VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MULT_Amp
  CLASS BLOCK ;
  FOREIGN MULT_Amp ;
  ORIGIN 0.000 0.050 ;
  SIZE 101.180 BY 158.870 ;
  PIN VDD
    ANTENNADIFFAREA 343.985596 ;
    PORT
      LAYER nwell ;
        RECT 18.615 111.070 81.715 138.270 ;
        RECT 29.340 84.755 70.390 90.960 ;
        RECT 31.140 84.750 69.230 84.755 ;
      LAYER li1 ;
        RECT 37.015 138.050 37.465 138.370 ;
        RECT 37.865 138.050 38.315 138.370 ;
        RECT 49.465 138.050 49.915 138.370 ;
        RECT 50.315 138.050 50.765 138.370 ;
        RECT 61.765 138.050 62.165 138.420 ;
        RECT 62.615 138.050 63.015 138.420 ;
        RECT 28.095 137.880 72.005 138.050 ;
        RECT 28.095 136.120 28.265 137.880 ;
        RECT 28.990 137.310 34.030 137.480 ;
        RECT 35.170 137.310 40.210 137.480 ;
        RECT 41.350 137.310 46.390 137.480 ;
        RECT 47.530 137.310 52.570 137.480 ;
        RECT 53.710 137.310 58.750 137.480 ;
        RECT 59.890 137.310 64.930 137.480 ;
        RECT 66.070 137.310 71.110 137.480 ;
        RECT 71.835 136.120 72.005 137.880 ;
        RECT 28.095 135.950 72.005 136.120 ;
        RECT 28.095 135.180 72.005 135.350 ;
        RECT 28.095 133.420 28.265 135.180 ;
        RECT 28.990 134.610 34.030 134.780 ;
        RECT 35.170 134.610 40.210 134.780 ;
        RECT 41.350 134.610 46.390 134.780 ;
        RECT 47.530 134.610 52.570 134.780 ;
        RECT 53.710 134.610 58.750 134.780 ;
        RECT 59.890 134.610 64.930 134.780 ;
        RECT 66.070 134.610 71.110 134.780 ;
        RECT 71.835 133.420 72.005 135.180 ;
        RECT 28.095 133.250 72.005 133.420 ;
        RECT 37.015 132.650 38.315 133.250 ;
        RECT 49.365 132.650 50.815 133.250 ;
        RECT 61.665 132.650 63.115 133.250 ;
        RECT 28.095 132.480 72.005 132.650 ;
        RECT 28.095 130.720 28.265 132.480 ;
        RECT 28.990 131.910 34.030 132.080 ;
        RECT 35.170 131.910 40.210 132.080 ;
        RECT 41.350 131.910 46.390 132.080 ;
        RECT 47.530 131.910 52.570 132.080 ;
        RECT 53.710 131.910 58.750 132.080 ;
        RECT 59.890 131.910 64.930 132.080 ;
        RECT 66.070 131.910 71.110 132.080 ;
        RECT 71.835 130.720 72.005 132.480 ;
        RECT 28.095 130.550 72.005 130.720 ;
        RECT 36.965 129.950 38.415 130.550 ;
        RECT 49.365 129.950 50.815 130.550 ;
        RECT 61.665 129.950 63.115 130.550 ;
        RECT 28.095 129.780 72.005 129.950 ;
        RECT 28.095 128.020 28.265 129.780 ;
        RECT 28.990 129.210 34.030 129.380 ;
        RECT 35.170 129.210 40.210 129.380 ;
        RECT 41.350 129.210 46.390 129.380 ;
        RECT 47.530 129.210 52.570 129.380 ;
        RECT 53.710 129.210 58.750 129.380 ;
        RECT 59.890 129.210 64.930 129.380 ;
        RECT 66.070 129.210 71.110 129.380 ;
        RECT 71.835 128.020 72.005 129.780 ;
        RECT 28.095 127.850 72.005 128.020 ;
        RECT 28.095 126.880 72.005 127.050 ;
        RECT 28.095 125.120 28.265 126.880 ;
        RECT 28.990 126.310 34.030 126.480 ;
        RECT 35.170 126.310 40.210 126.480 ;
        RECT 41.350 126.310 46.390 126.480 ;
        RECT 47.530 126.310 52.570 126.480 ;
        RECT 53.710 126.310 58.750 126.480 ;
        RECT 59.890 126.310 64.930 126.480 ;
        RECT 66.070 126.310 71.110 126.480 ;
        RECT 71.835 125.120 72.005 126.880 ;
        RECT 28.095 124.950 72.005 125.120 ;
        RECT 36.965 124.150 38.415 124.950 ;
        RECT 49.365 124.150 50.815 124.950 ;
        RECT 61.665 124.150 63.115 124.950 ;
        RECT 28.095 123.980 72.005 124.150 ;
        RECT 28.095 122.220 28.265 123.980 ;
        RECT 28.990 123.410 34.030 123.580 ;
        RECT 35.170 123.410 40.210 123.580 ;
        RECT 41.350 123.410 46.390 123.580 ;
        RECT 47.530 123.410 52.570 123.580 ;
        RECT 53.710 123.410 58.750 123.580 ;
        RECT 59.890 123.410 64.930 123.580 ;
        RECT 66.070 123.410 71.110 123.580 ;
        RECT 71.835 122.220 72.005 123.980 ;
        RECT 28.095 122.050 72.005 122.220 ;
        RECT 18.895 121.280 81.345 121.450 ;
        RECT 18.895 119.520 19.065 121.280 ;
        RECT 19.790 120.710 24.830 120.880 ;
        RECT 25.970 120.710 31.010 120.880 ;
        RECT 32.150 120.710 37.190 120.880 ;
        RECT 38.330 120.710 43.370 120.880 ;
        RECT 44.510 120.710 49.550 120.880 ;
        RECT 50.690 120.710 55.730 120.880 ;
        RECT 56.870 120.710 61.910 120.880 ;
        RECT 63.050 120.710 68.090 120.880 ;
        RECT 69.230 120.710 74.270 120.880 ;
        RECT 75.410 120.710 80.450 120.880 ;
        RECT 81.175 119.520 81.345 121.280 ;
        RECT 18.895 119.350 81.345 119.520 ;
        RECT 27.665 118.750 29.215 119.350 ;
        RECT 40.315 118.750 41.765 119.350 ;
        RECT 52.665 118.750 54.115 119.350 ;
        RECT 64.915 118.750 66.365 119.350 ;
        RECT 77.415 118.750 78.865 119.350 ;
        RECT 18.895 118.580 81.345 118.750 ;
        RECT 18.895 116.820 19.065 118.580 ;
        RECT 19.790 118.010 24.830 118.180 ;
        RECT 25.970 118.010 31.010 118.180 ;
        RECT 32.150 118.010 37.190 118.180 ;
        RECT 38.330 118.010 43.370 118.180 ;
        RECT 44.510 118.010 49.550 118.180 ;
        RECT 50.690 118.010 55.730 118.180 ;
        RECT 56.870 118.010 61.910 118.180 ;
        RECT 63.050 118.010 68.090 118.180 ;
        RECT 69.230 118.010 74.270 118.180 ;
        RECT 75.410 118.010 80.450 118.180 ;
        RECT 81.175 116.820 81.345 118.580 ;
        RECT 18.895 116.650 81.345 116.820 ;
        RECT 18.895 115.880 81.345 116.050 ;
        RECT 18.895 114.120 19.065 115.880 ;
        RECT 19.790 115.310 24.830 115.480 ;
        RECT 25.970 115.310 31.010 115.480 ;
        RECT 32.150 115.310 37.190 115.480 ;
        RECT 38.330 115.310 43.370 115.480 ;
        RECT 44.510 115.310 49.550 115.480 ;
        RECT 50.690 115.310 55.730 115.480 ;
        RECT 56.870 115.310 61.910 115.480 ;
        RECT 63.050 115.310 68.090 115.480 ;
        RECT 69.230 115.310 74.270 115.480 ;
        RECT 75.410 115.310 80.450 115.480 ;
        RECT 81.175 114.120 81.345 115.880 ;
        RECT 18.895 113.950 81.345 114.120 ;
        RECT 27.665 113.350 29.215 113.950 ;
        RECT 40.315 113.350 41.765 113.950 ;
        RECT 52.665 113.350 54.115 113.950 ;
        RECT 64.915 113.350 66.365 113.950 ;
        RECT 77.415 113.350 78.865 113.950 ;
        RECT 18.895 113.180 81.345 113.350 ;
        RECT 18.895 111.420 19.065 113.180 ;
        RECT 19.790 112.610 24.830 112.780 ;
        RECT 25.970 112.610 31.010 112.780 ;
        RECT 32.150 112.610 37.190 112.780 ;
        RECT 38.330 112.610 43.370 112.780 ;
        RECT 44.510 112.610 49.550 112.780 ;
        RECT 50.690 112.610 55.730 112.780 ;
        RECT 56.870 112.610 61.910 112.780 ;
        RECT 63.050 112.610 68.090 112.780 ;
        RECT 69.230 112.610 74.270 112.780 ;
        RECT 75.410 112.610 80.450 112.780 ;
        RECT 81.175 111.420 81.345 113.180 ;
        RECT 18.895 111.250 81.345 111.420 ;
        RECT 34.090 90.480 34.890 90.950 ;
        RECT 39.390 90.480 40.190 90.950 ;
        RECT 46.690 90.480 47.490 90.950 ;
        RECT 52.790 90.480 53.590 90.950 ;
        RECT 60.190 90.480 60.990 90.950 ;
        RECT 65.190 90.480 65.990 90.950 ;
        RECT 31.320 90.310 69.050 90.480 ;
        RECT 31.320 88.050 31.490 90.310 ;
        RECT 34.090 90.150 34.890 90.310 ;
        RECT 39.390 90.150 40.190 90.310 ;
        RECT 46.690 90.150 47.490 90.310 ;
        RECT 52.790 90.150 53.590 90.310 ;
        RECT 60.190 90.150 60.990 90.310 ;
        RECT 65.190 90.150 65.990 90.310 ;
        RECT 32.215 89.740 37.255 89.910 ;
        RECT 38.395 89.740 43.435 89.910 ;
        RECT 44.575 89.740 49.615 89.910 ;
        RECT 50.755 89.740 55.795 89.910 ;
        RECT 56.935 89.740 61.975 89.910 ;
        RECT 63.115 89.740 68.155 89.910 ;
        RECT 68.880 88.050 69.050 90.310 ;
        RECT 31.320 87.880 69.050 88.050 ;
        RECT 34.090 87.530 34.890 87.880 ;
        RECT 39.390 87.530 40.190 87.880 ;
        RECT 46.690 87.530 47.490 87.880 ;
        RECT 52.790 87.530 53.590 87.880 ;
        RECT 60.190 87.530 60.990 87.880 ;
        RECT 65.190 87.530 65.990 87.880 ;
        RECT 31.320 87.360 69.050 87.530 ;
        RECT 31.320 85.100 31.490 87.360 ;
        RECT 34.090 87.250 34.890 87.360 ;
        RECT 39.390 87.250 40.190 87.360 ;
        RECT 46.690 87.250 47.490 87.360 ;
        RECT 52.790 87.250 53.590 87.360 ;
        RECT 60.190 87.250 60.990 87.360 ;
        RECT 65.190 87.250 65.990 87.360 ;
        RECT 32.215 86.790 37.255 86.960 ;
        RECT 38.395 86.790 43.435 86.960 ;
        RECT 44.575 86.790 49.615 86.960 ;
        RECT 50.755 86.790 55.795 86.960 ;
        RECT 56.935 86.790 61.975 86.960 ;
        RECT 63.115 86.790 68.155 86.960 ;
        RECT 68.880 85.100 69.050 87.360 ;
        RECT 31.320 84.930 69.050 85.100 ;
      LAYER mcon ;
        RECT 37.155 138.110 37.325 138.280 ;
        RECT 38.005 138.110 38.175 138.280 ;
        RECT 49.605 138.110 49.775 138.280 ;
        RECT 50.455 138.110 50.625 138.280 ;
        RECT 61.880 138.135 62.050 138.305 ;
        RECT 62.730 138.135 62.900 138.305 ;
        RECT 29.085 137.310 29.255 137.480 ;
        RECT 29.445 137.310 29.615 137.480 ;
        RECT 29.805 137.310 29.975 137.480 ;
        RECT 30.165 137.310 30.335 137.480 ;
        RECT 30.525 137.310 30.695 137.480 ;
        RECT 30.885 137.310 31.055 137.480 ;
        RECT 31.245 137.310 31.415 137.480 ;
        RECT 31.605 137.310 31.775 137.480 ;
        RECT 31.965 137.310 32.135 137.480 ;
        RECT 32.325 137.310 32.495 137.480 ;
        RECT 32.685 137.310 32.855 137.480 ;
        RECT 33.045 137.310 33.215 137.480 ;
        RECT 33.405 137.310 33.575 137.480 ;
        RECT 33.765 137.310 33.935 137.480 ;
        RECT 35.265 137.310 35.435 137.480 ;
        RECT 35.625 137.310 35.795 137.480 ;
        RECT 35.985 137.310 36.155 137.480 ;
        RECT 36.345 137.310 36.515 137.480 ;
        RECT 36.705 137.310 36.875 137.480 ;
        RECT 37.065 137.310 37.235 137.480 ;
        RECT 37.425 137.310 37.595 137.480 ;
        RECT 37.785 137.310 37.955 137.480 ;
        RECT 38.145 137.310 38.315 137.480 ;
        RECT 38.505 137.310 38.675 137.480 ;
        RECT 38.865 137.310 39.035 137.480 ;
        RECT 39.225 137.310 39.395 137.480 ;
        RECT 39.585 137.310 39.755 137.480 ;
        RECT 39.945 137.310 40.115 137.480 ;
        RECT 41.445 137.310 41.615 137.480 ;
        RECT 41.805 137.310 41.975 137.480 ;
        RECT 42.165 137.310 42.335 137.480 ;
        RECT 42.525 137.310 42.695 137.480 ;
        RECT 42.885 137.310 43.055 137.480 ;
        RECT 43.245 137.310 43.415 137.480 ;
        RECT 43.605 137.310 43.775 137.480 ;
        RECT 43.965 137.310 44.135 137.480 ;
        RECT 44.325 137.310 44.495 137.480 ;
        RECT 44.685 137.310 44.855 137.480 ;
        RECT 45.045 137.310 45.215 137.480 ;
        RECT 45.405 137.310 45.575 137.480 ;
        RECT 45.765 137.310 45.935 137.480 ;
        RECT 46.125 137.310 46.295 137.480 ;
        RECT 47.625 137.310 47.795 137.480 ;
        RECT 47.985 137.310 48.155 137.480 ;
        RECT 48.345 137.310 48.515 137.480 ;
        RECT 48.705 137.310 48.875 137.480 ;
        RECT 49.065 137.310 49.235 137.480 ;
        RECT 49.425 137.310 49.595 137.480 ;
        RECT 49.785 137.310 49.955 137.480 ;
        RECT 50.145 137.310 50.315 137.480 ;
        RECT 50.505 137.310 50.675 137.480 ;
        RECT 50.865 137.310 51.035 137.480 ;
        RECT 51.225 137.310 51.395 137.480 ;
        RECT 51.585 137.310 51.755 137.480 ;
        RECT 51.945 137.310 52.115 137.480 ;
        RECT 52.305 137.310 52.475 137.480 ;
        RECT 53.805 137.310 53.975 137.480 ;
        RECT 54.165 137.310 54.335 137.480 ;
        RECT 54.525 137.310 54.695 137.480 ;
        RECT 54.885 137.310 55.055 137.480 ;
        RECT 55.245 137.310 55.415 137.480 ;
        RECT 55.605 137.310 55.775 137.480 ;
        RECT 55.965 137.310 56.135 137.480 ;
        RECT 56.325 137.310 56.495 137.480 ;
        RECT 56.685 137.310 56.855 137.480 ;
        RECT 57.045 137.310 57.215 137.480 ;
        RECT 57.405 137.310 57.575 137.480 ;
        RECT 57.765 137.310 57.935 137.480 ;
        RECT 58.125 137.310 58.295 137.480 ;
        RECT 58.485 137.310 58.655 137.480 ;
        RECT 59.985 137.310 60.155 137.480 ;
        RECT 60.345 137.310 60.515 137.480 ;
        RECT 60.705 137.310 60.875 137.480 ;
        RECT 61.065 137.310 61.235 137.480 ;
        RECT 61.425 137.310 61.595 137.480 ;
        RECT 61.785 137.310 61.955 137.480 ;
        RECT 62.145 137.310 62.315 137.480 ;
        RECT 62.505 137.310 62.675 137.480 ;
        RECT 62.865 137.310 63.035 137.480 ;
        RECT 63.225 137.310 63.395 137.480 ;
        RECT 63.585 137.310 63.755 137.480 ;
        RECT 63.945 137.310 64.115 137.480 ;
        RECT 64.305 137.310 64.475 137.480 ;
        RECT 64.665 137.310 64.835 137.480 ;
        RECT 66.165 137.310 66.335 137.480 ;
        RECT 66.525 137.310 66.695 137.480 ;
        RECT 66.885 137.310 67.055 137.480 ;
        RECT 67.245 137.310 67.415 137.480 ;
        RECT 67.605 137.310 67.775 137.480 ;
        RECT 67.965 137.310 68.135 137.480 ;
        RECT 68.325 137.310 68.495 137.480 ;
        RECT 68.685 137.310 68.855 137.480 ;
        RECT 69.045 137.310 69.215 137.480 ;
        RECT 69.405 137.310 69.575 137.480 ;
        RECT 69.765 137.310 69.935 137.480 ;
        RECT 70.125 137.310 70.295 137.480 ;
        RECT 70.485 137.310 70.655 137.480 ;
        RECT 70.845 137.310 71.015 137.480 ;
        RECT 29.085 134.610 29.255 134.780 ;
        RECT 29.445 134.610 29.615 134.780 ;
        RECT 29.805 134.610 29.975 134.780 ;
        RECT 30.165 134.610 30.335 134.780 ;
        RECT 30.525 134.610 30.695 134.780 ;
        RECT 30.885 134.610 31.055 134.780 ;
        RECT 31.245 134.610 31.415 134.780 ;
        RECT 31.605 134.610 31.775 134.780 ;
        RECT 31.965 134.610 32.135 134.780 ;
        RECT 32.325 134.610 32.495 134.780 ;
        RECT 32.685 134.610 32.855 134.780 ;
        RECT 33.045 134.610 33.215 134.780 ;
        RECT 33.405 134.610 33.575 134.780 ;
        RECT 33.765 134.610 33.935 134.780 ;
        RECT 35.265 134.610 35.435 134.780 ;
        RECT 35.625 134.610 35.795 134.780 ;
        RECT 35.985 134.610 36.155 134.780 ;
        RECT 36.345 134.610 36.515 134.780 ;
        RECT 36.705 134.610 36.875 134.780 ;
        RECT 37.065 134.610 37.235 134.780 ;
        RECT 37.425 134.610 37.595 134.780 ;
        RECT 37.785 134.610 37.955 134.780 ;
        RECT 38.145 134.610 38.315 134.780 ;
        RECT 38.505 134.610 38.675 134.780 ;
        RECT 38.865 134.610 39.035 134.780 ;
        RECT 39.225 134.610 39.395 134.780 ;
        RECT 39.585 134.610 39.755 134.780 ;
        RECT 39.945 134.610 40.115 134.780 ;
        RECT 41.445 134.610 41.615 134.780 ;
        RECT 41.805 134.610 41.975 134.780 ;
        RECT 42.165 134.610 42.335 134.780 ;
        RECT 42.525 134.610 42.695 134.780 ;
        RECT 42.885 134.610 43.055 134.780 ;
        RECT 43.245 134.610 43.415 134.780 ;
        RECT 43.605 134.610 43.775 134.780 ;
        RECT 43.965 134.610 44.135 134.780 ;
        RECT 44.325 134.610 44.495 134.780 ;
        RECT 44.685 134.610 44.855 134.780 ;
        RECT 45.045 134.610 45.215 134.780 ;
        RECT 45.405 134.610 45.575 134.780 ;
        RECT 45.765 134.610 45.935 134.780 ;
        RECT 46.125 134.610 46.295 134.780 ;
        RECT 47.625 134.610 47.795 134.780 ;
        RECT 47.985 134.610 48.155 134.780 ;
        RECT 48.345 134.610 48.515 134.780 ;
        RECT 48.705 134.610 48.875 134.780 ;
        RECT 49.065 134.610 49.235 134.780 ;
        RECT 49.425 134.610 49.595 134.780 ;
        RECT 49.785 134.610 49.955 134.780 ;
        RECT 50.145 134.610 50.315 134.780 ;
        RECT 50.505 134.610 50.675 134.780 ;
        RECT 50.865 134.610 51.035 134.780 ;
        RECT 51.225 134.610 51.395 134.780 ;
        RECT 51.585 134.610 51.755 134.780 ;
        RECT 51.945 134.610 52.115 134.780 ;
        RECT 52.305 134.610 52.475 134.780 ;
        RECT 53.805 134.610 53.975 134.780 ;
        RECT 54.165 134.610 54.335 134.780 ;
        RECT 54.525 134.610 54.695 134.780 ;
        RECT 54.885 134.610 55.055 134.780 ;
        RECT 55.245 134.610 55.415 134.780 ;
        RECT 55.605 134.610 55.775 134.780 ;
        RECT 55.965 134.610 56.135 134.780 ;
        RECT 56.325 134.610 56.495 134.780 ;
        RECT 56.685 134.610 56.855 134.780 ;
        RECT 57.045 134.610 57.215 134.780 ;
        RECT 57.405 134.610 57.575 134.780 ;
        RECT 57.765 134.610 57.935 134.780 ;
        RECT 58.125 134.610 58.295 134.780 ;
        RECT 58.485 134.610 58.655 134.780 ;
        RECT 59.985 134.610 60.155 134.780 ;
        RECT 60.345 134.610 60.515 134.780 ;
        RECT 60.705 134.610 60.875 134.780 ;
        RECT 61.065 134.610 61.235 134.780 ;
        RECT 61.425 134.610 61.595 134.780 ;
        RECT 61.785 134.610 61.955 134.780 ;
        RECT 62.145 134.610 62.315 134.780 ;
        RECT 62.505 134.610 62.675 134.780 ;
        RECT 62.865 134.610 63.035 134.780 ;
        RECT 63.225 134.610 63.395 134.780 ;
        RECT 63.585 134.610 63.755 134.780 ;
        RECT 63.945 134.610 64.115 134.780 ;
        RECT 64.305 134.610 64.475 134.780 ;
        RECT 64.665 134.610 64.835 134.780 ;
        RECT 66.165 134.610 66.335 134.780 ;
        RECT 66.525 134.610 66.695 134.780 ;
        RECT 66.885 134.610 67.055 134.780 ;
        RECT 67.245 134.610 67.415 134.780 ;
        RECT 67.605 134.610 67.775 134.780 ;
        RECT 67.965 134.610 68.135 134.780 ;
        RECT 68.325 134.610 68.495 134.780 ;
        RECT 68.685 134.610 68.855 134.780 ;
        RECT 69.045 134.610 69.215 134.780 ;
        RECT 69.405 134.610 69.575 134.780 ;
        RECT 69.765 134.610 69.935 134.780 ;
        RECT 70.125 134.610 70.295 134.780 ;
        RECT 70.485 134.610 70.655 134.780 ;
        RECT 70.845 134.610 71.015 134.780 ;
        RECT 37.205 132.860 37.375 133.030 ;
        RECT 37.905 132.860 38.075 133.030 ;
        RECT 49.605 132.860 49.775 133.030 ;
        RECT 50.405 132.910 50.575 133.080 ;
        RECT 61.880 132.910 62.050 133.080 ;
        RECT 62.730 132.910 62.900 133.080 ;
        RECT 29.085 131.910 29.255 132.080 ;
        RECT 29.445 131.910 29.615 132.080 ;
        RECT 29.805 131.910 29.975 132.080 ;
        RECT 30.165 131.910 30.335 132.080 ;
        RECT 30.525 131.910 30.695 132.080 ;
        RECT 30.885 131.910 31.055 132.080 ;
        RECT 31.245 131.910 31.415 132.080 ;
        RECT 31.605 131.910 31.775 132.080 ;
        RECT 31.965 131.910 32.135 132.080 ;
        RECT 32.325 131.910 32.495 132.080 ;
        RECT 32.685 131.910 32.855 132.080 ;
        RECT 33.045 131.910 33.215 132.080 ;
        RECT 33.405 131.910 33.575 132.080 ;
        RECT 33.765 131.910 33.935 132.080 ;
        RECT 35.265 131.910 35.435 132.080 ;
        RECT 35.625 131.910 35.795 132.080 ;
        RECT 35.985 131.910 36.155 132.080 ;
        RECT 36.345 131.910 36.515 132.080 ;
        RECT 36.705 131.910 36.875 132.080 ;
        RECT 37.065 131.910 37.235 132.080 ;
        RECT 37.425 131.910 37.595 132.080 ;
        RECT 37.785 131.910 37.955 132.080 ;
        RECT 38.145 131.910 38.315 132.080 ;
        RECT 38.505 131.910 38.675 132.080 ;
        RECT 38.865 131.910 39.035 132.080 ;
        RECT 39.225 131.910 39.395 132.080 ;
        RECT 39.585 131.910 39.755 132.080 ;
        RECT 39.945 131.910 40.115 132.080 ;
        RECT 41.445 131.910 41.615 132.080 ;
        RECT 41.805 131.910 41.975 132.080 ;
        RECT 42.165 131.910 42.335 132.080 ;
        RECT 42.525 131.910 42.695 132.080 ;
        RECT 42.885 131.910 43.055 132.080 ;
        RECT 43.245 131.910 43.415 132.080 ;
        RECT 43.605 131.910 43.775 132.080 ;
        RECT 43.965 131.910 44.135 132.080 ;
        RECT 44.325 131.910 44.495 132.080 ;
        RECT 44.685 131.910 44.855 132.080 ;
        RECT 45.045 131.910 45.215 132.080 ;
        RECT 45.405 131.910 45.575 132.080 ;
        RECT 45.765 131.910 45.935 132.080 ;
        RECT 46.125 131.910 46.295 132.080 ;
        RECT 47.625 131.910 47.795 132.080 ;
        RECT 47.985 131.910 48.155 132.080 ;
        RECT 48.345 131.910 48.515 132.080 ;
        RECT 48.705 131.910 48.875 132.080 ;
        RECT 49.065 131.910 49.235 132.080 ;
        RECT 49.425 131.910 49.595 132.080 ;
        RECT 49.785 131.910 49.955 132.080 ;
        RECT 50.145 131.910 50.315 132.080 ;
        RECT 50.505 131.910 50.675 132.080 ;
        RECT 50.865 131.910 51.035 132.080 ;
        RECT 51.225 131.910 51.395 132.080 ;
        RECT 51.585 131.910 51.755 132.080 ;
        RECT 51.945 131.910 52.115 132.080 ;
        RECT 52.305 131.910 52.475 132.080 ;
        RECT 53.805 131.910 53.975 132.080 ;
        RECT 54.165 131.910 54.335 132.080 ;
        RECT 54.525 131.910 54.695 132.080 ;
        RECT 54.885 131.910 55.055 132.080 ;
        RECT 55.245 131.910 55.415 132.080 ;
        RECT 55.605 131.910 55.775 132.080 ;
        RECT 55.965 131.910 56.135 132.080 ;
        RECT 56.325 131.910 56.495 132.080 ;
        RECT 56.685 131.910 56.855 132.080 ;
        RECT 57.045 131.910 57.215 132.080 ;
        RECT 57.405 131.910 57.575 132.080 ;
        RECT 57.765 131.910 57.935 132.080 ;
        RECT 58.125 131.910 58.295 132.080 ;
        RECT 58.485 131.910 58.655 132.080 ;
        RECT 59.985 131.910 60.155 132.080 ;
        RECT 60.345 131.910 60.515 132.080 ;
        RECT 60.705 131.910 60.875 132.080 ;
        RECT 61.065 131.910 61.235 132.080 ;
        RECT 61.425 131.910 61.595 132.080 ;
        RECT 61.785 131.910 61.955 132.080 ;
        RECT 62.145 131.910 62.315 132.080 ;
        RECT 62.505 131.910 62.675 132.080 ;
        RECT 62.865 131.910 63.035 132.080 ;
        RECT 63.225 131.910 63.395 132.080 ;
        RECT 63.585 131.910 63.755 132.080 ;
        RECT 63.945 131.910 64.115 132.080 ;
        RECT 64.305 131.910 64.475 132.080 ;
        RECT 64.665 131.910 64.835 132.080 ;
        RECT 66.165 131.910 66.335 132.080 ;
        RECT 66.525 131.910 66.695 132.080 ;
        RECT 66.885 131.910 67.055 132.080 ;
        RECT 67.245 131.910 67.415 132.080 ;
        RECT 67.605 131.910 67.775 132.080 ;
        RECT 67.965 131.910 68.135 132.080 ;
        RECT 68.325 131.910 68.495 132.080 ;
        RECT 68.685 131.910 68.855 132.080 ;
        RECT 69.045 131.910 69.215 132.080 ;
        RECT 69.405 131.910 69.575 132.080 ;
        RECT 69.765 131.910 69.935 132.080 ;
        RECT 70.125 131.910 70.295 132.080 ;
        RECT 70.485 131.910 70.655 132.080 ;
        RECT 70.845 131.910 71.015 132.080 ;
        RECT 37.180 130.185 37.350 130.355 ;
        RECT 38.030 130.185 38.200 130.355 ;
        RECT 49.580 130.185 49.750 130.355 ;
        RECT 50.430 130.185 50.600 130.355 ;
        RECT 61.880 130.185 62.050 130.355 ;
        RECT 62.730 130.185 62.900 130.355 ;
        RECT 29.085 129.210 29.255 129.380 ;
        RECT 29.445 129.210 29.615 129.380 ;
        RECT 29.805 129.210 29.975 129.380 ;
        RECT 30.165 129.210 30.335 129.380 ;
        RECT 30.525 129.210 30.695 129.380 ;
        RECT 30.885 129.210 31.055 129.380 ;
        RECT 31.245 129.210 31.415 129.380 ;
        RECT 31.605 129.210 31.775 129.380 ;
        RECT 31.965 129.210 32.135 129.380 ;
        RECT 32.325 129.210 32.495 129.380 ;
        RECT 32.685 129.210 32.855 129.380 ;
        RECT 33.045 129.210 33.215 129.380 ;
        RECT 33.405 129.210 33.575 129.380 ;
        RECT 33.765 129.210 33.935 129.380 ;
        RECT 35.265 129.210 35.435 129.380 ;
        RECT 35.625 129.210 35.795 129.380 ;
        RECT 35.985 129.210 36.155 129.380 ;
        RECT 36.345 129.210 36.515 129.380 ;
        RECT 36.705 129.210 36.875 129.380 ;
        RECT 37.065 129.210 37.235 129.380 ;
        RECT 37.425 129.210 37.595 129.380 ;
        RECT 37.785 129.210 37.955 129.380 ;
        RECT 38.145 129.210 38.315 129.380 ;
        RECT 38.505 129.210 38.675 129.380 ;
        RECT 38.865 129.210 39.035 129.380 ;
        RECT 39.225 129.210 39.395 129.380 ;
        RECT 39.585 129.210 39.755 129.380 ;
        RECT 39.945 129.210 40.115 129.380 ;
        RECT 41.445 129.210 41.615 129.380 ;
        RECT 41.805 129.210 41.975 129.380 ;
        RECT 42.165 129.210 42.335 129.380 ;
        RECT 42.525 129.210 42.695 129.380 ;
        RECT 42.885 129.210 43.055 129.380 ;
        RECT 43.245 129.210 43.415 129.380 ;
        RECT 43.605 129.210 43.775 129.380 ;
        RECT 43.965 129.210 44.135 129.380 ;
        RECT 44.325 129.210 44.495 129.380 ;
        RECT 44.685 129.210 44.855 129.380 ;
        RECT 45.045 129.210 45.215 129.380 ;
        RECT 45.405 129.210 45.575 129.380 ;
        RECT 45.765 129.210 45.935 129.380 ;
        RECT 46.125 129.210 46.295 129.380 ;
        RECT 47.625 129.210 47.795 129.380 ;
        RECT 47.985 129.210 48.155 129.380 ;
        RECT 48.345 129.210 48.515 129.380 ;
        RECT 48.705 129.210 48.875 129.380 ;
        RECT 49.065 129.210 49.235 129.380 ;
        RECT 49.425 129.210 49.595 129.380 ;
        RECT 49.785 129.210 49.955 129.380 ;
        RECT 50.145 129.210 50.315 129.380 ;
        RECT 50.505 129.210 50.675 129.380 ;
        RECT 50.865 129.210 51.035 129.380 ;
        RECT 51.225 129.210 51.395 129.380 ;
        RECT 51.585 129.210 51.755 129.380 ;
        RECT 51.945 129.210 52.115 129.380 ;
        RECT 52.305 129.210 52.475 129.380 ;
        RECT 53.805 129.210 53.975 129.380 ;
        RECT 54.165 129.210 54.335 129.380 ;
        RECT 54.525 129.210 54.695 129.380 ;
        RECT 54.885 129.210 55.055 129.380 ;
        RECT 55.245 129.210 55.415 129.380 ;
        RECT 55.605 129.210 55.775 129.380 ;
        RECT 55.965 129.210 56.135 129.380 ;
        RECT 56.325 129.210 56.495 129.380 ;
        RECT 56.685 129.210 56.855 129.380 ;
        RECT 57.045 129.210 57.215 129.380 ;
        RECT 57.405 129.210 57.575 129.380 ;
        RECT 57.765 129.210 57.935 129.380 ;
        RECT 58.125 129.210 58.295 129.380 ;
        RECT 58.485 129.210 58.655 129.380 ;
        RECT 59.985 129.210 60.155 129.380 ;
        RECT 60.345 129.210 60.515 129.380 ;
        RECT 60.705 129.210 60.875 129.380 ;
        RECT 61.065 129.210 61.235 129.380 ;
        RECT 61.425 129.210 61.595 129.380 ;
        RECT 61.785 129.210 61.955 129.380 ;
        RECT 62.145 129.210 62.315 129.380 ;
        RECT 62.505 129.210 62.675 129.380 ;
        RECT 62.865 129.210 63.035 129.380 ;
        RECT 63.225 129.210 63.395 129.380 ;
        RECT 63.585 129.210 63.755 129.380 ;
        RECT 63.945 129.210 64.115 129.380 ;
        RECT 64.305 129.210 64.475 129.380 ;
        RECT 64.665 129.210 64.835 129.380 ;
        RECT 66.165 129.210 66.335 129.380 ;
        RECT 66.525 129.210 66.695 129.380 ;
        RECT 66.885 129.210 67.055 129.380 ;
        RECT 67.245 129.210 67.415 129.380 ;
        RECT 67.605 129.210 67.775 129.380 ;
        RECT 67.965 129.210 68.135 129.380 ;
        RECT 68.325 129.210 68.495 129.380 ;
        RECT 68.685 129.210 68.855 129.380 ;
        RECT 69.045 129.210 69.215 129.380 ;
        RECT 69.405 129.210 69.575 129.380 ;
        RECT 69.765 129.210 69.935 129.380 ;
        RECT 70.125 129.210 70.295 129.380 ;
        RECT 70.485 129.210 70.655 129.380 ;
        RECT 70.845 129.210 71.015 129.380 ;
        RECT 29.085 126.310 29.255 126.480 ;
        RECT 29.445 126.310 29.615 126.480 ;
        RECT 29.805 126.310 29.975 126.480 ;
        RECT 30.165 126.310 30.335 126.480 ;
        RECT 30.525 126.310 30.695 126.480 ;
        RECT 30.885 126.310 31.055 126.480 ;
        RECT 31.245 126.310 31.415 126.480 ;
        RECT 31.605 126.310 31.775 126.480 ;
        RECT 31.965 126.310 32.135 126.480 ;
        RECT 32.325 126.310 32.495 126.480 ;
        RECT 32.685 126.310 32.855 126.480 ;
        RECT 33.045 126.310 33.215 126.480 ;
        RECT 33.405 126.310 33.575 126.480 ;
        RECT 33.765 126.310 33.935 126.480 ;
        RECT 35.265 126.310 35.435 126.480 ;
        RECT 35.625 126.310 35.795 126.480 ;
        RECT 35.985 126.310 36.155 126.480 ;
        RECT 36.345 126.310 36.515 126.480 ;
        RECT 36.705 126.310 36.875 126.480 ;
        RECT 37.065 126.310 37.235 126.480 ;
        RECT 37.425 126.310 37.595 126.480 ;
        RECT 37.785 126.310 37.955 126.480 ;
        RECT 38.145 126.310 38.315 126.480 ;
        RECT 38.505 126.310 38.675 126.480 ;
        RECT 38.865 126.310 39.035 126.480 ;
        RECT 39.225 126.310 39.395 126.480 ;
        RECT 39.585 126.310 39.755 126.480 ;
        RECT 39.945 126.310 40.115 126.480 ;
        RECT 41.445 126.310 41.615 126.480 ;
        RECT 41.805 126.310 41.975 126.480 ;
        RECT 42.165 126.310 42.335 126.480 ;
        RECT 42.525 126.310 42.695 126.480 ;
        RECT 42.885 126.310 43.055 126.480 ;
        RECT 43.245 126.310 43.415 126.480 ;
        RECT 43.605 126.310 43.775 126.480 ;
        RECT 43.965 126.310 44.135 126.480 ;
        RECT 44.325 126.310 44.495 126.480 ;
        RECT 44.685 126.310 44.855 126.480 ;
        RECT 45.045 126.310 45.215 126.480 ;
        RECT 45.405 126.310 45.575 126.480 ;
        RECT 45.765 126.310 45.935 126.480 ;
        RECT 46.125 126.310 46.295 126.480 ;
        RECT 47.625 126.310 47.795 126.480 ;
        RECT 47.985 126.310 48.155 126.480 ;
        RECT 48.345 126.310 48.515 126.480 ;
        RECT 48.705 126.310 48.875 126.480 ;
        RECT 49.065 126.310 49.235 126.480 ;
        RECT 49.425 126.310 49.595 126.480 ;
        RECT 49.785 126.310 49.955 126.480 ;
        RECT 50.145 126.310 50.315 126.480 ;
        RECT 50.505 126.310 50.675 126.480 ;
        RECT 50.865 126.310 51.035 126.480 ;
        RECT 51.225 126.310 51.395 126.480 ;
        RECT 51.585 126.310 51.755 126.480 ;
        RECT 51.945 126.310 52.115 126.480 ;
        RECT 52.305 126.310 52.475 126.480 ;
        RECT 53.805 126.310 53.975 126.480 ;
        RECT 54.165 126.310 54.335 126.480 ;
        RECT 54.525 126.310 54.695 126.480 ;
        RECT 54.885 126.310 55.055 126.480 ;
        RECT 55.245 126.310 55.415 126.480 ;
        RECT 55.605 126.310 55.775 126.480 ;
        RECT 55.965 126.310 56.135 126.480 ;
        RECT 56.325 126.310 56.495 126.480 ;
        RECT 56.685 126.310 56.855 126.480 ;
        RECT 57.045 126.310 57.215 126.480 ;
        RECT 57.405 126.310 57.575 126.480 ;
        RECT 57.765 126.310 57.935 126.480 ;
        RECT 58.125 126.310 58.295 126.480 ;
        RECT 58.485 126.310 58.655 126.480 ;
        RECT 59.985 126.310 60.155 126.480 ;
        RECT 60.345 126.310 60.515 126.480 ;
        RECT 60.705 126.310 60.875 126.480 ;
        RECT 61.065 126.310 61.235 126.480 ;
        RECT 61.425 126.310 61.595 126.480 ;
        RECT 61.785 126.310 61.955 126.480 ;
        RECT 62.145 126.310 62.315 126.480 ;
        RECT 62.505 126.310 62.675 126.480 ;
        RECT 62.865 126.310 63.035 126.480 ;
        RECT 63.225 126.310 63.395 126.480 ;
        RECT 63.585 126.310 63.755 126.480 ;
        RECT 63.945 126.310 64.115 126.480 ;
        RECT 64.305 126.310 64.475 126.480 ;
        RECT 64.665 126.310 64.835 126.480 ;
        RECT 66.165 126.310 66.335 126.480 ;
        RECT 66.525 126.310 66.695 126.480 ;
        RECT 66.885 126.310 67.055 126.480 ;
        RECT 67.245 126.310 67.415 126.480 ;
        RECT 67.605 126.310 67.775 126.480 ;
        RECT 67.965 126.310 68.135 126.480 ;
        RECT 68.325 126.310 68.495 126.480 ;
        RECT 68.685 126.310 68.855 126.480 ;
        RECT 69.045 126.310 69.215 126.480 ;
        RECT 69.405 126.310 69.575 126.480 ;
        RECT 69.765 126.310 69.935 126.480 ;
        RECT 70.125 126.310 70.295 126.480 ;
        RECT 70.485 126.310 70.655 126.480 ;
        RECT 70.845 126.310 71.015 126.480 ;
        RECT 37.205 124.385 37.375 124.555 ;
        RECT 38.005 124.385 38.175 124.555 ;
        RECT 49.580 124.360 49.750 124.530 ;
        RECT 50.430 124.360 50.600 124.530 ;
        RECT 61.880 124.360 62.050 124.530 ;
        RECT 62.730 124.360 62.900 124.530 ;
        RECT 29.085 123.410 29.255 123.580 ;
        RECT 29.445 123.410 29.615 123.580 ;
        RECT 29.805 123.410 29.975 123.580 ;
        RECT 30.165 123.410 30.335 123.580 ;
        RECT 30.525 123.410 30.695 123.580 ;
        RECT 30.885 123.410 31.055 123.580 ;
        RECT 31.245 123.410 31.415 123.580 ;
        RECT 31.605 123.410 31.775 123.580 ;
        RECT 31.965 123.410 32.135 123.580 ;
        RECT 32.325 123.410 32.495 123.580 ;
        RECT 32.685 123.410 32.855 123.580 ;
        RECT 33.045 123.410 33.215 123.580 ;
        RECT 33.405 123.410 33.575 123.580 ;
        RECT 33.765 123.410 33.935 123.580 ;
        RECT 35.265 123.410 35.435 123.580 ;
        RECT 35.625 123.410 35.795 123.580 ;
        RECT 35.985 123.410 36.155 123.580 ;
        RECT 36.345 123.410 36.515 123.580 ;
        RECT 36.705 123.410 36.875 123.580 ;
        RECT 37.065 123.410 37.235 123.580 ;
        RECT 37.425 123.410 37.595 123.580 ;
        RECT 37.785 123.410 37.955 123.580 ;
        RECT 38.145 123.410 38.315 123.580 ;
        RECT 38.505 123.410 38.675 123.580 ;
        RECT 38.865 123.410 39.035 123.580 ;
        RECT 39.225 123.410 39.395 123.580 ;
        RECT 39.585 123.410 39.755 123.580 ;
        RECT 39.945 123.410 40.115 123.580 ;
        RECT 41.445 123.410 41.615 123.580 ;
        RECT 41.805 123.410 41.975 123.580 ;
        RECT 42.165 123.410 42.335 123.580 ;
        RECT 42.525 123.410 42.695 123.580 ;
        RECT 42.885 123.410 43.055 123.580 ;
        RECT 43.245 123.410 43.415 123.580 ;
        RECT 43.605 123.410 43.775 123.580 ;
        RECT 43.965 123.410 44.135 123.580 ;
        RECT 44.325 123.410 44.495 123.580 ;
        RECT 44.685 123.410 44.855 123.580 ;
        RECT 45.045 123.410 45.215 123.580 ;
        RECT 45.405 123.410 45.575 123.580 ;
        RECT 45.765 123.410 45.935 123.580 ;
        RECT 46.125 123.410 46.295 123.580 ;
        RECT 47.625 123.410 47.795 123.580 ;
        RECT 47.985 123.410 48.155 123.580 ;
        RECT 48.345 123.410 48.515 123.580 ;
        RECT 48.705 123.410 48.875 123.580 ;
        RECT 49.065 123.410 49.235 123.580 ;
        RECT 49.425 123.410 49.595 123.580 ;
        RECT 49.785 123.410 49.955 123.580 ;
        RECT 50.145 123.410 50.315 123.580 ;
        RECT 50.505 123.410 50.675 123.580 ;
        RECT 50.865 123.410 51.035 123.580 ;
        RECT 51.225 123.410 51.395 123.580 ;
        RECT 51.585 123.410 51.755 123.580 ;
        RECT 51.945 123.410 52.115 123.580 ;
        RECT 52.305 123.410 52.475 123.580 ;
        RECT 53.805 123.410 53.975 123.580 ;
        RECT 54.165 123.410 54.335 123.580 ;
        RECT 54.525 123.410 54.695 123.580 ;
        RECT 54.885 123.410 55.055 123.580 ;
        RECT 55.245 123.410 55.415 123.580 ;
        RECT 55.605 123.410 55.775 123.580 ;
        RECT 55.965 123.410 56.135 123.580 ;
        RECT 56.325 123.410 56.495 123.580 ;
        RECT 56.685 123.410 56.855 123.580 ;
        RECT 57.045 123.410 57.215 123.580 ;
        RECT 57.405 123.410 57.575 123.580 ;
        RECT 57.765 123.410 57.935 123.580 ;
        RECT 58.125 123.410 58.295 123.580 ;
        RECT 58.485 123.410 58.655 123.580 ;
        RECT 59.985 123.410 60.155 123.580 ;
        RECT 60.345 123.410 60.515 123.580 ;
        RECT 60.705 123.410 60.875 123.580 ;
        RECT 61.065 123.410 61.235 123.580 ;
        RECT 61.425 123.410 61.595 123.580 ;
        RECT 61.785 123.410 61.955 123.580 ;
        RECT 62.145 123.410 62.315 123.580 ;
        RECT 62.505 123.410 62.675 123.580 ;
        RECT 62.865 123.410 63.035 123.580 ;
        RECT 63.225 123.410 63.395 123.580 ;
        RECT 63.585 123.410 63.755 123.580 ;
        RECT 63.945 123.410 64.115 123.580 ;
        RECT 64.305 123.410 64.475 123.580 ;
        RECT 64.665 123.410 64.835 123.580 ;
        RECT 66.165 123.410 66.335 123.580 ;
        RECT 66.525 123.410 66.695 123.580 ;
        RECT 66.885 123.410 67.055 123.580 ;
        RECT 67.245 123.410 67.415 123.580 ;
        RECT 67.605 123.410 67.775 123.580 ;
        RECT 67.965 123.410 68.135 123.580 ;
        RECT 68.325 123.410 68.495 123.580 ;
        RECT 68.685 123.410 68.855 123.580 ;
        RECT 69.045 123.410 69.215 123.580 ;
        RECT 69.405 123.410 69.575 123.580 ;
        RECT 69.765 123.410 69.935 123.580 ;
        RECT 70.125 123.410 70.295 123.580 ;
        RECT 70.485 123.410 70.655 123.580 ;
        RECT 70.845 123.410 71.015 123.580 ;
        RECT 19.885 120.710 20.055 120.880 ;
        RECT 20.245 120.710 20.415 120.880 ;
        RECT 20.605 120.710 20.775 120.880 ;
        RECT 20.965 120.710 21.135 120.880 ;
        RECT 21.325 120.710 21.495 120.880 ;
        RECT 21.685 120.710 21.855 120.880 ;
        RECT 22.045 120.710 22.215 120.880 ;
        RECT 22.405 120.710 22.575 120.880 ;
        RECT 22.765 120.710 22.935 120.880 ;
        RECT 23.125 120.710 23.295 120.880 ;
        RECT 23.485 120.710 23.655 120.880 ;
        RECT 23.845 120.710 24.015 120.880 ;
        RECT 24.205 120.710 24.375 120.880 ;
        RECT 24.565 120.710 24.735 120.880 ;
        RECT 26.065 120.710 26.235 120.880 ;
        RECT 26.425 120.710 26.595 120.880 ;
        RECT 26.785 120.710 26.955 120.880 ;
        RECT 27.145 120.710 27.315 120.880 ;
        RECT 27.505 120.710 27.675 120.880 ;
        RECT 27.865 120.710 28.035 120.880 ;
        RECT 28.225 120.710 28.395 120.880 ;
        RECT 28.585 120.710 28.755 120.880 ;
        RECT 28.945 120.710 29.115 120.880 ;
        RECT 29.305 120.710 29.475 120.880 ;
        RECT 29.665 120.710 29.835 120.880 ;
        RECT 30.025 120.710 30.195 120.880 ;
        RECT 30.385 120.710 30.555 120.880 ;
        RECT 30.745 120.710 30.915 120.880 ;
        RECT 32.245 120.710 32.415 120.880 ;
        RECT 32.605 120.710 32.775 120.880 ;
        RECT 32.965 120.710 33.135 120.880 ;
        RECT 33.325 120.710 33.495 120.880 ;
        RECT 33.685 120.710 33.855 120.880 ;
        RECT 34.045 120.710 34.215 120.880 ;
        RECT 34.405 120.710 34.575 120.880 ;
        RECT 34.765 120.710 34.935 120.880 ;
        RECT 35.125 120.710 35.295 120.880 ;
        RECT 35.485 120.710 35.655 120.880 ;
        RECT 35.845 120.710 36.015 120.880 ;
        RECT 36.205 120.710 36.375 120.880 ;
        RECT 36.565 120.710 36.735 120.880 ;
        RECT 36.925 120.710 37.095 120.880 ;
        RECT 38.425 120.710 38.595 120.880 ;
        RECT 38.785 120.710 38.955 120.880 ;
        RECT 39.145 120.710 39.315 120.880 ;
        RECT 39.505 120.710 39.675 120.880 ;
        RECT 39.865 120.710 40.035 120.880 ;
        RECT 40.225 120.710 40.395 120.880 ;
        RECT 40.585 120.710 40.755 120.880 ;
        RECT 40.945 120.710 41.115 120.880 ;
        RECT 41.305 120.710 41.475 120.880 ;
        RECT 41.665 120.710 41.835 120.880 ;
        RECT 42.025 120.710 42.195 120.880 ;
        RECT 42.385 120.710 42.555 120.880 ;
        RECT 42.745 120.710 42.915 120.880 ;
        RECT 43.105 120.710 43.275 120.880 ;
        RECT 44.605 120.710 44.775 120.880 ;
        RECT 44.965 120.710 45.135 120.880 ;
        RECT 45.325 120.710 45.495 120.880 ;
        RECT 45.685 120.710 45.855 120.880 ;
        RECT 46.045 120.710 46.215 120.880 ;
        RECT 46.405 120.710 46.575 120.880 ;
        RECT 46.765 120.710 46.935 120.880 ;
        RECT 47.125 120.710 47.295 120.880 ;
        RECT 47.485 120.710 47.655 120.880 ;
        RECT 47.845 120.710 48.015 120.880 ;
        RECT 48.205 120.710 48.375 120.880 ;
        RECT 48.565 120.710 48.735 120.880 ;
        RECT 48.925 120.710 49.095 120.880 ;
        RECT 49.285 120.710 49.455 120.880 ;
        RECT 50.785 120.710 50.955 120.880 ;
        RECT 51.145 120.710 51.315 120.880 ;
        RECT 51.505 120.710 51.675 120.880 ;
        RECT 51.865 120.710 52.035 120.880 ;
        RECT 52.225 120.710 52.395 120.880 ;
        RECT 52.585 120.710 52.755 120.880 ;
        RECT 52.945 120.710 53.115 120.880 ;
        RECT 53.305 120.710 53.475 120.880 ;
        RECT 53.665 120.710 53.835 120.880 ;
        RECT 54.025 120.710 54.195 120.880 ;
        RECT 54.385 120.710 54.555 120.880 ;
        RECT 54.745 120.710 54.915 120.880 ;
        RECT 55.105 120.710 55.275 120.880 ;
        RECT 55.465 120.710 55.635 120.880 ;
        RECT 56.965 120.710 57.135 120.880 ;
        RECT 57.325 120.710 57.495 120.880 ;
        RECT 57.685 120.710 57.855 120.880 ;
        RECT 58.045 120.710 58.215 120.880 ;
        RECT 58.405 120.710 58.575 120.880 ;
        RECT 58.765 120.710 58.935 120.880 ;
        RECT 59.125 120.710 59.295 120.880 ;
        RECT 59.485 120.710 59.655 120.880 ;
        RECT 59.845 120.710 60.015 120.880 ;
        RECT 60.205 120.710 60.375 120.880 ;
        RECT 60.565 120.710 60.735 120.880 ;
        RECT 60.925 120.710 61.095 120.880 ;
        RECT 61.285 120.710 61.455 120.880 ;
        RECT 61.645 120.710 61.815 120.880 ;
        RECT 63.145 120.710 63.315 120.880 ;
        RECT 63.505 120.710 63.675 120.880 ;
        RECT 63.865 120.710 64.035 120.880 ;
        RECT 64.225 120.710 64.395 120.880 ;
        RECT 64.585 120.710 64.755 120.880 ;
        RECT 64.945 120.710 65.115 120.880 ;
        RECT 65.305 120.710 65.475 120.880 ;
        RECT 65.665 120.710 65.835 120.880 ;
        RECT 66.025 120.710 66.195 120.880 ;
        RECT 66.385 120.710 66.555 120.880 ;
        RECT 66.745 120.710 66.915 120.880 ;
        RECT 67.105 120.710 67.275 120.880 ;
        RECT 67.465 120.710 67.635 120.880 ;
        RECT 67.825 120.710 67.995 120.880 ;
        RECT 69.325 120.710 69.495 120.880 ;
        RECT 69.685 120.710 69.855 120.880 ;
        RECT 70.045 120.710 70.215 120.880 ;
        RECT 70.405 120.710 70.575 120.880 ;
        RECT 70.765 120.710 70.935 120.880 ;
        RECT 71.125 120.710 71.295 120.880 ;
        RECT 71.485 120.710 71.655 120.880 ;
        RECT 71.845 120.710 72.015 120.880 ;
        RECT 72.205 120.710 72.375 120.880 ;
        RECT 72.565 120.710 72.735 120.880 ;
        RECT 72.925 120.710 73.095 120.880 ;
        RECT 73.285 120.710 73.455 120.880 ;
        RECT 73.645 120.710 73.815 120.880 ;
        RECT 74.005 120.710 74.175 120.880 ;
        RECT 75.505 120.710 75.675 120.880 ;
        RECT 75.865 120.710 76.035 120.880 ;
        RECT 76.225 120.710 76.395 120.880 ;
        RECT 76.585 120.710 76.755 120.880 ;
        RECT 76.945 120.710 77.115 120.880 ;
        RECT 77.305 120.710 77.475 120.880 ;
        RECT 77.665 120.710 77.835 120.880 ;
        RECT 78.025 120.710 78.195 120.880 ;
        RECT 78.385 120.710 78.555 120.880 ;
        RECT 78.745 120.710 78.915 120.880 ;
        RECT 79.105 120.710 79.275 120.880 ;
        RECT 79.465 120.710 79.635 120.880 ;
        RECT 79.825 120.710 79.995 120.880 ;
        RECT 80.185 120.710 80.355 120.880 ;
        RECT 27.905 118.985 28.075 119.155 ;
        RECT 28.805 118.985 28.975 119.155 ;
        RECT 40.555 118.985 40.725 119.155 ;
        RECT 41.355 118.985 41.525 119.155 ;
        RECT 52.905 118.985 53.075 119.155 ;
        RECT 53.705 118.985 53.875 119.155 ;
        RECT 65.155 118.985 65.325 119.155 ;
        RECT 65.955 118.985 66.125 119.155 ;
        RECT 77.655 118.985 77.825 119.155 ;
        RECT 78.455 118.985 78.625 119.155 ;
        RECT 19.885 118.010 20.055 118.180 ;
        RECT 20.245 118.010 20.415 118.180 ;
        RECT 20.605 118.010 20.775 118.180 ;
        RECT 20.965 118.010 21.135 118.180 ;
        RECT 21.325 118.010 21.495 118.180 ;
        RECT 21.685 118.010 21.855 118.180 ;
        RECT 22.045 118.010 22.215 118.180 ;
        RECT 22.405 118.010 22.575 118.180 ;
        RECT 22.765 118.010 22.935 118.180 ;
        RECT 23.125 118.010 23.295 118.180 ;
        RECT 23.485 118.010 23.655 118.180 ;
        RECT 23.845 118.010 24.015 118.180 ;
        RECT 24.205 118.010 24.375 118.180 ;
        RECT 24.565 118.010 24.735 118.180 ;
        RECT 26.065 118.010 26.235 118.180 ;
        RECT 26.425 118.010 26.595 118.180 ;
        RECT 26.785 118.010 26.955 118.180 ;
        RECT 27.145 118.010 27.315 118.180 ;
        RECT 27.505 118.010 27.675 118.180 ;
        RECT 27.865 118.010 28.035 118.180 ;
        RECT 28.225 118.010 28.395 118.180 ;
        RECT 28.585 118.010 28.755 118.180 ;
        RECT 28.945 118.010 29.115 118.180 ;
        RECT 29.305 118.010 29.475 118.180 ;
        RECT 29.665 118.010 29.835 118.180 ;
        RECT 30.025 118.010 30.195 118.180 ;
        RECT 30.385 118.010 30.555 118.180 ;
        RECT 30.745 118.010 30.915 118.180 ;
        RECT 32.245 118.010 32.415 118.180 ;
        RECT 32.605 118.010 32.775 118.180 ;
        RECT 32.965 118.010 33.135 118.180 ;
        RECT 33.325 118.010 33.495 118.180 ;
        RECT 33.685 118.010 33.855 118.180 ;
        RECT 34.045 118.010 34.215 118.180 ;
        RECT 34.405 118.010 34.575 118.180 ;
        RECT 34.765 118.010 34.935 118.180 ;
        RECT 35.125 118.010 35.295 118.180 ;
        RECT 35.485 118.010 35.655 118.180 ;
        RECT 35.845 118.010 36.015 118.180 ;
        RECT 36.205 118.010 36.375 118.180 ;
        RECT 36.565 118.010 36.735 118.180 ;
        RECT 36.925 118.010 37.095 118.180 ;
        RECT 38.425 118.010 38.595 118.180 ;
        RECT 38.785 118.010 38.955 118.180 ;
        RECT 39.145 118.010 39.315 118.180 ;
        RECT 39.505 118.010 39.675 118.180 ;
        RECT 39.865 118.010 40.035 118.180 ;
        RECT 40.225 118.010 40.395 118.180 ;
        RECT 40.585 118.010 40.755 118.180 ;
        RECT 40.945 118.010 41.115 118.180 ;
        RECT 41.305 118.010 41.475 118.180 ;
        RECT 41.665 118.010 41.835 118.180 ;
        RECT 42.025 118.010 42.195 118.180 ;
        RECT 42.385 118.010 42.555 118.180 ;
        RECT 42.745 118.010 42.915 118.180 ;
        RECT 43.105 118.010 43.275 118.180 ;
        RECT 44.605 118.010 44.775 118.180 ;
        RECT 44.965 118.010 45.135 118.180 ;
        RECT 45.325 118.010 45.495 118.180 ;
        RECT 45.685 118.010 45.855 118.180 ;
        RECT 46.045 118.010 46.215 118.180 ;
        RECT 46.405 118.010 46.575 118.180 ;
        RECT 46.765 118.010 46.935 118.180 ;
        RECT 47.125 118.010 47.295 118.180 ;
        RECT 47.485 118.010 47.655 118.180 ;
        RECT 47.845 118.010 48.015 118.180 ;
        RECT 48.205 118.010 48.375 118.180 ;
        RECT 48.565 118.010 48.735 118.180 ;
        RECT 48.925 118.010 49.095 118.180 ;
        RECT 49.285 118.010 49.455 118.180 ;
        RECT 50.785 118.010 50.955 118.180 ;
        RECT 51.145 118.010 51.315 118.180 ;
        RECT 51.505 118.010 51.675 118.180 ;
        RECT 51.865 118.010 52.035 118.180 ;
        RECT 52.225 118.010 52.395 118.180 ;
        RECT 52.585 118.010 52.755 118.180 ;
        RECT 52.945 118.010 53.115 118.180 ;
        RECT 53.305 118.010 53.475 118.180 ;
        RECT 53.665 118.010 53.835 118.180 ;
        RECT 54.025 118.010 54.195 118.180 ;
        RECT 54.385 118.010 54.555 118.180 ;
        RECT 54.745 118.010 54.915 118.180 ;
        RECT 55.105 118.010 55.275 118.180 ;
        RECT 55.465 118.010 55.635 118.180 ;
        RECT 56.965 118.010 57.135 118.180 ;
        RECT 57.325 118.010 57.495 118.180 ;
        RECT 57.685 118.010 57.855 118.180 ;
        RECT 58.045 118.010 58.215 118.180 ;
        RECT 58.405 118.010 58.575 118.180 ;
        RECT 58.765 118.010 58.935 118.180 ;
        RECT 59.125 118.010 59.295 118.180 ;
        RECT 59.485 118.010 59.655 118.180 ;
        RECT 59.845 118.010 60.015 118.180 ;
        RECT 60.205 118.010 60.375 118.180 ;
        RECT 60.565 118.010 60.735 118.180 ;
        RECT 60.925 118.010 61.095 118.180 ;
        RECT 61.285 118.010 61.455 118.180 ;
        RECT 61.645 118.010 61.815 118.180 ;
        RECT 63.145 118.010 63.315 118.180 ;
        RECT 63.505 118.010 63.675 118.180 ;
        RECT 63.865 118.010 64.035 118.180 ;
        RECT 64.225 118.010 64.395 118.180 ;
        RECT 64.585 118.010 64.755 118.180 ;
        RECT 64.945 118.010 65.115 118.180 ;
        RECT 65.305 118.010 65.475 118.180 ;
        RECT 65.665 118.010 65.835 118.180 ;
        RECT 66.025 118.010 66.195 118.180 ;
        RECT 66.385 118.010 66.555 118.180 ;
        RECT 66.745 118.010 66.915 118.180 ;
        RECT 67.105 118.010 67.275 118.180 ;
        RECT 67.465 118.010 67.635 118.180 ;
        RECT 67.825 118.010 67.995 118.180 ;
        RECT 69.325 118.010 69.495 118.180 ;
        RECT 69.685 118.010 69.855 118.180 ;
        RECT 70.045 118.010 70.215 118.180 ;
        RECT 70.405 118.010 70.575 118.180 ;
        RECT 70.765 118.010 70.935 118.180 ;
        RECT 71.125 118.010 71.295 118.180 ;
        RECT 71.485 118.010 71.655 118.180 ;
        RECT 71.845 118.010 72.015 118.180 ;
        RECT 72.205 118.010 72.375 118.180 ;
        RECT 72.565 118.010 72.735 118.180 ;
        RECT 72.925 118.010 73.095 118.180 ;
        RECT 73.285 118.010 73.455 118.180 ;
        RECT 73.645 118.010 73.815 118.180 ;
        RECT 74.005 118.010 74.175 118.180 ;
        RECT 75.505 118.010 75.675 118.180 ;
        RECT 75.865 118.010 76.035 118.180 ;
        RECT 76.225 118.010 76.395 118.180 ;
        RECT 76.585 118.010 76.755 118.180 ;
        RECT 76.945 118.010 77.115 118.180 ;
        RECT 77.305 118.010 77.475 118.180 ;
        RECT 77.665 118.010 77.835 118.180 ;
        RECT 78.025 118.010 78.195 118.180 ;
        RECT 78.385 118.010 78.555 118.180 ;
        RECT 78.745 118.010 78.915 118.180 ;
        RECT 79.105 118.010 79.275 118.180 ;
        RECT 79.465 118.010 79.635 118.180 ;
        RECT 79.825 118.010 79.995 118.180 ;
        RECT 80.185 118.010 80.355 118.180 ;
        RECT 19.885 115.310 20.055 115.480 ;
        RECT 20.245 115.310 20.415 115.480 ;
        RECT 20.605 115.310 20.775 115.480 ;
        RECT 20.965 115.310 21.135 115.480 ;
        RECT 21.325 115.310 21.495 115.480 ;
        RECT 21.685 115.310 21.855 115.480 ;
        RECT 22.045 115.310 22.215 115.480 ;
        RECT 22.405 115.310 22.575 115.480 ;
        RECT 22.765 115.310 22.935 115.480 ;
        RECT 23.125 115.310 23.295 115.480 ;
        RECT 23.485 115.310 23.655 115.480 ;
        RECT 23.845 115.310 24.015 115.480 ;
        RECT 24.205 115.310 24.375 115.480 ;
        RECT 24.565 115.310 24.735 115.480 ;
        RECT 26.065 115.310 26.235 115.480 ;
        RECT 26.425 115.310 26.595 115.480 ;
        RECT 26.785 115.310 26.955 115.480 ;
        RECT 27.145 115.310 27.315 115.480 ;
        RECT 27.505 115.310 27.675 115.480 ;
        RECT 27.865 115.310 28.035 115.480 ;
        RECT 28.225 115.310 28.395 115.480 ;
        RECT 28.585 115.310 28.755 115.480 ;
        RECT 28.945 115.310 29.115 115.480 ;
        RECT 29.305 115.310 29.475 115.480 ;
        RECT 29.665 115.310 29.835 115.480 ;
        RECT 30.025 115.310 30.195 115.480 ;
        RECT 30.385 115.310 30.555 115.480 ;
        RECT 30.745 115.310 30.915 115.480 ;
        RECT 32.245 115.310 32.415 115.480 ;
        RECT 32.605 115.310 32.775 115.480 ;
        RECT 32.965 115.310 33.135 115.480 ;
        RECT 33.325 115.310 33.495 115.480 ;
        RECT 33.685 115.310 33.855 115.480 ;
        RECT 34.045 115.310 34.215 115.480 ;
        RECT 34.405 115.310 34.575 115.480 ;
        RECT 34.765 115.310 34.935 115.480 ;
        RECT 35.125 115.310 35.295 115.480 ;
        RECT 35.485 115.310 35.655 115.480 ;
        RECT 35.845 115.310 36.015 115.480 ;
        RECT 36.205 115.310 36.375 115.480 ;
        RECT 36.565 115.310 36.735 115.480 ;
        RECT 36.925 115.310 37.095 115.480 ;
        RECT 38.425 115.310 38.595 115.480 ;
        RECT 38.785 115.310 38.955 115.480 ;
        RECT 39.145 115.310 39.315 115.480 ;
        RECT 39.505 115.310 39.675 115.480 ;
        RECT 39.865 115.310 40.035 115.480 ;
        RECT 40.225 115.310 40.395 115.480 ;
        RECT 40.585 115.310 40.755 115.480 ;
        RECT 40.945 115.310 41.115 115.480 ;
        RECT 41.305 115.310 41.475 115.480 ;
        RECT 41.665 115.310 41.835 115.480 ;
        RECT 42.025 115.310 42.195 115.480 ;
        RECT 42.385 115.310 42.555 115.480 ;
        RECT 42.745 115.310 42.915 115.480 ;
        RECT 43.105 115.310 43.275 115.480 ;
        RECT 44.605 115.310 44.775 115.480 ;
        RECT 44.965 115.310 45.135 115.480 ;
        RECT 45.325 115.310 45.495 115.480 ;
        RECT 45.685 115.310 45.855 115.480 ;
        RECT 46.045 115.310 46.215 115.480 ;
        RECT 46.405 115.310 46.575 115.480 ;
        RECT 46.765 115.310 46.935 115.480 ;
        RECT 47.125 115.310 47.295 115.480 ;
        RECT 47.485 115.310 47.655 115.480 ;
        RECT 47.845 115.310 48.015 115.480 ;
        RECT 48.205 115.310 48.375 115.480 ;
        RECT 48.565 115.310 48.735 115.480 ;
        RECT 48.925 115.310 49.095 115.480 ;
        RECT 49.285 115.310 49.455 115.480 ;
        RECT 50.785 115.310 50.955 115.480 ;
        RECT 51.145 115.310 51.315 115.480 ;
        RECT 51.505 115.310 51.675 115.480 ;
        RECT 51.865 115.310 52.035 115.480 ;
        RECT 52.225 115.310 52.395 115.480 ;
        RECT 52.585 115.310 52.755 115.480 ;
        RECT 52.945 115.310 53.115 115.480 ;
        RECT 53.305 115.310 53.475 115.480 ;
        RECT 53.665 115.310 53.835 115.480 ;
        RECT 54.025 115.310 54.195 115.480 ;
        RECT 54.385 115.310 54.555 115.480 ;
        RECT 54.745 115.310 54.915 115.480 ;
        RECT 55.105 115.310 55.275 115.480 ;
        RECT 55.465 115.310 55.635 115.480 ;
        RECT 56.965 115.310 57.135 115.480 ;
        RECT 57.325 115.310 57.495 115.480 ;
        RECT 57.685 115.310 57.855 115.480 ;
        RECT 58.045 115.310 58.215 115.480 ;
        RECT 58.405 115.310 58.575 115.480 ;
        RECT 58.765 115.310 58.935 115.480 ;
        RECT 59.125 115.310 59.295 115.480 ;
        RECT 59.485 115.310 59.655 115.480 ;
        RECT 59.845 115.310 60.015 115.480 ;
        RECT 60.205 115.310 60.375 115.480 ;
        RECT 60.565 115.310 60.735 115.480 ;
        RECT 60.925 115.310 61.095 115.480 ;
        RECT 61.285 115.310 61.455 115.480 ;
        RECT 61.645 115.310 61.815 115.480 ;
        RECT 63.145 115.310 63.315 115.480 ;
        RECT 63.505 115.310 63.675 115.480 ;
        RECT 63.865 115.310 64.035 115.480 ;
        RECT 64.225 115.310 64.395 115.480 ;
        RECT 64.585 115.310 64.755 115.480 ;
        RECT 64.945 115.310 65.115 115.480 ;
        RECT 65.305 115.310 65.475 115.480 ;
        RECT 65.665 115.310 65.835 115.480 ;
        RECT 66.025 115.310 66.195 115.480 ;
        RECT 66.385 115.310 66.555 115.480 ;
        RECT 66.745 115.310 66.915 115.480 ;
        RECT 67.105 115.310 67.275 115.480 ;
        RECT 67.465 115.310 67.635 115.480 ;
        RECT 67.825 115.310 67.995 115.480 ;
        RECT 69.325 115.310 69.495 115.480 ;
        RECT 69.685 115.310 69.855 115.480 ;
        RECT 70.045 115.310 70.215 115.480 ;
        RECT 70.405 115.310 70.575 115.480 ;
        RECT 70.765 115.310 70.935 115.480 ;
        RECT 71.125 115.310 71.295 115.480 ;
        RECT 71.485 115.310 71.655 115.480 ;
        RECT 71.845 115.310 72.015 115.480 ;
        RECT 72.205 115.310 72.375 115.480 ;
        RECT 72.565 115.310 72.735 115.480 ;
        RECT 72.925 115.310 73.095 115.480 ;
        RECT 73.285 115.310 73.455 115.480 ;
        RECT 73.645 115.310 73.815 115.480 ;
        RECT 74.005 115.310 74.175 115.480 ;
        RECT 75.505 115.310 75.675 115.480 ;
        RECT 75.865 115.310 76.035 115.480 ;
        RECT 76.225 115.310 76.395 115.480 ;
        RECT 76.585 115.310 76.755 115.480 ;
        RECT 76.945 115.310 77.115 115.480 ;
        RECT 77.305 115.310 77.475 115.480 ;
        RECT 77.665 115.310 77.835 115.480 ;
        RECT 78.025 115.310 78.195 115.480 ;
        RECT 78.385 115.310 78.555 115.480 ;
        RECT 78.745 115.310 78.915 115.480 ;
        RECT 79.105 115.310 79.275 115.480 ;
        RECT 79.465 115.310 79.635 115.480 ;
        RECT 79.825 115.310 79.995 115.480 ;
        RECT 80.185 115.310 80.355 115.480 ;
        RECT 27.905 113.585 28.075 113.755 ;
        RECT 28.805 113.635 28.975 113.805 ;
        RECT 40.555 113.585 40.725 113.755 ;
        RECT 41.355 113.585 41.525 113.755 ;
        RECT 52.905 113.585 53.075 113.755 ;
        RECT 53.705 113.585 53.875 113.755 ;
        RECT 65.155 113.585 65.325 113.755 ;
        RECT 65.955 113.585 66.125 113.755 ;
        RECT 77.655 113.585 77.825 113.755 ;
        RECT 78.455 113.585 78.625 113.755 ;
        RECT 19.885 112.610 20.055 112.780 ;
        RECT 20.245 112.610 20.415 112.780 ;
        RECT 20.605 112.610 20.775 112.780 ;
        RECT 20.965 112.610 21.135 112.780 ;
        RECT 21.325 112.610 21.495 112.780 ;
        RECT 21.685 112.610 21.855 112.780 ;
        RECT 22.045 112.610 22.215 112.780 ;
        RECT 22.405 112.610 22.575 112.780 ;
        RECT 22.765 112.610 22.935 112.780 ;
        RECT 23.125 112.610 23.295 112.780 ;
        RECT 23.485 112.610 23.655 112.780 ;
        RECT 23.845 112.610 24.015 112.780 ;
        RECT 24.205 112.610 24.375 112.780 ;
        RECT 24.565 112.610 24.735 112.780 ;
        RECT 26.065 112.610 26.235 112.780 ;
        RECT 26.425 112.610 26.595 112.780 ;
        RECT 26.785 112.610 26.955 112.780 ;
        RECT 27.145 112.610 27.315 112.780 ;
        RECT 27.505 112.610 27.675 112.780 ;
        RECT 27.865 112.610 28.035 112.780 ;
        RECT 28.225 112.610 28.395 112.780 ;
        RECT 28.585 112.610 28.755 112.780 ;
        RECT 28.945 112.610 29.115 112.780 ;
        RECT 29.305 112.610 29.475 112.780 ;
        RECT 29.665 112.610 29.835 112.780 ;
        RECT 30.025 112.610 30.195 112.780 ;
        RECT 30.385 112.610 30.555 112.780 ;
        RECT 30.745 112.610 30.915 112.780 ;
        RECT 32.245 112.610 32.415 112.780 ;
        RECT 32.605 112.610 32.775 112.780 ;
        RECT 32.965 112.610 33.135 112.780 ;
        RECT 33.325 112.610 33.495 112.780 ;
        RECT 33.685 112.610 33.855 112.780 ;
        RECT 34.045 112.610 34.215 112.780 ;
        RECT 34.405 112.610 34.575 112.780 ;
        RECT 34.765 112.610 34.935 112.780 ;
        RECT 35.125 112.610 35.295 112.780 ;
        RECT 35.485 112.610 35.655 112.780 ;
        RECT 35.845 112.610 36.015 112.780 ;
        RECT 36.205 112.610 36.375 112.780 ;
        RECT 36.565 112.610 36.735 112.780 ;
        RECT 36.925 112.610 37.095 112.780 ;
        RECT 38.425 112.610 38.595 112.780 ;
        RECT 38.785 112.610 38.955 112.780 ;
        RECT 39.145 112.610 39.315 112.780 ;
        RECT 39.505 112.610 39.675 112.780 ;
        RECT 39.865 112.610 40.035 112.780 ;
        RECT 40.225 112.610 40.395 112.780 ;
        RECT 40.585 112.610 40.755 112.780 ;
        RECT 40.945 112.610 41.115 112.780 ;
        RECT 41.305 112.610 41.475 112.780 ;
        RECT 41.665 112.610 41.835 112.780 ;
        RECT 42.025 112.610 42.195 112.780 ;
        RECT 42.385 112.610 42.555 112.780 ;
        RECT 42.745 112.610 42.915 112.780 ;
        RECT 43.105 112.610 43.275 112.780 ;
        RECT 44.605 112.610 44.775 112.780 ;
        RECT 44.965 112.610 45.135 112.780 ;
        RECT 45.325 112.610 45.495 112.780 ;
        RECT 45.685 112.610 45.855 112.780 ;
        RECT 46.045 112.610 46.215 112.780 ;
        RECT 46.405 112.610 46.575 112.780 ;
        RECT 46.765 112.610 46.935 112.780 ;
        RECT 47.125 112.610 47.295 112.780 ;
        RECT 47.485 112.610 47.655 112.780 ;
        RECT 47.845 112.610 48.015 112.780 ;
        RECT 48.205 112.610 48.375 112.780 ;
        RECT 48.565 112.610 48.735 112.780 ;
        RECT 48.925 112.610 49.095 112.780 ;
        RECT 49.285 112.610 49.455 112.780 ;
        RECT 50.785 112.610 50.955 112.780 ;
        RECT 51.145 112.610 51.315 112.780 ;
        RECT 51.505 112.610 51.675 112.780 ;
        RECT 51.865 112.610 52.035 112.780 ;
        RECT 52.225 112.610 52.395 112.780 ;
        RECT 52.585 112.610 52.755 112.780 ;
        RECT 52.945 112.610 53.115 112.780 ;
        RECT 53.305 112.610 53.475 112.780 ;
        RECT 53.665 112.610 53.835 112.780 ;
        RECT 54.025 112.610 54.195 112.780 ;
        RECT 54.385 112.610 54.555 112.780 ;
        RECT 54.745 112.610 54.915 112.780 ;
        RECT 55.105 112.610 55.275 112.780 ;
        RECT 55.465 112.610 55.635 112.780 ;
        RECT 56.965 112.610 57.135 112.780 ;
        RECT 57.325 112.610 57.495 112.780 ;
        RECT 57.685 112.610 57.855 112.780 ;
        RECT 58.045 112.610 58.215 112.780 ;
        RECT 58.405 112.610 58.575 112.780 ;
        RECT 58.765 112.610 58.935 112.780 ;
        RECT 59.125 112.610 59.295 112.780 ;
        RECT 59.485 112.610 59.655 112.780 ;
        RECT 59.845 112.610 60.015 112.780 ;
        RECT 60.205 112.610 60.375 112.780 ;
        RECT 60.565 112.610 60.735 112.780 ;
        RECT 60.925 112.610 61.095 112.780 ;
        RECT 61.285 112.610 61.455 112.780 ;
        RECT 61.645 112.610 61.815 112.780 ;
        RECT 63.145 112.610 63.315 112.780 ;
        RECT 63.505 112.610 63.675 112.780 ;
        RECT 63.865 112.610 64.035 112.780 ;
        RECT 64.225 112.610 64.395 112.780 ;
        RECT 64.585 112.610 64.755 112.780 ;
        RECT 64.945 112.610 65.115 112.780 ;
        RECT 65.305 112.610 65.475 112.780 ;
        RECT 65.665 112.610 65.835 112.780 ;
        RECT 66.025 112.610 66.195 112.780 ;
        RECT 66.385 112.610 66.555 112.780 ;
        RECT 66.745 112.610 66.915 112.780 ;
        RECT 67.105 112.610 67.275 112.780 ;
        RECT 67.465 112.610 67.635 112.780 ;
        RECT 67.825 112.610 67.995 112.780 ;
        RECT 69.325 112.610 69.495 112.780 ;
        RECT 69.685 112.610 69.855 112.780 ;
        RECT 70.045 112.610 70.215 112.780 ;
        RECT 70.405 112.610 70.575 112.780 ;
        RECT 70.765 112.610 70.935 112.780 ;
        RECT 71.125 112.610 71.295 112.780 ;
        RECT 71.485 112.610 71.655 112.780 ;
        RECT 71.845 112.610 72.015 112.780 ;
        RECT 72.205 112.610 72.375 112.780 ;
        RECT 72.565 112.610 72.735 112.780 ;
        RECT 72.925 112.610 73.095 112.780 ;
        RECT 73.285 112.610 73.455 112.780 ;
        RECT 73.645 112.610 73.815 112.780 ;
        RECT 74.005 112.610 74.175 112.780 ;
        RECT 75.505 112.610 75.675 112.780 ;
        RECT 75.865 112.610 76.035 112.780 ;
        RECT 76.225 112.610 76.395 112.780 ;
        RECT 76.585 112.610 76.755 112.780 ;
        RECT 76.945 112.610 77.115 112.780 ;
        RECT 77.305 112.610 77.475 112.780 ;
        RECT 77.665 112.610 77.835 112.780 ;
        RECT 78.025 112.610 78.195 112.780 ;
        RECT 78.385 112.610 78.555 112.780 ;
        RECT 78.745 112.610 78.915 112.780 ;
        RECT 79.105 112.610 79.275 112.780 ;
        RECT 79.465 112.610 79.635 112.780 ;
        RECT 79.825 112.610 79.995 112.780 ;
        RECT 80.185 112.610 80.355 112.780 ;
        RECT 34.225 90.285 34.755 90.815 ;
        RECT 39.525 90.285 40.055 90.815 ;
        RECT 46.825 90.285 47.355 90.815 ;
        RECT 52.925 90.285 53.455 90.815 ;
        RECT 60.325 90.285 60.855 90.815 ;
        RECT 65.325 90.285 65.855 90.815 ;
        RECT 32.310 89.740 32.480 89.910 ;
        RECT 32.670 89.740 32.840 89.910 ;
        RECT 33.030 89.740 33.200 89.910 ;
        RECT 33.390 89.740 33.560 89.910 ;
        RECT 33.750 89.740 33.920 89.910 ;
        RECT 34.110 89.740 34.280 89.910 ;
        RECT 34.470 89.740 34.640 89.910 ;
        RECT 34.830 89.740 35.000 89.910 ;
        RECT 35.190 89.740 35.360 89.910 ;
        RECT 35.550 89.740 35.720 89.910 ;
        RECT 35.910 89.740 36.080 89.910 ;
        RECT 36.270 89.740 36.440 89.910 ;
        RECT 36.630 89.740 36.800 89.910 ;
        RECT 36.990 89.740 37.160 89.910 ;
        RECT 38.490 89.740 38.660 89.910 ;
        RECT 38.850 89.740 39.020 89.910 ;
        RECT 39.210 89.740 39.380 89.910 ;
        RECT 39.570 89.740 39.740 89.910 ;
        RECT 39.930 89.740 40.100 89.910 ;
        RECT 40.290 89.740 40.460 89.910 ;
        RECT 40.650 89.740 40.820 89.910 ;
        RECT 41.010 89.740 41.180 89.910 ;
        RECT 41.370 89.740 41.540 89.910 ;
        RECT 41.730 89.740 41.900 89.910 ;
        RECT 42.090 89.740 42.260 89.910 ;
        RECT 42.450 89.740 42.620 89.910 ;
        RECT 42.810 89.740 42.980 89.910 ;
        RECT 43.170 89.740 43.340 89.910 ;
        RECT 44.670 89.740 44.840 89.910 ;
        RECT 45.030 89.740 45.200 89.910 ;
        RECT 45.390 89.740 45.560 89.910 ;
        RECT 45.750 89.740 45.920 89.910 ;
        RECT 46.110 89.740 46.280 89.910 ;
        RECT 46.470 89.740 46.640 89.910 ;
        RECT 46.830 89.740 47.000 89.910 ;
        RECT 47.190 89.740 47.360 89.910 ;
        RECT 47.550 89.740 47.720 89.910 ;
        RECT 47.910 89.740 48.080 89.910 ;
        RECT 48.270 89.740 48.440 89.910 ;
        RECT 48.630 89.740 48.800 89.910 ;
        RECT 48.990 89.740 49.160 89.910 ;
        RECT 49.350 89.740 49.520 89.910 ;
        RECT 50.850 89.740 51.020 89.910 ;
        RECT 51.210 89.740 51.380 89.910 ;
        RECT 51.570 89.740 51.740 89.910 ;
        RECT 51.930 89.740 52.100 89.910 ;
        RECT 52.290 89.740 52.460 89.910 ;
        RECT 52.650 89.740 52.820 89.910 ;
        RECT 53.010 89.740 53.180 89.910 ;
        RECT 53.370 89.740 53.540 89.910 ;
        RECT 53.730 89.740 53.900 89.910 ;
        RECT 54.090 89.740 54.260 89.910 ;
        RECT 54.450 89.740 54.620 89.910 ;
        RECT 54.810 89.740 54.980 89.910 ;
        RECT 55.170 89.740 55.340 89.910 ;
        RECT 55.530 89.740 55.700 89.910 ;
        RECT 57.030 89.740 57.200 89.910 ;
        RECT 57.390 89.740 57.560 89.910 ;
        RECT 57.750 89.740 57.920 89.910 ;
        RECT 58.110 89.740 58.280 89.910 ;
        RECT 58.470 89.740 58.640 89.910 ;
        RECT 58.830 89.740 59.000 89.910 ;
        RECT 59.190 89.740 59.360 89.910 ;
        RECT 59.550 89.740 59.720 89.910 ;
        RECT 59.910 89.740 60.080 89.910 ;
        RECT 60.270 89.740 60.440 89.910 ;
        RECT 60.630 89.740 60.800 89.910 ;
        RECT 60.990 89.740 61.160 89.910 ;
        RECT 61.350 89.740 61.520 89.910 ;
        RECT 61.710 89.740 61.880 89.910 ;
        RECT 63.210 89.740 63.380 89.910 ;
        RECT 63.570 89.740 63.740 89.910 ;
        RECT 63.930 89.740 64.100 89.910 ;
        RECT 64.290 89.740 64.460 89.910 ;
        RECT 64.650 89.740 64.820 89.910 ;
        RECT 65.010 89.740 65.180 89.910 ;
        RECT 65.370 89.740 65.540 89.910 ;
        RECT 65.730 89.740 65.900 89.910 ;
        RECT 66.090 89.740 66.260 89.910 ;
        RECT 66.450 89.740 66.620 89.910 ;
        RECT 66.810 89.740 66.980 89.910 ;
        RECT 67.170 89.740 67.340 89.910 ;
        RECT 67.530 89.740 67.700 89.910 ;
        RECT 67.890 89.740 68.060 89.910 ;
        RECT 34.225 87.385 34.755 87.915 ;
        RECT 39.525 87.385 40.055 87.915 ;
        RECT 46.825 87.385 47.355 87.915 ;
        RECT 52.925 87.385 53.455 87.915 ;
        RECT 60.325 87.385 60.855 87.915 ;
        RECT 65.325 87.385 65.855 87.915 ;
        RECT 32.310 86.790 32.480 86.960 ;
        RECT 32.670 86.790 32.840 86.960 ;
        RECT 33.030 86.790 33.200 86.960 ;
        RECT 33.390 86.790 33.560 86.960 ;
        RECT 33.750 86.790 33.920 86.960 ;
        RECT 34.110 86.790 34.280 86.960 ;
        RECT 34.470 86.790 34.640 86.960 ;
        RECT 34.830 86.790 35.000 86.960 ;
        RECT 35.190 86.790 35.360 86.960 ;
        RECT 35.550 86.790 35.720 86.960 ;
        RECT 35.910 86.790 36.080 86.960 ;
        RECT 36.270 86.790 36.440 86.960 ;
        RECT 36.630 86.790 36.800 86.960 ;
        RECT 36.990 86.790 37.160 86.960 ;
        RECT 38.490 86.790 38.660 86.960 ;
        RECT 38.850 86.790 39.020 86.960 ;
        RECT 39.210 86.790 39.380 86.960 ;
        RECT 39.570 86.790 39.740 86.960 ;
        RECT 39.930 86.790 40.100 86.960 ;
        RECT 40.290 86.790 40.460 86.960 ;
        RECT 40.650 86.790 40.820 86.960 ;
        RECT 41.010 86.790 41.180 86.960 ;
        RECT 41.370 86.790 41.540 86.960 ;
        RECT 41.730 86.790 41.900 86.960 ;
        RECT 42.090 86.790 42.260 86.960 ;
        RECT 42.450 86.790 42.620 86.960 ;
        RECT 42.810 86.790 42.980 86.960 ;
        RECT 43.170 86.790 43.340 86.960 ;
        RECT 44.670 86.790 44.840 86.960 ;
        RECT 45.030 86.790 45.200 86.960 ;
        RECT 45.390 86.790 45.560 86.960 ;
        RECT 45.750 86.790 45.920 86.960 ;
        RECT 46.110 86.790 46.280 86.960 ;
        RECT 46.470 86.790 46.640 86.960 ;
        RECT 46.830 86.790 47.000 86.960 ;
        RECT 47.190 86.790 47.360 86.960 ;
        RECT 47.550 86.790 47.720 86.960 ;
        RECT 47.910 86.790 48.080 86.960 ;
        RECT 48.270 86.790 48.440 86.960 ;
        RECT 48.630 86.790 48.800 86.960 ;
        RECT 48.990 86.790 49.160 86.960 ;
        RECT 49.350 86.790 49.520 86.960 ;
        RECT 50.850 86.790 51.020 86.960 ;
        RECT 51.210 86.790 51.380 86.960 ;
        RECT 51.570 86.790 51.740 86.960 ;
        RECT 51.930 86.790 52.100 86.960 ;
        RECT 52.290 86.790 52.460 86.960 ;
        RECT 52.650 86.790 52.820 86.960 ;
        RECT 53.010 86.790 53.180 86.960 ;
        RECT 53.370 86.790 53.540 86.960 ;
        RECT 53.730 86.790 53.900 86.960 ;
        RECT 54.090 86.790 54.260 86.960 ;
        RECT 54.450 86.790 54.620 86.960 ;
        RECT 54.810 86.790 54.980 86.960 ;
        RECT 55.170 86.790 55.340 86.960 ;
        RECT 55.530 86.790 55.700 86.960 ;
        RECT 57.030 86.790 57.200 86.960 ;
        RECT 57.390 86.790 57.560 86.960 ;
        RECT 57.750 86.790 57.920 86.960 ;
        RECT 58.110 86.790 58.280 86.960 ;
        RECT 58.470 86.790 58.640 86.960 ;
        RECT 58.830 86.790 59.000 86.960 ;
        RECT 59.190 86.790 59.360 86.960 ;
        RECT 59.550 86.790 59.720 86.960 ;
        RECT 59.910 86.790 60.080 86.960 ;
        RECT 60.270 86.790 60.440 86.960 ;
        RECT 60.630 86.790 60.800 86.960 ;
        RECT 60.990 86.790 61.160 86.960 ;
        RECT 61.350 86.790 61.520 86.960 ;
        RECT 61.710 86.790 61.880 86.960 ;
        RECT 63.210 86.790 63.380 86.960 ;
        RECT 63.570 86.790 63.740 86.960 ;
        RECT 63.930 86.790 64.100 86.960 ;
        RECT 64.290 86.790 64.460 86.960 ;
        RECT 64.650 86.790 64.820 86.960 ;
        RECT 65.010 86.790 65.180 86.960 ;
        RECT 65.370 86.790 65.540 86.960 ;
        RECT 65.730 86.790 65.900 86.960 ;
        RECT 66.090 86.790 66.260 86.960 ;
        RECT 66.450 86.790 66.620 86.960 ;
        RECT 66.810 86.790 66.980 86.960 ;
        RECT 67.170 86.790 67.340 86.960 ;
        RECT 67.530 86.790 67.700 86.960 ;
        RECT 67.890 86.790 68.060 86.960 ;
      LAYER met1 ;
        RECT 36.955 137.990 37.525 138.400 ;
        RECT 37.805 137.990 38.375 138.400 ;
        RECT 49.405 137.990 49.975 138.400 ;
        RECT 50.255 137.990 50.825 138.400 ;
        RECT 61.705 137.990 62.225 138.450 ;
        RECT 62.555 137.990 63.075 138.450 ;
        RECT 36.965 137.570 37.465 137.820 ;
        RECT 37.815 137.570 38.315 137.820 ;
        RECT 49.415 137.570 49.915 137.820 ;
        RECT 50.265 137.570 50.765 137.820 ;
        RECT 61.715 137.570 62.215 137.770 ;
        RECT 62.565 137.570 63.065 137.770 ;
        RECT 28.965 137.370 71.165 137.570 ;
        RECT 29.010 137.280 34.010 137.370 ;
        RECT 35.190 137.280 40.190 137.370 ;
        RECT 41.370 137.280 46.370 137.370 ;
        RECT 47.550 137.280 52.550 137.370 ;
        RECT 53.730 137.280 58.730 137.370 ;
        RECT 59.910 137.280 64.910 137.370 ;
        RECT 66.090 137.280 71.090 137.370 ;
        RECT 36.965 134.870 37.465 135.120 ;
        RECT 37.815 134.870 38.315 135.120 ;
        RECT 49.415 134.870 49.915 135.120 ;
        RECT 50.265 134.870 50.765 135.120 ;
        RECT 61.715 134.870 62.215 135.070 ;
        RECT 62.565 134.870 63.065 135.070 ;
        RECT 28.965 134.670 71.165 134.870 ;
        RECT 29.010 134.580 34.010 134.670 ;
        RECT 35.190 134.580 40.190 134.670 ;
        RECT 41.370 134.580 46.370 134.670 ;
        RECT 47.550 134.580 52.550 134.670 ;
        RECT 53.730 134.580 58.730 134.670 ;
        RECT 59.910 134.580 64.910 134.670 ;
        RECT 66.090 134.580 71.090 134.670 ;
        RECT 37.015 133.150 38.315 133.320 ;
        RECT 37.005 132.740 38.315 133.150 ;
        RECT 49.405 132.740 49.975 133.150 ;
        RECT 50.205 132.790 50.775 133.200 ;
        RECT 61.705 132.790 62.225 133.200 ;
        RECT 62.555 132.790 63.075 133.200 ;
        RECT 37.015 132.570 38.315 132.740 ;
        RECT 36.965 132.170 37.465 132.420 ;
        RECT 37.815 132.170 38.315 132.420 ;
        RECT 49.415 132.170 49.915 132.470 ;
        RECT 50.265 132.170 50.765 132.470 ;
        RECT 61.715 132.170 62.215 132.370 ;
        RECT 62.565 132.170 63.065 132.370 ;
        RECT 28.965 131.970 71.165 132.170 ;
        RECT 29.010 131.880 34.010 131.970 ;
        RECT 35.190 131.880 40.190 131.970 ;
        RECT 41.370 131.880 46.370 131.970 ;
        RECT 47.550 131.880 52.550 131.970 ;
        RECT 53.730 131.880 58.730 131.970 ;
        RECT 59.910 131.880 64.910 131.970 ;
        RECT 66.090 131.880 71.090 131.970 ;
        RECT 37.005 130.040 37.525 130.500 ;
        RECT 37.855 130.040 38.375 130.500 ;
        RECT 49.405 130.040 49.925 130.500 ;
        RECT 50.255 130.040 50.775 130.500 ;
        RECT 61.705 130.040 62.225 130.500 ;
        RECT 62.555 130.040 63.075 130.500 ;
        RECT 37.015 129.520 37.515 129.820 ;
        RECT 37.865 129.520 38.365 129.820 ;
        RECT 49.415 129.520 49.915 129.870 ;
        RECT 50.265 129.520 50.765 129.870 ;
        RECT 61.715 129.520 62.215 129.820 ;
        RECT 62.565 129.520 63.065 129.820 ;
        RECT 29.015 129.410 71.215 129.520 ;
        RECT 29.010 129.320 71.215 129.410 ;
        RECT 29.010 129.180 34.010 129.320 ;
        RECT 35.190 129.180 40.190 129.320 ;
        RECT 41.370 129.180 46.370 129.320 ;
        RECT 47.550 129.180 52.550 129.320 ;
        RECT 53.730 129.180 58.730 129.320 ;
        RECT 59.910 129.180 64.910 129.320 ;
        RECT 66.090 129.180 71.090 129.320 ;
        RECT 37.015 126.620 37.515 126.920 ;
        RECT 37.865 126.620 38.365 126.920 ;
        RECT 49.415 126.620 49.915 126.970 ;
        RECT 50.265 126.620 50.765 126.970 ;
        RECT 61.715 126.620 62.215 126.920 ;
        RECT 62.565 126.620 63.065 126.920 ;
        RECT 28.965 126.420 71.165 126.620 ;
        RECT 29.010 126.280 34.010 126.420 ;
        RECT 35.190 126.280 40.190 126.420 ;
        RECT 41.370 126.280 46.370 126.420 ;
        RECT 47.550 126.280 52.550 126.420 ;
        RECT 53.730 126.280 58.730 126.420 ;
        RECT 59.910 126.280 64.910 126.420 ;
        RECT 66.090 126.280 71.090 126.420 ;
        RECT 37.005 124.240 37.575 124.700 ;
        RECT 37.805 124.240 38.375 124.700 ;
        RECT 49.405 124.240 49.925 124.650 ;
        RECT 50.255 124.240 50.775 124.650 ;
        RECT 61.705 124.240 62.225 124.650 ;
        RECT 62.555 124.240 63.075 124.650 ;
        RECT 37.015 123.720 37.515 124.020 ;
        RECT 37.865 123.720 38.365 124.020 ;
        RECT 49.415 123.720 49.915 124.070 ;
        RECT 50.265 123.720 50.765 124.070 ;
        RECT 61.715 123.720 62.215 124.020 ;
        RECT 62.565 123.720 63.065 124.020 ;
        RECT 28.965 123.520 71.165 123.720 ;
        RECT 29.010 123.380 34.010 123.520 ;
        RECT 35.190 123.380 40.190 123.520 ;
        RECT 41.370 123.380 46.370 123.520 ;
        RECT 47.550 123.380 52.550 123.520 ;
        RECT 53.730 123.380 58.730 123.520 ;
        RECT 59.910 123.380 64.910 123.520 ;
        RECT 66.090 123.380 71.090 123.520 ;
        RECT 27.615 121.020 28.115 121.370 ;
        RECT 28.765 121.020 29.265 121.370 ;
        RECT 40.365 121.020 40.865 121.320 ;
        RECT 41.215 121.020 41.715 121.320 ;
        RECT 52.665 121.020 53.165 121.320 ;
        RECT 53.615 121.020 54.115 121.320 ;
        RECT 64.915 121.020 65.415 121.320 ;
        RECT 65.865 121.020 66.365 121.320 ;
        RECT 77.465 121.020 77.965 121.320 ;
        RECT 78.315 121.020 78.815 121.320 ;
        RECT 19.765 120.770 80.515 121.020 ;
        RECT 19.810 120.680 24.810 120.770 ;
        RECT 25.990 120.680 30.990 120.770 ;
        RECT 32.170 120.680 37.170 120.770 ;
        RECT 38.350 120.680 43.350 120.770 ;
        RECT 44.530 120.680 49.530 120.770 ;
        RECT 50.710 120.680 55.710 120.770 ;
        RECT 56.890 120.680 61.890 120.770 ;
        RECT 63.070 120.680 68.070 120.770 ;
        RECT 69.250 120.680 74.250 120.770 ;
        RECT 75.430 120.680 80.430 120.770 ;
        RECT 27.705 118.840 28.275 119.300 ;
        RECT 28.605 118.840 29.175 119.300 ;
        RECT 40.355 118.840 40.925 119.300 ;
        RECT 41.155 118.840 41.725 119.300 ;
        RECT 52.705 118.840 53.275 119.300 ;
        RECT 53.505 118.840 54.075 119.300 ;
        RECT 64.955 118.840 65.525 119.300 ;
        RECT 65.755 118.840 66.325 119.300 ;
        RECT 77.455 118.840 78.025 119.300 ;
        RECT 78.255 118.840 78.825 119.300 ;
        RECT 27.615 118.370 28.115 118.670 ;
        RECT 28.765 118.370 29.265 118.670 ;
        RECT 40.365 118.370 40.865 118.620 ;
        RECT 41.215 118.370 41.715 118.670 ;
        RECT 52.665 118.370 53.165 118.670 ;
        RECT 53.615 118.370 54.115 118.670 ;
        RECT 64.915 118.370 65.415 118.620 ;
        RECT 65.865 118.370 66.365 118.620 ;
        RECT 77.465 118.370 77.965 118.620 ;
        RECT 78.315 118.370 78.815 118.620 ;
        RECT 19.765 118.120 80.515 118.370 ;
        RECT 19.810 117.980 24.810 118.120 ;
        RECT 25.990 117.980 30.990 118.120 ;
        RECT 32.170 117.980 37.170 118.120 ;
        RECT 38.350 117.980 43.350 118.120 ;
        RECT 44.530 117.980 49.530 118.120 ;
        RECT 50.710 117.980 55.710 118.120 ;
        RECT 56.890 117.980 61.890 118.120 ;
        RECT 63.070 117.980 68.070 118.120 ;
        RECT 69.250 117.980 74.250 118.120 ;
        RECT 75.430 117.980 80.430 118.120 ;
        RECT 27.615 115.670 28.115 115.970 ;
        RECT 28.765 115.670 29.265 115.970 ;
        RECT 40.315 115.670 40.815 115.920 ;
        RECT 41.165 115.670 41.665 115.920 ;
        RECT 52.665 115.670 53.165 115.920 ;
        RECT 53.565 115.670 54.065 115.920 ;
        RECT 64.915 115.670 65.415 115.920 ;
        RECT 65.865 115.670 66.365 115.920 ;
        RECT 77.465 115.670 77.965 115.920 ;
        RECT 78.315 115.670 78.815 115.920 ;
        RECT 19.765 115.420 80.515 115.670 ;
        RECT 19.810 115.280 24.810 115.420 ;
        RECT 25.990 115.280 30.990 115.420 ;
        RECT 32.170 115.280 37.170 115.420 ;
        RECT 38.350 115.280 43.350 115.420 ;
        RECT 44.530 115.280 49.530 115.420 ;
        RECT 50.710 115.280 55.710 115.420 ;
        RECT 56.890 115.280 61.890 115.420 ;
        RECT 63.070 115.280 68.070 115.420 ;
        RECT 69.250 115.280 74.250 115.420 ;
        RECT 75.430 115.280 80.430 115.420 ;
        RECT 27.705 113.440 28.275 113.900 ;
        RECT 28.605 113.490 29.175 113.950 ;
        RECT 40.355 113.440 40.925 113.900 ;
        RECT 41.155 113.440 41.725 113.900 ;
        RECT 52.705 113.440 53.275 113.900 ;
        RECT 53.505 113.440 54.075 113.900 ;
        RECT 64.955 113.440 65.525 113.900 ;
        RECT 65.755 113.440 66.325 113.900 ;
        RECT 77.455 113.440 78.025 113.900 ;
        RECT 78.255 113.440 78.825 113.900 ;
        RECT 27.615 112.970 28.115 113.220 ;
        RECT 28.765 112.970 29.265 113.220 ;
        RECT 40.265 112.970 40.765 113.270 ;
        RECT 41.215 112.970 41.715 113.270 ;
        RECT 52.665 112.970 53.165 113.220 ;
        RECT 53.615 112.970 54.115 113.220 ;
        RECT 64.915 112.970 65.415 113.220 ;
        RECT 65.865 112.970 66.365 113.220 ;
        RECT 77.465 112.970 77.965 113.170 ;
        RECT 78.315 112.970 78.815 113.170 ;
        RECT 19.765 112.720 80.515 112.970 ;
        RECT 19.810 112.580 24.810 112.720 ;
        RECT 25.990 112.580 30.990 112.720 ;
        RECT 32.170 112.580 37.170 112.720 ;
        RECT 38.350 112.580 43.350 112.720 ;
        RECT 44.530 112.580 49.530 112.720 ;
        RECT 50.710 112.580 55.710 112.720 ;
        RECT 56.890 112.580 61.890 112.720 ;
        RECT 63.070 112.580 68.070 112.720 ;
        RECT 69.250 112.580 74.250 112.720 ;
        RECT 75.430 112.580 80.430 112.720 ;
        RECT 34.030 90.950 34.950 90.980 ;
        RECT 39.330 90.950 40.250 90.980 ;
        RECT 46.630 90.950 47.550 90.980 ;
        RECT 52.730 90.950 53.650 90.980 ;
        RECT 60.130 90.950 61.050 90.980 ;
        RECT 65.130 90.950 66.050 90.980 ;
        RECT 32.190 89.850 68.190 90.950 ;
        RECT 32.190 89.650 37.290 89.850 ;
        RECT 38.390 89.710 43.415 89.850 ;
        RECT 44.590 89.710 49.595 89.850 ;
        RECT 50.775 89.710 55.790 89.850 ;
        RECT 38.390 89.650 43.390 89.710 ;
        RECT 44.590 89.650 49.590 89.710 ;
        RECT 50.790 89.650 55.790 89.710 ;
        RECT 56.890 89.650 61.990 89.850 ;
        RECT 63.090 89.650 68.190 89.850 ;
        RECT 34.030 88.050 34.950 88.080 ;
        RECT 39.330 88.050 40.250 88.080 ;
        RECT 46.630 88.050 47.550 88.080 ;
        RECT 52.730 88.050 53.650 88.080 ;
        RECT 60.130 88.050 61.050 88.080 ;
        RECT 65.130 88.050 66.050 88.080 ;
        RECT 32.190 86.900 68.190 88.050 ;
        RECT 32.190 86.850 37.235 86.900 ;
        RECT 32.235 86.760 37.235 86.850 ;
        RECT 38.415 86.760 43.415 86.900 ;
        RECT 44.595 86.760 49.595 86.900 ;
        RECT 50.775 86.760 55.775 86.900 ;
        RECT 56.955 86.760 61.955 86.900 ;
        RECT 63.135 86.850 68.190 86.900 ;
        RECT 63.135 86.760 68.135 86.850 ;
      LAYER via ;
        RECT 37.110 138.065 37.370 138.325 ;
        RECT 37.960 138.065 38.220 138.325 ;
        RECT 49.560 138.065 49.820 138.325 ;
        RECT 50.410 138.065 50.670 138.325 ;
        RECT 61.835 138.090 62.095 138.350 ;
        RECT 62.685 138.090 62.945 138.350 ;
        RECT 37.085 137.490 37.345 137.750 ;
        RECT 37.935 137.490 38.195 137.750 ;
        RECT 49.535 137.490 49.795 137.750 ;
        RECT 50.385 137.490 50.645 137.750 ;
        RECT 61.835 137.440 62.095 137.700 ;
        RECT 62.685 137.440 62.945 137.700 ;
        RECT 37.085 134.790 37.345 135.050 ;
        RECT 37.935 134.790 38.195 135.050 ;
        RECT 49.535 134.790 49.795 135.050 ;
        RECT 50.385 134.790 50.645 135.050 ;
        RECT 61.835 134.740 62.095 135.000 ;
        RECT 62.685 134.740 62.945 135.000 ;
        RECT 37.160 132.815 37.420 133.075 ;
        RECT 37.860 132.815 38.120 133.075 ;
        RECT 49.560 132.815 49.820 133.075 ;
        RECT 50.360 132.865 50.620 133.125 ;
        RECT 61.835 132.865 62.095 133.125 ;
        RECT 62.685 132.865 62.945 133.125 ;
        RECT 37.085 132.090 37.345 132.350 ;
        RECT 37.935 132.090 38.195 132.350 ;
        RECT 49.535 132.140 49.795 132.400 ;
        RECT 50.385 132.140 50.645 132.400 ;
        RECT 61.835 132.040 62.095 132.300 ;
        RECT 62.685 132.040 62.945 132.300 ;
        RECT 37.135 130.140 37.395 130.400 ;
        RECT 37.985 130.140 38.245 130.400 ;
        RECT 49.535 130.140 49.795 130.400 ;
        RECT 50.385 130.140 50.645 130.400 ;
        RECT 61.835 130.140 62.095 130.400 ;
        RECT 62.685 130.140 62.945 130.400 ;
        RECT 37.135 129.490 37.395 129.750 ;
        RECT 37.985 129.490 38.245 129.750 ;
        RECT 49.535 129.540 49.795 129.800 ;
        RECT 50.385 129.540 50.645 129.800 ;
        RECT 61.835 129.490 62.095 129.750 ;
        RECT 62.685 129.490 62.945 129.750 ;
        RECT 37.135 126.590 37.395 126.850 ;
        RECT 37.985 126.590 38.245 126.850 ;
        RECT 49.535 126.640 49.795 126.900 ;
        RECT 50.385 126.640 50.645 126.900 ;
        RECT 61.835 126.590 62.095 126.850 ;
        RECT 62.685 126.590 62.945 126.850 ;
        RECT 37.160 124.340 37.420 124.600 ;
        RECT 37.960 124.340 38.220 124.600 ;
        RECT 49.535 124.315 49.795 124.575 ;
        RECT 50.385 124.315 50.645 124.575 ;
        RECT 61.835 124.315 62.095 124.575 ;
        RECT 62.685 124.315 62.945 124.575 ;
        RECT 37.135 123.690 37.395 123.950 ;
        RECT 37.985 123.690 38.245 123.950 ;
        RECT 49.535 123.740 49.795 124.000 ;
        RECT 50.385 123.740 50.645 124.000 ;
        RECT 61.835 123.690 62.095 123.950 ;
        RECT 62.685 123.690 62.945 123.950 ;
        RECT 27.735 121.040 27.995 121.300 ;
        RECT 28.885 121.040 29.145 121.300 ;
        RECT 40.485 120.990 40.745 121.250 ;
        RECT 41.335 120.990 41.595 121.250 ;
        RECT 52.785 120.990 53.045 121.250 ;
        RECT 53.735 120.990 53.995 121.250 ;
        RECT 65.035 120.990 65.295 121.250 ;
        RECT 65.985 120.990 66.245 121.250 ;
        RECT 77.585 120.990 77.845 121.250 ;
        RECT 78.435 120.990 78.695 121.250 ;
        RECT 27.860 118.940 28.120 119.200 ;
        RECT 28.760 118.940 29.020 119.200 ;
        RECT 40.510 118.940 40.770 119.200 ;
        RECT 41.310 118.940 41.570 119.200 ;
        RECT 52.860 118.940 53.120 119.200 ;
        RECT 53.660 118.940 53.920 119.200 ;
        RECT 65.110 118.940 65.370 119.200 ;
        RECT 65.910 118.940 66.170 119.200 ;
        RECT 77.610 118.940 77.870 119.200 ;
        RECT 78.410 118.940 78.670 119.200 ;
        RECT 27.735 118.340 27.995 118.600 ;
        RECT 28.885 118.340 29.145 118.600 ;
        RECT 40.485 118.290 40.745 118.550 ;
        RECT 41.335 118.340 41.595 118.600 ;
        RECT 52.785 118.340 53.045 118.600 ;
        RECT 53.735 118.340 53.995 118.600 ;
        RECT 65.035 118.290 65.295 118.550 ;
        RECT 65.985 118.290 66.245 118.550 ;
        RECT 77.585 118.290 77.845 118.550 ;
        RECT 78.435 118.290 78.695 118.550 ;
        RECT 27.735 115.640 27.995 115.900 ;
        RECT 28.885 115.640 29.145 115.900 ;
        RECT 40.435 115.590 40.695 115.850 ;
        RECT 41.285 115.590 41.545 115.850 ;
        RECT 52.785 115.590 53.045 115.850 ;
        RECT 53.685 115.590 53.945 115.850 ;
        RECT 65.035 115.590 65.295 115.850 ;
        RECT 65.985 115.590 66.245 115.850 ;
        RECT 77.585 115.590 77.845 115.850 ;
        RECT 78.435 115.590 78.695 115.850 ;
        RECT 27.860 113.540 28.120 113.800 ;
        RECT 28.760 113.590 29.020 113.850 ;
        RECT 40.510 113.540 40.770 113.800 ;
        RECT 41.310 113.540 41.570 113.800 ;
        RECT 52.860 113.540 53.120 113.800 ;
        RECT 53.660 113.540 53.920 113.800 ;
        RECT 65.110 113.540 65.370 113.800 ;
        RECT 65.910 113.540 66.170 113.800 ;
        RECT 77.610 113.540 77.870 113.800 ;
        RECT 78.410 113.540 78.670 113.800 ;
        RECT 27.735 112.890 27.995 113.150 ;
        RECT 28.885 112.890 29.145 113.150 ;
        RECT 40.385 112.940 40.645 113.200 ;
        RECT 41.335 112.940 41.595 113.200 ;
        RECT 52.785 112.890 53.045 113.150 ;
        RECT 53.735 112.890 53.995 113.150 ;
        RECT 65.035 112.890 65.295 113.150 ;
        RECT 65.985 112.890 66.245 113.150 ;
        RECT 77.585 112.840 77.845 113.100 ;
        RECT 78.435 112.840 78.695 113.100 ;
        RECT 34.200 90.260 34.780 90.840 ;
        RECT 39.500 90.260 40.080 90.840 ;
        RECT 46.800 90.260 47.380 90.840 ;
        RECT 52.900 90.260 53.480 90.840 ;
        RECT 60.300 90.260 60.880 90.840 ;
        RECT 65.300 90.260 65.880 90.840 ;
        RECT 34.200 87.360 34.780 87.940 ;
        RECT 39.500 87.360 40.080 87.940 ;
        RECT 46.800 87.360 47.380 87.940 ;
        RECT 52.900 87.360 53.480 87.940 ;
        RECT 60.300 87.360 60.880 87.940 ;
        RECT 65.300 87.360 65.880 87.940 ;
      LAYER met2 ;
        RECT 36.915 131.970 38.365 138.470 ;
        RECT 49.365 131.970 50.815 138.470 ;
        RECT 61.665 130.720 63.115 138.620 ;
        RECT 37.065 130.020 37.465 130.520 ;
        RECT 37.915 130.020 38.315 130.520 ;
        RECT 49.465 130.070 49.865 130.520 ;
        RECT 50.315 130.070 50.715 130.520 ;
        RECT 61.765 130.070 62.165 130.520 ;
        RECT 62.615 130.070 63.015 130.520 ;
        RECT 36.965 123.520 38.415 130.020 ;
        RECT 49.365 123.570 50.815 130.070 ;
        RECT 61.665 123.570 63.115 130.070 ;
        RECT 27.665 112.770 29.215 121.470 ;
        RECT 40.315 112.720 41.765 121.470 ;
        RECT 52.665 112.770 54.115 121.520 ;
        RECT 64.915 111.570 66.365 121.470 ;
        RECT 77.415 112.670 78.865 121.420 ;
        RECT 34.090 90.100 34.890 91.000 ;
        RECT 39.390 90.100 40.190 91.000 ;
        RECT 46.690 90.100 47.490 91.000 ;
        RECT 52.790 90.100 53.590 91.000 ;
        RECT 60.190 90.100 60.990 91.000 ;
        RECT 65.190 90.100 65.990 91.000 ;
        RECT 34.090 87.200 34.890 88.100 ;
        RECT 39.390 87.200 40.190 88.100 ;
        RECT 46.690 87.200 47.490 88.100 ;
        RECT 52.790 87.200 53.590 88.100 ;
        RECT 60.190 87.200 60.990 88.100 ;
        RECT 65.190 87.200 65.990 88.100 ;
      LAYER via2 ;
        RECT 37.100 138.055 37.380 138.335 ;
        RECT 37.950 138.055 38.230 138.335 ;
        RECT 37.150 132.805 37.430 133.085 ;
        RECT 37.850 132.805 38.130 133.085 ;
        RECT 49.550 138.055 49.830 138.335 ;
        RECT 50.400 138.055 50.680 138.335 ;
        RECT 49.550 132.805 49.830 133.085 ;
        RECT 50.350 132.855 50.630 133.135 ;
        RECT 61.825 138.080 62.105 138.360 ;
        RECT 62.675 138.080 62.955 138.360 ;
        RECT 61.825 132.855 62.105 133.135 ;
        RECT 62.675 132.855 62.955 133.135 ;
        RECT 37.125 130.130 37.405 130.410 ;
        RECT 37.975 130.130 38.255 130.410 ;
        RECT 49.525 130.130 49.805 130.410 ;
        RECT 50.375 130.130 50.655 130.410 ;
        RECT 61.825 130.130 62.105 130.410 ;
        RECT 62.675 130.130 62.955 130.410 ;
        RECT 37.150 124.330 37.430 124.610 ;
        RECT 37.950 124.330 38.230 124.610 ;
        RECT 49.525 124.305 49.805 124.585 ;
        RECT 50.375 124.305 50.655 124.585 ;
        RECT 61.825 124.305 62.105 124.585 ;
        RECT 62.675 124.305 62.955 124.585 ;
        RECT 27.850 118.930 28.130 119.210 ;
        RECT 28.750 118.930 29.030 119.210 ;
        RECT 27.850 113.530 28.130 113.810 ;
        RECT 28.750 113.580 29.030 113.860 ;
        RECT 40.500 118.930 40.780 119.210 ;
        RECT 41.300 118.930 41.580 119.210 ;
        RECT 40.500 113.530 40.780 113.810 ;
        RECT 41.300 113.530 41.580 113.810 ;
        RECT 52.850 118.930 53.130 119.210 ;
        RECT 53.650 118.930 53.930 119.210 ;
        RECT 52.850 113.530 53.130 113.810 ;
        RECT 53.650 113.530 53.930 113.810 ;
        RECT 65.100 118.930 65.380 119.210 ;
        RECT 65.900 118.930 66.180 119.210 ;
        RECT 65.100 113.530 65.380 113.810 ;
        RECT 65.900 113.530 66.180 113.810 ;
        RECT 77.600 118.930 77.880 119.210 ;
        RECT 78.400 118.930 78.680 119.210 ;
        RECT 77.600 113.530 77.880 113.810 ;
        RECT 78.400 113.530 78.680 113.810 ;
        RECT 34.150 90.210 34.830 90.890 ;
        RECT 39.450 90.210 40.130 90.890 ;
        RECT 46.750 90.210 47.430 90.890 ;
        RECT 52.850 90.210 53.530 90.890 ;
        RECT 60.250 90.210 60.930 90.890 ;
        RECT 65.250 90.210 65.930 90.890 ;
        RECT 34.150 87.310 34.830 87.990 ;
        RECT 39.450 87.310 40.130 87.990 ;
        RECT 46.750 87.310 47.430 87.990 ;
        RECT 52.850 87.310 53.530 87.990 ;
        RECT 60.250 87.310 60.930 87.990 ;
        RECT 65.250 87.310 65.930 87.990 ;
      LAYER met3 ;
        RECT 26.765 137.820 84.665 139.620 ;
        RECT 82.615 133.470 84.665 137.820 ;
        RECT 25.565 132.320 84.665 133.470 ;
        RECT 82.615 130.520 84.665 132.320 ;
        RECT 27.515 129.420 84.665 130.520 ;
        RECT 82.615 124.720 84.665 129.420 ;
        RECT 27.115 123.820 84.665 124.720 ;
        RECT 82.615 120.170 84.665 123.820 ;
        RECT 16.365 118.370 84.665 120.170 ;
        RECT 82.615 114.520 84.665 118.370 ;
        RECT 18.215 112.820 84.665 114.520 ;
        RECT 33.890 87.150 66.190 93.250 ;
      LAYER via3 ;
        RECT 83.025 113.240 84.145 113.960 ;
        RECT 64.385 88.740 64.705 89.060 ;
      LAYER met4 ;
        RECT 82.430 89.400 84.460 114.270 ;
        RECT 64.130 88.480 84.460 89.400 ;
        RECT 82.430 87.430 84.460 88.480 ;
    END
  END VDD
  PIN Vout
    ANTENNADIFFAREA 75.400002 ;
    PORT
      LAYER li1 ;
        RECT 19.790 119.920 24.830 120.090 ;
        RECT 25.970 119.920 31.010 120.090 ;
        RECT 32.150 119.920 37.190 120.090 ;
        RECT 38.330 119.920 43.370 120.090 ;
        RECT 44.510 119.920 49.550 120.090 ;
        RECT 50.690 119.920 55.730 120.090 ;
        RECT 56.870 119.920 61.910 120.090 ;
        RECT 63.050 119.920 68.090 120.090 ;
        RECT 69.230 119.920 74.270 120.090 ;
        RECT 75.410 119.920 80.450 120.090 ;
        RECT 19.790 117.220 24.830 117.390 ;
        RECT 25.970 117.220 31.010 117.390 ;
        RECT 32.150 117.220 37.190 117.390 ;
        RECT 38.330 117.220 43.370 117.390 ;
        RECT 44.510 117.220 49.550 117.390 ;
        RECT 50.690 117.220 55.730 117.390 ;
        RECT 56.870 117.220 61.910 117.390 ;
        RECT 63.050 117.220 68.090 117.390 ;
        RECT 69.230 117.220 74.270 117.390 ;
        RECT 75.410 117.220 80.450 117.390 ;
        RECT 19.790 114.520 24.830 114.690 ;
        RECT 25.970 114.520 31.010 114.690 ;
        RECT 32.150 114.520 37.190 114.690 ;
        RECT 38.330 114.520 43.370 114.690 ;
        RECT 44.510 114.520 49.550 114.690 ;
        RECT 50.690 114.520 55.730 114.690 ;
        RECT 56.870 114.520 61.910 114.690 ;
        RECT 63.050 114.520 68.090 114.690 ;
        RECT 69.230 114.520 74.270 114.690 ;
        RECT 75.410 114.520 80.450 114.690 ;
        RECT 19.790 111.820 24.830 111.990 ;
        RECT 25.970 111.820 31.010 111.990 ;
        RECT 32.150 111.820 37.190 111.990 ;
        RECT 38.330 111.820 43.370 111.990 ;
        RECT 44.510 111.820 49.550 111.990 ;
        RECT 50.690 111.820 55.730 111.990 ;
        RECT 56.870 111.820 61.910 111.990 ;
        RECT 63.050 111.820 68.090 111.990 ;
        RECT 69.230 111.820 74.270 111.990 ;
        RECT 75.410 111.820 80.450 111.990 ;
        RECT 32.245 103.710 37.285 103.880 ;
        RECT 38.335 103.710 43.375 103.880 ;
        RECT 44.425 103.710 49.465 103.880 ;
        RECT 50.515 103.710 55.555 103.880 ;
        RECT 56.605 103.710 61.645 103.880 ;
        RECT 62.695 103.710 67.735 103.880 ;
        RECT 32.245 100.610 37.285 100.780 ;
        RECT 38.335 100.610 43.375 100.780 ;
        RECT 44.425 100.610 49.465 100.780 ;
        RECT 50.515 100.610 55.555 100.780 ;
        RECT 56.605 100.610 61.645 100.780 ;
        RECT 62.695 100.610 67.735 100.780 ;
      LAYER mcon ;
        RECT 19.885 119.920 20.055 120.090 ;
        RECT 20.245 119.920 20.415 120.090 ;
        RECT 20.605 119.920 20.775 120.090 ;
        RECT 20.965 119.920 21.135 120.090 ;
        RECT 21.325 119.920 21.495 120.090 ;
        RECT 21.685 119.920 21.855 120.090 ;
        RECT 22.045 119.920 22.215 120.090 ;
        RECT 22.405 119.920 22.575 120.090 ;
        RECT 22.765 119.920 22.935 120.090 ;
        RECT 23.125 119.920 23.295 120.090 ;
        RECT 23.485 119.920 23.655 120.090 ;
        RECT 23.845 119.920 24.015 120.090 ;
        RECT 24.205 119.920 24.375 120.090 ;
        RECT 24.565 119.920 24.735 120.090 ;
        RECT 26.065 119.920 26.235 120.090 ;
        RECT 26.425 119.920 26.595 120.090 ;
        RECT 26.785 119.920 26.955 120.090 ;
        RECT 27.145 119.920 27.315 120.090 ;
        RECT 27.505 119.920 27.675 120.090 ;
        RECT 27.865 119.920 28.035 120.090 ;
        RECT 28.225 119.920 28.395 120.090 ;
        RECT 28.585 119.920 28.755 120.090 ;
        RECT 28.945 119.920 29.115 120.090 ;
        RECT 29.305 119.920 29.475 120.090 ;
        RECT 29.665 119.920 29.835 120.090 ;
        RECT 30.025 119.920 30.195 120.090 ;
        RECT 30.385 119.920 30.555 120.090 ;
        RECT 30.745 119.920 30.915 120.090 ;
        RECT 32.245 119.920 32.415 120.090 ;
        RECT 32.605 119.920 32.775 120.090 ;
        RECT 32.965 119.920 33.135 120.090 ;
        RECT 33.325 119.920 33.495 120.090 ;
        RECT 33.685 119.920 33.855 120.090 ;
        RECT 34.045 119.920 34.215 120.090 ;
        RECT 34.405 119.920 34.575 120.090 ;
        RECT 34.765 119.920 34.935 120.090 ;
        RECT 35.125 119.920 35.295 120.090 ;
        RECT 35.485 119.920 35.655 120.090 ;
        RECT 35.845 119.920 36.015 120.090 ;
        RECT 36.205 119.920 36.375 120.090 ;
        RECT 36.565 119.920 36.735 120.090 ;
        RECT 36.925 119.920 37.095 120.090 ;
        RECT 38.425 119.920 38.595 120.090 ;
        RECT 38.785 119.920 38.955 120.090 ;
        RECT 39.145 119.920 39.315 120.090 ;
        RECT 39.505 119.920 39.675 120.090 ;
        RECT 39.865 119.920 40.035 120.090 ;
        RECT 40.225 119.920 40.395 120.090 ;
        RECT 40.585 119.920 40.755 120.090 ;
        RECT 40.945 119.920 41.115 120.090 ;
        RECT 41.305 119.920 41.475 120.090 ;
        RECT 41.665 119.920 41.835 120.090 ;
        RECT 42.025 119.920 42.195 120.090 ;
        RECT 42.385 119.920 42.555 120.090 ;
        RECT 42.745 119.920 42.915 120.090 ;
        RECT 43.105 119.920 43.275 120.090 ;
        RECT 44.605 119.920 44.775 120.090 ;
        RECT 44.965 119.920 45.135 120.090 ;
        RECT 45.325 119.920 45.495 120.090 ;
        RECT 45.685 119.920 45.855 120.090 ;
        RECT 46.045 119.920 46.215 120.090 ;
        RECT 46.405 119.920 46.575 120.090 ;
        RECT 46.765 119.920 46.935 120.090 ;
        RECT 47.125 119.920 47.295 120.090 ;
        RECT 47.485 119.920 47.655 120.090 ;
        RECT 47.845 119.920 48.015 120.090 ;
        RECT 48.205 119.920 48.375 120.090 ;
        RECT 48.565 119.920 48.735 120.090 ;
        RECT 48.925 119.920 49.095 120.090 ;
        RECT 49.285 119.920 49.455 120.090 ;
        RECT 50.785 119.920 50.955 120.090 ;
        RECT 51.145 119.920 51.315 120.090 ;
        RECT 51.505 119.920 51.675 120.090 ;
        RECT 51.865 119.920 52.035 120.090 ;
        RECT 52.225 119.920 52.395 120.090 ;
        RECT 52.585 119.920 52.755 120.090 ;
        RECT 52.945 119.920 53.115 120.090 ;
        RECT 53.305 119.920 53.475 120.090 ;
        RECT 53.665 119.920 53.835 120.090 ;
        RECT 54.025 119.920 54.195 120.090 ;
        RECT 54.385 119.920 54.555 120.090 ;
        RECT 54.745 119.920 54.915 120.090 ;
        RECT 55.105 119.920 55.275 120.090 ;
        RECT 55.465 119.920 55.635 120.090 ;
        RECT 56.965 119.920 57.135 120.090 ;
        RECT 57.325 119.920 57.495 120.090 ;
        RECT 57.685 119.920 57.855 120.090 ;
        RECT 58.045 119.920 58.215 120.090 ;
        RECT 58.405 119.920 58.575 120.090 ;
        RECT 58.765 119.920 58.935 120.090 ;
        RECT 59.125 119.920 59.295 120.090 ;
        RECT 59.485 119.920 59.655 120.090 ;
        RECT 59.845 119.920 60.015 120.090 ;
        RECT 60.205 119.920 60.375 120.090 ;
        RECT 60.565 119.920 60.735 120.090 ;
        RECT 60.925 119.920 61.095 120.090 ;
        RECT 61.285 119.920 61.455 120.090 ;
        RECT 61.645 119.920 61.815 120.090 ;
        RECT 63.145 119.920 63.315 120.090 ;
        RECT 63.505 119.920 63.675 120.090 ;
        RECT 63.865 119.920 64.035 120.090 ;
        RECT 64.225 119.920 64.395 120.090 ;
        RECT 64.585 119.920 64.755 120.090 ;
        RECT 64.945 119.920 65.115 120.090 ;
        RECT 65.305 119.920 65.475 120.090 ;
        RECT 65.665 119.920 65.835 120.090 ;
        RECT 66.025 119.920 66.195 120.090 ;
        RECT 66.385 119.920 66.555 120.090 ;
        RECT 66.745 119.920 66.915 120.090 ;
        RECT 67.105 119.920 67.275 120.090 ;
        RECT 67.465 119.920 67.635 120.090 ;
        RECT 67.825 119.920 67.995 120.090 ;
        RECT 69.325 119.920 69.495 120.090 ;
        RECT 69.685 119.920 69.855 120.090 ;
        RECT 70.045 119.920 70.215 120.090 ;
        RECT 70.405 119.920 70.575 120.090 ;
        RECT 70.765 119.920 70.935 120.090 ;
        RECT 71.125 119.920 71.295 120.090 ;
        RECT 71.485 119.920 71.655 120.090 ;
        RECT 71.845 119.920 72.015 120.090 ;
        RECT 72.205 119.920 72.375 120.090 ;
        RECT 72.565 119.920 72.735 120.090 ;
        RECT 72.925 119.920 73.095 120.090 ;
        RECT 73.285 119.920 73.455 120.090 ;
        RECT 73.645 119.920 73.815 120.090 ;
        RECT 74.005 119.920 74.175 120.090 ;
        RECT 75.505 119.920 75.675 120.090 ;
        RECT 75.865 119.920 76.035 120.090 ;
        RECT 76.225 119.920 76.395 120.090 ;
        RECT 76.585 119.920 76.755 120.090 ;
        RECT 76.945 119.920 77.115 120.090 ;
        RECT 77.305 119.920 77.475 120.090 ;
        RECT 77.665 119.920 77.835 120.090 ;
        RECT 78.025 119.920 78.195 120.090 ;
        RECT 78.385 119.920 78.555 120.090 ;
        RECT 78.745 119.920 78.915 120.090 ;
        RECT 79.105 119.920 79.275 120.090 ;
        RECT 79.465 119.920 79.635 120.090 ;
        RECT 79.825 119.920 79.995 120.090 ;
        RECT 80.185 119.920 80.355 120.090 ;
        RECT 19.885 117.220 20.055 117.390 ;
        RECT 20.245 117.220 20.415 117.390 ;
        RECT 20.605 117.220 20.775 117.390 ;
        RECT 20.965 117.220 21.135 117.390 ;
        RECT 21.325 117.220 21.495 117.390 ;
        RECT 21.685 117.220 21.855 117.390 ;
        RECT 22.045 117.220 22.215 117.390 ;
        RECT 22.405 117.220 22.575 117.390 ;
        RECT 22.765 117.220 22.935 117.390 ;
        RECT 23.125 117.220 23.295 117.390 ;
        RECT 23.485 117.220 23.655 117.390 ;
        RECT 23.845 117.220 24.015 117.390 ;
        RECT 24.205 117.220 24.375 117.390 ;
        RECT 24.565 117.220 24.735 117.390 ;
        RECT 26.065 117.220 26.235 117.390 ;
        RECT 26.425 117.220 26.595 117.390 ;
        RECT 26.785 117.220 26.955 117.390 ;
        RECT 27.145 117.220 27.315 117.390 ;
        RECT 27.505 117.220 27.675 117.390 ;
        RECT 27.865 117.220 28.035 117.390 ;
        RECT 28.225 117.220 28.395 117.390 ;
        RECT 28.585 117.220 28.755 117.390 ;
        RECT 28.945 117.220 29.115 117.390 ;
        RECT 29.305 117.220 29.475 117.390 ;
        RECT 29.665 117.220 29.835 117.390 ;
        RECT 30.025 117.220 30.195 117.390 ;
        RECT 30.385 117.220 30.555 117.390 ;
        RECT 30.745 117.220 30.915 117.390 ;
        RECT 32.245 117.220 32.415 117.390 ;
        RECT 32.605 117.220 32.775 117.390 ;
        RECT 32.965 117.220 33.135 117.390 ;
        RECT 33.325 117.220 33.495 117.390 ;
        RECT 33.685 117.220 33.855 117.390 ;
        RECT 34.045 117.220 34.215 117.390 ;
        RECT 34.405 117.220 34.575 117.390 ;
        RECT 34.765 117.220 34.935 117.390 ;
        RECT 35.125 117.220 35.295 117.390 ;
        RECT 35.485 117.220 35.655 117.390 ;
        RECT 35.845 117.220 36.015 117.390 ;
        RECT 36.205 117.220 36.375 117.390 ;
        RECT 36.565 117.220 36.735 117.390 ;
        RECT 36.925 117.220 37.095 117.390 ;
        RECT 38.425 117.220 38.595 117.390 ;
        RECT 38.785 117.220 38.955 117.390 ;
        RECT 39.145 117.220 39.315 117.390 ;
        RECT 39.505 117.220 39.675 117.390 ;
        RECT 39.865 117.220 40.035 117.390 ;
        RECT 40.225 117.220 40.395 117.390 ;
        RECT 40.585 117.220 40.755 117.390 ;
        RECT 40.945 117.220 41.115 117.390 ;
        RECT 41.305 117.220 41.475 117.390 ;
        RECT 41.665 117.220 41.835 117.390 ;
        RECT 42.025 117.220 42.195 117.390 ;
        RECT 42.385 117.220 42.555 117.390 ;
        RECT 42.745 117.220 42.915 117.390 ;
        RECT 43.105 117.220 43.275 117.390 ;
        RECT 44.605 117.220 44.775 117.390 ;
        RECT 44.965 117.220 45.135 117.390 ;
        RECT 45.325 117.220 45.495 117.390 ;
        RECT 45.685 117.220 45.855 117.390 ;
        RECT 46.045 117.220 46.215 117.390 ;
        RECT 46.405 117.220 46.575 117.390 ;
        RECT 46.765 117.220 46.935 117.390 ;
        RECT 47.125 117.220 47.295 117.390 ;
        RECT 47.485 117.220 47.655 117.390 ;
        RECT 47.845 117.220 48.015 117.390 ;
        RECT 48.205 117.220 48.375 117.390 ;
        RECT 48.565 117.220 48.735 117.390 ;
        RECT 48.925 117.220 49.095 117.390 ;
        RECT 49.285 117.220 49.455 117.390 ;
        RECT 50.785 117.220 50.955 117.390 ;
        RECT 51.145 117.220 51.315 117.390 ;
        RECT 51.505 117.220 51.675 117.390 ;
        RECT 51.865 117.220 52.035 117.390 ;
        RECT 52.225 117.220 52.395 117.390 ;
        RECT 52.585 117.220 52.755 117.390 ;
        RECT 52.945 117.220 53.115 117.390 ;
        RECT 53.305 117.220 53.475 117.390 ;
        RECT 53.665 117.220 53.835 117.390 ;
        RECT 54.025 117.220 54.195 117.390 ;
        RECT 54.385 117.220 54.555 117.390 ;
        RECT 54.745 117.220 54.915 117.390 ;
        RECT 55.105 117.220 55.275 117.390 ;
        RECT 55.465 117.220 55.635 117.390 ;
        RECT 56.965 117.220 57.135 117.390 ;
        RECT 57.325 117.220 57.495 117.390 ;
        RECT 57.685 117.220 57.855 117.390 ;
        RECT 58.045 117.220 58.215 117.390 ;
        RECT 58.405 117.220 58.575 117.390 ;
        RECT 58.765 117.220 58.935 117.390 ;
        RECT 59.125 117.220 59.295 117.390 ;
        RECT 59.485 117.220 59.655 117.390 ;
        RECT 59.845 117.220 60.015 117.390 ;
        RECT 60.205 117.220 60.375 117.390 ;
        RECT 60.565 117.220 60.735 117.390 ;
        RECT 60.925 117.220 61.095 117.390 ;
        RECT 61.285 117.220 61.455 117.390 ;
        RECT 61.645 117.220 61.815 117.390 ;
        RECT 63.145 117.220 63.315 117.390 ;
        RECT 63.505 117.220 63.675 117.390 ;
        RECT 63.865 117.220 64.035 117.390 ;
        RECT 64.225 117.220 64.395 117.390 ;
        RECT 64.585 117.220 64.755 117.390 ;
        RECT 64.945 117.220 65.115 117.390 ;
        RECT 65.305 117.220 65.475 117.390 ;
        RECT 65.665 117.220 65.835 117.390 ;
        RECT 66.025 117.220 66.195 117.390 ;
        RECT 66.385 117.220 66.555 117.390 ;
        RECT 66.745 117.220 66.915 117.390 ;
        RECT 67.105 117.220 67.275 117.390 ;
        RECT 67.465 117.220 67.635 117.390 ;
        RECT 67.825 117.220 67.995 117.390 ;
        RECT 69.325 117.220 69.495 117.390 ;
        RECT 69.685 117.220 69.855 117.390 ;
        RECT 70.045 117.220 70.215 117.390 ;
        RECT 70.405 117.220 70.575 117.390 ;
        RECT 70.765 117.220 70.935 117.390 ;
        RECT 71.125 117.220 71.295 117.390 ;
        RECT 71.485 117.220 71.655 117.390 ;
        RECT 71.845 117.220 72.015 117.390 ;
        RECT 72.205 117.220 72.375 117.390 ;
        RECT 72.565 117.220 72.735 117.390 ;
        RECT 72.925 117.220 73.095 117.390 ;
        RECT 73.285 117.220 73.455 117.390 ;
        RECT 73.645 117.220 73.815 117.390 ;
        RECT 74.005 117.220 74.175 117.390 ;
        RECT 75.505 117.220 75.675 117.390 ;
        RECT 75.865 117.220 76.035 117.390 ;
        RECT 76.225 117.220 76.395 117.390 ;
        RECT 76.585 117.220 76.755 117.390 ;
        RECT 76.945 117.220 77.115 117.390 ;
        RECT 77.305 117.220 77.475 117.390 ;
        RECT 77.665 117.220 77.835 117.390 ;
        RECT 78.025 117.220 78.195 117.390 ;
        RECT 78.385 117.220 78.555 117.390 ;
        RECT 78.745 117.220 78.915 117.390 ;
        RECT 79.105 117.220 79.275 117.390 ;
        RECT 79.465 117.220 79.635 117.390 ;
        RECT 79.825 117.220 79.995 117.390 ;
        RECT 80.185 117.220 80.355 117.390 ;
        RECT 19.885 114.520 20.055 114.690 ;
        RECT 20.245 114.520 20.415 114.690 ;
        RECT 20.605 114.520 20.775 114.690 ;
        RECT 20.965 114.520 21.135 114.690 ;
        RECT 21.325 114.520 21.495 114.690 ;
        RECT 21.685 114.520 21.855 114.690 ;
        RECT 22.045 114.520 22.215 114.690 ;
        RECT 22.405 114.520 22.575 114.690 ;
        RECT 22.765 114.520 22.935 114.690 ;
        RECT 23.125 114.520 23.295 114.690 ;
        RECT 23.485 114.520 23.655 114.690 ;
        RECT 23.845 114.520 24.015 114.690 ;
        RECT 24.205 114.520 24.375 114.690 ;
        RECT 24.565 114.520 24.735 114.690 ;
        RECT 26.065 114.520 26.235 114.690 ;
        RECT 26.425 114.520 26.595 114.690 ;
        RECT 26.785 114.520 26.955 114.690 ;
        RECT 27.145 114.520 27.315 114.690 ;
        RECT 27.505 114.520 27.675 114.690 ;
        RECT 27.865 114.520 28.035 114.690 ;
        RECT 28.225 114.520 28.395 114.690 ;
        RECT 28.585 114.520 28.755 114.690 ;
        RECT 28.945 114.520 29.115 114.690 ;
        RECT 29.305 114.520 29.475 114.690 ;
        RECT 29.665 114.520 29.835 114.690 ;
        RECT 30.025 114.520 30.195 114.690 ;
        RECT 30.385 114.520 30.555 114.690 ;
        RECT 30.745 114.520 30.915 114.690 ;
        RECT 32.245 114.520 32.415 114.690 ;
        RECT 32.605 114.520 32.775 114.690 ;
        RECT 32.965 114.520 33.135 114.690 ;
        RECT 33.325 114.520 33.495 114.690 ;
        RECT 33.685 114.520 33.855 114.690 ;
        RECT 34.045 114.520 34.215 114.690 ;
        RECT 34.405 114.520 34.575 114.690 ;
        RECT 34.765 114.520 34.935 114.690 ;
        RECT 35.125 114.520 35.295 114.690 ;
        RECT 35.485 114.520 35.655 114.690 ;
        RECT 35.845 114.520 36.015 114.690 ;
        RECT 36.205 114.520 36.375 114.690 ;
        RECT 36.565 114.520 36.735 114.690 ;
        RECT 36.925 114.520 37.095 114.690 ;
        RECT 38.425 114.520 38.595 114.690 ;
        RECT 38.785 114.520 38.955 114.690 ;
        RECT 39.145 114.520 39.315 114.690 ;
        RECT 39.505 114.520 39.675 114.690 ;
        RECT 39.865 114.520 40.035 114.690 ;
        RECT 40.225 114.520 40.395 114.690 ;
        RECT 40.585 114.520 40.755 114.690 ;
        RECT 40.945 114.520 41.115 114.690 ;
        RECT 41.305 114.520 41.475 114.690 ;
        RECT 41.665 114.520 41.835 114.690 ;
        RECT 42.025 114.520 42.195 114.690 ;
        RECT 42.385 114.520 42.555 114.690 ;
        RECT 42.745 114.520 42.915 114.690 ;
        RECT 43.105 114.520 43.275 114.690 ;
        RECT 44.605 114.520 44.775 114.690 ;
        RECT 44.965 114.520 45.135 114.690 ;
        RECT 45.325 114.520 45.495 114.690 ;
        RECT 45.685 114.520 45.855 114.690 ;
        RECT 46.045 114.520 46.215 114.690 ;
        RECT 46.405 114.520 46.575 114.690 ;
        RECT 46.765 114.520 46.935 114.690 ;
        RECT 47.125 114.520 47.295 114.690 ;
        RECT 47.485 114.520 47.655 114.690 ;
        RECT 47.845 114.520 48.015 114.690 ;
        RECT 48.205 114.520 48.375 114.690 ;
        RECT 48.565 114.520 48.735 114.690 ;
        RECT 48.925 114.520 49.095 114.690 ;
        RECT 49.285 114.520 49.455 114.690 ;
        RECT 50.785 114.520 50.955 114.690 ;
        RECT 51.145 114.520 51.315 114.690 ;
        RECT 51.505 114.520 51.675 114.690 ;
        RECT 51.865 114.520 52.035 114.690 ;
        RECT 52.225 114.520 52.395 114.690 ;
        RECT 52.585 114.520 52.755 114.690 ;
        RECT 52.945 114.520 53.115 114.690 ;
        RECT 53.305 114.520 53.475 114.690 ;
        RECT 53.665 114.520 53.835 114.690 ;
        RECT 54.025 114.520 54.195 114.690 ;
        RECT 54.385 114.520 54.555 114.690 ;
        RECT 54.745 114.520 54.915 114.690 ;
        RECT 55.105 114.520 55.275 114.690 ;
        RECT 55.465 114.520 55.635 114.690 ;
        RECT 56.965 114.520 57.135 114.690 ;
        RECT 57.325 114.520 57.495 114.690 ;
        RECT 57.685 114.520 57.855 114.690 ;
        RECT 58.045 114.520 58.215 114.690 ;
        RECT 58.405 114.520 58.575 114.690 ;
        RECT 58.765 114.520 58.935 114.690 ;
        RECT 59.125 114.520 59.295 114.690 ;
        RECT 59.485 114.520 59.655 114.690 ;
        RECT 59.845 114.520 60.015 114.690 ;
        RECT 60.205 114.520 60.375 114.690 ;
        RECT 60.565 114.520 60.735 114.690 ;
        RECT 60.925 114.520 61.095 114.690 ;
        RECT 61.285 114.520 61.455 114.690 ;
        RECT 61.645 114.520 61.815 114.690 ;
        RECT 63.145 114.520 63.315 114.690 ;
        RECT 63.505 114.520 63.675 114.690 ;
        RECT 63.865 114.520 64.035 114.690 ;
        RECT 64.225 114.520 64.395 114.690 ;
        RECT 64.585 114.520 64.755 114.690 ;
        RECT 64.945 114.520 65.115 114.690 ;
        RECT 65.305 114.520 65.475 114.690 ;
        RECT 65.665 114.520 65.835 114.690 ;
        RECT 66.025 114.520 66.195 114.690 ;
        RECT 66.385 114.520 66.555 114.690 ;
        RECT 66.745 114.520 66.915 114.690 ;
        RECT 67.105 114.520 67.275 114.690 ;
        RECT 67.465 114.520 67.635 114.690 ;
        RECT 67.825 114.520 67.995 114.690 ;
        RECT 69.325 114.520 69.495 114.690 ;
        RECT 69.685 114.520 69.855 114.690 ;
        RECT 70.045 114.520 70.215 114.690 ;
        RECT 70.405 114.520 70.575 114.690 ;
        RECT 70.765 114.520 70.935 114.690 ;
        RECT 71.125 114.520 71.295 114.690 ;
        RECT 71.485 114.520 71.655 114.690 ;
        RECT 71.845 114.520 72.015 114.690 ;
        RECT 72.205 114.520 72.375 114.690 ;
        RECT 72.565 114.520 72.735 114.690 ;
        RECT 72.925 114.520 73.095 114.690 ;
        RECT 73.285 114.520 73.455 114.690 ;
        RECT 73.645 114.520 73.815 114.690 ;
        RECT 74.005 114.520 74.175 114.690 ;
        RECT 75.505 114.520 75.675 114.690 ;
        RECT 75.865 114.520 76.035 114.690 ;
        RECT 76.225 114.520 76.395 114.690 ;
        RECT 76.585 114.520 76.755 114.690 ;
        RECT 76.945 114.520 77.115 114.690 ;
        RECT 77.305 114.520 77.475 114.690 ;
        RECT 77.665 114.520 77.835 114.690 ;
        RECT 78.025 114.520 78.195 114.690 ;
        RECT 78.385 114.520 78.555 114.690 ;
        RECT 78.745 114.520 78.915 114.690 ;
        RECT 79.105 114.520 79.275 114.690 ;
        RECT 79.465 114.520 79.635 114.690 ;
        RECT 79.825 114.520 79.995 114.690 ;
        RECT 80.185 114.520 80.355 114.690 ;
        RECT 19.885 111.820 20.055 111.990 ;
        RECT 20.245 111.820 20.415 111.990 ;
        RECT 20.605 111.820 20.775 111.990 ;
        RECT 20.965 111.820 21.135 111.990 ;
        RECT 21.325 111.820 21.495 111.990 ;
        RECT 21.685 111.820 21.855 111.990 ;
        RECT 22.045 111.820 22.215 111.990 ;
        RECT 22.405 111.820 22.575 111.990 ;
        RECT 22.765 111.820 22.935 111.990 ;
        RECT 23.125 111.820 23.295 111.990 ;
        RECT 23.485 111.820 23.655 111.990 ;
        RECT 23.845 111.820 24.015 111.990 ;
        RECT 24.205 111.820 24.375 111.990 ;
        RECT 24.565 111.820 24.735 111.990 ;
        RECT 26.065 111.820 26.235 111.990 ;
        RECT 26.425 111.820 26.595 111.990 ;
        RECT 26.785 111.820 26.955 111.990 ;
        RECT 27.145 111.820 27.315 111.990 ;
        RECT 27.505 111.820 27.675 111.990 ;
        RECT 27.865 111.820 28.035 111.990 ;
        RECT 28.225 111.820 28.395 111.990 ;
        RECT 28.585 111.820 28.755 111.990 ;
        RECT 28.945 111.820 29.115 111.990 ;
        RECT 29.305 111.820 29.475 111.990 ;
        RECT 29.665 111.820 29.835 111.990 ;
        RECT 30.025 111.820 30.195 111.990 ;
        RECT 30.385 111.820 30.555 111.990 ;
        RECT 30.745 111.820 30.915 111.990 ;
        RECT 32.245 111.820 32.415 111.990 ;
        RECT 32.605 111.820 32.775 111.990 ;
        RECT 32.965 111.820 33.135 111.990 ;
        RECT 33.325 111.820 33.495 111.990 ;
        RECT 33.685 111.820 33.855 111.990 ;
        RECT 34.045 111.820 34.215 111.990 ;
        RECT 34.405 111.820 34.575 111.990 ;
        RECT 34.765 111.820 34.935 111.990 ;
        RECT 35.125 111.820 35.295 111.990 ;
        RECT 35.485 111.820 35.655 111.990 ;
        RECT 35.845 111.820 36.015 111.990 ;
        RECT 36.205 111.820 36.375 111.990 ;
        RECT 36.565 111.820 36.735 111.990 ;
        RECT 36.925 111.820 37.095 111.990 ;
        RECT 38.425 111.820 38.595 111.990 ;
        RECT 38.785 111.820 38.955 111.990 ;
        RECT 39.145 111.820 39.315 111.990 ;
        RECT 39.505 111.820 39.675 111.990 ;
        RECT 39.865 111.820 40.035 111.990 ;
        RECT 40.225 111.820 40.395 111.990 ;
        RECT 40.585 111.820 40.755 111.990 ;
        RECT 40.945 111.820 41.115 111.990 ;
        RECT 41.305 111.820 41.475 111.990 ;
        RECT 41.665 111.820 41.835 111.990 ;
        RECT 42.025 111.820 42.195 111.990 ;
        RECT 42.385 111.820 42.555 111.990 ;
        RECT 42.745 111.820 42.915 111.990 ;
        RECT 43.105 111.820 43.275 111.990 ;
        RECT 44.605 111.820 44.775 111.990 ;
        RECT 44.965 111.820 45.135 111.990 ;
        RECT 45.325 111.820 45.495 111.990 ;
        RECT 45.685 111.820 45.855 111.990 ;
        RECT 46.045 111.820 46.215 111.990 ;
        RECT 46.405 111.820 46.575 111.990 ;
        RECT 46.765 111.820 46.935 111.990 ;
        RECT 47.125 111.820 47.295 111.990 ;
        RECT 47.485 111.820 47.655 111.990 ;
        RECT 47.845 111.820 48.015 111.990 ;
        RECT 48.205 111.820 48.375 111.990 ;
        RECT 48.565 111.820 48.735 111.990 ;
        RECT 48.925 111.820 49.095 111.990 ;
        RECT 49.285 111.820 49.455 111.990 ;
        RECT 50.785 111.820 50.955 111.990 ;
        RECT 51.145 111.820 51.315 111.990 ;
        RECT 51.505 111.820 51.675 111.990 ;
        RECT 51.865 111.820 52.035 111.990 ;
        RECT 52.225 111.820 52.395 111.990 ;
        RECT 52.585 111.820 52.755 111.990 ;
        RECT 52.945 111.820 53.115 111.990 ;
        RECT 53.305 111.820 53.475 111.990 ;
        RECT 53.665 111.820 53.835 111.990 ;
        RECT 54.025 111.820 54.195 111.990 ;
        RECT 54.385 111.820 54.555 111.990 ;
        RECT 54.745 111.820 54.915 111.990 ;
        RECT 55.105 111.820 55.275 111.990 ;
        RECT 55.465 111.820 55.635 111.990 ;
        RECT 56.965 111.820 57.135 111.990 ;
        RECT 57.325 111.820 57.495 111.990 ;
        RECT 57.685 111.820 57.855 111.990 ;
        RECT 58.045 111.820 58.215 111.990 ;
        RECT 58.405 111.820 58.575 111.990 ;
        RECT 58.765 111.820 58.935 111.990 ;
        RECT 59.125 111.820 59.295 111.990 ;
        RECT 59.485 111.820 59.655 111.990 ;
        RECT 59.845 111.820 60.015 111.990 ;
        RECT 60.205 111.820 60.375 111.990 ;
        RECT 60.565 111.820 60.735 111.990 ;
        RECT 60.925 111.820 61.095 111.990 ;
        RECT 61.285 111.820 61.455 111.990 ;
        RECT 61.645 111.820 61.815 111.990 ;
        RECT 63.145 111.820 63.315 111.990 ;
        RECT 63.505 111.820 63.675 111.990 ;
        RECT 63.865 111.820 64.035 111.990 ;
        RECT 64.225 111.820 64.395 111.990 ;
        RECT 64.585 111.820 64.755 111.990 ;
        RECT 64.945 111.820 65.115 111.990 ;
        RECT 65.305 111.820 65.475 111.990 ;
        RECT 65.665 111.820 65.835 111.990 ;
        RECT 66.025 111.820 66.195 111.990 ;
        RECT 66.385 111.820 66.555 111.990 ;
        RECT 66.745 111.820 66.915 111.990 ;
        RECT 67.105 111.820 67.275 111.990 ;
        RECT 67.465 111.820 67.635 111.990 ;
        RECT 67.825 111.820 67.995 111.990 ;
        RECT 69.325 111.820 69.495 111.990 ;
        RECT 69.685 111.820 69.855 111.990 ;
        RECT 70.045 111.820 70.215 111.990 ;
        RECT 70.405 111.820 70.575 111.990 ;
        RECT 70.765 111.820 70.935 111.990 ;
        RECT 71.125 111.820 71.295 111.990 ;
        RECT 71.485 111.820 71.655 111.990 ;
        RECT 71.845 111.820 72.015 111.990 ;
        RECT 72.205 111.820 72.375 111.990 ;
        RECT 72.565 111.820 72.735 111.990 ;
        RECT 72.925 111.820 73.095 111.990 ;
        RECT 73.285 111.820 73.455 111.990 ;
        RECT 73.645 111.820 73.815 111.990 ;
        RECT 74.005 111.820 74.175 111.990 ;
        RECT 75.505 111.820 75.675 111.990 ;
        RECT 75.865 111.820 76.035 111.990 ;
        RECT 76.225 111.820 76.395 111.990 ;
        RECT 76.585 111.820 76.755 111.990 ;
        RECT 76.945 111.820 77.115 111.990 ;
        RECT 77.305 111.820 77.475 111.990 ;
        RECT 77.665 111.820 77.835 111.990 ;
        RECT 78.025 111.820 78.195 111.990 ;
        RECT 78.385 111.820 78.555 111.990 ;
        RECT 78.745 111.820 78.915 111.990 ;
        RECT 79.105 111.820 79.275 111.990 ;
        RECT 79.465 111.820 79.635 111.990 ;
        RECT 79.825 111.820 79.995 111.990 ;
        RECT 80.185 111.820 80.355 111.990 ;
        RECT 32.340 103.710 32.510 103.880 ;
        RECT 32.700 103.710 32.870 103.880 ;
        RECT 33.060 103.710 33.230 103.880 ;
        RECT 33.420 103.710 33.590 103.880 ;
        RECT 33.780 103.710 33.950 103.880 ;
        RECT 34.140 103.710 34.310 103.880 ;
        RECT 34.500 103.710 34.670 103.880 ;
        RECT 34.860 103.710 35.030 103.880 ;
        RECT 35.220 103.710 35.390 103.880 ;
        RECT 35.580 103.710 35.750 103.880 ;
        RECT 35.940 103.710 36.110 103.880 ;
        RECT 36.300 103.710 36.470 103.880 ;
        RECT 36.660 103.710 36.830 103.880 ;
        RECT 37.020 103.710 37.190 103.880 ;
        RECT 38.430 103.710 38.600 103.880 ;
        RECT 38.790 103.710 38.960 103.880 ;
        RECT 39.150 103.710 39.320 103.880 ;
        RECT 39.510 103.710 39.680 103.880 ;
        RECT 39.870 103.710 40.040 103.880 ;
        RECT 40.230 103.710 40.400 103.880 ;
        RECT 40.590 103.710 40.760 103.880 ;
        RECT 40.950 103.710 41.120 103.880 ;
        RECT 41.310 103.710 41.480 103.880 ;
        RECT 41.670 103.710 41.840 103.880 ;
        RECT 42.030 103.710 42.200 103.880 ;
        RECT 42.390 103.710 42.560 103.880 ;
        RECT 42.750 103.710 42.920 103.880 ;
        RECT 43.110 103.710 43.280 103.880 ;
        RECT 44.520 103.710 44.690 103.880 ;
        RECT 44.880 103.710 45.050 103.880 ;
        RECT 45.240 103.710 45.410 103.880 ;
        RECT 45.600 103.710 45.770 103.880 ;
        RECT 45.960 103.710 46.130 103.880 ;
        RECT 46.320 103.710 46.490 103.880 ;
        RECT 46.680 103.710 46.850 103.880 ;
        RECT 47.040 103.710 47.210 103.880 ;
        RECT 47.400 103.710 47.570 103.880 ;
        RECT 47.760 103.710 47.930 103.880 ;
        RECT 48.120 103.710 48.290 103.880 ;
        RECT 48.480 103.710 48.650 103.880 ;
        RECT 48.840 103.710 49.010 103.880 ;
        RECT 49.200 103.710 49.370 103.880 ;
        RECT 50.610 103.710 50.780 103.880 ;
        RECT 50.970 103.710 51.140 103.880 ;
        RECT 51.330 103.710 51.500 103.880 ;
        RECT 51.690 103.710 51.860 103.880 ;
        RECT 52.050 103.710 52.220 103.880 ;
        RECT 52.410 103.710 52.580 103.880 ;
        RECT 52.770 103.710 52.940 103.880 ;
        RECT 53.130 103.710 53.300 103.880 ;
        RECT 53.490 103.710 53.660 103.880 ;
        RECT 53.850 103.710 54.020 103.880 ;
        RECT 54.210 103.710 54.380 103.880 ;
        RECT 54.570 103.710 54.740 103.880 ;
        RECT 54.930 103.710 55.100 103.880 ;
        RECT 55.290 103.710 55.460 103.880 ;
        RECT 56.700 103.710 56.870 103.880 ;
        RECT 57.060 103.710 57.230 103.880 ;
        RECT 57.420 103.710 57.590 103.880 ;
        RECT 57.780 103.710 57.950 103.880 ;
        RECT 58.140 103.710 58.310 103.880 ;
        RECT 58.500 103.710 58.670 103.880 ;
        RECT 58.860 103.710 59.030 103.880 ;
        RECT 59.220 103.710 59.390 103.880 ;
        RECT 59.580 103.710 59.750 103.880 ;
        RECT 59.940 103.710 60.110 103.880 ;
        RECT 60.300 103.710 60.470 103.880 ;
        RECT 60.660 103.710 60.830 103.880 ;
        RECT 61.020 103.710 61.190 103.880 ;
        RECT 61.380 103.710 61.550 103.880 ;
        RECT 62.790 103.710 62.960 103.880 ;
        RECT 63.150 103.710 63.320 103.880 ;
        RECT 63.510 103.710 63.680 103.880 ;
        RECT 63.870 103.710 64.040 103.880 ;
        RECT 64.230 103.710 64.400 103.880 ;
        RECT 64.590 103.710 64.760 103.880 ;
        RECT 64.950 103.710 65.120 103.880 ;
        RECT 65.310 103.710 65.480 103.880 ;
        RECT 65.670 103.710 65.840 103.880 ;
        RECT 66.030 103.710 66.200 103.880 ;
        RECT 66.390 103.710 66.560 103.880 ;
        RECT 66.750 103.710 66.920 103.880 ;
        RECT 67.110 103.710 67.280 103.880 ;
        RECT 67.470 103.710 67.640 103.880 ;
        RECT 32.340 100.610 32.510 100.780 ;
        RECT 32.700 100.610 32.870 100.780 ;
        RECT 33.060 100.610 33.230 100.780 ;
        RECT 33.420 100.610 33.590 100.780 ;
        RECT 33.780 100.610 33.950 100.780 ;
        RECT 34.140 100.610 34.310 100.780 ;
        RECT 34.500 100.610 34.670 100.780 ;
        RECT 34.860 100.610 35.030 100.780 ;
        RECT 35.220 100.610 35.390 100.780 ;
        RECT 35.580 100.610 35.750 100.780 ;
        RECT 35.940 100.610 36.110 100.780 ;
        RECT 36.300 100.610 36.470 100.780 ;
        RECT 36.660 100.610 36.830 100.780 ;
        RECT 37.020 100.610 37.190 100.780 ;
        RECT 38.430 100.610 38.600 100.780 ;
        RECT 38.790 100.610 38.960 100.780 ;
        RECT 39.150 100.610 39.320 100.780 ;
        RECT 39.510 100.610 39.680 100.780 ;
        RECT 39.870 100.610 40.040 100.780 ;
        RECT 40.230 100.610 40.400 100.780 ;
        RECT 40.590 100.610 40.760 100.780 ;
        RECT 40.950 100.610 41.120 100.780 ;
        RECT 41.310 100.610 41.480 100.780 ;
        RECT 41.670 100.610 41.840 100.780 ;
        RECT 42.030 100.610 42.200 100.780 ;
        RECT 42.390 100.610 42.560 100.780 ;
        RECT 42.750 100.610 42.920 100.780 ;
        RECT 43.110 100.610 43.280 100.780 ;
        RECT 44.520 100.610 44.690 100.780 ;
        RECT 44.880 100.610 45.050 100.780 ;
        RECT 45.240 100.610 45.410 100.780 ;
        RECT 45.600 100.610 45.770 100.780 ;
        RECT 45.960 100.610 46.130 100.780 ;
        RECT 46.320 100.610 46.490 100.780 ;
        RECT 46.680 100.610 46.850 100.780 ;
        RECT 47.040 100.610 47.210 100.780 ;
        RECT 47.400 100.610 47.570 100.780 ;
        RECT 47.760 100.610 47.930 100.780 ;
        RECT 48.120 100.610 48.290 100.780 ;
        RECT 48.480 100.610 48.650 100.780 ;
        RECT 48.840 100.610 49.010 100.780 ;
        RECT 49.200 100.610 49.370 100.780 ;
        RECT 50.610 100.610 50.780 100.780 ;
        RECT 50.970 100.610 51.140 100.780 ;
        RECT 51.330 100.610 51.500 100.780 ;
        RECT 51.690 100.610 51.860 100.780 ;
        RECT 52.050 100.610 52.220 100.780 ;
        RECT 52.410 100.610 52.580 100.780 ;
        RECT 52.770 100.610 52.940 100.780 ;
        RECT 53.130 100.610 53.300 100.780 ;
        RECT 53.490 100.610 53.660 100.780 ;
        RECT 53.850 100.610 54.020 100.780 ;
        RECT 54.210 100.610 54.380 100.780 ;
        RECT 54.570 100.610 54.740 100.780 ;
        RECT 54.930 100.610 55.100 100.780 ;
        RECT 55.290 100.610 55.460 100.780 ;
        RECT 56.700 100.610 56.870 100.780 ;
        RECT 57.060 100.610 57.230 100.780 ;
        RECT 57.420 100.610 57.590 100.780 ;
        RECT 57.780 100.610 57.950 100.780 ;
        RECT 58.140 100.610 58.310 100.780 ;
        RECT 58.500 100.610 58.670 100.780 ;
        RECT 58.860 100.610 59.030 100.780 ;
        RECT 59.220 100.610 59.390 100.780 ;
        RECT 59.580 100.610 59.750 100.780 ;
        RECT 59.940 100.610 60.110 100.780 ;
        RECT 60.300 100.610 60.470 100.780 ;
        RECT 60.660 100.610 60.830 100.780 ;
        RECT 61.020 100.610 61.190 100.780 ;
        RECT 61.380 100.610 61.550 100.780 ;
        RECT 62.790 100.610 62.960 100.780 ;
        RECT 63.150 100.610 63.320 100.780 ;
        RECT 63.510 100.610 63.680 100.780 ;
        RECT 63.870 100.610 64.040 100.780 ;
        RECT 64.230 100.610 64.400 100.780 ;
        RECT 64.590 100.610 64.760 100.780 ;
        RECT 64.950 100.610 65.120 100.780 ;
        RECT 65.310 100.610 65.480 100.780 ;
        RECT 65.670 100.610 65.840 100.780 ;
        RECT 66.030 100.610 66.200 100.780 ;
        RECT 66.390 100.610 66.560 100.780 ;
        RECT 66.750 100.610 66.920 100.780 ;
        RECT 67.110 100.610 67.280 100.780 ;
        RECT 67.470 100.610 67.640 100.780 ;
      LAYER met1 ;
        RECT 19.810 120.020 24.810 120.120 ;
        RECT 25.990 120.020 30.990 120.120 ;
        RECT 32.170 120.020 37.170 120.120 ;
        RECT 38.350 120.020 43.350 120.120 ;
        RECT 44.530 120.020 49.530 120.120 ;
        RECT 50.710 120.020 55.710 120.120 ;
        RECT 56.890 120.020 61.890 120.120 ;
        RECT 63.070 120.020 68.070 120.120 ;
        RECT 69.250 120.020 74.250 120.120 ;
        RECT 75.430 120.020 80.430 120.120 ;
        RECT 19.765 119.770 80.515 120.020 ;
        RECT 21.365 119.570 21.865 119.770 ;
        RECT 22.415 119.570 22.915 119.770 ;
        RECT 33.765 119.570 34.265 119.770 ;
        RECT 34.865 119.570 35.365 119.770 ;
        RECT 46.415 119.570 46.915 119.770 ;
        RECT 47.315 119.570 47.815 119.770 ;
        RECT 58.715 119.520 59.215 119.770 ;
        RECT 59.615 119.520 60.115 119.770 ;
        RECT 71.115 119.520 71.615 119.770 ;
        RECT 71.965 119.520 72.465 119.770 ;
        RECT 19.810 117.320 24.810 117.420 ;
        RECT 25.990 117.320 30.990 117.420 ;
        RECT 32.170 117.320 37.170 117.420 ;
        RECT 38.350 117.320 43.350 117.420 ;
        RECT 44.530 117.320 49.530 117.420 ;
        RECT 50.710 117.320 55.710 117.420 ;
        RECT 56.890 117.320 61.890 117.420 ;
        RECT 63.070 117.320 68.070 117.420 ;
        RECT 69.250 117.320 74.250 117.420 ;
        RECT 75.430 117.320 80.430 117.420 ;
        RECT 19.765 117.070 80.515 117.320 ;
        RECT 21.365 116.870 21.865 117.070 ;
        RECT 22.415 116.870 22.915 117.070 ;
        RECT 33.765 116.870 34.265 117.070 ;
        RECT 34.865 116.870 35.365 117.070 ;
        RECT 46.415 116.870 46.915 117.070 ;
        RECT 47.365 116.870 47.865 117.070 ;
        RECT 58.715 116.820 59.215 117.070 ;
        RECT 59.615 116.820 60.115 117.070 ;
        RECT 71.115 116.820 71.615 117.070 ;
        RECT 71.965 116.820 72.465 117.070 ;
        RECT 19.810 114.620 24.810 114.720 ;
        RECT 25.990 114.620 30.990 114.720 ;
        RECT 32.170 114.620 37.170 114.720 ;
        RECT 38.350 114.620 43.350 114.720 ;
        RECT 44.530 114.620 49.530 114.720 ;
        RECT 50.710 114.620 55.710 114.720 ;
        RECT 56.890 114.620 61.890 114.720 ;
        RECT 63.070 114.620 68.070 114.720 ;
        RECT 69.250 114.620 74.250 114.720 ;
        RECT 75.430 114.620 80.430 114.720 ;
        RECT 19.765 114.370 80.515 114.620 ;
        RECT 21.365 114.170 21.865 114.370 ;
        RECT 22.415 114.170 22.915 114.370 ;
        RECT 33.715 114.170 34.215 114.370 ;
        RECT 34.915 114.170 35.415 114.370 ;
        RECT 46.415 114.170 46.915 114.370 ;
        RECT 47.315 114.170 47.815 114.370 ;
        RECT 58.765 114.120 59.265 114.370 ;
        RECT 59.615 114.120 60.115 114.370 ;
        RECT 71.115 114.120 71.615 114.370 ;
        RECT 71.965 114.120 72.465 114.370 ;
        RECT 19.810 111.920 24.810 112.020 ;
        RECT 25.990 111.920 30.990 112.020 ;
        RECT 32.170 111.920 37.170 112.020 ;
        RECT 38.350 111.920 43.350 112.020 ;
        RECT 44.530 111.920 49.530 112.020 ;
        RECT 50.710 111.920 55.710 112.020 ;
        RECT 56.890 111.920 61.890 112.020 ;
        RECT 63.070 111.920 68.070 112.020 ;
        RECT 69.250 111.920 74.250 112.020 ;
        RECT 75.430 111.920 80.430 112.020 ;
        RECT 19.765 111.670 80.515 111.920 ;
        RECT 21.365 111.470 21.865 111.670 ;
        RECT 22.415 111.470 22.915 111.670 ;
        RECT 33.715 111.420 34.215 111.670 ;
        RECT 34.915 111.420 35.415 111.670 ;
        RECT 46.415 111.470 46.915 111.670 ;
        RECT 47.365 111.470 47.865 111.670 ;
        RECT 58.715 111.420 59.215 111.670 ;
        RECT 59.665 111.420 60.165 111.670 ;
        RECT 71.115 111.370 71.615 111.670 ;
        RECT 71.965 111.370 72.465 111.670 ;
        RECT 34.415 104.270 35.965 104.420 ;
        RECT 33.815 103.970 35.965 104.270 ;
        RECT 46.865 103.970 47.365 104.120 ;
        RECT 59.115 103.970 60.215 104.270 ;
        RECT 65.115 103.970 65.615 104.170 ;
        RECT 32.215 103.770 67.815 103.970 ;
        RECT 32.265 103.680 37.265 103.770 ;
        RECT 38.355 103.680 43.355 103.770 ;
        RECT 44.445 103.680 49.445 103.770 ;
        RECT 50.535 103.680 55.535 103.770 ;
        RECT 56.625 103.680 61.625 103.770 ;
        RECT 62.715 103.680 67.715 103.770 ;
        RECT 46.865 100.870 47.365 101.020 ;
        RECT 65.115 100.870 65.615 101.070 ;
        RECT 32.215 100.670 67.815 100.870 ;
        RECT 32.265 100.580 37.265 100.670 ;
        RECT 38.355 100.580 43.355 100.670 ;
        RECT 44.445 100.580 49.445 100.670 ;
        RECT 50.535 100.580 55.535 100.670 ;
        RECT 56.625 100.580 61.625 100.670 ;
        RECT 62.715 100.580 67.715 100.670 ;
      LAYER via ;
        RECT 21.485 119.640 21.745 119.900 ;
        RECT 22.535 119.640 22.795 119.900 ;
        RECT 33.885 119.640 34.145 119.900 ;
        RECT 34.985 119.640 35.245 119.900 ;
        RECT 46.535 119.640 46.795 119.900 ;
        RECT 47.435 119.640 47.695 119.900 ;
        RECT 58.835 119.590 59.095 119.850 ;
        RECT 59.735 119.590 59.995 119.850 ;
        RECT 71.235 119.590 71.495 119.850 ;
        RECT 72.085 119.590 72.345 119.850 ;
        RECT 21.485 116.940 21.745 117.200 ;
        RECT 22.535 116.940 22.795 117.200 ;
        RECT 33.885 116.940 34.145 117.200 ;
        RECT 34.985 116.940 35.245 117.200 ;
        RECT 46.535 116.940 46.795 117.200 ;
        RECT 47.485 116.940 47.745 117.200 ;
        RECT 58.835 116.890 59.095 117.150 ;
        RECT 59.735 116.890 59.995 117.150 ;
        RECT 71.235 116.890 71.495 117.150 ;
        RECT 72.085 116.890 72.345 117.150 ;
        RECT 21.485 114.240 21.745 114.500 ;
        RECT 22.535 114.240 22.795 114.500 ;
        RECT 33.835 114.240 34.095 114.500 ;
        RECT 35.035 114.240 35.295 114.500 ;
        RECT 46.535 114.240 46.795 114.500 ;
        RECT 47.435 114.240 47.695 114.500 ;
        RECT 58.885 114.190 59.145 114.450 ;
        RECT 59.735 114.190 59.995 114.450 ;
        RECT 71.235 114.190 71.495 114.450 ;
        RECT 72.085 114.190 72.345 114.450 ;
        RECT 21.485 111.540 21.745 111.800 ;
        RECT 22.535 111.540 22.795 111.800 ;
        RECT 33.835 111.490 34.095 111.750 ;
        RECT 35.035 111.490 35.295 111.750 ;
        RECT 46.535 111.540 46.795 111.800 ;
        RECT 47.485 111.540 47.745 111.800 ;
        RECT 58.835 111.490 59.095 111.750 ;
        RECT 59.785 111.490 60.045 111.750 ;
        RECT 71.235 111.440 71.495 111.700 ;
        RECT 72.085 111.440 72.345 111.700 ;
        RECT 34.935 103.940 35.195 104.200 ;
        RECT 35.485 103.940 35.745 104.200 ;
        RECT 46.985 103.790 47.245 104.050 ;
        RECT 59.235 103.890 59.495 104.150 ;
        RECT 59.835 103.890 60.095 104.150 ;
        RECT 65.235 103.840 65.495 104.100 ;
        RECT 46.985 100.690 47.245 100.950 ;
        RECT 65.235 100.740 65.495 101.000 ;
      LAYER met2 ;
        RECT 21.415 111.420 22.865 122.220 ;
        RECT 33.765 112.220 35.365 120.120 ;
        RECT 33.765 110.920 35.815 112.220 ;
        RECT 34.865 104.420 35.815 110.920 ;
        RECT 34.415 103.770 35.965 104.420 ;
        RECT 46.415 103.870 47.865 120.420 ;
        RECT 58.715 112.320 60.165 120.420 ;
        RECT 58.715 111.320 60.215 112.320 ;
        RECT 71.065 111.320 72.515 121.770 ;
        RECT 46.915 100.570 47.315 103.870 ;
        RECT 59.115 103.770 60.215 111.320 ;
        RECT 64.915 103.970 66.365 104.220 ;
        RECT 65.165 100.620 65.565 103.970 ;
      LAYER via2 ;
        RECT 21.600 121.405 21.880 121.685 ;
        RECT 22.400 121.405 22.680 121.685 ;
        RECT 71.225 121.230 71.505 121.510 ;
        RECT 72.075 121.230 72.355 121.510 ;
      LAYER met3 ;
        RECT 21.415 121.220 22.865 121.920 ;
        RECT 71.065 121.130 72.525 121.620 ;
      LAYER via3 ;
        RECT 21.580 121.385 21.900 121.705 ;
        RECT 22.380 121.385 22.700 121.705 ;
        RECT 71.205 121.210 71.525 121.530 ;
        RECT 72.055 121.210 72.375 121.530 ;
      LAYER met4 ;
        RECT 13.710 151.320 29.320 157.075 ;
        RECT 32.710 151.320 48.320 157.075 ;
        RECT 51.710 151.320 67.320 157.075 ;
        RECT 70.710 151.320 86.320 157.075 ;
        RECT 13.710 149.520 86.320 151.320 ;
        RECT 13.710 141.465 29.320 149.520 ;
        RECT 30.415 140.420 31.265 149.520 ;
        RECT 32.710 141.465 48.320 149.520 ;
        RECT 51.710 141.465 67.320 149.520 ;
        RECT 21.415 139.470 31.265 140.420 ;
        RECT 68.615 140.520 69.415 149.520 ;
        RECT 70.710 141.465 86.320 149.520 ;
        RECT 68.615 139.870 72.515 140.520 ;
        RECT 21.415 120.170 22.865 139.470 ;
        RECT 71.065 119.120 72.515 139.870 ;
    END
  END Vout
  PIN VSS
    ANTENNADIFFAREA 183.797394 ;
    PORT
      LAYER pwell ;
        RECT 0.000 123.765 15.880 124.195 ;
        RECT 0.000 117.335 0.430 123.765 ;
        RECT 15.450 117.335 15.880 123.765 ;
        RECT 0.000 116.905 15.880 117.335 ;
        RECT 85.300 123.765 101.180 124.195 ;
        RECT 85.300 117.335 85.730 123.765 ;
        RECT 100.750 117.335 101.180 123.765 ;
        RECT 85.300 116.905 101.180 117.335 ;
        RECT 0.000 116.415 15.880 116.845 ;
        RECT 0.000 109.985 0.430 116.415 ;
        RECT 15.450 109.985 15.880 116.415 ;
        RECT 0.000 109.555 15.880 109.985 ;
        RECT 85.300 116.415 101.180 116.845 ;
        RECT 85.300 109.985 85.730 116.415 ;
        RECT 100.750 109.985 101.180 116.415 ;
        RECT 28.465 107.220 72.005 109.580 ;
        RECT 85.300 109.555 101.180 109.985 ;
        RECT 28.465 104.720 72.005 107.080 ;
        RECT 31.265 101.720 68.715 104.580 ;
        RECT 31.265 98.620 68.715 101.480 ;
        RECT 28.465 95.620 72.005 98.480 ;
        RECT 28.465 92.620 72.005 95.480 ;
        RECT 45.040 80.850 55.310 83.710 ;
        RECT 46.140 77.960 54.230 80.850 ;
        RECT 31.465 75.100 68.915 77.960 ;
        RECT 33.860 68.000 34.720 69.100 ;
        RECT 65.710 68.000 66.570 69.100 ;
        RECT 33.860 53.000 34.720 54.100 ;
        RECT 65.710 53.000 66.570 54.100 ;
        RECT 33.860 38.000 34.720 39.100 ;
        RECT 65.710 38.000 66.570 39.100 ;
        RECT 33.860 23.000 34.720 24.100 ;
        RECT 65.710 23.000 66.570 24.100 ;
        RECT 33.860 8.000 34.720 9.100 ;
        RECT 65.710 8.000 66.570 9.100 ;
      LAYER li1 ;
        RECT 0.130 123.895 15.750 124.065 ;
        RECT 0.130 117.205 0.300 123.895 ;
        RECT 6.065 117.205 6.515 117.270 ;
        RECT 15.580 117.205 15.750 123.895 ;
        RECT 0.130 117.035 15.750 117.205 ;
        RECT 85.430 123.895 101.050 124.065 ;
        RECT 85.430 117.205 85.600 123.895 ;
        RECT 100.880 117.205 101.050 123.895 ;
        RECT 85.430 117.035 101.050 117.205 ;
        RECT 6.065 116.715 6.515 117.035 ;
        RECT 92.315 116.715 93.015 117.035 ;
        RECT 0.130 116.545 15.750 116.715 ;
        RECT 0.130 109.855 0.300 116.545 ;
        RECT 15.580 109.855 15.750 116.545 ;
        RECT 0.130 109.685 15.750 109.855 ;
        RECT 85.430 116.545 101.050 116.715 ;
        RECT 85.430 109.855 85.600 116.545 ;
        RECT 100.880 109.855 101.050 116.545 ;
        RECT 85.430 109.685 101.050 109.855 ;
        RECT 5.965 109.170 6.415 109.685 ;
        RECT 7.015 109.170 7.465 109.685 ;
        RECT 28.595 109.280 71.875 109.450 ;
        RECT 92.515 109.320 92.865 109.685 ;
        RECT 93.315 109.320 93.665 109.685 ;
        RECT 28.595 107.520 28.765 109.280 ;
        RECT 71.705 107.520 71.875 109.280 ;
        RECT 28.595 107.350 71.875 107.520 ;
        RECT 38.565 106.950 39.115 107.350 ;
        RECT 42.865 106.950 43.415 107.350 ;
        RECT 48.915 106.950 49.465 107.350 ;
        RECT 53.165 106.950 53.715 107.350 ;
        RECT 61.015 106.950 61.565 107.350 ;
        RECT 65.415 106.950 65.965 107.350 ;
        RECT 28.595 106.780 71.875 106.950 ;
        RECT 28.595 105.020 28.765 106.780 ;
        RECT 71.705 105.020 71.875 106.780 ;
        RECT 28.595 104.850 71.875 105.020 ;
        RECT 31.395 104.280 68.585 104.450 ;
        RECT 31.395 102.020 31.565 104.280 ;
        RECT 32.245 102.420 37.285 102.590 ;
        RECT 38.335 102.420 43.375 102.590 ;
        RECT 44.425 102.420 49.465 102.590 ;
        RECT 50.515 102.420 55.555 102.590 ;
        RECT 56.605 102.420 61.645 102.590 ;
        RECT 62.695 102.420 67.735 102.590 ;
        RECT 68.415 102.020 68.585 104.280 ;
        RECT 31.395 101.850 68.585 102.020 ;
        RECT 34.865 101.350 35.715 101.850 ;
        RECT 59.415 101.350 60.265 101.850 ;
        RECT 31.395 101.180 68.585 101.350 ;
        RECT 31.395 98.920 31.565 101.180 ;
        RECT 32.245 99.320 37.285 99.490 ;
        RECT 38.335 99.320 43.375 99.490 ;
        RECT 44.425 99.320 49.465 99.490 ;
        RECT 50.515 99.320 55.555 99.490 ;
        RECT 56.605 99.320 61.645 99.490 ;
        RECT 62.695 99.320 67.735 99.490 ;
        RECT 68.415 98.920 68.585 101.180 ;
        RECT 31.395 98.750 68.585 98.920 ;
        RECT 28.595 98.180 71.875 98.350 ;
        RECT 28.595 95.920 28.765 98.180 ;
        RECT 29.445 97.610 34.485 97.780 ;
        RECT 35.535 97.610 40.575 97.780 ;
        RECT 41.625 97.610 46.665 97.780 ;
        RECT 47.715 97.610 52.755 97.780 ;
        RECT 53.805 97.610 58.845 97.780 ;
        RECT 59.895 97.610 64.935 97.780 ;
        RECT 65.985 97.610 71.025 97.780 ;
        RECT 71.705 95.920 71.875 98.180 ;
        RECT 28.595 95.750 71.875 95.920 ;
        RECT 34.715 95.350 35.315 95.750 ;
        RECT 40.815 95.350 41.415 95.750 ;
        RECT 46.865 95.350 47.465 95.750 ;
        RECT 52.965 95.350 53.565 95.750 ;
        RECT 59.115 95.350 59.715 95.750 ;
        RECT 65.165 95.350 65.765 95.750 ;
        RECT 28.595 95.180 71.875 95.350 ;
        RECT 28.595 92.920 28.765 95.180 ;
        RECT 29.445 94.610 34.485 94.780 ;
        RECT 35.535 94.610 40.575 94.780 ;
        RECT 41.625 94.610 46.665 94.780 ;
        RECT 47.715 94.610 52.755 94.780 ;
        RECT 53.805 94.610 58.845 94.780 ;
        RECT 59.895 94.610 64.935 94.780 ;
        RECT 65.985 94.610 71.025 94.780 ;
        RECT 71.705 92.920 71.875 95.180 ;
        RECT 28.595 92.750 71.875 92.920 ;
        RECT 45.170 83.410 55.180 83.580 ;
        RECT 45.170 81.150 45.340 83.410 ;
        RECT 46.020 81.550 47.310 81.720 ;
        RECT 48.360 81.550 49.650 81.720 ;
        RECT 50.700 81.550 51.990 81.720 ;
        RECT 53.040 81.550 54.330 81.720 ;
        RECT 55.010 81.150 55.180 83.410 ;
        RECT 45.170 80.980 55.180 81.150 ;
        RECT 45.990 80.455 47.090 80.980 ;
        RECT 48.590 80.455 49.690 80.980 ;
        RECT 50.690 80.455 51.790 80.980 ;
        RECT 53.440 80.455 54.540 80.980 ;
        RECT 45.990 80.400 54.540 80.455 ;
        RECT 46.270 80.285 54.100 80.400 ;
        RECT 46.270 78.525 46.440 80.285 ;
        RECT 53.930 78.525 54.100 80.285 ;
        RECT 34.190 77.830 35.090 78.350 ;
        RECT 39.890 77.830 40.790 78.350 ;
        RECT 44.790 77.830 45.690 78.400 ;
        RECT 46.270 78.355 54.100 78.525 ;
        RECT 48.640 77.830 49.540 78.355 ;
        RECT 50.840 77.830 51.740 78.355 ;
        RECT 54.440 77.830 55.340 78.350 ;
        RECT 59.790 77.830 60.690 78.400 ;
        RECT 64.790 77.830 65.690 78.400 ;
        RECT 31.595 77.660 68.785 77.830 ;
        RECT 31.595 75.400 31.765 77.660 ;
        RECT 68.615 75.400 68.785 77.660 ;
        RECT 31.595 75.230 68.785 75.400 ;
        RECT 33.990 68.170 34.590 68.930 ;
        RECT 65.840 68.170 66.440 68.930 ;
        RECT 33.990 53.170 34.590 53.930 ;
        RECT 65.840 53.170 66.440 53.930 ;
        RECT 33.990 38.170 34.590 38.930 ;
        RECT 65.840 38.170 66.440 38.930 ;
        RECT 33.990 23.170 34.590 23.930 ;
        RECT 65.840 23.170 66.440 23.930 ;
        RECT 33.990 8.170 34.590 8.930 ;
        RECT 65.840 8.170 66.440 8.930 ;
        RECT 35.975 0.250 41.705 2.410 ;
        RECT 43.575 0.250 49.305 2.410 ;
        RECT 51.125 0.280 56.855 2.440 ;
        RECT 58.675 0.280 64.405 2.440 ;
      LAYER mcon ;
        RECT 6.105 109.590 6.275 109.760 ;
        RECT 6.105 109.230 6.275 109.400 ;
        RECT 7.155 109.590 7.325 109.760 ;
        RECT 92.605 109.460 92.775 109.630 ;
        RECT 7.155 109.230 7.325 109.400 ;
        RECT 93.405 109.460 93.575 109.630 ;
        RECT 38.575 106.880 39.105 107.410 ;
        RECT 42.875 106.880 43.405 107.410 ;
        RECT 48.925 106.880 49.455 107.410 ;
        RECT 53.175 106.880 53.705 107.410 ;
        RECT 61.025 106.880 61.555 107.410 ;
        RECT 65.425 106.880 65.955 107.410 ;
        RECT 32.340 102.420 32.510 102.590 ;
        RECT 32.700 102.420 32.870 102.590 ;
        RECT 33.060 102.420 33.230 102.590 ;
        RECT 33.420 102.420 33.590 102.590 ;
        RECT 33.780 102.420 33.950 102.590 ;
        RECT 34.140 102.420 34.310 102.590 ;
        RECT 34.500 102.420 34.670 102.590 ;
        RECT 34.860 102.420 35.030 102.590 ;
        RECT 35.220 102.420 35.390 102.590 ;
        RECT 35.580 102.420 35.750 102.590 ;
        RECT 35.940 102.420 36.110 102.590 ;
        RECT 36.300 102.420 36.470 102.590 ;
        RECT 36.660 102.420 36.830 102.590 ;
        RECT 37.020 102.420 37.190 102.590 ;
        RECT 38.430 102.420 38.600 102.590 ;
        RECT 38.790 102.420 38.960 102.590 ;
        RECT 39.150 102.420 39.320 102.590 ;
        RECT 39.510 102.420 39.680 102.590 ;
        RECT 39.870 102.420 40.040 102.590 ;
        RECT 40.230 102.420 40.400 102.590 ;
        RECT 40.590 102.420 40.760 102.590 ;
        RECT 40.950 102.420 41.120 102.590 ;
        RECT 41.310 102.420 41.480 102.590 ;
        RECT 41.670 102.420 41.840 102.590 ;
        RECT 42.030 102.420 42.200 102.590 ;
        RECT 42.390 102.420 42.560 102.590 ;
        RECT 42.750 102.420 42.920 102.590 ;
        RECT 43.110 102.420 43.280 102.590 ;
        RECT 44.520 102.420 44.690 102.590 ;
        RECT 44.880 102.420 45.050 102.590 ;
        RECT 45.240 102.420 45.410 102.590 ;
        RECT 45.600 102.420 45.770 102.590 ;
        RECT 45.960 102.420 46.130 102.590 ;
        RECT 46.320 102.420 46.490 102.590 ;
        RECT 46.680 102.420 46.850 102.590 ;
        RECT 47.040 102.420 47.210 102.590 ;
        RECT 47.400 102.420 47.570 102.590 ;
        RECT 47.760 102.420 47.930 102.590 ;
        RECT 48.120 102.420 48.290 102.590 ;
        RECT 48.480 102.420 48.650 102.590 ;
        RECT 48.840 102.420 49.010 102.590 ;
        RECT 49.200 102.420 49.370 102.590 ;
        RECT 50.610 102.420 50.780 102.590 ;
        RECT 50.970 102.420 51.140 102.590 ;
        RECT 51.330 102.420 51.500 102.590 ;
        RECT 51.690 102.420 51.860 102.590 ;
        RECT 52.050 102.420 52.220 102.590 ;
        RECT 52.410 102.420 52.580 102.590 ;
        RECT 52.770 102.420 52.940 102.590 ;
        RECT 53.130 102.420 53.300 102.590 ;
        RECT 53.490 102.420 53.660 102.590 ;
        RECT 53.850 102.420 54.020 102.590 ;
        RECT 54.210 102.420 54.380 102.590 ;
        RECT 54.570 102.420 54.740 102.590 ;
        RECT 54.930 102.420 55.100 102.590 ;
        RECT 55.290 102.420 55.460 102.590 ;
        RECT 56.700 102.420 56.870 102.590 ;
        RECT 57.060 102.420 57.230 102.590 ;
        RECT 57.420 102.420 57.590 102.590 ;
        RECT 57.780 102.420 57.950 102.590 ;
        RECT 58.140 102.420 58.310 102.590 ;
        RECT 58.500 102.420 58.670 102.590 ;
        RECT 58.860 102.420 59.030 102.590 ;
        RECT 59.220 102.420 59.390 102.590 ;
        RECT 59.580 102.420 59.750 102.590 ;
        RECT 59.940 102.420 60.110 102.590 ;
        RECT 60.300 102.420 60.470 102.590 ;
        RECT 60.660 102.420 60.830 102.590 ;
        RECT 61.020 102.420 61.190 102.590 ;
        RECT 61.380 102.420 61.550 102.590 ;
        RECT 62.790 102.420 62.960 102.590 ;
        RECT 63.150 102.420 63.320 102.590 ;
        RECT 63.510 102.420 63.680 102.590 ;
        RECT 63.870 102.420 64.040 102.590 ;
        RECT 64.230 102.420 64.400 102.590 ;
        RECT 64.590 102.420 64.760 102.590 ;
        RECT 64.950 102.420 65.120 102.590 ;
        RECT 65.310 102.420 65.480 102.590 ;
        RECT 65.670 102.420 65.840 102.590 ;
        RECT 66.030 102.420 66.200 102.590 ;
        RECT 66.390 102.420 66.560 102.590 ;
        RECT 66.750 102.420 66.920 102.590 ;
        RECT 67.110 102.420 67.280 102.590 ;
        RECT 67.470 102.420 67.640 102.590 ;
        RECT 35.025 101.510 35.195 101.680 ;
        RECT 35.385 101.510 35.555 101.680 ;
        RECT 59.575 101.510 59.745 101.680 ;
        RECT 59.935 101.510 60.105 101.680 ;
        RECT 32.340 99.320 32.510 99.490 ;
        RECT 32.700 99.320 32.870 99.490 ;
        RECT 33.060 99.320 33.230 99.490 ;
        RECT 33.420 99.320 33.590 99.490 ;
        RECT 33.780 99.320 33.950 99.490 ;
        RECT 34.140 99.320 34.310 99.490 ;
        RECT 34.500 99.320 34.670 99.490 ;
        RECT 34.860 99.320 35.030 99.490 ;
        RECT 35.220 99.320 35.390 99.490 ;
        RECT 35.580 99.320 35.750 99.490 ;
        RECT 35.940 99.320 36.110 99.490 ;
        RECT 36.300 99.320 36.470 99.490 ;
        RECT 36.660 99.320 36.830 99.490 ;
        RECT 37.020 99.320 37.190 99.490 ;
        RECT 38.430 99.320 38.600 99.490 ;
        RECT 38.790 99.320 38.960 99.490 ;
        RECT 39.150 99.320 39.320 99.490 ;
        RECT 39.510 99.320 39.680 99.490 ;
        RECT 39.870 99.320 40.040 99.490 ;
        RECT 40.230 99.320 40.400 99.490 ;
        RECT 40.590 99.320 40.760 99.490 ;
        RECT 40.950 99.320 41.120 99.490 ;
        RECT 41.310 99.320 41.480 99.490 ;
        RECT 41.670 99.320 41.840 99.490 ;
        RECT 42.030 99.320 42.200 99.490 ;
        RECT 42.390 99.320 42.560 99.490 ;
        RECT 42.750 99.320 42.920 99.490 ;
        RECT 43.110 99.320 43.280 99.490 ;
        RECT 44.520 99.320 44.690 99.490 ;
        RECT 44.880 99.320 45.050 99.490 ;
        RECT 45.240 99.320 45.410 99.490 ;
        RECT 45.600 99.320 45.770 99.490 ;
        RECT 45.960 99.320 46.130 99.490 ;
        RECT 46.320 99.320 46.490 99.490 ;
        RECT 46.680 99.320 46.850 99.490 ;
        RECT 47.040 99.320 47.210 99.490 ;
        RECT 47.400 99.320 47.570 99.490 ;
        RECT 47.760 99.320 47.930 99.490 ;
        RECT 48.120 99.320 48.290 99.490 ;
        RECT 48.480 99.320 48.650 99.490 ;
        RECT 48.840 99.320 49.010 99.490 ;
        RECT 49.200 99.320 49.370 99.490 ;
        RECT 50.610 99.320 50.780 99.490 ;
        RECT 50.970 99.320 51.140 99.490 ;
        RECT 51.330 99.320 51.500 99.490 ;
        RECT 51.690 99.320 51.860 99.490 ;
        RECT 52.050 99.320 52.220 99.490 ;
        RECT 52.410 99.320 52.580 99.490 ;
        RECT 52.770 99.320 52.940 99.490 ;
        RECT 53.130 99.320 53.300 99.490 ;
        RECT 53.490 99.320 53.660 99.490 ;
        RECT 53.850 99.320 54.020 99.490 ;
        RECT 54.210 99.320 54.380 99.490 ;
        RECT 54.570 99.320 54.740 99.490 ;
        RECT 54.930 99.320 55.100 99.490 ;
        RECT 55.290 99.320 55.460 99.490 ;
        RECT 56.700 99.320 56.870 99.490 ;
        RECT 57.060 99.320 57.230 99.490 ;
        RECT 57.420 99.320 57.590 99.490 ;
        RECT 57.780 99.320 57.950 99.490 ;
        RECT 58.140 99.320 58.310 99.490 ;
        RECT 58.500 99.320 58.670 99.490 ;
        RECT 58.860 99.320 59.030 99.490 ;
        RECT 59.220 99.320 59.390 99.490 ;
        RECT 59.580 99.320 59.750 99.490 ;
        RECT 59.940 99.320 60.110 99.490 ;
        RECT 60.300 99.320 60.470 99.490 ;
        RECT 60.660 99.320 60.830 99.490 ;
        RECT 61.020 99.320 61.190 99.490 ;
        RECT 61.380 99.320 61.550 99.490 ;
        RECT 62.790 99.320 62.960 99.490 ;
        RECT 63.150 99.320 63.320 99.490 ;
        RECT 63.510 99.320 63.680 99.490 ;
        RECT 63.870 99.320 64.040 99.490 ;
        RECT 64.230 99.320 64.400 99.490 ;
        RECT 64.590 99.320 64.760 99.490 ;
        RECT 64.950 99.320 65.120 99.490 ;
        RECT 65.310 99.320 65.480 99.490 ;
        RECT 65.670 99.320 65.840 99.490 ;
        RECT 66.030 99.320 66.200 99.490 ;
        RECT 66.390 99.320 66.560 99.490 ;
        RECT 66.750 99.320 66.920 99.490 ;
        RECT 67.110 99.320 67.280 99.490 ;
        RECT 67.470 99.320 67.640 99.490 ;
        RECT 29.540 97.610 29.710 97.780 ;
        RECT 29.900 97.610 30.070 97.780 ;
        RECT 30.260 97.610 30.430 97.780 ;
        RECT 30.620 97.610 30.790 97.780 ;
        RECT 30.980 97.610 31.150 97.780 ;
        RECT 31.340 97.610 31.510 97.780 ;
        RECT 31.700 97.610 31.870 97.780 ;
        RECT 32.060 97.610 32.230 97.780 ;
        RECT 32.420 97.610 32.590 97.780 ;
        RECT 32.780 97.610 32.950 97.780 ;
        RECT 33.140 97.610 33.310 97.780 ;
        RECT 33.500 97.610 33.670 97.780 ;
        RECT 33.860 97.610 34.030 97.780 ;
        RECT 34.220 97.610 34.390 97.780 ;
        RECT 35.630 97.610 35.800 97.780 ;
        RECT 35.990 97.610 36.160 97.780 ;
        RECT 36.350 97.610 36.520 97.780 ;
        RECT 36.710 97.610 36.880 97.780 ;
        RECT 37.070 97.610 37.240 97.780 ;
        RECT 37.430 97.610 37.600 97.780 ;
        RECT 37.790 97.610 37.960 97.780 ;
        RECT 38.150 97.610 38.320 97.780 ;
        RECT 38.510 97.610 38.680 97.780 ;
        RECT 38.870 97.610 39.040 97.780 ;
        RECT 39.230 97.610 39.400 97.780 ;
        RECT 39.590 97.610 39.760 97.780 ;
        RECT 39.950 97.610 40.120 97.780 ;
        RECT 40.310 97.610 40.480 97.780 ;
        RECT 41.720 97.610 41.890 97.780 ;
        RECT 42.080 97.610 42.250 97.780 ;
        RECT 42.440 97.610 42.610 97.780 ;
        RECT 42.800 97.610 42.970 97.780 ;
        RECT 43.160 97.610 43.330 97.780 ;
        RECT 43.520 97.610 43.690 97.780 ;
        RECT 43.880 97.610 44.050 97.780 ;
        RECT 44.240 97.610 44.410 97.780 ;
        RECT 44.600 97.610 44.770 97.780 ;
        RECT 44.960 97.610 45.130 97.780 ;
        RECT 45.320 97.610 45.490 97.780 ;
        RECT 45.680 97.610 45.850 97.780 ;
        RECT 46.040 97.610 46.210 97.780 ;
        RECT 46.400 97.610 46.570 97.780 ;
        RECT 47.810 97.610 47.980 97.780 ;
        RECT 48.170 97.610 48.340 97.780 ;
        RECT 48.530 97.610 48.700 97.780 ;
        RECT 48.890 97.610 49.060 97.780 ;
        RECT 49.250 97.610 49.420 97.780 ;
        RECT 49.610 97.610 49.780 97.780 ;
        RECT 49.970 97.610 50.140 97.780 ;
        RECT 50.330 97.610 50.500 97.780 ;
        RECT 50.690 97.610 50.860 97.780 ;
        RECT 51.050 97.610 51.220 97.780 ;
        RECT 51.410 97.610 51.580 97.780 ;
        RECT 51.770 97.610 51.940 97.780 ;
        RECT 52.130 97.610 52.300 97.780 ;
        RECT 52.490 97.610 52.660 97.780 ;
        RECT 53.900 97.610 54.070 97.780 ;
        RECT 54.260 97.610 54.430 97.780 ;
        RECT 54.620 97.610 54.790 97.780 ;
        RECT 54.980 97.610 55.150 97.780 ;
        RECT 55.340 97.610 55.510 97.780 ;
        RECT 55.700 97.610 55.870 97.780 ;
        RECT 56.060 97.610 56.230 97.780 ;
        RECT 56.420 97.610 56.590 97.780 ;
        RECT 56.780 97.610 56.950 97.780 ;
        RECT 57.140 97.610 57.310 97.780 ;
        RECT 57.500 97.610 57.670 97.780 ;
        RECT 57.860 97.610 58.030 97.780 ;
        RECT 58.220 97.610 58.390 97.780 ;
        RECT 58.580 97.610 58.750 97.780 ;
        RECT 59.990 97.610 60.160 97.780 ;
        RECT 60.350 97.610 60.520 97.780 ;
        RECT 60.710 97.610 60.880 97.780 ;
        RECT 61.070 97.610 61.240 97.780 ;
        RECT 61.430 97.610 61.600 97.780 ;
        RECT 61.790 97.610 61.960 97.780 ;
        RECT 62.150 97.610 62.320 97.780 ;
        RECT 62.510 97.610 62.680 97.780 ;
        RECT 62.870 97.610 63.040 97.780 ;
        RECT 63.230 97.610 63.400 97.780 ;
        RECT 63.590 97.610 63.760 97.780 ;
        RECT 63.950 97.610 64.120 97.780 ;
        RECT 64.310 97.610 64.480 97.780 ;
        RECT 64.670 97.610 64.840 97.780 ;
        RECT 66.080 97.610 66.250 97.780 ;
        RECT 66.440 97.610 66.610 97.780 ;
        RECT 66.800 97.610 66.970 97.780 ;
        RECT 67.160 97.610 67.330 97.780 ;
        RECT 67.520 97.610 67.690 97.780 ;
        RECT 67.880 97.610 68.050 97.780 ;
        RECT 68.240 97.610 68.410 97.780 ;
        RECT 68.600 97.610 68.770 97.780 ;
        RECT 68.960 97.610 69.130 97.780 ;
        RECT 69.320 97.610 69.490 97.780 ;
        RECT 69.680 97.610 69.850 97.780 ;
        RECT 70.040 97.610 70.210 97.780 ;
        RECT 70.400 97.610 70.570 97.780 ;
        RECT 70.760 97.610 70.930 97.780 ;
        RECT 34.750 95.485 34.920 95.655 ;
        RECT 35.110 95.485 35.280 95.655 ;
        RECT 40.850 95.485 41.020 95.655 ;
        RECT 41.210 95.485 41.380 95.655 ;
        RECT 46.900 95.485 47.070 95.655 ;
        RECT 47.260 95.485 47.430 95.655 ;
        RECT 53.000 95.485 53.170 95.655 ;
        RECT 53.360 95.485 53.530 95.655 ;
        RECT 59.150 95.435 59.320 95.605 ;
        RECT 59.510 95.435 59.680 95.605 ;
        RECT 65.200 95.485 65.370 95.655 ;
        RECT 65.560 95.485 65.730 95.655 ;
        RECT 29.540 94.610 29.710 94.780 ;
        RECT 29.900 94.610 30.070 94.780 ;
        RECT 30.260 94.610 30.430 94.780 ;
        RECT 30.620 94.610 30.790 94.780 ;
        RECT 30.980 94.610 31.150 94.780 ;
        RECT 31.340 94.610 31.510 94.780 ;
        RECT 31.700 94.610 31.870 94.780 ;
        RECT 32.060 94.610 32.230 94.780 ;
        RECT 32.420 94.610 32.590 94.780 ;
        RECT 32.780 94.610 32.950 94.780 ;
        RECT 33.140 94.610 33.310 94.780 ;
        RECT 33.500 94.610 33.670 94.780 ;
        RECT 33.860 94.610 34.030 94.780 ;
        RECT 34.220 94.610 34.390 94.780 ;
        RECT 35.630 94.610 35.800 94.780 ;
        RECT 35.990 94.610 36.160 94.780 ;
        RECT 36.350 94.610 36.520 94.780 ;
        RECT 36.710 94.610 36.880 94.780 ;
        RECT 37.070 94.610 37.240 94.780 ;
        RECT 37.430 94.610 37.600 94.780 ;
        RECT 37.790 94.610 37.960 94.780 ;
        RECT 38.150 94.610 38.320 94.780 ;
        RECT 38.510 94.610 38.680 94.780 ;
        RECT 38.870 94.610 39.040 94.780 ;
        RECT 39.230 94.610 39.400 94.780 ;
        RECT 39.590 94.610 39.760 94.780 ;
        RECT 39.950 94.610 40.120 94.780 ;
        RECT 40.310 94.610 40.480 94.780 ;
        RECT 41.720 94.610 41.890 94.780 ;
        RECT 42.080 94.610 42.250 94.780 ;
        RECT 42.440 94.610 42.610 94.780 ;
        RECT 42.800 94.610 42.970 94.780 ;
        RECT 43.160 94.610 43.330 94.780 ;
        RECT 43.520 94.610 43.690 94.780 ;
        RECT 43.880 94.610 44.050 94.780 ;
        RECT 44.240 94.610 44.410 94.780 ;
        RECT 44.600 94.610 44.770 94.780 ;
        RECT 44.960 94.610 45.130 94.780 ;
        RECT 45.320 94.610 45.490 94.780 ;
        RECT 45.680 94.610 45.850 94.780 ;
        RECT 46.040 94.610 46.210 94.780 ;
        RECT 46.400 94.610 46.570 94.780 ;
        RECT 47.810 94.610 47.980 94.780 ;
        RECT 48.170 94.610 48.340 94.780 ;
        RECT 48.530 94.610 48.700 94.780 ;
        RECT 48.890 94.610 49.060 94.780 ;
        RECT 49.250 94.610 49.420 94.780 ;
        RECT 49.610 94.610 49.780 94.780 ;
        RECT 49.970 94.610 50.140 94.780 ;
        RECT 50.330 94.610 50.500 94.780 ;
        RECT 50.690 94.610 50.860 94.780 ;
        RECT 51.050 94.610 51.220 94.780 ;
        RECT 51.410 94.610 51.580 94.780 ;
        RECT 51.770 94.610 51.940 94.780 ;
        RECT 52.130 94.610 52.300 94.780 ;
        RECT 52.490 94.610 52.660 94.780 ;
        RECT 53.900 94.610 54.070 94.780 ;
        RECT 54.260 94.610 54.430 94.780 ;
        RECT 54.620 94.610 54.790 94.780 ;
        RECT 54.980 94.610 55.150 94.780 ;
        RECT 55.340 94.610 55.510 94.780 ;
        RECT 55.700 94.610 55.870 94.780 ;
        RECT 56.060 94.610 56.230 94.780 ;
        RECT 56.420 94.610 56.590 94.780 ;
        RECT 56.780 94.610 56.950 94.780 ;
        RECT 57.140 94.610 57.310 94.780 ;
        RECT 57.500 94.610 57.670 94.780 ;
        RECT 57.860 94.610 58.030 94.780 ;
        RECT 58.220 94.610 58.390 94.780 ;
        RECT 58.580 94.610 58.750 94.780 ;
        RECT 59.990 94.610 60.160 94.780 ;
        RECT 60.350 94.610 60.520 94.780 ;
        RECT 60.710 94.610 60.880 94.780 ;
        RECT 61.070 94.610 61.240 94.780 ;
        RECT 61.430 94.610 61.600 94.780 ;
        RECT 61.790 94.610 61.960 94.780 ;
        RECT 62.150 94.610 62.320 94.780 ;
        RECT 62.510 94.610 62.680 94.780 ;
        RECT 62.870 94.610 63.040 94.780 ;
        RECT 63.230 94.610 63.400 94.780 ;
        RECT 63.590 94.610 63.760 94.780 ;
        RECT 63.950 94.610 64.120 94.780 ;
        RECT 64.310 94.610 64.480 94.780 ;
        RECT 64.670 94.610 64.840 94.780 ;
        RECT 66.080 94.610 66.250 94.780 ;
        RECT 66.440 94.610 66.610 94.780 ;
        RECT 66.800 94.610 66.970 94.780 ;
        RECT 67.160 94.610 67.330 94.780 ;
        RECT 67.520 94.610 67.690 94.780 ;
        RECT 67.880 94.610 68.050 94.780 ;
        RECT 68.240 94.610 68.410 94.780 ;
        RECT 68.600 94.610 68.770 94.780 ;
        RECT 68.960 94.610 69.130 94.780 ;
        RECT 69.320 94.610 69.490 94.780 ;
        RECT 69.680 94.610 69.850 94.780 ;
        RECT 70.040 94.610 70.210 94.780 ;
        RECT 70.400 94.610 70.570 94.780 ;
        RECT 70.760 94.610 70.930 94.780 ;
        RECT 46.220 81.550 46.390 81.720 ;
        RECT 46.580 81.550 46.750 81.720 ;
        RECT 46.940 81.550 47.110 81.720 ;
        RECT 48.560 81.550 48.730 81.720 ;
        RECT 48.920 81.550 49.090 81.720 ;
        RECT 49.280 81.550 49.450 81.720 ;
        RECT 50.900 81.550 51.070 81.720 ;
        RECT 51.260 81.550 51.430 81.720 ;
        RECT 51.620 81.550 51.790 81.720 ;
        RECT 53.240 81.550 53.410 81.720 ;
        RECT 53.600 81.550 53.770 81.720 ;
        RECT 53.960 81.550 54.130 81.720 ;
        RECT 46.095 80.510 46.985 81.040 ;
        RECT 48.695 80.510 49.585 81.040 ;
        RECT 50.795 80.510 51.685 81.040 ;
        RECT 53.545 80.510 54.435 81.040 ;
        RECT 34.195 77.760 35.085 78.290 ;
        RECT 39.895 77.760 40.785 78.290 ;
        RECT 44.795 77.810 45.685 78.340 ;
        RECT 48.645 77.810 49.535 78.340 ;
        RECT 50.845 77.810 51.735 78.340 ;
        RECT 54.445 77.760 55.335 78.290 ;
        RECT 59.795 77.810 60.685 78.340 ;
        RECT 64.795 77.810 65.685 78.340 ;
        RECT 34.025 68.285 34.555 68.815 ;
        RECT 65.875 68.285 66.405 68.815 ;
        RECT 34.025 53.285 34.555 53.815 ;
        RECT 65.875 53.285 66.405 53.815 ;
        RECT 34.025 38.285 34.555 38.815 ;
        RECT 65.875 38.285 66.405 38.815 ;
        RECT 34.025 23.285 34.555 23.815 ;
        RECT 65.875 23.285 66.405 23.815 ;
        RECT 34.025 8.285 34.555 8.815 ;
        RECT 65.875 8.285 66.405 8.815 ;
        RECT 36.055 0.345 41.625 2.315 ;
        RECT 43.655 0.345 49.225 2.315 ;
        RECT 51.205 0.375 56.775 2.345 ;
        RECT 58.755 0.375 64.325 2.345 ;
      LAYER met1 ;
        RECT 5.935 109.820 6.445 109.880 ;
        RECT 6.985 109.820 7.495 109.880 ;
        RECT 5.915 109.170 6.465 109.820 ;
        RECT 6.965 109.170 7.515 109.820 ;
        RECT 92.485 109.770 92.895 109.830 ;
        RECT 93.285 109.770 93.695 109.830 ;
        RECT 92.465 109.320 92.915 109.770 ;
        RECT 93.265 109.320 93.715 109.770 ;
        RECT 92.485 109.260 92.895 109.320 ;
        RECT 93.285 109.260 93.695 109.320 ;
        RECT 5.935 109.110 6.445 109.170 ;
        RECT 6.985 109.110 7.495 109.170 ;
        RECT 38.505 106.840 39.175 107.450 ;
        RECT 42.805 106.840 43.475 107.450 ;
        RECT 48.855 106.840 49.525 107.450 ;
        RECT 53.105 106.840 53.775 107.450 ;
        RECT 60.955 106.840 61.625 107.450 ;
        RECT 65.355 106.840 66.025 107.450 ;
        RECT 32.265 102.470 37.265 102.620 ;
        RECT 38.355 102.470 43.355 102.620 ;
        RECT 44.445 102.470 49.445 102.620 ;
        RECT 50.535 102.470 55.535 102.620 ;
        RECT 56.625 102.470 61.625 102.620 ;
        RECT 62.715 102.470 67.715 102.620 ;
        RECT 32.215 102.270 67.815 102.470 ;
        RECT 34.415 102.070 34.915 102.270 ;
        RECT 58.865 102.070 59.365 102.270 ;
        RECT 34.955 101.340 35.625 101.850 ;
        RECT 59.505 101.340 60.175 101.850 ;
        RECT 32.265 99.370 37.265 99.520 ;
        RECT 38.355 99.370 43.355 99.520 ;
        RECT 44.445 99.370 49.445 99.520 ;
        RECT 50.535 99.370 55.535 99.520 ;
        RECT 56.625 99.370 61.625 99.520 ;
        RECT 62.715 99.370 67.715 99.520 ;
        RECT 32.215 99.170 67.815 99.370 ;
        RECT 34.415 98.970 34.915 99.170 ;
        RECT 58.865 98.970 59.365 99.170 ;
        RECT 43.815 97.970 44.365 98.120 ;
        RECT 68.215 97.970 68.765 98.220 ;
        RECT 29.415 97.770 71.015 97.970 ;
        RECT 29.465 97.580 34.465 97.770 ;
        RECT 35.555 97.580 40.555 97.770 ;
        RECT 41.645 97.580 46.645 97.770 ;
        RECT 47.735 97.580 52.735 97.770 ;
        RECT 53.825 97.580 58.825 97.770 ;
        RECT 59.915 97.580 64.915 97.770 ;
        RECT 66.005 97.580 71.005 97.770 ;
        RECT 34.615 94.970 35.415 95.870 ;
        RECT 40.715 94.970 41.515 95.870 ;
        RECT 43.815 94.970 44.365 95.120 ;
        RECT 46.765 94.970 47.565 95.870 ;
        RECT 52.905 95.820 53.625 95.850 ;
        RECT 65.105 95.820 65.825 95.850 ;
        RECT 52.865 94.970 53.665 95.820 ;
        RECT 59.055 95.770 59.775 95.800 ;
        RECT 59.015 94.970 59.815 95.770 ;
        RECT 65.065 94.970 65.865 95.820 ;
        RECT 68.215 94.970 68.765 95.220 ;
        RECT 29.415 94.770 71.015 94.970 ;
        RECT 29.465 94.580 34.465 94.770 ;
        RECT 35.555 94.580 40.555 94.770 ;
        RECT 41.645 94.580 46.645 94.770 ;
        RECT 47.735 94.580 52.735 94.770 ;
        RECT 53.825 94.580 58.825 94.770 ;
        RECT 59.915 94.580 64.915 94.770 ;
        RECT 66.005 94.580 71.005 94.770 ;
        RECT 46.040 81.650 47.290 81.750 ;
        RECT 48.380 81.650 49.630 81.750 ;
        RECT 50.720 81.650 51.970 81.750 ;
        RECT 53.060 81.650 54.310 81.750 ;
        RECT 45.990 81.450 54.340 81.650 ;
        RECT 45.990 81.180 54.540 81.450 ;
        RECT 45.930 81.100 54.600 81.180 ;
        RECT 45.930 80.370 47.150 81.100 ;
        RECT 48.530 80.370 49.750 81.100 ;
        RECT 50.630 80.370 51.850 81.100 ;
        RECT 53.380 80.370 54.600 81.100 ;
        RECT 34.130 77.670 35.150 78.380 ;
        RECT 39.830 77.670 40.850 78.380 ;
        RECT 44.730 77.720 45.750 78.430 ;
        RECT 48.580 77.720 49.600 78.430 ;
        RECT 50.780 77.720 51.800 78.430 ;
        RECT 54.380 77.670 55.400 78.380 ;
        RECT 59.730 77.720 60.750 78.430 ;
        RECT 64.730 77.720 65.750 78.430 ;
        RECT 33.930 68.220 34.650 68.880 ;
        RECT 65.780 68.220 66.500 68.880 ;
        RECT 33.930 53.220 34.650 53.880 ;
        RECT 65.780 53.220 66.500 53.880 ;
        RECT 33.930 38.220 34.650 38.880 ;
        RECT 65.780 38.220 66.500 38.880 ;
        RECT 33.930 23.220 34.650 23.880 ;
        RECT 65.780 23.220 66.500 23.880 ;
        RECT 33.930 8.220 34.650 8.880 ;
        RECT 65.780 8.220 66.500 8.880 ;
        RECT 35.190 0.050 65.190 2.550 ;
      LAYER via ;
        RECT 6.060 109.525 6.320 109.785 ;
        RECT 6.060 109.205 6.320 109.465 ;
        RECT 7.110 109.525 7.370 109.785 ;
        RECT 7.110 109.205 7.370 109.465 ;
        RECT 92.560 109.415 92.820 109.675 ;
        RECT 93.360 109.415 93.620 109.675 ;
        RECT 38.710 107.015 38.970 107.275 ;
        RECT 43.010 107.015 43.270 107.275 ;
        RECT 49.060 107.015 49.320 107.275 ;
        RECT 53.310 107.015 53.570 107.275 ;
        RECT 61.160 107.015 61.420 107.275 ;
        RECT 65.560 107.015 65.820 107.275 ;
        RECT 34.535 102.140 34.795 102.400 ;
        RECT 58.985 102.140 59.245 102.400 ;
        RECT 35.160 101.465 35.420 101.725 ;
        RECT 59.710 101.465 59.970 101.725 ;
        RECT 34.535 99.040 34.795 99.300 ;
        RECT 58.985 99.040 59.245 99.300 ;
        RECT 43.960 97.790 44.220 98.050 ;
        RECT 68.360 97.890 68.620 98.150 ;
        RECT 34.725 95.440 34.985 95.700 ;
        RECT 35.045 95.440 35.305 95.700 ;
        RECT 40.825 95.440 41.085 95.700 ;
        RECT 41.145 95.440 41.405 95.700 ;
        RECT 46.875 95.440 47.135 95.700 ;
        RECT 47.195 95.440 47.455 95.700 ;
        RECT 43.960 94.790 44.220 95.050 ;
        RECT 52.975 95.440 53.235 95.700 ;
        RECT 53.295 95.440 53.555 95.700 ;
        RECT 59.125 95.390 59.385 95.650 ;
        RECT 59.445 95.390 59.705 95.650 ;
        RECT 65.175 95.440 65.435 95.700 ;
        RECT 65.495 95.440 65.755 95.700 ;
        RECT 68.360 94.890 68.620 95.150 ;
        RECT 46.090 80.485 46.990 81.065 ;
        RECT 48.690 80.485 49.590 81.065 ;
        RECT 50.790 80.485 51.690 81.065 ;
        RECT 53.540 80.485 54.440 81.065 ;
        RECT 34.190 77.735 35.090 78.315 ;
        RECT 39.890 77.735 40.790 78.315 ;
        RECT 44.790 77.785 45.690 78.365 ;
        RECT 48.640 77.785 49.540 78.365 ;
        RECT 50.840 77.785 51.740 78.365 ;
        RECT 54.440 77.735 55.340 78.315 ;
        RECT 59.790 77.785 60.690 78.365 ;
        RECT 64.790 77.785 65.690 78.365 ;
        RECT 34.000 68.260 34.580 68.840 ;
        RECT 65.850 68.260 66.430 68.840 ;
        RECT 34.000 53.260 34.580 53.840 ;
        RECT 65.850 53.260 66.430 53.840 ;
        RECT 34.000 38.260 34.580 38.840 ;
        RECT 65.850 38.260 66.430 38.840 ;
        RECT 34.000 23.260 34.580 23.840 ;
        RECT 65.850 23.260 66.430 23.840 ;
        RECT 34.000 8.260 34.580 8.840 ;
        RECT 65.850 8.260 66.430 8.840 ;
        RECT 35.965 0.245 41.665 2.105 ;
        RECT 43.515 0.245 49.215 2.105 ;
        RECT 51.115 0.245 56.815 2.105 ;
        RECT 58.715 0.295 64.415 2.155 ;
      LAYER met2 ;
        RECT 5.965 109.120 6.415 109.870 ;
        RECT 7.015 109.120 7.465 109.870 ;
        RECT 92.515 109.270 92.865 109.820 ;
        RECT 93.315 109.270 93.665 109.820 ;
        RECT 38.565 106.820 39.115 107.470 ;
        RECT 42.865 106.820 43.415 107.470 ;
        RECT 48.915 106.820 49.465 107.470 ;
        RECT 53.165 106.820 53.715 107.470 ;
        RECT 61.015 106.820 61.565 107.470 ;
        RECT 65.415 106.820 65.965 107.470 ;
        RECT 34.465 102.020 34.865 102.620 ;
        RECT 58.915 102.020 59.315 102.620 ;
        RECT 34.465 101.170 35.765 102.020 ;
        RECT 58.915 101.170 60.265 102.020 ;
        RECT 34.465 98.920 34.865 101.170 ;
        RECT 58.915 98.920 59.315 101.170 ;
        RECT 34.715 95.270 35.315 95.870 ;
        RECT 40.815 95.270 41.415 95.870 ;
        RECT 43.865 94.670 44.315 98.270 ;
        RECT 46.865 95.270 47.465 95.870 ;
        RECT 52.965 95.270 53.565 95.870 ;
        RECT 59.115 95.220 59.715 95.820 ;
        RECT 65.165 95.270 65.765 95.870 ;
        RECT 68.265 94.770 68.715 98.370 ;
        RECT 45.990 80.350 47.090 81.200 ;
        RECT 48.590 80.350 49.690 81.200 ;
        RECT 50.690 80.350 51.790 81.200 ;
        RECT 53.440 80.350 54.540 81.200 ;
        RECT 34.190 77.650 35.090 78.400 ;
        RECT 39.890 77.650 40.790 78.400 ;
        RECT 44.790 77.700 45.690 78.450 ;
        RECT 48.640 77.700 49.540 78.450 ;
        RECT 50.840 77.700 51.740 78.450 ;
        RECT 54.440 77.650 55.340 78.400 ;
        RECT 59.790 77.700 60.690 78.450 ;
        RECT 64.790 77.700 65.690 78.450 ;
        RECT 33.990 68.200 34.590 68.900 ;
        RECT 65.840 68.200 66.440 68.900 ;
        RECT 33.990 53.200 34.590 53.900 ;
        RECT 65.840 53.200 66.440 53.900 ;
        RECT 33.990 38.200 34.590 38.900 ;
        RECT 65.840 38.200 66.440 38.900 ;
        RECT 33.990 23.200 34.590 23.900 ;
        RECT 65.840 23.200 66.440 23.900 ;
        RECT 33.990 8.200 34.590 8.900 ;
        RECT 65.840 8.200 66.440 8.900 ;
        RECT 35.890 0.100 41.740 2.250 ;
        RECT 43.440 0.100 49.290 2.250 ;
        RECT 51.040 0.100 56.890 2.250 ;
        RECT 58.640 0.150 64.490 2.300 ;
      LAYER via2 ;
        RECT 6.050 109.355 6.330 109.635 ;
        RECT 7.100 109.355 7.380 109.635 ;
        RECT 92.550 109.405 92.830 109.685 ;
        RECT 93.350 109.405 93.630 109.685 ;
        RECT 38.700 107.005 38.980 107.285 ;
        RECT 43.000 107.005 43.280 107.285 ;
        RECT 49.050 107.005 49.330 107.285 ;
        RECT 53.300 107.005 53.580 107.285 ;
        RECT 61.150 107.005 61.430 107.285 ;
        RECT 65.550 107.005 65.830 107.285 ;
        RECT 35.150 101.455 35.430 101.735 ;
        RECT 59.700 101.455 59.980 101.735 ;
        RECT 34.875 95.430 35.155 95.710 ;
        RECT 40.975 95.430 41.255 95.710 ;
        RECT 47.025 95.430 47.305 95.710 ;
        RECT 53.125 95.430 53.405 95.710 ;
        RECT 65.325 95.430 65.605 95.710 ;
        RECT 46.000 80.435 47.080 81.115 ;
        RECT 48.600 80.435 49.680 81.115 ;
        RECT 50.700 80.435 51.780 81.115 ;
        RECT 53.450 80.435 54.530 81.115 ;
        RECT 34.300 77.885 34.580 78.165 ;
        RECT 34.700 77.885 34.980 78.165 ;
        RECT 40.000 77.885 40.280 78.165 ;
        RECT 40.400 77.885 40.680 78.165 ;
        RECT 44.900 77.935 45.180 78.215 ;
        RECT 45.300 77.935 45.580 78.215 ;
        RECT 48.750 77.935 49.030 78.215 ;
        RECT 49.150 77.935 49.430 78.215 ;
        RECT 50.950 77.935 51.230 78.215 ;
        RECT 51.350 77.935 51.630 78.215 ;
        RECT 54.550 77.885 54.830 78.165 ;
        RECT 54.950 77.885 55.230 78.165 ;
        RECT 59.900 77.935 60.180 78.215 ;
        RECT 60.300 77.935 60.580 78.215 ;
        RECT 64.900 77.935 65.180 78.215 ;
        RECT 65.300 77.935 65.580 78.215 ;
        RECT 34.150 68.410 34.430 68.690 ;
        RECT 66.000 68.410 66.280 68.690 ;
        RECT 34.150 53.410 34.430 53.690 ;
        RECT 66.000 53.410 66.280 53.690 ;
        RECT 34.150 38.410 34.430 38.690 ;
        RECT 66.000 38.410 66.280 38.690 ;
        RECT 34.150 23.410 34.430 23.690 ;
        RECT 66.000 23.410 66.280 23.690 ;
        RECT 34.150 8.410 34.430 8.690 ;
        RECT 66.000 8.410 66.280 8.690 ;
        RECT 36.075 0.235 41.555 2.115 ;
        RECT 43.625 0.235 49.105 2.115 ;
        RECT 51.225 0.235 56.705 2.115 ;
        RECT 58.825 0.285 64.305 2.165 ;
      LAYER met3 ;
        RECT 5.865 108.170 7.615 109.870 ;
        RECT 3.365 108.120 26.715 108.170 ;
        RECT 92.465 108.120 93.765 109.820 ;
        RECT 3.365 107.020 99.415 108.120 ;
        RECT 25.315 106.320 99.415 107.020 ;
        RECT 25.315 102.820 26.715 106.320 ;
        RECT 74.165 106.270 99.415 106.320 ;
        RECT 74.515 102.820 75.615 106.270 ;
        RECT 25.315 100.520 75.615 102.820 ;
        RECT 25.315 96.920 26.715 100.520 ;
        RECT 74.515 96.920 75.615 100.520 ;
        RECT 25.315 95.610 75.615 96.920 ;
        RECT 25.315 94.620 77.680 95.610 ;
        RECT 73.000 81.450 77.680 94.620 ;
        RECT 31.640 81.190 66.740 81.350 ;
        RECT 72.320 81.190 77.680 81.450 ;
        RECT 31.640 80.450 77.680 81.190 ;
        RECT 33.640 78.500 77.680 80.450 ;
        RECT 33.640 77.550 66.740 78.500 ;
        RECT 72.320 78.210 77.680 78.500 ;
        RECT 72.320 78.060 74.270 78.210 ;
        RECT 33.640 2.350 35.240 77.550 ;
        RECT 65.140 2.350 66.740 77.550 ;
        RECT 33.640 -0.050 66.740 2.350 ;
      LAYER via3 ;
        RECT 59.255 95.360 59.575 95.680 ;
      LAYER met4 ;
        RECT 59.110 95.265 59.720 95.775 ;
    END
  END VSS
  PIN Vp
    ANTENNAGATEAREA 17.500000 ;
    PORT
      LAYER li1 ;
        RECT 29.105 108.150 29.275 108.650 ;
        RECT 34.655 108.150 34.825 108.650 ;
        RECT 35.195 108.150 35.365 108.650 ;
        RECT 40.745 108.150 40.915 108.650 ;
        RECT 41.285 108.150 41.455 108.650 ;
        RECT 46.835 108.150 47.005 108.650 ;
        RECT 47.375 108.150 47.545 108.650 ;
        RECT 52.925 108.150 53.095 108.650 ;
        RECT 53.465 108.150 53.635 108.650 ;
        RECT 59.015 108.150 59.185 108.650 ;
        RECT 59.555 108.150 59.725 108.650 ;
        RECT 65.105 108.150 65.275 108.650 ;
        RECT 65.645 108.150 65.815 108.650 ;
        RECT 71.195 108.150 71.365 108.650 ;
      LAYER mcon ;
        RECT 29.105 108.315 29.275 108.485 ;
        RECT 34.655 108.315 34.825 108.485 ;
        RECT 35.195 108.315 35.365 108.485 ;
        RECT 40.745 108.315 40.915 108.485 ;
        RECT 41.285 108.315 41.455 108.485 ;
        RECT 46.835 108.315 47.005 108.485 ;
        RECT 47.375 108.315 47.545 108.485 ;
        RECT 52.925 108.315 53.095 108.485 ;
        RECT 53.465 108.315 53.635 108.485 ;
        RECT 59.015 108.315 59.185 108.485 ;
        RECT 59.555 108.315 59.725 108.485 ;
        RECT 65.105 108.315 65.275 108.485 ;
        RECT 65.645 108.315 65.815 108.485 ;
        RECT 71.195 108.315 71.365 108.485 ;
      LAYER met1 ;
        RECT 29.075 108.520 29.305 108.630 ;
        RECT 34.625 108.520 34.855 108.630 ;
        RECT 35.165 108.520 35.395 108.630 ;
        RECT 40.715 108.570 40.945 108.630 ;
        RECT 41.255 108.570 41.485 108.630 ;
        RECT 40.715 108.520 41.485 108.570 ;
        RECT 46.805 108.570 47.035 108.630 ;
        RECT 47.345 108.570 47.575 108.630 ;
        RECT 46.805 108.520 47.575 108.570 ;
        RECT 52.895 108.570 53.125 108.630 ;
        RECT 53.435 108.570 53.665 108.630 ;
        RECT 52.895 108.520 53.665 108.570 ;
        RECT 58.985 108.570 59.215 108.630 ;
        RECT 59.525 108.570 59.755 108.630 ;
        RECT 65.075 108.570 65.305 108.630 ;
        RECT 65.615 108.570 65.845 108.630 ;
        RECT 58.985 108.520 59.765 108.570 ;
        RECT 65.065 108.520 65.845 108.570 ;
        RECT 71.165 108.520 71.395 108.630 ;
        RECT 29.065 108.320 71.395 108.520 ;
        RECT 29.075 108.170 29.305 108.320 ;
        RECT 34.625 108.170 34.855 108.320 ;
        RECT 35.165 108.170 35.395 108.320 ;
        RECT 40.715 108.220 41.485 108.320 ;
        RECT 40.715 108.170 40.945 108.220 ;
        RECT 41.255 108.170 41.485 108.220 ;
        RECT 46.805 108.220 47.575 108.320 ;
        RECT 46.805 108.170 47.035 108.220 ;
        RECT 47.345 108.170 47.575 108.220 ;
        RECT 52.895 108.220 53.665 108.320 ;
        RECT 52.895 108.170 53.125 108.220 ;
        RECT 53.435 108.170 53.665 108.220 ;
        RECT 58.985 108.220 59.765 108.320 ;
        RECT 65.065 108.220 65.845 108.320 ;
        RECT 58.985 108.170 59.215 108.220 ;
        RECT 59.525 108.170 59.755 108.220 ;
        RECT 65.075 108.170 65.305 108.220 ;
        RECT 65.615 108.170 65.845 108.220 ;
        RECT 71.165 108.170 71.395 108.320 ;
    END
  END Vp
  PIN Vn
    ANTENNAGATEAREA 17.500000 ;
    PORT
      LAYER li1 ;
        RECT 29.105 105.650 29.275 106.150 ;
        RECT 34.655 105.650 34.825 106.150 ;
        RECT 35.195 105.650 35.365 106.150 ;
        RECT 40.745 105.650 40.915 106.150 ;
        RECT 41.285 105.650 41.455 106.150 ;
        RECT 46.835 105.650 47.005 106.150 ;
        RECT 47.375 105.650 47.545 106.150 ;
        RECT 52.925 105.650 53.095 106.150 ;
        RECT 53.465 105.650 53.635 106.150 ;
        RECT 59.015 105.650 59.185 106.150 ;
        RECT 59.555 105.650 59.725 106.150 ;
        RECT 65.105 105.650 65.275 106.150 ;
        RECT 65.645 105.650 65.815 106.150 ;
        RECT 71.195 105.650 71.365 106.150 ;
      LAYER mcon ;
        RECT 29.105 105.815 29.275 105.985 ;
        RECT 34.655 105.815 34.825 105.985 ;
        RECT 35.195 105.815 35.365 105.985 ;
        RECT 40.745 105.815 40.915 105.985 ;
        RECT 41.285 105.815 41.455 105.985 ;
        RECT 46.835 105.815 47.005 105.985 ;
        RECT 47.375 105.815 47.545 105.985 ;
        RECT 52.925 105.815 53.095 105.985 ;
        RECT 53.465 105.815 53.635 105.985 ;
        RECT 59.015 105.815 59.185 105.985 ;
        RECT 59.555 105.815 59.725 105.985 ;
        RECT 65.105 105.815 65.275 105.985 ;
        RECT 65.645 105.815 65.815 105.985 ;
        RECT 71.195 105.815 71.365 105.985 ;
      LAYER met1 ;
        RECT 29.075 106.020 29.305 106.130 ;
        RECT 34.625 106.020 34.855 106.130 ;
        RECT 35.165 106.020 35.395 106.130 ;
        RECT 40.715 106.070 40.945 106.130 ;
        RECT 41.255 106.070 41.485 106.130 ;
        RECT 40.715 106.020 41.485 106.070 ;
        RECT 46.805 106.070 47.035 106.130 ;
        RECT 47.345 106.070 47.575 106.130 ;
        RECT 46.805 106.020 47.575 106.070 ;
        RECT 52.895 106.070 53.125 106.130 ;
        RECT 53.435 106.070 53.665 106.130 ;
        RECT 52.895 106.020 53.665 106.070 ;
        RECT 58.985 106.070 59.215 106.130 ;
        RECT 59.525 106.070 59.755 106.130 ;
        RECT 65.075 106.070 65.305 106.130 ;
        RECT 65.615 106.070 65.845 106.130 ;
        RECT 58.985 106.020 59.765 106.070 ;
        RECT 65.065 106.020 65.845 106.070 ;
        RECT 71.165 106.020 71.395 106.130 ;
        RECT 29.075 105.820 71.415 106.020 ;
        RECT 29.075 105.670 29.305 105.820 ;
        RECT 34.625 105.670 34.855 105.820 ;
        RECT 35.165 105.670 35.395 105.820 ;
        RECT 40.715 105.720 41.485 105.820 ;
        RECT 40.715 105.670 40.945 105.720 ;
        RECT 41.255 105.670 41.485 105.720 ;
        RECT 46.805 105.720 47.575 105.820 ;
        RECT 46.805 105.670 47.035 105.720 ;
        RECT 47.345 105.670 47.575 105.720 ;
        RECT 52.895 105.720 53.665 105.820 ;
        RECT 52.895 105.670 53.125 105.720 ;
        RECT 53.435 105.670 53.665 105.720 ;
        RECT 58.985 105.720 59.765 105.820 ;
        RECT 65.065 105.720 65.845 105.820 ;
        RECT 58.985 105.670 59.215 105.720 ;
        RECT 59.525 105.670 59.755 105.720 ;
        RECT 65.075 105.670 65.305 105.720 ;
        RECT 65.615 105.670 65.845 105.720 ;
        RECT 71.165 105.670 71.395 105.820 ;
    END
  END Vn
  OBS
      LAYER li1 ;
        RECT 28.605 136.750 28.775 137.250 ;
        RECT 34.245 136.750 34.415 137.250 ;
        RECT 34.785 136.750 34.955 137.250 ;
        RECT 40.425 136.750 40.595 137.250 ;
        RECT 40.965 136.750 41.135 137.250 ;
        RECT 46.605 136.750 46.775 137.250 ;
        RECT 47.145 136.750 47.315 137.250 ;
        RECT 52.785 136.750 52.955 137.250 ;
        RECT 53.325 136.750 53.495 137.250 ;
        RECT 58.965 136.750 59.135 137.250 ;
        RECT 59.505 136.750 59.675 137.250 ;
        RECT 65.145 136.750 65.315 137.250 ;
        RECT 65.685 136.750 65.855 137.250 ;
        RECT 71.325 136.750 71.495 137.250 ;
        RECT 28.990 136.520 34.030 136.690 ;
        RECT 35.170 136.520 40.210 136.690 ;
        RECT 41.350 136.520 46.390 136.690 ;
        RECT 47.530 136.520 52.570 136.690 ;
        RECT 53.710 136.520 58.750 136.690 ;
        RECT 59.890 136.520 64.930 136.690 ;
        RECT 66.070 136.520 71.110 136.690 ;
        RECT 28.605 134.050 28.775 134.550 ;
        RECT 34.245 134.050 34.415 134.550 ;
        RECT 34.785 134.050 34.955 134.550 ;
        RECT 40.425 134.050 40.595 134.550 ;
        RECT 40.965 134.050 41.135 134.550 ;
        RECT 46.605 134.050 46.775 134.550 ;
        RECT 47.145 134.050 47.315 134.550 ;
        RECT 52.785 134.050 52.955 134.550 ;
        RECT 53.325 134.050 53.495 134.550 ;
        RECT 58.965 134.050 59.135 134.550 ;
        RECT 59.505 134.050 59.675 134.550 ;
        RECT 65.145 134.050 65.315 134.550 ;
        RECT 65.685 134.050 65.855 134.550 ;
        RECT 71.325 134.050 71.495 134.550 ;
        RECT 28.990 133.820 34.030 133.990 ;
        RECT 35.170 133.820 40.210 133.990 ;
        RECT 41.350 133.820 46.390 133.990 ;
        RECT 47.530 133.820 52.570 133.990 ;
        RECT 53.710 133.820 58.750 133.990 ;
        RECT 59.890 133.820 64.930 133.990 ;
        RECT 66.070 133.820 71.110 133.990 ;
        RECT 28.605 131.350 28.775 131.850 ;
        RECT 34.245 131.350 34.415 131.850 ;
        RECT 34.785 131.350 34.955 131.850 ;
        RECT 40.425 131.350 40.595 131.850 ;
        RECT 40.965 131.350 41.135 131.850 ;
        RECT 46.605 131.350 46.775 131.850 ;
        RECT 47.145 131.350 47.315 131.850 ;
        RECT 52.785 131.350 52.955 131.850 ;
        RECT 53.325 131.350 53.495 131.850 ;
        RECT 58.965 131.350 59.135 131.850 ;
        RECT 59.505 131.350 59.675 131.850 ;
        RECT 65.145 131.350 65.315 131.850 ;
        RECT 65.685 131.350 65.855 131.850 ;
        RECT 71.325 131.350 71.495 131.850 ;
        RECT 28.990 131.120 34.030 131.290 ;
        RECT 35.170 131.120 40.210 131.290 ;
        RECT 41.350 131.120 46.390 131.290 ;
        RECT 47.530 131.120 52.570 131.290 ;
        RECT 53.710 131.120 58.750 131.290 ;
        RECT 59.890 131.120 64.930 131.290 ;
        RECT 66.070 131.120 71.110 131.290 ;
        RECT 28.605 128.650 28.775 129.150 ;
        RECT 34.245 128.650 34.415 129.150 ;
        RECT 34.785 128.650 34.955 129.150 ;
        RECT 40.425 128.650 40.595 129.150 ;
        RECT 40.965 128.650 41.135 129.150 ;
        RECT 46.605 128.650 46.775 129.150 ;
        RECT 47.145 128.650 47.315 129.150 ;
        RECT 52.785 128.650 52.955 129.150 ;
        RECT 53.325 128.650 53.495 129.150 ;
        RECT 58.965 128.650 59.135 129.150 ;
        RECT 59.505 128.650 59.675 129.150 ;
        RECT 65.145 128.650 65.315 129.150 ;
        RECT 65.685 128.650 65.855 129.150 ;
        RECT 71.325 128.650 71.495 129.150 ;
        RECT 28.990 128.420 34.030 128.590 ;
        RECT 35.170 128.420 40.210 128.590 ;
        RECT 41.350 128.420 46.390 128.590 ;
        RECT 47.530 128.420 52.570 128.590 ;
        RECT 53.710 128.420 58.750 128.590 ;
        RECT 59.890 128.420 64.930 128.590 ;
        RECT 66.070 128.420 71.110 128.590 ;
        RECT 28.605 125.750 28.775 126.250 ;
        RECT 34.245 125.750 34.415 126.250 ;
        RECT 34.785 125.750 34.955 126.250 ;
        RECT 40.425 125.750 40.595 126.250 ;
        RECT 40.965 125.750 41.135 126.250 ;
        RECT 46.605 125.750 46.775 126.250 ;
        RECT 47.145 125.750 47.315 126.250 ;
        RECT 52.785 125.750 52.955 126.250 ;
        RECT 53.325 125.750 53.495 126.250 ;
        RECT 58.965 125.750 59.135 126.250 ;
        RECT 59.505 125.750 59.675 126.250 ;
        RECT 65.145 125.750 65.315 126.250 ;
        RECT 65.685 125.750 65.855 126.250 ;
        RECT 71.325 125.750 71.495 126.250 ;
        RECT 28.990 125.520 34.030 125.690 ;
        RECT 35.170 125.520 40.210 125.690 ;
        RECT 41.350 125.520 46.390 125.690 ;
        RECT 47.530 125.520 52.570 125.690 ;
        RECT 53.710 125.520 58.750 125.690 ;
        RECT 59.890 125.520 64.930 125.690 ;
        RECT 66.070 125.520 71.110 125.690 ;
        RECT 0.780 117.685 2.940 123.415 ;
        RECT 12.940 117.685 15.100 123.415 ;
        RECT 28.605 122.850 28.775 123.350 ;
        RECT 34.245 122.850 34.415 123.350 ;
        RECT 34.785 122.850 34.955 123.350 ;
        RECT 40.425 122.850 40.595 123.350 ;
        RECT 40.965 122.850 41.135 123.350 ;
        RECT 46.605 122.850 46.775 123.350 ;
        RECT 47.145 122.850 47.315 123.350 ;
        RECT 52.785 122.850 52.955 123.350 ;
        RECT 53.325 122.850 53.495 123.350 ;
        RECT 58.965 122.850 59.135 123.350 ;
        RECT 59.505 122.850 59.675 123.350 ;
        RECT 65.145 122.850 65.315 123.350 ;
        RECT 65.685 122.850 65.855 123.350 ;
        RECT 71.325 122.850 71.495 123.350 ;
        RECT 28.990 122.620 34.030 122.790 ;
        RECT 35.170 122.620 40.210 122.790 ;
        RECT 41.350 122.620 46.390 122.790 ;
        RECT 47.530 122.620 52.570 122.790 ;
        RECT 53.710 122.620 58.750 122.790 ;
        RECT 59.890 122.620 64.930 122.790 ;
        RECT 66.070 122.620 71.110 122.790 ;
        RECT 19.405 120.150 19.575 120.650 ;
        RECT 25.045 120.150 25.215 120.650 ;
        RECT 25.585 120.150 25.755 120.650 ;
        RECT 31.225 120.150 31.395 120.650 ;
        RECT 31.765 120.150 31.935 120.650 ;
        RECT 37.405 120.150 37.575 120.650 ;
        RECT 37.945 120.150 38.115 120.650 ;
        RECT 43.585 120.150 43.755 120.650 ;
        RECT 44.125 120.150 44.295 120.650 ;
        RECT 49.765 120.150 49.935 120.650 ;
        RECT 50.305 120.150 50.475 120.650 ;
        RECT 55.945 120.150 56.115 120.650 ;
        RECT 56.485 120.150 56.655 120.650 ;
        RECT 62.125 120.150 62.295 120.650 ;
        RECT 62.665 120.150 62.835 120.650 ;
        RECT 68.305 120.150 68.475 120.650 ;
        RECT 68.845 120.150 69.015 120.650 ;
        RECT 74.485 120.150 74.655 120.650 ;
        RECT 75.025 120.150 75.195 120.650 ;
        RECT 80.665 120.150 80.835 120.650 ;
        RECT 19.405 117.450 19.575 117.950 ;
        RECT 25.045 117.450 25.215 117.950 ;
        RECT 25.585 117.450 25.755 117.950 ;
        RECT 31.225 117.450 31.395 117.950 ;
        RECT 31.765 117.450 31.935 117.950 ;
        RECT 37.405 117.450 37.575 117.950 ;
        RECT 37.945 117.450 38.115 117.950 ;
        RECT 43.585 117.450 43.755 117.950 ;
        RECT 44.125 117.450 44.295 117.950 ;
        RECT 49.765 117.450 49.935 117.950 ;
        RECT 50.305 117.450 50.475 117.950 ;
        RECT 55.945 117.450 56.115 117.950 ;
        RECT 56.485 117.450 56.655 117.950 ;
        RECT 62.125 117.450 62.295 117.950 ;
        RECT 62.665 117.450 62.835 117.950 ;
        RECT 68.305 117.450 68.475 117.950 ;
        RECT 68.845 117.450 69.015 117.950 ;
        RECT 74.485 117.450 74.655 117.950 ;
        RECT 75.025 117.450 75.195 117.950 ;
        RECT 80.665 117.450 80.835 117.950 ;
        RECT 86.080 117.685 88.240 123.415 ;
        RECT 98.240 117.685 100.400 123.415 ;
        RECT 0.780 110.335 2.940 116.065 ;
        RECT 12.940 110.335 15.100 116.065 ;
        RECT 19.405 114.750 19.575 115.250 ;
        RECT 25.045 114.750 25.215 115.250 ;
        RECT 25.585 114.750 25.755 115.250 ;
        RECT 31.225 114.750 31.395 115.250 ;
        RECT 31.765 114.750 31.935 115.250 ;
        RECT 37.405 114.750 37.575 115.250 ;
        RECT 37.945 114.750 38.115 115.250 ;
        RECT 43.585 114.750 43.755 115.250 ;
        RECT 44.125 114.750 44.295 115.250 ;
        RECT 49.765 114.750 49.935 115.250 ;
        RECT 50.305 114.750 50.475 115.250 ;
        RECT 55.945 114.750 56.115 115.250 ;
        RECT 56.485 114.750 56.655 115.250 ;
        RECT 62.125 114.750 62.295 115.250 ;
        RECT 62.665 114.750 62.835 115.250 ;
        RECT 68.305 114.750 68.475 115.250 ;
        RECT 68.845 114.750 69.015 115.250 ;
        RECT 74.485 114.750 74.655 115.250 ;
        RECT 75.025 114.750 75.195 115.250 ;
        RECT 80.665 114.750 80.835 115.250 ;
        RECT 19.405 112.050 19.575 112.550 ;
        RECT 25.045 112.050 25.215 112.550 ;
        RECT 25.585 112.050 25.755 112.550 ;
        RECT 31.225 112.050 31.395 112.550 ;
        RECT 31.765 112.050 31.935 112.550 ;
        RECT 37.405 112.050 37.575 112.550 ;
        RECT 37.945 112.050 38.115 112.550 ;
        RECT 43.585 112.050 43.755 112.550 ;
        RECT 44.125 112.050 44.295 112.550 ;
        RECT 49.765 112.050 49.935 112.550 ;
        RECT 50.305 112.050 50.475 112.550 ;
        RECT 55.945 112.050 56.115 112.550 ;
        RECT 56.485 112.050 56.655 112.550 ;
        RECT 62.125 112.050 62.295 112.550 ;
        RECT 62.665 112.050 62.835 112.550 ;
        RECT 68.305 112.050 68.475 112.550 ;
        RECT 68.845 112.050 69.015 112.550 ;
        RECT 74.485 112.050 74.655 112.550 ;
        RECT 75.025 112.050 75.195 112.550 ;
        RECT 80.665 112.050 80.835 112.550 ;
        RECT 86.080 110.335 88.240 116.065 ;
        RECT 98.240 110.335 100.400 116.065 ;
        RECT 29.445 108.710 34.485 108.880 ;
        RECT 35.535 108.710 40.575 108.880 ;
        RECT 41.625 108.710 46.665 108.880 ;
        RECT 47.715 108.710 52.755 108.880 ;
        RECT 53.805 108.710 58.845 108.880 ;
        RECT 59.895 108.710 64.935 108.880 ;
        RECT 65.985 108.710 71.025 108.880 ;
        RECT 29.445 107.920 34.485 108.090 ;
        RECT 35.535 107.920 40.575 108.090 ;
        RECT 41.625 107.920 46.665 108.090 ;
        RECT 47.715 107.920 52.755 108.090 ;
        RECT 53.805 107.920 58.845 108.090 ;
        RECT 59.895 107.920 64.935 108.090 ;
        RECT 65.985 107.920 71.025 108.090 ;
        RECT 29.445 106.210 34.485 106.380 ;
        RECT 35.535 106.210 40.575 106.380 ;
        RECT 41.625 106.210 46.665 106.380 ;
        RECT 47.715 106.210 52.755 106.380 ;
        RECT 53.805 106.210 58.845 106.380 ;
        RECT 59.895 106.210 64.935 106.380 ;
        RECT 65.985 106.210 71.025 106.380 ;
        RECT 29.445 105.420 34.485 105.590 ;
        RECT 35.535 105.420 40.575 105.590 ;
        RECT 41.625 105.420 46.665 105.590 ;
        RECT 47.715 105.420 52.755 105.590 ;
        RECT 53.805 105.420 58.845 105.590 ;
        RECT 59.895 105.420 64.935 105.590 ;
        RECT 65.985 105.420 71.025 105.590 ;
        RECT 31.905 102.650 32.075 103.650 ;
        RECT 37.455 102.650 37.625 103.650 ;
        RECT 37.995 102.650 38.165 103.650 ;
        RECT 43.545 102.650 43.715 103.650 ;
        RECT 44.085 102.650 44.255 103.650 ;
        RECT 49.635 102.650 49.805 103.650 ;
        RECT 50.175 102.650 50.345 103.650 ;
        RECT 55.725 102.650 55.895 103.650 ;
        RECT 56.265 102.650 56.435 103.650 ;
        RECT 61.815 102.650 61.985 103.650 ;
        RECT 62.355 102.650 62.525 103.650 ;
        RECT 67.905 102.650 68.075 103.650 ;
        RECT 31.905 99.550 32.075 100.550 ;
        RECT 37.455 99.550 37.625 100.550 ;
        RECT 37.995 99.550 38.165 100.550 ;
        RECT 43.545 99.550 43.715 100.550 ;
        RECT 44.085 99.550 44.255 100.550 ;
        RECT 49.635 99.550 49.805 100.550 ;
        RECT 50.175 99.550 50.345 100.550 ;
        RECT 55.725 99.550 55.895 100.550 ;
        RECT 56.265 99.550 56.435 100.550 ;
        RECT 61.815 99.550 61.985 100.550 ;
        RECT 62.355 99.550 62.525 100.550 ;
        RECT 67.905 99.550 68.075 100.550 ;
        RECT 29.105 96.550 29.275 97.550 ;
        RECT 34.655 96.550 34.825 97.550 ;
        RECT 35.195 96.550 35.365 97.550 ;
        RECT 40.745 96.550 40.915 97.550 ;
        RECT 41.285 96.550 41.455 97.550 ;
        RECT 46.835 96.550 47.005 97.550 ;
        RECT 47.375 96.550 47.545 97.550 ;
        RECT 52.925 96.550 53.095 97.550 ;
        RECT 53.465 96.550 53.635 97.550 ;
        RECT 59.015 96.550 59.185 97.550 ;
        RECT 59.555 96.550 59.725 97.550 ;
        RECT 65.105 96.550 65.275 97.550 ;
        RECT 65.645 96.550 65.815 97.550 ;
        RECT 71.195 96.550 71.365 97.550 ;
        RECT 29.445 96.320 34.485 96.490 ;
        RECT 35.535 96.320 40.575 96.490 ;
        RECT 41.625 96.320 46.665 96.490 ;
        RECT 47.715 96.320 52.755 96.490 ;
        RECT 53.805 96.320 58.845 96.490 ;
        RECT 59.895 96.320 64.935 96.490 ;
        RECT 65.985 96.320 71.025 96.490 ;
        RECT 29.105 93.550 29.275 94.550 ;
        RECT 34.655 93.550 34.825 94.550 ;
        RECT 35.195 93.550 35.365 94.550 ;
        RECT 40.745 93.550 40.915 94.550 ;
        RECT 41.285 93.550 41.455 94.550 ;
        RECT 46.835 93.550 47.005 94.550 ;
        RECT 47.375 93.550 47.545 94.550 ;
        RECT 52.925 93.550 53.095 94.550 ;
        RECT 53.465 93.550 53.635 94.550 ;
        RECT 59.015 93.550 59.185 94.550 ;
        RECT 59.555 93.550 59.725 94.550 ;
        RECT 65.105 93.550 65.275 94.550 ;
        RECT 65.645 93.550 65.815 94.550 ;
        RECT 71.195 93.550 71.365 94.550 ;
        RECT 29.445 93.320 34.485 93.490 ;
        RECT 35.535 93.320 40.575 93.490 ;
        RECT 41.625 93.320 46.665 93.490 ;
        RECT 47.715 93.320 52.755 93.490 ;
        RECT 53.805 93.320 58.845 93.490 ;
        RECT 59.895 93.320 64.935 93.490 ;
        RECT 65.985 93.320 71.025 93.490 ;
        RECT 31.830 88.680 32.000 89.680 ;
        RECT 37.470 88.680 37.640 89.680 ;
        RECT 38.010 88.680 38.180 89.680 ;
        RECT 43.650 88.680 43.820 89.680 ;
        RECT 44.190 88.680 44.360 89.680 ;
        RECT 49.830 88.680 50.000 89.680 ;
        RECT 50.370 88.680 50.540 89.680 ;
        RECT 56.010 88.680 56.180 89.680 ;
        RECT 56.550 88.680 56.720 89.680 ;
        RECT 62.190 88.680 62.360 89.680 ;
        RECT 62.730 88.680 62.900 89.680 ;
        RECT 68.370 88.680 68.540 89.680 ;
        RECT 32.215 88.450 37.255 88.620 ;
        RECT 38.395 88.450 43.435 88.620 ;
        RECT 44.575 88.450 49.615 88.620 ;
        RECT 50.755 88.450 55.795 88.620 ;
        RECT 56.935 88.450 61.975 88.620 ;
        RECT 63.115 88.450 68.155 88.620 ;
        RECT 31.830 85.730 32.000 86.730 ;
        RECT 37.470 85.730 37.640 86.730 ;
        RECT 38.010 85.730 38.180 86.730 ;
        RECT 43.650 85.730 43.820 86.730 ;
        RECT 44.190 85.730 44.360 86.730 ;
        RECT 49.830 85.730 50.000 86.730 ;
        RECT 50.370 85.730 50.540 86.730 ;
        RECT 56.010 85.730 56.180 86.730 ;
        RECT 56.550 85.730 56.720 86.730 ;
        RECT 62.190 85.730 62.360 86.730 ;
        RECT 62.730 85.730 62.900 86.730 ;
        RECT 68.370 85.730 68.540 86.730 ;
        RECT 32.215 85.500 37.255 85.670 ;
        RECT 38.395 85.500 43.435 85.670 ;
        RECT 44.575 85.500 49.615 85.670 ;
        RECT 50.755 85.500 55.795 85.670 ;
        RECT 56.935 85.500 61.975 85.670 ;
        RECT 63.115 85.500 68.155 85.670 ;
        RECT 46.020 82.840 47.310 83.010 ;
        RECT 48.360 82.840 49.650 83.010 ;
        RECT 50.700 82.840 51.990 83.010 ;
        RECT 53.040 82.840 54.330 83.010 ;
        RECT 45.680 81.780 45.850 82.780 ;
        RECT 47.480 81.780 47.650 82.780 ;
        RECT 48.020 81.780 48.190 82.780 ;
        RECT 49.820 81.780 49.990 82.780 ;
        RECT 50.360 81.780 50.530 82.780 ;
        RECT 52.160 81.780 52.330 82.780 ;
        RECT 52.700 81.780 52.870 82.780 ;
        RECT 54.500 81.780 54.670 82.780 ;
        RECT 47.120 79.715 49.660 79.885 ;
        RECT 50.710 79.715 53.250 79.885 ;
        RECT 46.780 79.155 46.950 79.655 ;
        RECT 49.830 79.155 50.000 79.655 ;
        RECT 50.370 79.155 50.540 79.655 ;
        RECT 53.420 79.155 53.590 79.655 ;
        RECT 47.120 78.925 49.660 79.095 ;
        RECT 50.710 78.925 53.250 79.095 ;
        RECT 32.445 77.090 37.485 77.260 ;
        RECT 38.535 77.090 43.575 77.260 ;
        RECT 44.625 77.090 49.665 77.260 ;
        RECT 50.715 77.090 55.755 77.260 ;
        RECT 56.805 77.090 61.845 77.260 ;
        RECT 62.895 77.090 67.935 77.260 ;
        RECT 32.105 76.030 32.275 77.030 ;
        RECT 37.655 76.030 37.825 77.030 ;
        RECT 38.195 76.030 38.365 77.030 ;
        RECT 43.745 76.030 43.915 77.030 ;
        RECT 44.285 76.030 44.455 77.030 ;
        RECT 49.835 76.030 50.005 77.030 ;
        RECT 50.375 76.030 50.545 77.030 ;
        RECT 55.925 76.030 56.095 77.030 ;
        RECT 56.465 76.030 56.635 77.030 ;
        RECT 62.015 76.030 62.185 77.030 ;
        RECT 62.555 76.030 62.725 77.030 ;
        RECT 68.105 76.030 68.275 77.030 ;
        RECT 32.445 75.800 37.485 75.970 ;
        RECT 38.535 75.800 43.575 75.970 ;
        RECT 44.625 75.800 49.665 75.970 ;
        RECT 50.715 75.800 55.755 75.970 ;
        RECT 56.805 75.800 61.845 75.970 ;
        RECT 62.895 75.800 67.935 75.970 ;
        RECT 35.975 71.410 41.705 73.570 ;
        RECT 43.575 71.410 49.305 73.570 ;
        RECT 51.125 71.440 56.855 73.600 ;
        RECT 58.675 71.440 64.405 73.600 ;
      LAYER mcon ;
        RECT 28.605 136.915 28.775 137.085 ;
        RECT 34.245 136.915 34.415 137.085 ;
        RECT 34.785 136.915 34.955 137.085 ;
        RECT 40.425 136.915 40.595 137.085 ;
        RECT 40.965 136.915 41.135 137.085 ;
        RECT 46.605 136.915 46.775 137.085 ;
        RECT 47.145 136.915 47.315 137.085 ;
        RECT 52.785 136.915 52.955 137.085 ;
        RECT 53.325 136.915 53.495 137.085 ;
        RECT 58.965 136.915 59.135 137.085 ;
        RECT 59.505 136.915 59.675 137.085 ;
        RECT 65.145 136.915 65.315 137.085 ;
        RECT 65.685 136.915 65.855 137.085 ;
        RECT 71.325 136.915 71.495 137.085 ;
        RECT 29.085 136.520 29.255 136.690 ;
        RECT 29.445 136.520 29.615 136.690 ;
        RECT 29.805 136.520 29.975 136.690 ;
        RECT 30.165 136.520 30.335 136.690 ;
        RECT 30.525 136.520 30.695 136.690 ;
        RECT 30.885 136.520 31.055 136.690 ;
        RECT 31.245 136.520 31.415 136.690 ;
        RECT 31.605 136.520 31.775 136.690 ;
        RECT 31.965 136.520 32.135 136.690 ;
        RECT 32.325 136.520 32.495 136.690 ;
        RECT 32.685 136.520 32.855 136.690 ;
        RECT 33.045 136.520 33.215 136.690 ;
        RECT 33.405 136.520 33.575 136.690 ;
        RECT 33.765 136.520 33.935 136.690 ;
        RECT 35.265 136.520 35.435 136.690 ;
        RECT 35.625 136.520 35.795 136.690 ;
        RECT 35.985 136.520 36.155 136.690 ;
        RECT 36.345 136.520 36.515 136.690 ;
        RECT 36.705 136.520 36.875 136.690 ;
        RECT 37.065 136.520 37.235 136.690 ;
        RECT 37.425 136.520 37.595 136.690 ;
        RECT 37.785 136.520 37.955 136.690 ;
        RECT 38.145 136.520 38.315 136.690 ;
        RECT 38.505 136.520 38.675 136.690 ;
        RECT 38.865 136.520 39.035 136.690 ;
        RECT 39.225 136.520 39.395 136.690 ;
        RECT 39.585 136.520 39.755 136.690 ;
        RECT 39.945 136.520 40.115 136.690 ;
        RECT 41.445 136.520 41.615 136.690 ;
        RECT 41.805 136.520 41.975 136.690 ;
        RECT 42.165 136.520 42.335 136.690 ;
        RECT 42.525 136.520 42.695 136.690 ;
        RECT 42.885 136.520 43.055 136.690 ;
        RECT 43.245 136.520 43.415 136.690 ;
        RECT 43.605 136.520 43.775 136.690 ;
        RECT 43.965 136.520 44.135 136.690 ;
        RECT 44.325 136.520 44.495 136.690 ;
        RECT 44.685 136.520 44.855 136.690 ;
        RECT 45.045 136.520 45.215 136.690 ;
        RECT 45.405 136.520 45.575 136.690 ;
        RECT 45.765 136.520 45.935 136.690 ;
        RECT 46.125 136.520 46.295 136.690 ;
        RECT 47.625 136.520 47.795 136.690 ;
        RECT 47.985 136.520 48.155 136.690 ;
        RECT 48.345 136.520 48.515 136.690 ;
        RECT 48.705 136.520 48.875 136.690 ;
        RECT 49.065 136.520 49.235 136.690 ;
        RECT 49.425 136.520 49.595 136.690 ;
        RECT 49.785 136.520 49.955 136.690 ;
        RECT 50.145 136.520 50.315 136.690 ;
        RECT 50.505 136.520 50.675 136.690 ;
        RECT 50.865 136.520 51.035 136.690 ;
        RECT 51.225 136.520 51.395 136.690 ;
        RECT 51.585 136.520 51.755 136.690 ;
        RECT 51.945 136.520 52.115 136.690 ;
        RECT 52.305 136.520 52.475 136.690 ;
        RECT 53.805 136.520 53.975 136.690 ;
        RECT 54.165 136.520 54.335 136.690 ;
        RECT 54.525 136.520 54.695 136.690 ;
        RECT 54.885 136.520 55.055 136.690 ;
        RECT 55.245 136.520 55.415 136.690 ;
        RECT 55.605 136.520 55.775 136.690 ;
        RECT 55.965 136.520 56.135 136.690 ;
        RECT 56.325 136.520 56.495 136.690 ;
        RECT 56.685 136.520 56.855 136.690 ;
        RECT 57.045 136.520 57.215 136.690 ;
        RECT 57.405 136.520 57.575 136.690 ;
        RECT 57.765 136.520 57.935 136.690 ;
        RECT 58.125 136.520 58.295 136.690 ;
        RECT 58.485 136.520 58.655 136.690 ;
        RECT 59.985 136.520 60.155 136.690 ;
        RECT 60.345 136.520 60.515 136.690 ;
        RECT 60.705 136.520 60.875 136.690 ;
        RECT 61.065 136.520 61.235 136.690 ;
        RECT 61.425 136.520 61.595 136.690 ;
        RECT 61.785 136.520 61.955 136.690 ;
        RECT 62.145 136.520 62.315 136.690 ;
        RECT 62.505 136.520 62.675 136.690 ;
        RECT 62.865 136.520 63.035 136.690 ;
        RECT 63.225 136.520 63.395 136.690 ;
        RECT 63.585 136.520 63.755 136.690 ;
        RECT 63.945 136.520 64.115 136.690 ;
        RECT 64.305 136.520 64.475 136.690 ;
        RECT 64.665 136.520 64.835 136.690 ;
        RECT 66.165 136.520 66.335 136.690 ;
        RECT 66.525 136.520 66.695 136.690 ;
        RECT 66.885 136.520 67.055 136.690 ;
        RECT 67.245 136.520 67.415 136.690 ;
        RECT 67.605 136.520 67.775 136.690 ;
        RECT 67.965 136.520 68.135 136.690 ;
        RECT 68.325 136.520 68.495 136.690 ;
        RECT 68.685 136.520 68.855 136.690 ;
        RECT 69.045 136.520 69.215 136.690 ;
        RECT 69.405 136.520 69.575 136.690 ;
        RECT 69.765 136.520 69.935 136.690 ;
        RECT 70.125 136.520 70.295 136.690 ;
        RECT 70.485 136.520 70.655 136.690 ;
        RECT 70.845 136.520 71.015 136.690 ;
        RECT 28.605 134.215 28.775 134.385 ;
        RECT 34.245 134.215 34.415 134.385 ;
        RECT 34.785 134.215 34.955 134.385 ;
        RECT 40.425 134.215 40.595 134.385 ;
        RECT 40.965 134.215 41.135 134.385 ;
        RECT 46.605 134.215 46.775 134.385 ;
        RECT 47.145 134.215 47.315 134.385 ;
        RECT 52.785 134.215 52.955 134.385 ;
        RECT 53.325 134.215 53.495 134.385 ;
        RECT 58.965 134.215 59.135 134.385 ;
        RECT 59.505 134.215 59.675 134.385 ;
        RECT 65.145 134.215 65.315 134.385 ;
        RECT 65.685 134.215 65.855 134.385 ;
        RECT 71.325 134.215 71.495 134.385 ;
        RECT 29.085 133.820 29.255 133.990 ;
        RECT 29.445 133.820 29.615 133.990 ;
        RECT 29.805 133.820 29.975 133.990 ;
        RECT 30.165 133.820 30.335 133.990 ;
        RECT 30.525 133.820 30.695 133.990 ;
        RECT 30.885 133.820 31.055 133.990 ;
        RECT 31.245 133.820 31.415 133.990 ;
        RECT 31.605 133.820 31.775 133.990 ;
        RECT 31.965 133.820 32.135 133.990 ;
        RECT 32.325 133.820 32.495 133.990 ;
        RECT 32.685 133.820 32.855 133.990 ;
        RECT 33.045 133.820 33.215 133.990 ;
        RECT 33.405 133.820 33.575 133.990 ;
        RECT 33.765 133.820 33.935 133.990 ;
        RECT 35.265 133.820 35.435 133.990 ;
        RECT 35.625 133.820 35.795 133.990 ;
        RECT 35.985 133.820 36.155 133.990 ;
        RECT 36.345 133.820 36.515 133.990 ;
        RECT 36.705 133.820 36.875 133.990 ;
        RECT 37.065 133.820 37.235 133.990 ;
        RECT 37.425 133.820 37.595 133.990 ;
        RECT 37.785 133.820 37.955 133.990 ;
        RECT 38.145 133.820 38.315 133.990 ;
        RECT 38.505 133.820 38.675 133.990 ;
        RECT 38.865 133.820 39.035 133.990 ;
        RECT 39.225 133.820 39.395 133.990 ;
        RECT 39.585 133.820 39.755 133.990 ;
        RECT 39.945 133.820 40.115 133.990 ;
        RECT 41.445 133.820 41.615 133.990 ;
        RECT 41.805 133.820 41.975 133.990 ;
        RECT 42.165 133.820 42.335 133.990 ;
        RECT 42.525 133.820 42.695 133.990 ;
        RECT 42.885 133.820 43.055 133.990 ;
        RECT 43.245 133.820 43.415 133.990 ;
        RECT 43.605 133.820 43.775 133.990 ;
        RECT 43.965 133.820 44.135 133.990 ;
        RECT 44.325 133.820 44.495 133.990 ;
        RECT 44.685 133.820 44.855 133.990 ;
        RECT 45.045 133.820 45.215 133.990 ;
        RECT 45.405 133.820 45.575 133.990 ;
        RECT 45.765 133.820 45.935 133.990 ;
        RECT 46.125 133.820 46.295 133.990 ;
        RECT 47.625 133.820 47.795 133.990 ;
        RECT 47.985 133.820 48.155 133.990 ;
        RECT 48.345 133.820 48.515 133.990 ;
        RECT 48.705 133.820 48.875 133.990 ;
        RECT 49.065 133.820 49.235 133.990 ;
        RECT 49.425 133.820 49.595 133.990 ;
        RECT 49.785 133.820 49.955 133.990 ;
        RECT 50.145 133.820 50.315 133.990 ;
        RECT 50.505 133.820 50.675 133.990 ;
        RECT 50.865 133.820 51.035 133.990 ;
        RECT 51.225 133.820 51.395 133.990 ;
        RECT 51.585 133.820 51.755 133.990 ;
        RECT 51.945 133.820 52.115 133.990 ;
        RECT 52.305 133.820 52.475 133.990 ;
        RECT 53.805 133.820 53.975 133.990 ;
        RECT 54.165 133.820 54.335 133.990 ;
        RECT 54.525 133.820 54.695 133.990 ;
        RECT 54.885 133.820 55.055 133.990 ;
        RECT 55.245 133.820 55.415 133.990 ;
        RECT 55.605 133.820 55.775 133.990 ;
        RECT 55.965 133.820 56.135 133.990 ;
        RECT 56.325 133.820 56.495 133.990 ;
        RECT 56.685 133.820 56.855 133.990 ;
        RECT 57.045 133.820 57.215 133.990 ;
        RECT 57.405 133.820 57.575 133.990 ;
        RECT 57.765 133.820 57.935 133.990 ;
        RECT 58.125 133.820 58.295 133.990 ;
        RECT 58.485 133.820 58.655 133.990 ;
        RECT 59.985 133.820 60.155 133.990 ;
        RECT 60.345 133.820 60.515 133.990 ;
        RECT 60.705 133.820 60.875 133.990 ;
        RECT 61.065 133.820 61.235 133.990 ;
        RECT 61.425 133.820 61.595 133.990 ;
        RECT 61.785 133.820 61.955 133.990 ;
        RECT 62.145 133.820 62.315 133.990 ;
        RECT 62.505 133.820 62.675 133.990 ;
        RECT 62.865 133.820 63.035 133.990 ;
        RECT 63.225 133.820 63.395 133.990 ;
        RECT 63.585 133.820 63.755 133.990 ;
        RECT 63.945 133.820 64.115 133.990 ;
        RECT 64.305 133.820 64.475 133.990 ;
        RECT 64.665 133.820 64.835 133.990 ;
        RECT 66.165 133.820 66.335 133.990 ;
        RECT 66.525 133.820 66.695 133.990 ;
        RECT 66.885 133.820 67.055 133.990 ;
        RECT 67.245 133.820 67.415 133.990 ;
        RECT 67.605 133.820 67.775 133.990 ;
        RECT 67.965 133.820 68.135 133.990 ;
        RECT 68.325 133.820 68.495 133.990 ;
        RECT 68.685 133.820 68.855 133.990 ;
        RECT 69.045 133.820 69.215 133.990 ;
        RECT 69.405 133.820 69.575 133.990 ;
        RECT 69.765 133.820 69.935 133.990 ;
        RECT 70.125 133.820 70.295 133.990 ;
        RECT 70.485 133.820 70.655 133.990 ;
        RECT 70.845 133.820 71.015 133.990 ;
        RECT 28.605 131.515 28.775 131.685 ;
        RECT 34.245 131.515 34.415 131.685 ;
        RECT 34.785 131.515 34.955 131.685 ;
        RECT 40.425 131.515 40.595 131.685 ;
        RECT 40.965 131.515 41.135 131.685 ;
        RECT 46.605 131.515 46.775 131.685 ;
        RECT 47.145 131.515 47.315 131.685 ;
        RECT 52.785 131.515 52.955 131.685 ;
        RECT 53.325 131.515 53.495 131.685 ;
        RECT 58.965 131.515 59.135 131.685 ;
        RECT 59.505 131.515 59.675 131.685 ;
        RECT 65.145 131.515 65.315 131.685 ;
        RECT 65.685 131.515 65.855 131.685 ;
        RECT 71.325 131.515 71.495 131.685 ;
        RECT 29.085 131.120 29.255 131.290 ;
        RECT 29.445 131.120 29.615 131.290 ;
        RECT 29.805 131.120 29.975 131.290 ;
        RECT 30.165 131.120 30.335 131.290 ;
        RECT 30.525 131.120 30.695 131.290 ;
        RECT 30.885 131.120 31.055 131.290 ;
        RECT 31.245 131.120 31.415 131.290 ;
        RECT 31.605 131.120 31.775 131.290 ;
        RECT 31.965 131.120 32.135 131.290 ;
        RECT 32.325 131.120 32.495 131.290 ;
        RECT 32.685 131.120 32.855 131.290 ;
        RECT 33.045 131.120 33.215 131.290 ;
        RECT 33.405 131.120 33.575 131.290 ;
        RECT 33.765 131.120 33.935 131.290 ;
        RECT 35.265 131.120 35.435 131.290 ;
        RECT 35.625 131.120 35.795 131.290 ;
        RECT 35.985 131.120 36.155 131.290 ;
        RECT 36.345 131.120 36.515 131.290 ;
        RECT 36.705 131.120 36.875 131.290 ;
        RECT 37.065 131.120 37.235 131.290 ;
        RECT 37.425 131.120 37.595 131.290 ;
        RECT 37.785 131.120 37.955 131.290 ;
        RECT 38.145 131.120 38.315 131.290 ;
        RECT 38.505 131.120 38.675 131.290 ;
        RECT 38.865 131.120 39.035 131.290 ;
        RECT 39.225 131.120 39.395 131.290 ;
        RECT 39.585 131.120 39.755 131.290 ;
        RECT 39.945 131.120 40.115 131.290 ;
        RECT 41.445 131.120 41.615 131.290 ;
        RECT 41.805 131.120 41.975 131.290 ;
        RECT 42.165 131.120 42.335 131.290 ;
        RECT 42.525 131.120 42.695 131.290 ;
        RECT 42.885 131.120 43.055 131.290 ;
        RECT 43.245 131.120 43.415 131.290 ;
        RECT 43.605 131.120 43.775 131.290 ;
        RECT 43.965 131.120 44.135 131.290 ;
        RECT 44.325 131.120 44.495 131.290 ;
        RECT 44.685 131.120 44.855 131.290 ;
        RECT 45.045 131.120 45.215 131.290 ;
        RECT 45.405 131.120 45.575 131.290 ;
        RECT 45.765 131.120 45.935 131.290 ;
        RECT 46.125 131.120 46.295 131.290 ;
        RECT 47.625 131.120 47.795 131.290 ;
        RECT 47.985 131.120 48.155 131.290 ;
        RECT 48.345 131.120 48.515 131.290 ;
        RECT 48.705 131.120 48.875 131.290 ;
        RECT 49.065 131.120 49.235 131.290 ;
        RECT 49.425 131.120 49.595 131.290 ;
        RECT 49.785 131.120 49.955 131.290 ;
        RECT 50.145 131.120 50.315 131.290 ;
        RECT 50.505 131.120 50.675 131.290 ;
        RECT 50.865 131.120 51.035 131.290 ;
        RECT 51.225 131.120 51.395 131.290 ;
        RECT 51.585 131.120 51.755 131.290 ;
        RECT 51.945 131.120 52.115 131.290 ;
        RECT 52.305 131.120 52.475 131.290 ;
        RECT 53.805 131.120 53.975 131.290 ;
        RECT 54.165 131.120 54.335 131.290 ;
        RECT 54.525 131.120 54.695 131.290 ;
        RECT 54.885 131.120 55.055 131.290 ;
        RECT 55.245 131.120 55.415 131.290 ;
        RECT 55.605 131.120 55.775 131.290 ;
        RECT 55.965 131.120 56.135 131.290 ;
        RECT 56.325 131.120 56.495 131.290 ;
        RECT 56.685 131.120 56.855 131.290 ;
        RECT 57.045 131.120 57.215 131.290 ;
        RECT 57.405 131.120 57.575 131.290 ;
        RECT 57.765 131.120 57.935 131.290 ;
        RECT 58.125 131.120 58.295 131.290 ;
        RECT 58.485 131.120 58.655 131.290 ;
        RECT 59.985 131.120 60.155 131.290 ;
        RECT 60.345 131.120 60.515 131.290 ;
        RECT 60.705 131.120 60.875 131.290 ;
        RECT 61.065 131.120 61.235 131.290 ;
        RECT 61.425 131.120 61.595 131.290 ;
        RECT 61.785 131.120 61.955 131.290 ;
        RECT 62.145 131.120 62.315 131.290 ;
        RECT 62.505 131.120 62.675 131.290 ;
        RECT 62.865 131.120 63.035 131.290 ;
        RECT 63.225 131.120 63.395 131.290 ;
        RECT 63.585 131.120 63.755 131.290 ;
        RECT 63.945 131.120 64.115 131.290 ;
        RECT 64.305 131.120 64.475 131.290 ;
        RECT 64.665 131.120 64.835 131.290 ;
        RECT 66.165 131.120 66.335 131.290 ;
        RECT 66.525 131.120 66.695 131.290 ;
        RECT 66.885 131.120 67.055 131.290 ;
        RECT 67.245 131.120 67.415 131.290 ;
        RECT 67.605 131.120 67.775 131.290 ;
        RECT 67.965 131.120 68.135 131.290 ;
        RECT 68.325 131.120 68.495 131.290 ;
        RECT 68.685 131.120 68.855 131.290 ;
        RECT 69.045 131.120 69.215 131.290 ;
        RECT 69.405 131.120 69.575 131.290 ;
        RECT 69.765 131.120 69.935 131.290 ;
        RECT 70.125 131.120 70.295 131.290 ;
        RECT 70.485 131.120 70.655 131.290 ;
        RECT 70.845 131.120 71.015 131.290 ;
        RECT 28.605 128.815 28.775 128.985 ;
        RECT 34.245 128.815 34.415 128.985 ;
        RECT 34.785 128.815 34.955 128.985 ;
        RECT 40.425 128.815 40.595 128.985 ;
        RECT 40.965 128.815 41.135 128.985 ;
        RECT 46.605 128.815 46.775 128.985 ;
        RECT 47.145 128.815 47.315 128.985 ;
        RECT 52.785 128.815 52.955 128.985 ;
        RECT 53.325 128.815 53.495 128.985 ;
        RECT 58.965 128.815 59.135 128.985 ;
        RECT 59.505 128.815 59.675 128.985 ;
        RECT 65.145 128.815 65.315 128.985 ;
        RECT 65.685 128.815 65.855 128.985 ;
        RECT 71.325 128.815 71.495 128.985 ;
        RECT 29.085 128.420 29.255 128.590 ;
        RECT 29.445 128.420 29.615 128.590 ;
        RECT 29.805 128.420 29.975 128.590 ;
        RECT 30.165 128.420 30.335 128.590 ;
        RECT 30.525 128.420 30.695 128.590 ;
        RECT 30.885 128.420 31.055 128.590 ;
        RECT 31.245 128.420 31.415 128.590 ;
        RECT 31.605 128.420 31.775 128.590 ;
        RECT 31.965 128.420 32.135 128.590 ;
        RECT 32.325 128.420 32.495 128.590 ;
        RECT 32.685 128.420 32.855 128.590 ;
        RECT 33.045 128.420 33.215 128.590 ;
        RECT 33.405 128.420 33.575 128.590 ;
        RECT 33.765 128.420 33.935 128.590 ;
        RECT 35.265 128.420 35.435 128.590 ;
        RECT 35.625 128.420 35.795 128.590 ;
        RECT 35.985 128.420 36.155 128.590 ;
        RECT 36.345 128.420 36.515 128.590 ;
        RECT 36.705 128.420 36.875 128.590 ;
        RECT 37.065 128.420 37.235 128.590 ;
        RECT 37.425 128.420 37.595 128.590 ;
        RECT 37.785 128.420 37.955 128.590 ;
        RECT 38.145 128.420 38.315 128.590 ;
        RECT 38.505 128.420 38.675 128.590 ;
        RECT 38.865 128.420 39.035 128.590 ;
        RECT 39.225 128.420 39.395 128.590 ;
        RECT 39.585 128.420 39.755 128.590 ;
        RECT 39.945 128.420 40.115 128.590 ;
        RECT 41.445 128.420 41.615 128.590 ;
        RECT 41.805 128.420 41.975 128.590 ;
        RECT 42.165 128.420 42.335 128.590 ;
        RECT 42.525 128.420 42.695 128.590 ;
        RECT 42.885 128.420 43.055 128.590 ;
        RECT 43.245 128.420 43.415 128.590 ;
        RECT 43.605 128.420 43.775 128.590 ;
        RECT 43.965 128.420 44.135 128.590 ;
        RECT 44.325 128.420 44.495 128.590 ;
        RECT 44.685 128.420 44.855 128.590 ;
        RECT 45.045 128.420 45.215 128.590 ;
        RECT 45.405 128.420 45.575 128.590 ;
        RECT 45.765 128.420 45.935 128.590 ;
        RECT 46.125 128.420 46.295 128.590 ;
        RECT 47.625 128.420 47.795 128.590 ;
        RECT 47.985 128.420 48.155 128.590 ;
        RECT 48.345 128.420 48.515 128.590 ;
        RECT 48.705 128.420 48.875 128.590 ;
        RECT 49.065 128.420 49.235 128.590 ;
        RECT 49.425 128.420 49.595 128.590 ;
        RECT 49.785 128.420 49.955 128.590 ;
        RECT 50.145 128.420 50.315 128.590 ;
        RECT 50.505 128.420 50.675 128.590 ;
        RECT 50.865 128.420 51.035 128.590 ;
        RECT 51.225 128.420 51.395 128.590 ;
        RECT 51.585 128.420 51.755 128.590 ;
        RECT 51.945 128.420 52.115 128.590 ;
        RECT 52.305 128.420 52.475 128.590 ;
        RECT 53.805 128.420 53.975 128.590 ;
        RECT 54.165 128.420 54.335 128.590 ;
        RECT 54.525 128.420 54.695 128.590 ;
        RECT 54.885 128.420 55.055 128.590 ;
        RECT 55.245 128.420 55.415 128.590 ;
        RECT 55.605 128.420 55.775 128.590 ;
        RECT 55.965 128.420 56.135 128.590 ;
        RECT 56.325 128.420 56.495 128.590 ;
        RECT 56.685 128.420 56.855 128.590 ;
        RECT 57.045 128.420 57.215 128.590 ;
        RECT 57.405 128.420 57.575 128.590 ;
        RECT 57.765 128.420 57.935 128.590 ;
        RECT 58.125 128.420 58.295 128.590 ;
        RECT 58.485 128.420 58.655 128.590 ;
        RECT 59.985 128.420 60.155 128.590 ;
        RECT 60.345 128.420 60.515 128.590 ;
        RECT 60.705 128.420 60.875 128.590 ;
        RECT 61.065 128.420 61.235 128.590 ;
        RECT 61.425 128.420 61.595 128.590 ;
        RECT 61.785 128.420 61.955 128.590 ;
        RECT 62.145 128.420 62.315 128.590 ;
        RECT 62.505 128.420 62.675 128.590 ;
        RECT 62.865 128.420 63.035 128.590 ;
        RECT 63.225 128.420 63.395 128.590 ;
        RECT 63.585 128.420 63.755 128.590 ;
        RECT 63.945 128.420 64.115 128.590 ;
        RECT 64.305 128.420 64.475 128.590 ;
        RECT 64.665 128.420 64.835 128.590 ;
        RECT 66.165 128.420 66.335 128.590 ;
        RECT 66.525 128.420 66.695 128.590 ;
        RECT 66.885 128.420 67.055 128.590 ;
        RECT 67.245 128.420 67.415 128.590 ;
        RECT 67.605 128.420 67.775 128.590 ;
        RECT 67.965 128.420 68.135 128.590 ;
        RECT 68.325 128.420 68.495 128.590 ;
        RECT 68.685 128.420 68.855 128.590 ;
        RECT 69.045 128.420 69.215 128.590 ;
        RECT 69.405 128.420 69.575 128.590 ;
        RECT 69.765 128.420 69.935 128.590 ;
        RECT 70.125 128.420 70.295 128.590 ;
        RECT 70.485 128.420 70.655 128.590 ;
        RECT 70.845 128.420 71.015 128.590 ;
        RECT 28.605 125.915 28.775 126.085 ;
        RECT 34.245 125.915 34.415 126.085 ;
        RECT 34.785 125.915 34.955 126.085 ;
        RECT 40.425 125.915 40.595 126.085 ;
        RECT 40.965 125.915 41.135 126.085 ;
        RECT 46.605 125.915 46.775 126.085 ;
        RECT 47.145 125.915 47.315 126.085 ;
        RECT 52.785 125.915 52.955 126.085 ;
        RECT 53.325 125.915 53.495 126.085 ;
        RECT 58.965 125.915 59.135 126.085 ;
        RECT 59.505 125.915 59.675 126.085 ;
        RECT 65.145 125.915 65.315 126.085 ;
        RECT 65.685 125.915 65.855 126.085 ;
        RECT 71.325 125.915 71.495 126.085 ;
        RECT 29.085 125.520 29.255 125.690 ;
        RECT 29.445 125.520 29.615 125.690 ;
        RECT 29.805 125.520 29.975 125.690 ;
        RECT 30.165 125.520 30.335 125.690 ;
        RECT 30.525 125.520 30.695 125.690 ;
        RECT 30.885 125.520 31.055 125.690 ;
        RECT 31.245 125.520 31.415 125.690 ;
        RECT 31.605 125.520 31.775 125.690 ;
        RECT 31.965 125.520 32.135 125.690 ;
        RECT 32.325 125.520 32.495 125.690 ;
        RECT 32.685 125.520 32.855 125.690 ;
        RECT 33.045 125.520 33.215 125.690 ;
        RECT 33.405 125.520 33.575 125.690 ;
        RECT 33.765 125.520 33.935 125.690 ;
        RECT 35.265 125.520 35.435 125.690 ;
        RECT 35.625 125.520 35.795 125.690 ;
        RECT 35.985 125.520 36.155 125.690 ;
        RECT 36.345 125.520 36.515 125.690 ;
        RECT 36.705 125.520 36.875 125.690 ;
        RECT 37.065 125.520 37.235 125.690 ;
        RECT 37.425 125.520 37.595 125.690 ;
        RECT 37.785 125.520 37.955 125.690 ;
        RECT 38.145 125.520 38.315 125.690 ;
        RECT 38.505 125.520 38.675 125.690 ;
        RECT 38.865 125.520 39.035 125.690 ;
        RECT 39.225 125.520 39.395 125.690 ;
        RECT 39.585 125.520 39.755 125.690 ;
        RECT 39.945 125.520 40.115 125.690 ;
        RECT 41.445 125.520 41.615 125.690 ;
        RECT 41.805 125.520 41.975 125.690 ;
        RECT 42.165 125.520 42.335 125.690 ;
        RECT 42.525 125.520 42.695 125.690 ;
        RECT 42.885 125.520 43.055 125.690 ;
        RECT 43.245 125.520 43.415 125.690 ;
        RECT 43.605 125.520 43.775 125.690 ;
        RECT 43.965 125.520 44.135 125.690 ;
        RECT 44.325 125.520 44.495 125.690 ;
        RECT 44.685 125.520 44.855 125.690 ;
        RECT 45.045 125.520 45.215 125.690 ;
        RECT 45.405 125.520 45.575 125.690 ;
        RECT 45.765 125.520 45.935 125.690 ;
        RECT 46.125 125.520 46.295 125.690 ;
        RECT 47.625 125.520 47.795 125.690 ;
        RECT 47.985 125.520 48.155 125.690 ;
        RECT 48.345 125.520 48.515 125.690 ;
        RECT 48.705 125.520 48.875 125.690 ;
        RECT 49.065 125.520 49.235 125.690 ;
        RECT 49.425 125.520 49.595 125.690 ;
        RECT 49.785 125.520 49.955 125.690 ;
        RECT 50.145 125.520 50.315 125.690 ;
        RECT 50.505 125.520 50.675 125.690 ;
        RECT 50.865 125.520 51.035 125.690 ;
        RECT 51.225 125.520 51.395 125.690 ;
        RECT 51.585 125.520 51.755 125.690 ;
        RECT 51.945 125.520 52.115 125.690 ;
        RECT 52.305 125.520 52.475 125.690 ;
        RECT 53.805 125.520 53.975 125.690 ;
        RECT 54.165 125.520 54.335 125.690 ;
        RECT 54.525 125.520 54.695 125.690 ;
        RECT 54.885 125.520 55.055 125.690 ;
        RECT 55.245 125.520 55.415 125.690 ;
        RECT 55.605 125.520 55.775 125.690 ;
        RECT 55.965 125.520 56.135 125.690 ;
        RECT 56.325 125.520 56.495 125.690 ;
        RECT 56.685 125.520 56.855 125.690 ;
        RECT 57.045 125.520 57.215 125.690 ;
        RECT 57.405 125.520 57.575 125.690 ;
        RECT 57.765 125.520 57.935 125.690 ;
        RECT 58.125 125.520 58.295 125.690 ;
        RECT 58.485 125.520 58.655 125.690 ;
        RECT 59.985 125.520 60.155 125.690 ;
        RECT 60.345 125.520 60.515 125.690 ;
        RECT 60.705 125.520 60.875 125.690 ;
        RECT 61.065 125.520 61.235 125.690 ;
        RECT 61.425 125.520 61.595 125.690 ;
        RECT 61.785 125.520 61.955 125.690 ;
        RECT 62.145 125.520 62.315 125.690 ;
        RECT 62.505 125.520 62.675 125.690 ;
        RECT 62.865 125.520 63.035 125.690 ;
        RECT 63.225 125.520 63.395 125.690 ;
        RECT 63.585 125.520 63.755 125.690 ;
        RECT 63.945 125.520 64.115 125.690 ;
        RECT 64.305 125.520 64.475 125.690 ;
        RECT 64.665 125.520 64.835 125.690 ;
        RECT 66.165 125.520 66.335 125.690 ;
        RECT 66.525 125.520 66.695 125.690 ;
        RECT 66.885 125.520 67.055 125.690 ;
        RECT 67.245 125.520 67.415 125.690 ;
        RECT 67.605 125.520 67.775 125.690 ;
        RECT 67.965 125.520 68.135 125.690 ;
        RECT 68.325 125.520 68.495 125.690 ;
        RECT 68.685 125.520 68.855 125.690 ;
        RECT 69.045 125.520 69.215 125.690 ;
        RECT 69.405 125.520 69.575 125.690 ;
        RECT 69.765 125.520 69.935 125.690 ;
        RECT 70.125 125.520 70.295 125.690 ;
        RECT 70.485 125.520 70.655 125.690 ;
        RECT 70.845 125.520 71.015 125.690 ;
        RECT 0.875 117.765 2.845 123.335 ;
        RECT 13.030 117.765 15.000 123.335 ;
        RECT 28.605 123.015 28.775 123.185 ;
        RECT 34.245 123.015 34.415 123.185 ;
        RECT 34.785 123.015 34.955 123.185 ;
        RECT 40.425 123.015 40.595 123.185 ;
        RECT 40.965 123.015 41.135 123.185 ;
        RECT 46.605 123.015 46.775 123.185 ;
        RECT 47.145 123.015 47.315 123.185 ;
        RECT 52.785 123.015 52.955 123.185 ;
        RECT 53.325 123.015 53.495 123.185 ;
        RECT 58.965 123.015 59.135 123.185 ;
        RECT 59.505 123.015 59.675 123.185 ;
        RECT 65.145 123.015 65.315 123.185 ;
        RECT 65.685 123.015 65.855 123.185 ;
        RECT 71.325 123.015 71.495 123.185 ;
        RECT 29.085 122.620 29.255 122.790 ;
        RECT 29.445 122.620 29.615 122.790 ;
        RECT 29.805 122.620 29.975 122.790 ;
        RECT 30.165 122.620 30.335 122.790 ;
        RECT 30.525 122.620 30.695 122.790 ;
        RECT 30.885 122.620 31.055 122.790 ;
        RECT 31.245 122.620 31.415 122.790 ;
        RECT 31.605 122.620 31.775 122.790 ;
        RECT 31.965 122.620 32.135 122.790 ;
        RECT 32.325 122.620 32.495 122.790 ;
        RECT 32.685 122.620 32.855 122.790 ;
        RECT 33.045 122.620 33.215 122.790 ;
        RECT 33.405 122.620 33.575 122.790 ;
        RECT 33.765 122.620 33.935 122.790 ;
        RECT 35.265 122.620 35.435 122.790 ;
        RECT 35.625 122.620 35.795 122.790 ;
        RECT 35.985 122.620 36.155 122.790 ;
        RECT 36.345 122.620 36.515 122.790 ;
        RECT 36.705 122.620 36.875 122.790 ;
        RECT 37.065 122.620 37.235 122.790 ;
        RECT 37.425 122.620 37.595 122.790 ;
        RECT 37.785 122.620 37.955 122.790 ;
        RECT 38.145 122.620 38.315 122.790 ;
        RECT 38.505 122.620 38.675 122.790 ;
        RECT 38.865 122.620 39.035 122.790 ;
        RECT 39.225 122.620 39.395 122.790 ;
        RECT 39.585 122.620 39.755 122.790 ;
        RECT 39.945 122.620 40.115 122.790 ;
        RECT 41.445 122.620 41.615 122.790 ;
        RECT 41.805 122.620 41.975 122.790 ;
        RECT 42.165 122.620 42.335 122.790 ;
        RECT 42.525 122.620 42.695 122.790 ;
        RECT 42.885 122.620 43.055 122.790 ;
        RECT 43.245 122.620 43.415 122.790 ;
        RECT 43.605 122.620 43.775 122.790 ;
        RECT 43.965 122.620 44.135 122.790 ;
        RECT 44.325 122.620 44.495 122.790 ;
        RECT 44.685 122.620 44.855 122.790 ;
        RECT 45.045 122.620 45.215 122.790 ;
        RECT 45.405 122.620 45.575 122.790 ;
        RECT 45.765 122.620 45.935 122.790 ;
        RECT 46.125 122.620 46.295 122.790 ;
        RECT 47.625 122.620 47.795 122.790 ;
        RECT 47.985 122.620 48.155 122.790 ;
        RECT 48.345 122.620 48.515 122.790 ;
        RECT 48.705 122.620 48.875 122.790 ;
        RECT 49.065 122.620 49.235 122.790 ;
        RECT 49.425 122.620 49.595 122.790 ;
        RECT 49.785 122.620 49.955 122.790 ;
        RECT 50.145 122.620 50.315 122.790 ;
        RECT 50.505 122.620 50.675 122.790 ;
        RECT 50.865 122.620 51.035 122.790 ;
        RECT 51.225 122.620 51.395 122.790 ;
        RECT 51.585 122.620 51.755 122.790 ;
        RECT 51.945 122.620 52.115 122.790 ;
        RECT 52.305 122.620 52.475 122.790 ;
        RECT 53.805 122.620 53.975 122.790 ;
        RECT 54.165 122.620 54.335 122.790 ;
        RECT 54.525 122.620 54.695 122.790 ;
        RECT 54.885 122.620 55.055 122.790 ;
        RECT 55.245 122.620 55.415 122.790 ;
        RECT 55.605 122.620 55.775 122.790 ;
        RECT 55.965 122.620 56.135 122.790 ;
        RECT 56.325 122.620 56.495 122.790 ;
        RECT 56.685 122.620 56.855 122.790 ;
        RECT 57.045 122.620 57.215 122.790 ;
        RECT 57.405 122.620 57.575 122.790 ;
        RECT 57.765 122.620 57.935 122.790 ;
        RECT 58.125 122.620 58.295 122.790 ;
        RECT 58.485 122.620 58.655 122.790 ;
        RECT 59.985 122.620 60.155 122.790 ;
        RECT 60.345 122.620 60.515 122.790 ;
        RECT 60.705 122.620 60.875 122.790 ;
        RECT 61.065 122.620 61.235 122.790 ;
        RECT 61.425 122.620 61.595 122.790 ;
        RECT 61.785 122.620 61.955 122.790 ;
        RECT 62.145 122.620 62.315 122.790 ;
        RECT 62.505 122.620 62.675 122.790 ;
        RECT 62.865 122.620 63.035 122.790 ;
        RECT 63.225 122.620 63.395 122.790 ;
        RECT 63.585 122.620 63.755 122.790 ;
        RECT 63.945 122.620 64.115 122.790 ;
        RECT 64.305 122.620 64.475 122.790 ;
        RECT 64.665 122.620 64.835 122.790 ;
        RECT 66.165 122.620 66.335 122.790 ;
        RECT 66.525 122.620 66.695 122.790 ;
        RECT 66.885 122.620 67.055 122.790 ;
        RECT 67.245 122.620 67.415 122.790 ;
        RECT 67.605 122.620 67.775 122.790 ;
        RECT 67.965 122.620 68.135 122.790 ;
        RECT 68.325 122.620 68.495 122.790 ;
        RECT 68.685 122.620 68.855 122.790 ;
        RECT 69.045 122.620 69.215 122.790 ;
        RECT 69.405 122.620 69.575 122.790 ;
        RECT 69.765 122.620 69.935 122.790 ;
        RECT 70.125 122.620 70.295 122.790 ;
        RECT 70.485 122.620 70.655 122.790 ;
        RECT 70.845 122.620 71.015 122.790 ;
        RECT 19.405 120.315 19.575 120.485 ;
        RECT 25.045 120.315 25.215 120.485 ;
        RECT 25.585 120.315 25.755 120.485 ;
        RECT 31.225 120.315 31.395 120.485 ;
        RECT 31.765 120.315 31.935 120.485 ;
        RECT 37.405 120.315 37.575 120.485 ;
        RECT 37.945 120.315 38.115 120.485 ;
        RECT 43.585 120.315 43.755 120.485 ;
        RECT 44.125 120.315 44.295 120.485 ;
        RECT 49.765 120.315 49.935 120.485 ;
        RECT 50.305 120.315 50.475 120.485 ;
        RECT 55.945 120.315 56.115 120.485 ;
        RECT 56.485 120.315 56.655 120.485 ;
        RECT 62.125 120.315 62.295 120.485 ;
        RECT 62.665 120.315 62.835 120.485 ;
        RECT 68.305 120.315 68.475 120.485 ;
        RECT 68.845 120.315 69.015 120.485 ;
        RECT 74.485 120.315 74.655 120.485 ;
        RECT 75.025 120.315 75.195 120.485 ;
        RECT 80.665 120.315 80.835 120.485 ;
        RECT 19.405 117.615 19.575 117.785 ;
        RECT 25.045 117.615 25.215 117.785 ;
        RECT 25.585 117.615 25.755 117.785 ;
        RECT 31.225 117.615 31.395 117.785 ;
        RECT 31.765 117.615 31.935 117.785 ;
        RECT 37.405 117.615 37.575 117.785 ;
        RECT 37.945 117.615 38.115 117.785 ;
        RECT 43.585 117.615 43.755 117.785 ;
        RECT 44.125 117.615 44.295 117.785 ;
        RECT 49.765 117.615 49.935 117.785 ;
        RECT 50.305 117.615 50.475 117.785 ;
        RECT 55.945 117.615 56.115 117.785 ;
        RECT 56.485 117.615 56.655 117.785 ;
        RECT 62.125 117.615 62.295 117.785 ;
        RECT 62.665 117.615 62.835 117.785 ;
        RECT 68.305 117.615 68.475 117.785 ;
        RECT 68.845 117.615 69.015 117.785 ;
        RECT 74.485 117.615 74.655 117.785 ;
        RECT 75.025 117.615 75.195 117.785 ;
        RECT 80.665 117.615 80.835 117.785 ;
        RECT 86.175 117.765 88.145 123.335 ;
        RECT 98.330 117.765 100.300 123.335 ;
        RECT 0.875 110.415 2.845 115.985 ;
        RECT 13.030 110.415 15.000 115.985 ;
        RECT 19.405 114.915 19.575 115.085 ;
        RECT 25.045 114.915 25.215 115.085 ;
        RECT 25.585 114.915 25.755 115.085 ;
        RECT 31.225 114.915 31.395 115.085 ;
        RECT 31.765 114.915 31.935 115.085 ;
        RECT 37.405 114.915 37.575 115.085 ;
        RECT 37.945 114.915 38.115 115.085 ;
        RECT 43.585 114.915 43.755 115.085 ;
        RECT 44.125 114.915 44.295 115.085 ;
        RECT 49.765 114.915 49.935 115.085 ;
        RECT 50.305 114.915 50.475 115.085 ;
        RECT 55.945 114.915 56.115 115.085 ;
        RECT 56.485 114.915 56.655 115.085 ;
        RECT 62.125 114.915 62.295 115.085 ;
        RECT 62.665 114.915 62.835 115.085 ;
        RECT 68.305 114.915 68.475 115.085 ;
        RECT 68.845 114.915 69.015 115.085 ;
        RECT 74.485 114.915 74.655 115.085 ;
        RECT 75.025 114.915 75.195 115.085 ;
        RECT 80.665 114.915 80.835 115.085 ;
        RECT 19.405 112.215 19.575 112.385 ;
        RECT 25.045 112.215 25.215 112.385 ;
        RECT 25.585 112.215 25.755 112.385 ;
        RECT 31.225 112.215 31.395 112.385 ;
        RECT 31.765 112.215 31.935 112.385 ;
        RECT 37.405 112.215 37.575 112.385 ;
        RECT 37.945 112.215 38.115 112.385 ;
        RECT 43.585 112.215 43.755 112.385 ;
        RECT 44.125 112.215 44.295 112.385 ;
        RECT 49.765 112.215 49.935 112.385 ;
        RECT 50.305 112.215 50.475 112.385 ;
        RECT 55.945 112.215 56.115 112.385 ;
        RECT 56.485 112.215 56.655 112.385 ;
        RECT 62.125 112.215 62.295 112.385 ;
        RECT 62.665 112.215 62.835 112.385 ;
        RECT 68.305 112.215 68.475 112.385 ;
        RECT 68.845 112.215 69.015 112.385 ;
        RECT 74.485 112.215 74.655 112.385 ;
        RECT 75.025 112.215 75.195 112.385 ;
        RECT 80.665 112.215 80.835 112.385 ;
        RECT 86.175 110.415 88.145 115.985 ;
        RECT 98.330 110.415 100.300 115.985 ;
        RECT 29.540 108.710 29.710 108.880 ;
        RECT 29.900 108.710 30.070 108.880 ;
        RECT 30.260 108.710 30.430 108.880 ;
        RECT 30.620 108.710 30.790 108.880 ;
        RECT 30.980 108.710 31.150 108.880 ;
        RECT 31.340 108.710 31.510 108.880 ;
        RECT 31.700 108.710 31.870 108.880 ;
        RECT 32.060 108.710 32.230 108.880 ;
        RECT 32.420 108.710 32.590 108.880 ;
        RECT 32.780 108.710 32.950 108.880 ;
        RECT 33.140 108.710 33.310 108.880 ;
        RECT 33.500 108.710 33.670 108.880 ;
        RECT 33.860 108.710 34.030 108.880 ;
        RECT 34.220 108.710 34.390 108.880 ;
        RECT 35.630 108.710 35.800 108.880 ;
        RECT 35.990 108.710 36.160 108.880 ;
        RECT 36.350 108.710 36.520 108.880 ;
        RECT 36.710 108.710 36.880 108.880 ;
        RECT 37.070 108.710 37.240 108.880 ;
        RECT 37.430 108.710 37.600 108.880 ;
        RECT 37.790 108.710 37.960 108.880 ;
        RECT 38.150 108.710 38.320 108.880 ;
        RECT 38.510 108.710 38.680 108.880 ;
        RECT 38.870 108.710 39.040 108.880 ;
        RECT 39.230 108.710 39.400 108.880 ;
        RECT 39.590 108.710 39.760 108.880 ;
        RECT 39.950 108.710 40.120 108.880 ;
        RECT 40.310 108.710 40.480 108.880 ;
        RECT 41.720 108.710 41.890 108.880 ;
        RECT 42.080 108.710 42.250 108.880 ;
        RECT 42.440 108.710 42.610 108.880 ;
        RECT 42.800 108.710 42.970 108.880 ;
        RECT 43.160 108.710 43.330 108.880 ;
        RECT 43.520 108.710 43.690 108.880 ;
        RECT 43.880 108.710 44.050 108.880 ;
        RECT 44.240 108.710 44.410 108.880 ;
        RECT 44.600 108.710 44.770 108.880 ;
        RECT 44.960 108.710 45.130 108.880 ;
        RECT 45.320 108.710 45.490 108.880 ;
        RECT 45.680 108.710 45.850 108.880 ;
        RECT 46.040 108.710 46.210 108.880 ;
        RECT 46.400 108.710 46.570 108.880 ;
        RECT 47.810 108.710 47.980 108.880 ;
        RECT 48.170 108.710 48.340 108.880 ;
        RECT 48.530 108.710 48.700 108.880 ;
        RECT 48.890 108.710 49.060 108.880 ;
        RECT 49.250 108.710 49.420 108.880 ;
        RECT 49.610 108.710 49.780 108.880 ;
        RECT 49.970 108.710 50.140 108.880 ;
        RECT 50.330 108.710 50.500 108.880 ;
        RECT 50.690 108.710 50.860 108.880 ;
        RECT 51.050 108.710 51.220 108.880 ;
        RECT 51.410 108.710 51.580 108.880 ;
        RECT 51.770 108.710 51.940 108.880 ;
        RECT 52.130 108.710 52.300 108.880 ;
        RECT 52.490 108.710 52.660 108.880 ;
        RECT 53.900 108.710 54.070 108.880 ;
        RECT 54.260 108.710 54.430 108.880 ;
        RECT 54.620 108.710 54.790 108.880 ;
        RECT 54.980 108.710 55.150 108.880 ;
        RECT 55.340 108.710 55.510 108.880 ;
        RECT 55.700 108.710 55.870 108.880 ;
        RECT 56.060 108.710 56.230 108.880 ;
        RECT 56.420 108.710 56.590 108.880 ;
        RECT 56.780 108.710 56.950 108.880 ;
        RECT 57.140 108.710 57.310 108.880 ;
        RECT 57.500 108.710 57.670 108.880 ;
        RECT 57.860 108.710 58.030 108.880 ;
        RECT 58.220 108.710 58.390 108.880 ;
        RECT 58.580 108.710 58.750 108.880 ;
        RECT 59.990 108.710 60.160 108.880 ;
        RECT 60.350 108.710 60.520 108.880 ;
        RECT 60.710 108.710 60.880 108.880 ;
        RECT 61.070 108.710 61.240 108.880 ;
        RECT 61.430 108.710 61.600 108.880 ;
        RECT 61.790 108.710 61.960 108.880 ;
        RECT 62.150 108.710 62.320 108.880 ;
        RECT 62.510 108.710 62.680 108.880 ;
        RECT 62.870 108.710 63.040 108.880 ;
        RECT 63.230 108.710 63.400 108.880 ;
        RECT 63.590 108.710 63.760 108.880 ;
        RECT 63.950 108.710 64.120 108.880 ;
        RECT 64.310 108.710 64.480 108.880 ;
        RECT 64.670 108.710 64.840 108.880 ;
        RECT 66.080 108.710 66.250 108.880 ;
        RECT 66.440 108.710 66.610 108.880 ;
        RECT 66.800 108.710 66.970 108.880 ;
        RECT 67.160 108.710 67.330 108.880 ;
        RECT 67.520 108.710 67.690 108.880 ;
        RECT 67.880 108.710 68.050 108.880 ;
        RECT 68.240 108.710 68.410 108.880 ;
        RECT 68.600 108.710 68.770 108.880 ;
        RECT 68.960 108.710 69.130 108.880 ;
        RECT 69.320 108.710 69.490 108.880 ;
        RECT 69.680 108.710 69.850 108.880 ;
        RECT 70.040 108.710 70.210 108.880 ;
        RECT 70.400 108.710 70.570 108.880 ;
        RECT 70.760 108.710 70.930 108.880 ;
        RECT 29.540 107.920 29.710 108.090 ;
        RECT 29.900 107.920 30.070 108.090 ;
        RECT 30.260 107.920 30.430 108.090 ;
        RECT 30.620 107.920 30.790 108.090 ;
        RECT 30.980 107.920 31.150 108.090 ;
        RECT 31.340 107.920 31.510 108.090 ;
        RECT 31.700 107.920 31.870 108.090 ;
        RECT 32.060 107.920 32.230 108.090 ;
        RECT 32.420 107.920 32.590 108.090 ;
        RECT 32.780 107.920 32.950 108.090 ;
        RECT 33.140 107.920 33.310 108.090 ;
        RECT 33.500 107.920 33.670 108.090 ;
        RECT 33.860 107.920 34.030 108.090 ;
        RECT 34.220 107.920 34.390 108.090 ;
        RECT 35.630 107.920 35.800 108.090 ;
        RECT 35.990 107.920 36.160 108.090 ;
        RECT 36.350 107.920 36.520 108.090 ;
        RECT 36.710 107.920 36.880 108.090 ;
        RECT 37.070 107.920 37.240 108.090 ;
        RECT 37.430 107.920 37.600 108.090 ;
        RECT 37.790 107.920 37.960 108.090 ;
        RECT 38.150 107.920 38.320 108.090 ;
        RECT 38.510 107.920 38.680 108.090 ;
        RECT 38.870 107.920 39.040 108.090 ;
        RECT 39.230 107.920 39.400 108.090 ;
        RECT 39.590 107.920 39.760 108.090 ;
        RECT 39.950 107.920 40.120 108.090 ;
        RECT 40.310 107.920 40.480 108.090 ;
        RECT 41.720 107.920 41.890 108.090 ;
        RECT 42.080 107.920 42.250 108.090 ;
        RECT 42.440 107.920 42.610 108.090 ;
        RECT 42.800 107.920 42.970 108.090 ;
        RECT 43.160 107.920 43.330 108.090 ;
        RECT 43.520 107.920 43.690 108.090 ;
        RECT 43.880 107.920 44.050 108.090 ;
        RECT 44.240 107.920 44.410 108.090 ;
        RECT 44.600 107.920 44.770 108.090 ;
        RECT 44.960 107.920 45.130 108.090 ;
        RECT 45.320 107.920 45.490 108.090 ;
        RECT 45.680 107.920 45.850 108.090 ;
        RECT 46.040 107.920 46.210 108.090 ;
        RECT 46.400 107.920 46.570 108.090 ;
        RECT 47.810 107.920 47.980 108.090 ;
        RECT 48.170 107.920 48.340 108.090 ;
        RECT 48.530 107.920 48.700 108.090 ;
        RECT 48.890 107.920 49.060 108.090 ;
        RECT 49.250 107.920 49.420 108.090 ;
        RECT 49.610 107.920 49.780 108.090 ;
        RECT 49.970 107.920 50.140 108.090 ;
        RECT 50.330 107.920 50.500 108.090 ;
        RECT 50.690 107.920 50.860 108.090 ;
        RECT 51.050 107.920 51.220 108.090 ;
        RECT 51.410 107.920 51.580 108.090 ;
        RECT 51.770 107.920 51.940 108.090 ;
        RECT 52.130 107.920 52.300 108.090 ;
        RECT 52.490 107.920 52.660 108.090 ;
        RECT 53.900 107.920 54.070 108.090 ;
        RECT 54.260 107.920 54.430 108.090 ;
        RECT 54.620 107.920 54.790 108.090 ;
        RECT 54.980 107.920 55.150 108.090 ;
        RECT 55.340 107.920 55.510 108.090 ;
        RECT 55.700 107.920 55.870 108.090 ;
        RECT 56.060 107.920 56.230 108.090 ;
        RECT 56.420 107.920 56.590 108.090 ;
        RECT 56.780 107.920 56.950 108.090 ;
        RECT 57.140 107.920 57.310 108.090 ;
        RECT 57.500 107.920 57.670 108.090 ;
        RECT 57.860 107.920 58.030 108.090 ;
        RECT 58.220 107.920 58.390 108.090 ;
        RECT 58.580 107.920 58.750 108.090 ;
        RECT 59.990 107.920 60.160 108.090 ;
        RECT 60.350 107.920 60.520 108.090 ;
        RECT 60.710 107.920 60.880 108.090 ;
        RECT 61.070 107.920 61.240 108.090 ;
        RECT 61.430 107.920 61.600 108.090 ;
        RECT 61.790 107.920 61.960 108.090 ;
        RECT 62.150 107.920 62.320 108.090 ;
        RECT 62.510 107.920 62.680 108.090 ;
        RECT 62.870 107.920 63.040 108.090 ;
        RECT 63.230 107.920 63.400 108.090 ;
        RECT 63.590 107.920 63.760 108.090 ;
        RECT 63.950 107.920 64.120 108.090 ;
        RECT 64.310 107.920 64.480 108.090 ;
        RECT 64.670 107.920 64.840 108.090 ;
        RECT 66.080 107.920 66.250 108.090 ;
        RECT 66.440 107.920 66.610 108.090 ;
        RECT 66.800 107.920 66.970 108.090 ;
        RECT 67.160 107.920 67.330 108.090 ;
        RECT 67.520 107.920 67.690 108.090 ;
        RECT 67.880 107.920 68.050 108.090 ;
        RECT 68.240 107.920 68.410 108.090 ;
        RECT 68.600 107.920 68.770 108.090 ;
        RECT 68.960 107.920 69.130 108.090 ;
        RECT 69.320 107.920 69.490 108.090 ;
        RECT 69.680 107.920 69.850 108.090 ;
        RECT 70.040 107.920 70.210 108.090 ;
        RECT 70.400 107.920 70.570 108.090 ;
        RECT 70.760 107.920 70.930 108.090 ;
        RECT 29.540 106.210 29.710 106.380 ;
        RECT 29.900 106.210 30.070 106.380 ;
        RECT 30.260 106.210 30.430 106.380 ;
        RECT 30.620 106.210 30.790 106.380 ;
        RECT 30.980 106.210 31.150 106.380 ;
        RECT 31.340 106.210 31.510 106.380 ;
        RECT 31.700 106.210 31.870 106.380 ;
        RECT 32.060 106.210 32.230 106.380 ;
        RECT 32.420 106.210 32.590 106.380 ;
        RECT 32.780 106.210 32.950 106.380 ;
        RECT 33.140 106.210 33.310 106.380 ;
        RECT 33.500 106.210 33.670 106.380 ;
        RECT 33.860 106.210 34.030 106.380 ;
        RECT 34.220 106.210 34.390 106.380 ;
        RECT 35.630 106.210 35.800 106.380 ;
        RECT 35.990 106.210 36.160 106.380 ;
        RECT 36.350 106.210 36.520 106.380 ;
        RECT 36.710 106.210 36.880 106.380 ;
        RECT 37.070 106.210 37.240 106.380 ;
        RECT 37.430 106.210 37.600 106.380 ;
        RECT 37.790 106.210 37.960 106.380 ;
        RECT 38.150 106.210 38.320 106.380 ;
        RECT 38.510 106.210 38.680 106.380 ;
        RECT 38.870 106.210 39.040 106.380 ;
        RECT 39.230 106.210 39.400 106.380 ;
        RECT 39.590 106.210 39.760 106.380 ;
        RECT 39.950 106.210 40.120 106.380 ;
        RECT 40.310 106.210 40.480 106.380 ;
        RECT 41.720 106.210 41.890 106.380 ;
        RECT 42.080 106.210 42.250 106.380 ;
        RECT 42.440 106.210 42.610 106.380 ;
        RECT 42.800 106.210 42.970 106.380 ;
        RECT 43.160 106.210 43.330 106.380 ;
        RECT 43.520 106.210 43.690 106.380 ;
        RECT 43.880 106.210 44.050 106.380 ;
        RECT 44.240 106.210 44.410 106.380 ;
        RECT 44.600 106.210 44.770 106.380 ;
        RECT 44.960 106.210 45.130 106.380 ;
        RECT 45.320 106.210 45.490 106.380 ;
        RECT 45.680 106.210 45.850 106.380 ;
        RECT 46.040 106.210 46.210 106.380 ;
        RECT 46.400 106.210 46.570 106.380 ;
        RECT 47.810 106.210 47.980 106.380 ;
        RECT 48.170 106.210 48.340 106.380 ;
        RECT 48.530 106.210 48.700 106.380 ;
        RECT 48.890 106.210 49.060 106.380 ;
        RECT 49.250 106.210 49.420 106.380 ;
        RECT 49.610 106.210 49.780 106.380 ;
        RECT 49.970 106.210 50.140 106.380 ;
        RECT 50.330 106.210 50.500 106.380 ;
        RECT 50.690 106.210 50.860 106.380 ;
        RECT 51.050 106.210 51.220 106.380 ;
        RECT 51.410 106.210 51.580 106.380 ;
        RECT 51.770 106.210 51.940 106.380 ;
        RECT 52.130 106.210 52.300 106.380 ;
        RECT 52.490 106.210 52.660 106.380 ;
        RECT 53.900 106.210 54.070 106.380 ;
        RECT 54.260 106.210 54.430 106.380 ;
        RECT 54.620 106.210 54.790 106.380 ;
        RECT 54.980 106.210 55.150 106.380 ;
        RECT 55.340 106.210 55.510 106.380 ;
        RECT 55.700 106.210 55.870 106.380 ;
        RECT 56.060 106.210 56.230 106.380 ;
        RECT 56.420 106.210 56.590 106.380 ;
        RECT 56.780 106.210 56.950 106.380 ;
        RECT 57.140 106.210 57.310 106.380 ;
        RECT 57.500 106.210 57.670 106.380 ;
        RECT 57.860 106.210 58.030 106.380 ;
        RECT 58.220 106.210 58.390 106.380 ;
        RECT 58.580 106.210 58.750 106.380 ;
        RECT 59.990 106.210 60.160 106.380 ;
        RECT 60.350 106.210 60.520 106.380 ;
        RECT 60.710 106.210 60.880 106.380 ;
        RECT 61.070 106.210 61.240 106.380 ;
        RECT 61.430 106.210 61.600 106.380 ;
        RECT 61.790 106.210 61.960 106.380 ;
        RECT 62.150 106.210 62.320 106.380 ;
        RECT 62.510 106.210 62.680 106.380 ;
        RECT 62.870 106.210 63.040 106.380 ;
        RECT 63.230 106.210 63.400 106.380 ;
        RECT 63.590 106.210 63.760 106.380 ;
        RECT 63.950 106.210 64.120 106.380 ;
        RECT 64.310 106.210 64.480 106.380 ;
        RECT 64.670 106.210 64.840 106.380 ;
        RECT 66.080 106.210 66.250 106.380 ;
        RECT 66.440 106.210 66.610 106.380 ;
        RECT 66.800 106.210 66.970 106.380 ;
        RECT 67.160 106.210 67.330 106.380 ;
        RECT 67.520 106.210 67.690 106.380 ;
        RECT 67.880 106.210 68.050 106.380 ;
        RECT 68.240 106.210 68.410 106.380 ;
        RECT 68.600 106.210 68.770 106.380 ;
        RECT 68.960 106.210 69.130 106.380 ;
        RECT 69.320 106.210 69.490 106.380 ;
        RECT 69.680 106.210 69.850 106.380 ;
        RECT 70.040 106.210 70.210 106.380 ;
        RECT 70.400 106.210 70.570 106.380 ;
        RECT 70.760 106.210 70.930 106.380 ;
        RECT 29.540 105.420 29.710 105.590 ;
        RECT 29.900 105.420 30.070 105.590 ;
        RECT 30.260 105.420 30.430 105.590 ;
        RECT 30.620 105.420 30.790 105.590 ;
        RECT 30.980 105.420 31.150 105.590 ;
        RECT 31.340 105.420 31.510 105.590 ;
        RECT 31.700 105.420 31.870 105.590 ;
        RECT 32.060 105.420 32.230 105.590 ;
        RECT 32.420 105.420 32.590 105.590 ;
        RECT 32.780 105.420 32.950 105.590 ;
        RECT 33.140 105.420 33.310 105.590 ;
        RECT 33.500 105.420 33.670 105.590 ;
        RECT 33.860 105.420 34.030 105.590 ;
        RECT 34.220 105.420 34.390 105.590 ;
        RECT 35.630 105.420 35.800 105.590 ;
        RECT 35.990 105.420 36.160 105.590 ;
        RECT 36.350 105.420 36.520 105.590 ;
        RECT 36.710 105.420 36.880 105.590 ;
        RECT 37.070 105.420 37.240 105.590 ;
        RECT 37.430 105.420 37.600 105.590 ;
        RECT 37.790 105.420 37.960 105.590 ;
        RECT 38.150 105.420 38.320 105.590 ;
        RECT 38.510 105.420 38.680 105.590 ;
        RECT 38.870 105.420 39.040 105.590 ;
        RECT 39.230 105.420 39.400 105.590 ;
        RECT 39.590 105.420 39.760 105.590 ;
        RECT 39.950 105.420 40.120 105.590 ;
        RECT 40.310 105.420 40.480 105.590 ;
        RECT 41.720 105.420 41.890 105.590 ;
        RECT 42.080 105.420 42.250 105.590 ;
        RECT 42.440 105.420 42.610 105.590 ;
        RECT 42.800 105.420 42.970 105.590 ;
        RECT 43.160 105.420 43.330 105.590 ;
        RECT 43.520 105.420 43.690 105.590 ;
        RECT 43.880 105.420 44.050 105.590 ;
        RECT 44.240 105.420 44.410 105.590 ;
        RECT 44.600 105.420 44.770 105.590 ;
        RECT 44.960 105.420 45.130 105.590 ;
        RECT 45.320 105.420 45.490 105.590 ;
        RECT 45.680 105.420 45.850 105.590 ;
        RECT 46.040 105.420 46.210 105.590 ;
        RECT 46.400 105.420 46.570 105.590 ;
        RECT 47.810 105.420 47.980 105.590 ;
        RECT 48.170 105.420 48.340 105.590 ;
        RECT 48.530 105.420 48.700 105.590 ;
        RECT 48.890 105.420 49.060 105.590 ;
        RECT 49.250 105.420 49.420 105.590 ;
        RECT 49.610 105.420 49.780 105.590 ;
        RECT 49.970 105.420 50.140 105.590 ;
        RECT 50.330 105.420 50.500 105.590 ;
        RECT 50.690 105.420 50.860 105.590 ;
        RECT 51.050 105.420 51.220 105.590 ;
        RECT 51.410 105.420 51.580 105.590 ;
        RECT 51.770 105.420 51.940 105.590 ;
        RECT 52.130 105.420 52.300 105.590 ;
        RECT 52.490 105.420 52.660 105.590 ;
        RECT 53.900 105.420 54.070 105.590 ;
        RECT 54.260 105.420 54.430 105.590 ;
        RECT 54.620 105.420 54.790 105.590 ;
        RECT 54.980 105.420 55.150 105.590 ;
        RECT 55.340 105.420 55.510 105.590 ;
        RECT 55.700 105.420 55.870 105.590 ;
        RECT 56.060 105.420 56.230 105.590 ;
        RECT 56.420 105.420 56.590 105.590 ;
        RECT 56.780 105.420 56.950 105.590 ;
        RECT 57.140 105.420 57.310 105.590 ;
        RECT 57.500 105.420 57.670 105.590 ;
        RECT 57.860 105.420 58.030 105.590 ;
        RECT 58.220 105.420 58.390 105.590 ;
        RECT 58.580 105.420 58.750 105.590 ;
        RECT 59.990 105.420 60.160 105.590 ;
        RECT 60.350 105.420 60.520 105.590 ;
        RECT 60.710 105.420 60.880 105.590 ;
        RECT 61.070 105.420 61.240 105.590 ;
        RECT 61.430 105.420 61.600 105.590 ;
        RECT 61.790 105.420 61.960 105.590 ;
        RECT 62.150 105.420 62.320 105.590 ;
        RECT 62.510 105.420 62.680 105.590 ;
        RECT 62.870 105.420 63.040 105.590 ;
        RECT 63.230 105.420 63.400 105.590 ;
        RECT 63.590 105.420 63.760 105.590 ;
        RECT 63.950 105.420 64.120 105.590 ;
        RECT 64.310 105.420 64.480 105.590 ;
        RECT 64.670 105.420 64.840 105.590 ;
        RECT 66.080 105.420 66.250 105.590 ;
        RECT 66.440 105.420 66.610 105.590 ;
        RECT 66.800 105.420 66.970 105.590 ;
        RECT 67.160 105.420 67.330 105.590 ;
        RECT 67.520 105.420 67.690 105.590 ;
        RECT 67.880 105.420 68.050 105.590 ;
        RECT 68.240 105.420 68.410 105.590 ;
        RECT 68.600 105.420 68.770 105.590 ;
        RECT 68.960 105.420 69.130 105.590 ;
        RECT 69.320 105.420 69.490 105.590 ;
        RECT 69.680 105.420 69.850 105.590 ;
        RECT 70.040 105.420 70.210 105.590 ;
        RECT 70.400 105.420 70.570 105.590 ;
        RECT 70.760 105.420 70.930 105.590 ;
        RECT 31.905 103.245 32.075 103.415 ;
        RECT 31.905 102.885 32.075 103.055 ;
        RECT 37.455 103.245 37.625 103.415 ;
        RECT 37.455 102.885 37.625 103.055 ;
        RECT 37.995 103.245 38.165 103.415 ;
        RECT 37.995 102.885 38.165 103.055 ;
        RECT 43.545 103.245 43.715 103.415 ;
        RECT 43.545 102.885 43.715 103.055 ;
        RECT 44.085 103.245 44.255 103.415 ;
        RECT 44.085 102.885 44.255 103.055 ;
        RECT 49.635 103.245 49.805 103.415 ;
        RECT 49.635 102.885 49.805 103.055 ;
        RECT 50.175 103.245 50.345 103.415 ;
        RECT 50.175 102.885 50.345 103.055 ;
        RECT 55.725 103.245 55.895 103.415 ;
        RECT 55.725 102.885 55.895 103.055 ;
        RECT 56.265 103.245 56.435 103.415 ;
        RECT 56.265 102.885 56.435 103.055 ;
        RECT 61.815 103.245 61.985 103.415 ;
        RECT 61.815 102.885 61.985 103.055 ;
        RECT 62.355 103.245 62.525 103.415 ;
        RECT 62.355 102.885 62.525 103.055 ;
        RECT 67.905 103.245 68.075 103.415 ;
        RECT 67.905 102.885 68.075 103.055 ;
        RECT 31.905 100.145 32.075 100.315 ;
        RECT 31.905 99.785 32.075 99.955 ;
        RECT 37.455 100.145 37.625 100.315 ;
        RECT 37.455 99.785 37.625 99.955 ;
        RECT 37.995 100.145 38.165 100.315 ;
        RECT 37.995 99.785 38.165 99.955 ;
        RECT 43.545 100.145 43.715 100.315 ;
        RECT 43.545 99.785 43.715 99.955 ;
        RECT 44.085 100.145 44.255 100.315 ;
        RECT 44.085 99.785 44.255 99.955 ;
        RECT 49.635 100.145 49.805 100.315 ;
        RECT 49.635 99.785 49.805 99.955 ;
        RECT 50.175 100.145 50.345 100.315 ;
        RECT 50.175 99.785 50.345 99.955 ;
        RECT 55.725 100.145 55.895 100.315 ;
        RECT 55.725 99.785 55.895 99.955 ;
        RECT 56.265 100.145 56.435 100.315 ;
        RECT 56.265 99.785 56.435 99.955 ;
        RECT 61.815 100.145 61.985 100.315 ;
        RECT 61.815 99.785 61.985 99.955 ;
        RECT 62.355 100.145 62.525 100.315 ;
        RECT 62.355 99.785 62.525 99.955 ;
        RECT 67.905 100.145 68.075 100.315 ;
        RECT 67.905 99.785 68.075 99.955 ;
        RECT 29.105 97.145 29.275 97.315 ;
        RECT 29.105 96.785 29.275 96.955 ;
        RECT 34.655 97.145 34.825 97.315 ;
        RECT 34.655 96.785 34.825 96.955 ;
        RECT 35.195 97.145 35.365 97.315 ;
        RECT 35.195 96.785 35.365 96.955 ;
        RECT 40.745 97.145 40.915 97.315 ;
        RECT 40.745 96.785 40.915 96.955 ;
        RECT 41.285 97.145 41.455 97.315 ;
        RECT 41.285 96.785 41.455 96.955 ;
        RECT 46.835 97.145 47.005 97.315 ;
        RECT 46.835 96.785 47.005 96.955 ;
        RECT 47.375 97.145 47.545 97.315 ;
        RECT 47.375 96.785 47.545 96.955 ;
        RECT 52.925 97.145 53.095 97.315 ;
        RECT 52.925 96.785 53.095 96.955 ;
        RECT 53.465 97.145 53.635 97.315 ;
        RECT 53.465 96.785 53.635 96.955 ;
        RECT 59.015 97.145 59.185 97.315 ;
        RECT 59.015 96.785 59.185 96.955 ;
        RECT 59.555 97.145 59.725 97.315 ;
        RECT 59.555 96.785 59.725 96.955 ;
        RECT 65.105 97.145 65.275 97.315 ;
        RECT 65.105 96.785 65.275 96.955 ;
        RECT 65.645 97.145 65.815 97.315 ;
        RECT 65.645 96.785 65.815 96.955 ;
        RECT 71.195 97.145 71.365 97.315 ;
        RECT 71.195 96.785 71.365 96.955 ;
        RECT 29.540 96.320 29.710 96.490 ;
        RECT 29.900 96.320 30.070 96.490 ;
        RECT 30.260 96.320 30.430 96.490 ;
        RECT 30.620 96.320 30.790 96.490 ;
        RECT 30.980 96.320 31.150 96.490 ;
        RECT 31.340 96.320 31.510 96.490 ;
        RECT 31.700 96.320 31.870 96.490 ;
        RECT 32.060 96.320 32.230 96.490 ;
        RECT 32.420 96.320 32.590 96.490 ;
        RECT 32.780 96.320 32.950 96.490 ;
        RECT 33.140 96.320 33.310 96.490 ;
        RECT 33.500 96.320 33.670 96.490 ;
        RECT 33.860 96.320 34.030 96.490 ;
        RECT 34.220 96.320 34.390 96.490 ;
        RECT 35.630 96.320 35.800 96.490 ;
        RECT 35.990 96.320 36.160 96.490 ;
        RECT 36.350 96.320 36.520 96.490 ;
        RECT 36.710 96.320 36.880 96.490 ;
        RECT 37.070 96.320 37.240 96.490 ;
        RECT 37.430 96.320 37.600 96.490 ;
        RECT 37.790 96.320 37.960 96.490 ;
        RECT 38.150 96.320 38.320 96.490 ;
        RECT 38.510 96.320 38.680 96.490 ;
        RECT 38.870 96.320 39.040 96.490 ;
        RECT 39.230 96.320 39.400 96.490 ;
        RECT 39.590 96.320 39.760 96.490 ;
        RECT 39.950 96.320 40.120 96.490 ;
        RECT 40.310 96.320 40.480 96.490 ;
        RECT 41.720 96.320 41.890 96.490 ;
        RECT 42.080 96.320 42.250 96.490 ;
        RECT 42.440 96.320 42.610 96.490 ;
        RECT 42.800 96.320 42.970 96.490 ;
        RECT 43.160 96.320 43.330 96.490 ;
        RECT 43.520 96.320 43.690 96.490 ;
        RECT 43.880 96.320 44.050 96.490 ;
        RECT 44.240 96.320 44.410 96.490 ;
        RECT 44.600 96.320 44.770 96.490 ;
        RECT 44.960 96.320 45.130 96.490 ;
        RECT 45.320 96.320 45.490 96.490 ;
        RECT 45.680 96.320 45.850 96.490 ;
        RECT 46.040 96.320 46.210 96.490 ;
        RECT 46.400 96.320 46.570 96.490 ;
        RECT 47.810 96.320 47.980 96.490 ;
        RECT 48.170 96.320 48.340 96.490 ;
        RECT 48.530 96.320 48.700 96.490 ;
        RECT 48.890 96.320 49.060 96.490 ;
        RECT 49.250 96.320 49.420 96.490 ;
        RECT 49.610 96.320 49.780 96.490 ;
        RECT 49.970 96.320 50.140 96.490 ;
        RECT 50.330 96.320 50.500 96.490 ;
        RECT 50.690 96.320 50.860 96.490 ;
        RECT 51.050 96.320 51.220 96.490 ;
        RECT 51.410 96.320 51.580 96.490 ;
        RECT 51.770 96.320 51.940 96.490 ;
        RECT 52.130 96.320 52.300 96.490 ;
        RECT 52.490 96.320 52.660 96.490 ;
        RECT 53.900 96.320 54.070 96.490 ;
        RECT 54.260 96.320 54.430 96.490 ;
        RECT 54.620 96.320 54.790 96.490 ;
        RECT 54.980 96.320 55.150 96.490 ;
        RECT 55.340 96.320 55.510 96.490 ;
        RECT 55.700 96.320 55.870 96.490 ;
        RECT 56.060 96.320 56.230 96.490 ;
        RECT 56.420 96.320 56.590 96.490 ;
        RECT 56.780 96.320 56.950 96.490 ;
        RECT 57.140 96.320 57.310 96.490 ;
        RECT 57.500 96.320 57.670 96.490 ;
        RECT 57.860 96.320 58.030 96.490 ;
        RECT 58.220 96.320 58.390 96.490 ;
        RECT 58.580 96.320 58.750 96.490 ;
        RECT 59.990 96.320 60.160 96.490 ;
        RECT 60.350 96.320 60.520 96.490 ;
        RECT 60.710 96.320 60.880 96.490 ;
        RECT 61.070 96.320 61.240 96.490 ;
        RECT 61.430 96.320 61.600 96.490 ;
        RECT 61.790 96.320 61.960 96.490 ;
        RECT 62.150 96.320 62.320 96.490 ;
        RECT 62.510 96.320 62.680 96.490 ;
        RECT 62.870 96.320 63.040 96.490 ;
        RECT 63.230 96.320 63.400 96.490 ;
        RECT 63.590 96.320 63.760 96.490 ;
        RECT 63.950 96.320 64.120 96.490 ;
        RECT 64.310 96.320 64.480 96.490 ;
        RECT 64.670 96.320 64.840 96.490 ;
        RECT 66.080 96.320 66.250 96.490 ;
        RECT 66.440 96.320 66.610 96.490 ;
        RECT 66.800 96.320 66.970 96.490 ;
        RECT 67.160 96.320 67.330 96.490 ;
        RECT 67.520 96.320 67.690 96.490 ;
        RECT 67.880 96.320 68.050 96.490 ;
        RECT 68.240 96.320 68.410 96.490 ;
        RECT 68.600 96.320 68.770 96.490 ;
        RECT 68.960 96.320 69.130 96.490 ;
        RECT 69.320 96.320 69.490 96.490 ;
        RECT 69.680 96.320 69.850 96.490 ;
        RECT 70.040 96.320 70.210 96.490 ;
        RECT 70.400 96.320 70.570 96.490 ;
        RECT 70.760 96.320 70.930 96.490 ;
        RECT 29.105 94.145 29.275 94.315 ;
        RECT 29.105 93.785 29.275 93.955 ;
        RECT 34.655 94.145 34.825 94.315 ;
        RECT 34.655 93.785 34.825 93.955 ;
        RECT 35.195 94.145 35.365 94.315 ;
        RECT 35.195 93.785 35.365 93.955 ;
        RECT 40.745 94.145 40.915 94.315 ;
        RECT 40.745 93.785 40.915 93.955 ;
        RECT 41.285 94.145 41.455 94.315 ;
        RECT 41.285 93.785 41.455 93.955 ;
        RECT 46.835 94.145 47.005 94.315 ;
        RECT 46.835 93.785 47.005 93.955 ;
        RECT 47.375 94.145 47.545 94.315 ;
        RECT 47.375 93.785 47.545 93.955 ;
        RECT 52.925 94.145 53.095 94.315 ;
        RECT 52.925 93.785 53.095 93.955 ;
        RECT 53.465 94.145 53.635 94.315 ;
        RECT 53.465 93.785 53.635 93.955 ;
        RECT 59.015 94.145 59.185 94.315 ;
        RECT 59.015 93.785 59.185 93.955 ;
        RECT 59.555 94.145 59.725 94.315 ;
        RECT 59.555 93.785 59.725 93.955 ;
        RECT 65.105 94.145 65.275 94.315 ;
        RECT 65.105 93.785 65.275 93.955 ;
        RECT 65.645 94.145 65.815 94.315 ;
        RECT 65.645 93.785 65.815 93.955 ;
        RECT 71.195 94.145 71.365 94.315 ;
        RECT 71.195 93.785 71.365 93.955 ;
        RECT 29.540 93.320 29.710 93.490 ;
        RECT 29.900 93.320 30.070 93.490 ;
        RECT 30.260 93.320 30.430 93.490 ;
        RECT 30.620 93.320 30.790 93.490 ;
        RECT 30.980 93.320 31.150 93.490 ;
        RECT 31.340 93.320 31.510 93.490 ;
        RECT 31.700 93.320 31.870 93.490 ;
        RECT 32.060 93.320 32.230 93.490 ;
        RECT 32.420 93.320 32.590 93.490 ;
        RECT 32.780 93.320 32.950 93.490 ;
        RECT 33.140 93.320 33.310 93.490 ;
        RECT 33.500 93.320 33.670 93.490 ;
        RECT 33.860 93.320 34.030 93.490 ;
        RECT 34.220 93.320 34.390 93.490 ;
        RECT 35.630 93.320 35.800 93.490 ;
        RECT 35.990 93.320 36.160 93.490 ;
        RECT 36.350 93.320 36.520 93.490 ;
        RECT 36.710 93.320 36.880 93.490 ;
        RECT 37.070 93.320 37.240 93.490 ;
        RECT 37.430 93.320 37.600 93.490 ;
        RECT 37.790 93.320 37.960 93.490 ;
        RECT 38.150 93.320 38.320 93.490 ;
        RECT 38.510 93.320 38.680 93.490 ;
        RECT 38.870 93.320 39.040 93.490 ;
        RECT 39.230 93.320 39.400 93.490 ;
        RECT 39.590 93.320 39.760 93.490 ;
        RECT 39.950 93.320 40.120 93.490 ;
        RECT 40.310 93.320 40.480 93.490 ;
        RECT 41.720 93.320 41.890 93.490 ;
        RECT 42.080 93.320 42.250 93.490 ;
        RECT 42.440 93.320 42.610 93.490 ;
        RECT 42.800 93.320 42.970 93.490 ;
        RECT 43.160 93.320 43.330 93.490 ;
        RECT 43.520 93.320 43.690 93.490 ;
        RECT 43.880 93.320 44.050 93.490 ;
        RECT 44.240 93.320 44.410 93.490 ;
        RECT 44.600 93.320 44.770 93.490 ;
        RECT 44.960 93.320 45.130 93.490 ;
        RECT 45.320 93.320 45.490 93.490 ;
        RECT 45.680 93.320 45.850 93.490 ;
        RECT 46.040 93.320 46.210 93.490 ;
        RECT 46.400 93.320 46.570 93.490 ;
        RECT 47.810 93.320 47.980 93.490 ;
        RECT 48.170 93.320 48.340 93.490 ;
        RECT 48.530 93.320 48.700 93.490 ;
        RECT 48.890 93.320 49.060 93.490 ;
        RECT 49.250 93.320 49.420 93.490 ;
        RECT 49.610 93.320 49.780 93.490 ;
        RECT 49.970 93.320 50.140 93.490 ;
        RECT 50.330 93.320 50.500 93.490 ;
        RECT 50.690 93.320 50.860 93.490 ;
        RECT 51.050 93.320 51.220 93.490 ;
        RECT 51.410 93.320 51.580 93.490 ;
        RECT 51.770 93.320 51.940 93.490 ;
        RECT 52.130 93.320 52.300 93.490 ;
        RECT 52.490 93.320 52.660 93.490 ;
        RECT 53.900 93.320 54.070 93.490 ;
        RECT 54.260 93.320 54.430 93.490 ;
        RECT 54.620 93.320 54.790 93.490 ;
        RECT 54.980 93.320 55.150 93.490 ;
        RECT 55.340 93.320 55.510 93.490 ;
        RECT 55.700 93.320 55.870 93.490 ;
        RECT 56.060 93.320 56.230 93.490 ;
        RECT 56.420 93.320 56.590 93.490 ;
        RECT 56.780 93.320 56.950 93.490 ;
        RECT 57.140 93.320 57.310 93.490 ;
        RECT 57.500 93.320 57.670 93.490 ;
        RECT 57.860 93.320 58.030 93.490 ;
        RECT 58.220 93.320 58.390 93.490 ;
        RECT 58.580 93.320 58.750 93.490 ;
        RECT 59.990 93.320 60.160 93.490 ;
        RECT 60.350 93.320 60.520 93.490 ;
        RECT 60.710 93.320 60.880 93.490 ;
        RECT 61.070 93.320 61.240 93.490 ;
        RECT 61.430 93.320 61.600 93.490 ;
        RECT 61.790 93.320 61.960 93.490 ;
        RECT 62.150 93.320 62.320 93.490 ;
        RECT 62.510 93.320 62.680 93.490 ;
        RECT 62.870 93.320 63.040 93.490 ;
        RECT 63.230 93.320 63.400 93.490 ;
        RECT 63.590 93.320 63.760 93.490 ;
        RECT 63.950 93.320 64.120 93.490 ;
        RECT 64.310 93.320 64.480 93.490 ;
        RECT 64.670 93.320 64.840 93.490 ;
        RECT 66.080 93.320 66.250 93.490 ;
        RECT 66.440 93.320 66.610 93.490 ;
        RECT 66.800 93.320 66.970 93.490 ;
        RECT 67.160 93.320 67.330 93.490 ;
        RECT 67.520 93.320 67.690 93.490 ;
        RECT 67.880 93.320 68.050 93.490 ;
        RECT 68.240 93.320 68.410 93.490 ;
        RECT 68.600 93.320 68.770 93.490 ;
        RECT 68.960 93.320 69.130 93.490 ;
        RECT 69.320 93.320 69.490 93.490 ;
        RECT 69.680 93.320 69.850 93.490 ;
        RECT 70.040 93.320 70.210 93.490 ;
        RECT 70.400 93.320 70.570 93.490 ;
        RECT 70.760 93.320 70.930 93.490 ;
        RECT 31.830 89.275 32.000 89.445 ;
        RECT 31.830 88.915 32.000 89.085 ;
        RECT 37.470 89.275 37.640 89.445 ;
        RECT 37.470 88.915 37.640 89.085 ;
        RECT 38.010 89.275 38.180 89.445 ;
        RECT 38.010 88.915 38.180 89.085 ;
        RECT 43.650 89.275 43.820 89.445 ;
        RECT 43.650 88.915 43.820 89.085 ;
        RECT 44.190 89.275 44.360 89.445 ;
        RECT 44.190 88.915 44.360 89.085 ;
        RECT 49.830 89.275 50.000 89.445 ;
        RECT 49.830 88.915 50.000 89.085 ;
        RECT 50.370 89.275 50.540 89.445 ;
        RECT 50.370 88.915 50.540 89.085 ;
        RECT 56.010 89.275 56.180 89.445 ;
        RECT 56.010 88.915 56.180 89.085 ;
        RECT 56.550 89.275 56.720 89.445 ;
        RECT 56.550 88.915 56.720 89.085 ;
        RECT 62.190 89.275 62.360 89.445 ;
        RECT 62.190 88.915 62.360 89.085 ;
        RECT 62.730 89.275 62.900 89.445 ;
        RECT 62.730 88.915 62.900 89.085 ;
        RECT 68.370 89.275 68.540 89.445 ;
        RECT 68.370 88.915 68.540 89.085 ;
        RECT 32.310 88.450 32.480 88.620 ;
        RECT 32.670 88.450 32.840 88.620 ;
        RECT 33.030 88.450 33.200 88.620 ;
        RECT 33.390 88.450 33.560 88.620 ;
        RECT 33.750 88.450 33.920 88.620 ;
        RECT 34.110 88.450 34.280 88.620 ;
        RECT 34.470 88.450 34.640 88.620 ;
        RECT 34.830 88.450 35.000 88.620 ;
        RECT 35.190 88.450 35.360 88.620 ;
        RECT 35.550 88.450 35.720 88.620 ;
        RECT 35.910 88.450 36.080 88.620 ;
        RECT 36.270 88.450 36.440 88.620 ;
        RECT 36.630 88.450 36.800 88.620 ;
        RECT 36.990 88.450 37.160 88.620 ;
        RECT 38.490 88.450 38.660 88.620 ;
        RECT 38.850 88.450 39.020 88.620 ;
        RECT 39.210 88.450 39.380 88.620 ;
        RECT 39.570 88.450 39.740 88.620 ;
        RECT 39.930 88.450 40.100 88.620 ;
        RECT 40.290 88.450 40.460 88.620 ;
        RECT 40.650 88.450 40.820 88.620 ;
        RECT 41.010 88.450 41.180 88.620 ;
        RECT 41.370 88.450 41.540 88.620 ;
        RECT 41.730 88.450 41.900 88.620 ;
        RECT 42.090 88.450 42.260 88.620 ;
        RECT 42.450 88.450 42.620 88.620 ;
        RECT 42.810 88.450 42.980 88.620 ;
        RECT 43.170 88.450 43.340 88.620 ;
        RECT 44.670 88.450 44.840 88.620 ;
        RECT 45.030 88.450 45.200 88.620 ;
        RECT 45.390 88.450 45.560 88.620 ;
        RECT 45.750 88.450 45.920 88.620 ;
        RECT 46.110 88.450 46.280 88.620 ;
        RECT 46.470 88.450 46.640 88.620 ;
        RECT 46.830 88.450 47.000 88.620 ;
        RECT 47.190 88.450 47.360 88.620 ;
        RECT 47.550 88.450 47.720 88.620 ;
        RECT 47.910 88.450 48.080 88.620 ;
        RECT 48.270 88.450 48.440 88.620 ;
        RECT 48.630 88.450 48.800 88.620 ;
        RECT 48.990 88.450 49.160 88.620 ;
        RECT 49.350 88.450 49.520 88.620 ;
        RECT 50.850 88.450 51.020 88.620 ;
        RECT 51.210 88.450 51.380 88.620 ;
        RECT 51.570 88.450 51.740 88.620 ;
        RECT 51.930 88.450 52.100 88.620 ;
        RECT 52.290 88.450 52.460 88.620 ;
        RECT 52.650 88.450 52.820 88.620 ;
        RECT 53.010 88.450 53.180 88.620 ;
        RECT 53.370 88.450 53.540 88.620 ;
        RECT 53.730 88.450 53.900 88.620 ;
        RECT 54.090 88.450 54.260 88.620 ;
        RECT 54.450 88.450 54.620 88.620 ;
        RECT 54.810 88.450 54.980 88.620 ;
        RECT 55.170 88.450 55.340 88.620 ;
        RECT 55.530 88.450 55.700 88.620 ;
        RECT 57.030 88.450 57.200 88.620 ;
        RECT 57.390 88.450 57.560 88.620 ;
        RECT 57.750 88.450 57.920 88.620 ;
        RECT 58.110 88.450 58.280 88.620 ;
        RECT 58.470 88.450 58.640 88.620 ;
        RECT 58.830 88.450 59.000 88.620 ;
        RECT 59.190 88.450 59.360 88.620 ;
        RECT 59.550 88.450 59.720 88.620 ;
        RECT 59.910 88.450 60.080 88.620 ;
        RECT 60.270 88.450 60.440 88.620 ;
        RECT 60.630 88.450 60.800 88.620 ;
        RECT 60.990 88.450 61.160 88.620 ;
        RECT 61.350 88.450 61.520 88.620 ;
        RECT 61.710 88.450 61.880 88.620 ;
        RECT 63.210 88.450 63.380 88.620 ;
        RECT 63.570 88.450 63.740 88.620 ;
        RECT 63.930 88.450 64.100 88.620 ;
        RECT 64.290 88.450 64.460 88.620 ;
        RECT 64.650 88.450 64.820 88.620 ;
        RECT 65.010 88.450 65.180 88.620 ;
        RECT 65.370 88.450 65.540 88.620 ;
        RECT 65.730 88.450 65.900 88.620 ;
        RECT 66.090 88.450 66.260 88.620 ;
        RECT 66.450 88.450 66.620 88.620 ;
        RECT 66.810 88.450 66.980 88.620 ;
        RECT 67.170 88.450 67.340 88.620 ;
        RECT 67.530 88.450 67.700 88.620 ;
        RECT 67.890 88.450 68.060 88.620 ;
        RECT 31.830 86.325 32.000 86.495 ;
        RECT 31.830 85.965 32.000 86.135 ;
        RECT 37.470 86.325 37.640 86.495 ;
        RECT 37.470 85.965 37.640 86.135 ;
        RECT 38.010 86.325 38.180 86.495 ;
        RECT 38.010 85.965 38.180 86.135 ;
        RECT 43.650 86.325 43.820 86.495 ;
        RECT 43.650 85.965 43.820 86.135 ;
        RECT 44.190 86.325 44.360 86.495 ;
        RECT 44.190 85.965 44.360 86.135 ;
        RECT 49.830 86.325 50.000 86.495 ;
        RECT 49.830 85.965 50.000 86.135 ;
        RECT 50.370 86.325 50.540 86.495 ;
        RECT 50.370 85.965 50.540 86.135 ;
        RECT 56.010 86.325 56.180 86.495 ;
        RECT 56.010 85.965 56.180 86.135 ;
        RECT 56.550 86.325 56.720 86.495 ;
        RECT 56.550 85.965 56.720 86.135 ;
        RECT 62.190 86.325 62.360 86.495 ;
        RECT 62.190 85.965 62.360 86.135 ;
        RECT 62.730 86.325 62.900 86.495 ;
        RECT 62.730 85.965 62.900 86.135 ;
        RECT 68.370 86.325 68.540 86.495 ;
        RECT 68.370 85.965 68.540 86.135 ;
        RECT 32.310 85.500 32.480 85.670 ;
        RECT 32.670 85.500 32.840 85.670 ;
        RECT 33.030 85.500 33.200 85.670 ;
        RECT 33.390 85.500 33.560 85.670 ;
        RECT 33.750 85.500 33.920 85.670 ;
        RECT 34.110 85.500 34.280 85.670 ;
        RECT 34.470 85.500 34.640 85.670 ;
        RECT 34.830 85.500 35.000 85.670 ;
        RECT 35.190 85.500 35.360 85.670 ;
        RECT 35.550 85.500 35.720 85.670 ;
        RECT 35.910 85.500 36.080 85.670 ;
        RECT 36.270 85.500 36.440 85.670 ;
        RECT 36.630 85.500 36.800 85.670 ;
        RECT 36.990 85.500 37.160 85.670 ;
        RECT 38.490 85.500 38.660 85.670 ;
        RECT 38.850 85.500 39.020 85.670 ;
        RECT 39.210 85.500 39.380 85.670 ;
        RECT 39.570 85.500 39.740 85.670 ;
        RECT 39.930 85.500 40.100 85.670 ;
        RECT 40.290 85.500 40.460 85.670 ;
        RECT 40.650 85.500 40.820 85.670 ;
        RECT 41.010 85.500 41.180 85.670 ;
        RECT 41.370 85.500 41.540 85.670 ;
        RECT 41.730 85.500 41.900 85.670 ;
        RECT 42.090 85.500 42.260 85.670 ;
        RECT 42.450 85.500 42.620 85.670 ;
        RECT 42.810 85.500 42.980 85.670 ;
        RECT 43.170 85.500 43.340 85.670 ;
        RECT 44.670 85.500 44.840 85.670 ;
        RECT 45.030 85.500 45.200 85.670 ;
        RECT 45.390 85.500 45.560 85.670 ;
        RECT 45.750 85.500 45.920 85.670 ;
        RECT 46.110 85.500 46.280 85.670 ;
        RECT 46.470 85.500 46.640 85.670 ;
        RECT 46.830 85.500 47.000 85.670 ;
        RECT 47.190 85.500 47.360 85.670 ;
        RECT 47.550 85.500 47.720 85.670 ;
        RECT 47.910 85.500 48.080 85.670 ;
        RECT 48.270 85.500 48.440 85.670 ;
        RECT 48.630 85.500 48.800 85.670 ;
        RECT 48.990 85.500 49.160 85.670 ;
        RECT 49.350 85.500 49.520 85.670 ;
        RECT 50.850 85.500 51.020 85.670 ;
        RECT 51.210 85.500 51.380 85.670 ;
        RECT 51.570 85.500 51.740 85.670 ;
        RECT 51.930 85.500 52.100 85.670 ;
        RECT 52.290 85.500 52.460 85.670 ;
        RECT 52.650 85.500 52.820 85.670 ;
        RECT 53.010 85.500 53.180 85.670 ;
        RECT 53.370 85.500 53.540 85.670 ;
        RECT 53.730 85.500 53.900 85.670 ;
        RECT 54.090 85.500 54.260 85.670 ;
        RECT 54.450 85.500 54.620 85.670 ;
        RECT 54.810 85.500 54.980 85.670 ;
        RECT 55.170 85.500 55.340 85.670 ;
        RECT 55.530 85.500 55.700 85.670 ;
        RECT 57.030 85.500 57.200 85.670 ;
        RECT 57.390 85.500 57.560 85.670 ;
        RECT 57.750 85.500 57.920 85.670 ;
        RECT 58.110 85.500 58.280 85.670 ;
        RECT 58.470 85.500 58.640 85.670 ;
        RECT 58.830 85.500 59.000 85.670 ;
        RECT 59.190 85.500 59.360 85.670 ;
        RECT 59.550 85.500 59.720 85.670 ;
        RECT 59.910 85.500 60.080 85.670 ;
        RECT 60.270 85.500 60.440 85.670 ;
        RECT 60.630 85.500 60.800 85.670 ;
        RECT 60.990 85.500 61.160 85.670 ;
        RECT 61.350 85.500 61.520 85.670 ;
        RECT 61.710 85.500 61.880 85.670 ;
        RECT 63.210 85.500 63.380 85.670 ;
        RECT 63.570 85.500 63.740 85.670 ;
        RECT 63.930 85.500 64.100 85.670 ;
        RECT 64.290 85.500 64.460 85.670 ;
        RECT 64.650 85.500 64.820 85.670 ;
        RECT 65.010 85.500 65.180 85.670 ;
        RECT 65.370 85.500 65.540 85.670 ;
        RECT 65.730 85.500 65.900 85.670 ;
        RECT 66.090 85.500 66.260 85.670 ;
        RECT 66.450 85.500 66.620 85.670 ;
        RECT 66.810 85.500 66.980 85.670 ;
        RECT 67.170 85.500 67.340 85.670 ;
        RECT 67.530 85.500 67.700 85.670 ;
        RECT 67.890 85.500 68.060 85.670 ;
        RECT 46.220 82.840 46.390 83.010 ;
        RECT 46.580 82.840 46.750 83.010 ;
        RECT 46.940 82.840 47.110 83.010 ;
        RECT 48.560 82.840 48.730 83.010 ;
        RECT 48.920 82.840 49.090 83.010 ;
        RECT 49.280 82.840 49.450 83.010 ;
        RECT 50.900 82.840 51.070 83.010 ;
        RECT 51.260 82.840 51.430 83.010 ;
        RECT 51.620 82.840 51.790 83.010 ;
        RECT 53.240 82.840 53.410 83.010 ;
        RECT 53.600 82.840 53.770 83.010 ;
        RECT 53.960 82.840 54.130 83.010 ;
        RECT 45.680 82.375 45.850 82.545 ;
        RECT 45.680 82.015 45.850 82.185 ;
        RECT 47.480 82.375 47.650 82.545 ;
        RECT 47.480 82.015 47.650 82.185 ;
        RECT 48.020 82.375 48.190 82.545 ;
        RECT 48.020 82.015 48.190 82.185 ;
        RECT 49.820 82.375 49.990 82.545 ;
        RECT 49.820 82.015 49.990 82.185 ;
        RECT 50.360 82.375 50.530 82.545 ;
        RECT 50.360 82.015 50.530 82.185 ;
        RECT 52.160 82.375 52.330 82.545 ;
        RECT 52.160 82.015 52.330 82.185 ;
        RECT 52.700 82.375 52.870 82.545 ;
        RECT 52.700 82.015 52.870 82.185 ;
        RECT 54.500 82.375 54.670 82.545 ;
        RECT 54.500 82.015 54.670 82.185 ;
        RECT 47.225 79.715 47.395 79.885 ;
        RECT 47.585 79.715 47.755 79.885 ;
        RECT 47.945 79.715 48.115 79.885 ;
        RECT 48.305 79.715 48.475 79.885 ;
        RECT 48.665 79.715 48.835 79.885 ;
        RECT 49.025 79.715 49.195 79.885 ;
        RECT 49.385 79.715 49.555 79.885 ;
        RECT 50.815 79.715 50.985 79.885 ;
        RECT 51.175 79.715 51.345 79.885 ;
        RECT 51.535 79.715 51.705 79.885 ;
        RECT 51.895 79.715 52.065 79.885 ;
        RECT 52.255 79.715 52.425 79.885 ;
        RECT 52.615 79.715 52.785 79.885 ;
        RECT 52.975 79.715 53.145 79.885 ;
        RECT 46.780 79.320 46.950 79.490 ;
        RECT 49.830 79.320 50.000 79.490 ;
        RECT 50.370 79.320 50.540 79.490 ;
        RECT 53.420 79.320 53.590 79.490 ;
        RECT 47.225 78.925 47.395 79.095 ;
        RECT 47.585 78.925 47.755 79.095 ;
        RECT 47.945 78.925 48.115 79.095 ;
        RECT 48.305 78.925 48.475 79.095 ;
        RECT 48.665 78.925 48.835 79.095 ;
        RECT 49.025 78.925 49.195 79.095 ;
        RECT 49.385 78.925 49.555 79.095 ;
        RECT 50.815 78.925 50.985 79.095 ;
        RECT 51.175 78.925 51.345 79.095 ;
        RECT 51.535 78.925 51.705 79.095 ;
        RECT 51.895 78.925 52.065 79.095 ;
        RECT 52.255 78.925 52.425 79.095 ;
        RECT 52.615 78.925 52.785 79.095 ;
        RECT 52.975 78.925 53.145 79.095 ;
        RECT 32.540 77.090 32.710 77.260 ;
        RECT 32.900 77.090 33.070 77.260 ;
        RECT 33.260 77.090 33.430 77.260 ;
        RECT 33.620 77.090 33.790 77.260 ;
        RECT 33.980 77.090 34.150 77.260 ;
        RECT 34.340 77.090 34.510 77.260 ;
        RECT 34.700 77.090 34.870 77.260 ;
        RECT 35.060 77.090 35.230 77.260 ;
        RECT 35.420 77.090 35.590 77.260 ;
        RECT 35.780 77.090 35.950 77.260 ;
        RECT 36.140 77.090 36.310 77.260 ;
        RECT 36.500 77.090 36.670 77.260 ;
        RECT 36.860 77.090 37.030 77.260 ;
        RECT 37.220 77.090 37.390 77.260 ;
        RECT 38.630 77.090 38.800 77.260 ;
        RECT 38.990 77.090 39.160 77.260 ;
        RECT 39.350 77.090 39.520 77.260 ;
        RECT 39.710 77.090 39.880 77.260 ;
        RECT 40.070 77.090 40.240 77.260 ;
        RECT 40.430 77.090 40.600 77.260 ;
        RECT 40.790 77.090 40.960 77.260 ;
        RECT 41.150 77.090 41.320 77.260 ;
        RECT 41.510 77.090 41.680 77.260 ;
        RECT 41.870 77.090 42.040 77.260 ;
        RECT 42.230 77.090 42.400 77.260 ;
        RECT 42.590 77.090 42.760 77.260 ;
        RECT 42.950 77.090 43.120 77.260 ;
        RECT 43.310 77.090 43.480 77.260 ;
        RECT 44.720 77.090 44.890 77.260 ;
        RECT 45.080 77.090 45.250 77.260 ;
        RECT 45.440 77.090 45.610 77.260 ;
        RECT 45.800 77.090 45.970 77.260 ;
        RECT 46.160 77.090 46.330 77.260 ;
        RECT 46.520 77.090 46.690 77.260 ;
        RECT 46.880 77.090 47.050 77.260 ;
        RECT 47.240 77.090 47.410 77.260 ;
        RECT 47.600 77.090 47.770 77.260 ;
        RECT 47.960 77.090 48.130 77.260 ;
        RECT 48.320 77.090 48.490 77.260 ;
        RECT 48.680 77.090 48.850 77.260 ;
        RECT 49.040 77.090 49.210 77.260 ;
        RECT 49.400 77.090 49.570 77.260 ;
        RECT 50.810 77.090 50.980 77.260 ;
        RECT 51.170 77.090 51.340 77.260 ;
        RECT 51.530 77.090 51.700 77.260 ;
        RECT 51.890 77.090 52.060 77.260 ;
        RECT 52.250 77.090 52.420 77.260 ;
        RECT 52.610 77.090 52.780 77.260 ;
        RECT 52.970 77.090 53.140 77.260 ;
        RECT 53.330 77.090 53.500 77.260 ;
        RECT 53.690 77.090 53.860 77.260 ;
        RECT 54.050 77.090 54.220 77.260 ;
        RECT 54.410 77.090 54.580 77.260 ;
        RECT 54.770 77.090 54.940 77.260 ;
        RECT 55.130 77.090 55.300 77.260 ;
        RECT 55.490 77.090 55.660 77.260 ;
        RECT 56.900 77.090 57.070 77.260 ;
        RECT 57.260 77.090 57.430 77.260 ;
        RECT 57.620 77.090 57.790 77.260 ;
        RECT 57.980 77.090 58.150 77.260 ;
        RECT 58.340 77.090 58.510 77.260 ;
        RECT 58.700 77.090 58.870 77.260 ;
        RECT 59.060 77.090 59.230 77.260 ;
        RECT 59.420 77.090 59.590 77.260 ;
        RECT 59.780 77.090 59.950 77.260 ;
        RECT 60.140 77.090 60.310 77.260 ;
        RECT 60.500 77.090 60.670 77.260 ;
        RECT 60.860 77.090 61.030 77.260 ;
        RECT 61.220 77.090 61.390 77.260 ;
        RECT 61.580 77.090 61.750 77.260 ;
        RECT 62.990 77.090 63.160 77.260 ;
        RECT 63.350 77.090 63.520 77.260 ;
        RECT 63.710 77.090 63.880 77.260 ;
        RECT 64.070 77.090 64.240 77.260 ;
        RECT 64.430 77.090 64.600 77.260 ;
        RECT 64.790 77.090 64.960 77.260 ;
        RECT 65.150 77.090 65.320 77.260 ;
        RECT 65.510 77.090 65.680 77.260 ;
        RECT 65.870 77.090 66.040 77.260 ;
        RECT 66.230 77.090 66.400 77.260 ;
        RECT 66.590 77.090 66.760 77.260 ;
        RECT 66.950 77.090 67.120 77.260 ;
        RECT 67.310 77.090 67.480 77.260 ;
        RECT 67.670 77.090 67.840 77.260 ;
        RECT 32.105 76.625 32.275 76.795 ;
        RECT 32.105 76.265 32.275 76.435 ;
        RECT 37.655 76.625 37.825 76.795 ;
        RECT 37.655 76.265 37.825 76.435 ;
        RECT 38.195 76.625 38.365 76.795 ;
        RECT 38.195 76.265 38.365 76.435 ;
        RECT 43.745 76.625 43.915 76.795 ;
        RECT 43.745 76.265 43.915 76.435 ;
        RECT 44.285 76.625 44.455 76.795 ;
        RECT 44.285 76.265 44.455 76.435 ;
        RECT 49.835 76.625 50.005 76.795 ;
        RECT 49.835 76.265 50.005 76.435 ;
        RECT 50.375 76.625 50.545 76.795 ;
        RECT 50.375 76.265 50.545 76.435 ;
        RECT 55.925 76.625 56.095 76.795 ;
        RECT 55.925 76.265 56.095 76.435 ;
        RECT 56.465 76.625 56.635 76.795 ;
        RECT 56.465 76.265 56.635 76.435 ;
        RECT 62.015 76.625 62.185 76.795 ;
        RECT 62.015 76.265 62.185 76.435 ;
        RECT 62.555 76.625 62.725 76.795 ;
        RECT 62.555 76.265 62.725 76.435 ;
        RECT 68.105 76.625 68.275 76.795 ;
        RECT 68.105 76.265 68.275 76.435 ;
        RECT 32.540 75.800 32.710 75.970 ;
        RECT 32.900 75.800 33.070 75.970 ;
        RECT 33.260 75.800 33.430 75.970 ;
        RECT 33.620 75.800 33.790 75.970 ;
        RECT 33.980 75.800 34.150 75.970 ;
        RECT 34.340 75.800 34.510 75.970 ;
        RECT 34.700 75.800 34.870 75.970 ;
        RECT 35.060 75.800 35.230 75.970 ;
        RECT 35.420 75.800 35.590 75.970 ;
        RECT 35.780 75.800 35.950 75.970 ;
        RECT 36.140 75.800 36.310 75.970 ;
        RECT 36.500 75.800 36.670 75.970 ;
        RECT 36.860 75.800 37.030 75.970 ;
        RECT 37.220 75.800 37.390 75.970 ;
        RECT 38.630 75.800 38.800 75.970 ;
        RECT 38.990 75.800 39.160 75.970 ;
        RECT 39.350 75.800 39.520 75.970 ;
        RECT 39.710 75.800 39.880 75.970 ;
        RECT 40.070 75.800 40.240 75.970 ;
        RECT 40.430 75.800 40.600 75.970 ;
        RECT 40.790 75.800 40.960 75.970 ;
        RECT 41.150 75.800 41.320 75.970 ;
        RECT 41.510 75.800 41.680 75.970 ;
        RECT 41.870 75.800 42.040 75.970 ;
        RECT 42.230 75.800 42.400 75.970 ;
        RECT 42.590 75.800 42.760 75.970 ;
        RECT 42.950 75.800 43.120 75.970 ;
        RECT 43.310 75.800 43.480 75.970 ;
        RECT 44.720 75.800 44.890 75.970 ;
        RECT 45.080 75.800 45.250 75.970 ;
        RECT 45.440 75.800 45.610 75.970 ;
        RECT 45.800 75.800 45.970 75.970 ;
        RECT 46.160 75.800 46.330 75.970 ;
        RECT 46.520 75.800 46.690 75.970 ;
        RECT 46.880 75.800 47.050 75.970 ;
        RECT 47.240 75.800 47.410 75.970 ;
        RECT 47.600 75.800 47.770 75.970 ;
        RECT 47.960 75.800 48.130 75.970 ;
        RECT 48.320 75.800 48.490 75.970 ;
        RECT 48.680 75.800 48.850 75.970 ;
        RECT 49.040 75.800 49.210 75.970 ;
        RECT 49.400 75.800 49.570 75.970 ;
        RECT 50.810 75.800 50.980 75.970 ;
        RECT 51.170 75.800 51.340 75.970 ;
        RECT 51.530 75.800 51.700 75.970 ;
        RECT 51.890 75.800 52.060 75.970 ;
        RECT 52.250 75.800 52.420 75.970 ;
        RECT 52.610 75.800 52.780 75.970 ;
        RECT 52.970 75.800 53.140 75.970 ;
        RECT 53.330 75.800 53.500 75.970 ;
        RECT 53.690 75.800 53.860 75.970 ;
        RECT 54.050 75.800 54.220 75.970 ;
        RECT 54.410 75.800 54.580 75.970 ;
        RECT 54.770 75.800 54.940 75.970 ;
        RECT 55.130 75.800 55.300 75.970 ;
        RECT 55.490 75.800 55.660 75.970 ;
        RECT 56.900 75.800 57.070 75.970 ;
        RECT 57.260 75.800 57.430 75.970 ;
        RECT 57.620 75.800 57.790 75.970 ;
        RECT 57.980 75.800 58.150 75.970 ;
        RECT 58.340 75.800 58.510 75.970 ;
        RECT 58.700 75.800 58.870 75.970 ;
        RECT 59.060 75.800 59.230 75.970 ;
        RECT 59.420 75.800 59.590 75.970 ;
        RECT 59.780 75.800 59.950 75.970 ;
        RECT 60.140 75.800 60.310 75.970 ;
        RECT 60.500 75.800 60.670 75.970 ;
        RECT 60.860 75.800 61.030 75.970 ;
        RECT 61.220 75.800 61.390 75.970 ;
        RECT 61.580 75.800 61.750 75.970 ;
        RECT 62.990 75.800 63.160 75.970 ;
        RECT 63.350 75.800 63.520 75.970 ;
        RECT 63.710 75.800 63.880 75.970 ;
        RECT 64.070 75.800 64.240 75.970 ;
        RECT 64.430 75.800 64.600 75.970 ;
        RECT 64.790 75.800 64.960 75.970 ;
        RECT 65.150 75.800 65.320 75.970 ;
        RECT 65.510 75.800 65.680 75.970 ;
        RECT 65.870 75.800 66.040 75.970 ;
        RECT 66.230 75.800 66.400 75.970 ;
        RECT 66.590 75.800 66.760 75.970 ;
        RECT 66.950 75.800 67.120 75.970 ;
        RECT 67.310 75.800 67.480 75.970 ;
        RECT 67.670 75.800 67.840 75.970 ;
        RECT 36.055 71.500 41.625 73.470 ;
        RECT 43.655 71.500 49.225 73.470 ;
        RECT 51.205 71.530 56.775 73.500 ;
        RECT 58.755 71.530 64.325 73.500 ;
      LAYER met1 ;
        RECT 28.575 137.120 28.805 137.230 ;
        RECT 34.215 137.170 34.445 137.230 ;
        RECT 34.755 137.170 34.985 137.230 ;
        RECT 34.215 137.120 34.985 137.170 ;
        RECT 40.395 137.170 40.625 137.230 ;
        RECT 40.935 137.170 41.165 137.230 ;
        RECT 46.575 137.170 46.805 137.230 ;
        RECT 47.115 137.170 47.345 137.230 ;
        RECT 40.395 137.120 41.165 137.170 ;
        RECT 46.565 137.120 47.345 137.170 ;
        RECT 52.755 137.170 52.985 137.230 ;
        RECT 53.295 137.170 53.525 137.230 ;
        RECT 52.755 137.120 53.525 137.170 ;
        RECT 58.935 137.170 59.165 137.230 ;
        RECT 59.475 137.170 59.705 137.230 ;
        RECT 65.115 137.170 65.345 137.230 ;
        RECT 65.655 137.170 65.885 137.230 ;
        RECT 58.935 137.120 59.715 137.170 ;
        RECT 65.115 137.120 65.885 137.170 ;
        RECT 71.295 137.120 71.525 137.230 ;
        RECT 28.575 136.920 71.525 137.120 ;
        RECT 28.515 136.420 71.565 136.920 ;
        RECT 30.615 136.220 31.115 136.420 ;
        RECT 31.465 136.220 31.965 136.420 ;
        RECT 43.215 136.220 43.715 136.420 ;
        RECT 44.065 136.220 44.565 136.420 ;
        RECT 55.665 136.220 56.165 136.420 ;
        RECT 56.515 136.220 57.015 136.420 ;
        RECT 67.915 136.220 68.415 136.420 ;
        RECT 68.765 136.220 69.265 136.420 ;
        RECT 28.575 134.420 28.805 134.530 ;
        RECT 34.215 134.470 34.445 134.530 ;
        RECT 34.755 134.470 34.985 134.530 ;
        RECT 34.215 134.420 34.985 134.470 ;
        RECT 40.395 134.470 40.625 134.530 ;
        RECT 40.935 134.470 41.165 134.530 ;
        RECT 46.575 134.470 46.805 134.530 ;
        RECT 47.115 134.470 47.345 134.530 ;
        RECT 40.395 134.420 41.165 134.470 ;
        RECT 46.565 134.420 47.345 134.470 ;
        RECT 52.755 134.470 52.985 134.530 ;
        RECT 53.295 134.470 53.525 134.530 ;
        RECT 52.755 134.420 53.525 134.470 ;
        RECT 58.935 134.470 59.165 134.530 ;
        RECT 59.475 134.470 59.705 134.530 ;
        RECT 65.115 134.470 65.345 134.530 ;
        RECT 65.655 134.470 65.885 134.530 ;
        RECT 58.935 134.420 59.715 134.470 ;
        RECT 65.115 134.420 65.885 134.470 ;
        RECT 71.295 134.420 71.525 134.530 ;
        RECT 28.575 134.220 71.525 134.420 ;
        RECT 28.565 134.070 71.525 134.220 ;
        RECT 28.565 133.720 71.465 134.070 ;
        RECT 30.615 133.520 31.115 133.720 ;
        RECT 31.465 133.520 31.965 133.720 ;
        RECT 43.215 133.520 43.715 133.720 ;
        RECT 44.065 133.520 44.565 133.720 ;
        RECT 55.665 133.520 56.165 133.720 ;
        RECT 56.515 133.520 57.015 133.720 ;
        RECT 67.915 133.470 68.415 133.720 ;
        RECT 68.765 133.470 69.265 133.720 ;
        RECT 28.575 131.720 28.805 131.830 ;
        RECT 34.215 131.770 34.445 131.830 ;
        RECT 34.755 131.770 34.985 131.830 ;
        RECT 34.215 131.720 34.985 131.770 ;
        RECT 40.395 131.770 40.625 131.830 ;
        RECT 40.935 131.770 41.165 131.830 ;
        RECT 46.575 131.770 46.805 131.830 ;
        RECT 47.115 131.770 47.345 131.830 ;
        RECT 40.395 131.720 41.165 131.770 ;
        RECT 46.565 131.720 47.345 131.770 ;
        RECT 52.755 131.770 52.985 131.830 ;
        RECT 53.295 131.770 53.525 131.830 ;
        RECT 52.755 131.720 53.525 131.770 ;
        RECT 58.935 131.770 59.165 131.830 ;
        RECT 59.475 131.770 59.705 131.830 ;
        RECT 65.115 131.770 65.345 131.830 ;
        RECT 65.655 131.770 65.885 131.830 ;
        RECT 58.935 131.720 59.715 131.770 ;
        RECT 65.115 131.720 65.885 131.770 ;
        RECT 71.295 131.720 71.525 131.830 ;
        RECT 28.575 131.370 71.525 131.720 ;
        RECT 28.615 131.020 71.515 131.370 ;
        RECT 30.615 130.820 31.115 131.020 ;
        RECT 31.465 130.820 31.965 131.020 ;
        RECT 43.215 130.820 43.715 131.020 ;
        RECT 44.065 130.820 44.565 131.020 ;
        RECT 55.665 130.770 56.165 131.020 ;
        RECT 56.515 130.770 57.015 131.020 ;
        RECT 67.915 130.820 68.415 131.020 ;
        RECT 68.765 130.820 69.265 131.020 ;
        RECT 28.575 129.020 28.805 129.130 ;
        RECT 34.215 129.070 34.445 129.130 ;
        RECT 34.755 129.070 34.985 129.130 ;
        RECT 34.215 129.020 34.985 129.070 ;
        RECT 40.395 129.070 40.625 129.130 ;
        RECT 40.935 129.070 41.165 129.130 ;
        RECT 46.575 129.070 46.805 129.130 ;
        RECT 47.115 129.070 47.345 129.130 ;
        RECT 40.395 129.020 41.165 129.070 ;
        RECT 46.565 129.020 47.345 129.070 ;
        RECT 52.755 129.070 52.985 129.130 ;
        RECT 53.295 129.070 53.525 129.130 ;
        RECT 58.935 129.070 59.165 129.130 ;
        RECT 59.475 129.070 59.705 129.130 ;
        RECT 52.755 129.020 53.525 129.070 ;
        RECT 58.915 129.020 59.705 129.070 ;
        RECT 65.115 129.070 65.345 129.130 ;
        RECT 65.655 129.070 65.885 129.130 ;
        RECT 65.115 129.020 65.885 129.070 ;
        RECT 71.295 129.020 71.525 129.130 ;
        RECT 28.575 128.770 71.525 129.020 ;
        RECT 28.575 128.670 28.805 128.770 ;
        RECT 34.215 128.720 34.985 128.770 ;
        RECT 34.215 128.670 34.445 128.720 ;
        RECT 34.755 128.670 34.985 128.720 ;
        RECT 40.395 128.720 41.165 128.770 ;
        RECT 46.565 128.720 47.345 128.770 ;
        RECT 40.395 128.670 40.625 128.720 ;
        RECT 40.935 128.670 41.165 128.720 ;
        RECT 46.575 128.670 46.805 128.720 ;
        RECT 47.115 128.670 47.345 128.720 ;
        RECT 52.755 128.720 53.525 128.770 ;
        RECT 58.915 128.720 59.705 128.770 ;
        RECT 52.755 128.670 52.985 128.720 ;
        RECT 53.295 128.670 53.525 128.720 ;
        RECT 58.935 128.670 59.165 128.720 ;
        RECT 59.475 128.670 59.705 128.720 ;
        RECT 65.115 128.720 65.885 128.770 ;
        RECT 65.115 128.670 65.345 128.720 ;
        RECT 65.655 128.670 65.885 128.720 ;
        RECT 71.295 128.670 71.525 128.770 ;
        RECT 29.010 128.520 34.010 128.620 ;
        RECT 35.190 128.520 40.190 128.620 ;
        RECT 41.370 128.520 46.370 128.620 ;
        RECT 47.550 128.520 52.550 128.620 ;
        RECT 53.730 128.520 58.730 128.620 ;
        RECT 59.910 128.520 64.910 128.620 ;
        RECT 66.090 128.520 71.090 128.620 ;
        RECT 28.965 128.320 71.165 128.520 ;
        RECT 30.615 128.120 31.115 128.320 ;
        RECT 31.465 128.120 31.965 128.320 ;
        RECT 38.965 128.020 40.115 128.320 ;
        RECT 43.165 128.120 43.665 128.320 ;
        RECT 44.015 128.120 44.515 128.320 ;
        RECT 51.015 128.120 52.165 128.320 ;
        RECT 55.615 128.120 56.115 128.320 ;
        RECT 56.465 128.120 56.965 128.320 ;
        RECT 63.315 128.020 64.465 128.320 ;
        RECT 68.065 128.120 68.565 128.320 ;
        RECT 68.915 128.120 69.415 128.320 ;
        RECT 28.575 126.120 28.805 126.230 ;
        RECT 34.215 126.170 34.445 126.230 ;
        RECT 34.755 126.170 34.985 126.230 ;
        RECT 34.215 126.120 34.985 126.170 ;
        RECT 40.395 126.170 40.625 126.230 ;
        RECT 40.935 126.170 41.165 126.230 ;
        RECT 40.395 126.120 41.165 126.170 ;
        RECT 46.575 126.170 46.805 126.230 ;
        RECT 47.115 126.170 47.345 126.230 ;
        RECT 52.755 126.170 52.985 126.230 ;
        RECT 53.295 126.170 53.525 126.230 ;
        RECT 58.935 126.170 59.165 126.230 ;
        RECT 59.475 126.170 59.705 126.230 ;
        RECT 46.575 126.120 47.365 126.170 ;
        RECT 52.755 126.120 53.525 126.170 ;
        RECT 58.915 126.120 59.705 126.170 ;
        RECT 65.115 126.170 65.345 126.230 ;
        RECT 65.655 126.170 65.885 126.230 ;
        RECT 65.115 126.120 65.885 126.170 ;
        RECT 71.295 126.120 71.525 126.230 ;
        RECT 28.575 125.870 71.525 126.120 ;
        RECT 28.575 125.770 28.805 125.870 ;
        RECT 34.215 125.820 34.985 125.870 ;
        RECT 34.215 125.770 34.445 125.820 ;
        RECT 34.755 125.770 34.985 125.820 ;
        RECT 40.395 125.820 41.165 125.870 ;
        RECT 40.395 125.770 40.625 125.820 ;
        RECT 40.935 125.770 41.165 125.820 ;
        RECT 46.575 125.820 47.365 125.870 ;
        RECT 52.755 125.820 53.525 125.870 ;
        RECT 58.915 125.820 59.705 125.870 ;
        RECT 46.575 125.770 46.805 125.820 ;
        RECT 47.115 125.770 47.345 125.820 ;
        RECT 52.755 125.770 52.985 125.820 ;
        RECT 53.295 125.770 53.525 125.820 ;
        RECT 58.935 125.770 59.165 125.820 ;
        RECT 59.475 125.770 59.705 125.820 ;
        RECT 65.115 125.820 65.885 125.870 ;
        RECT 65.115 125.770 65.345 125.820 ;
        RECT 65.655 125.770 65.885 125.820 ;
        RECT 71.295 125.770 71.525 125.870 ;
        RECT 29.010 125.620 34.010 125.720 ;
        RECT 35.190 125.620 40.190 125.720 ;
        RECT 41.370 125.620 46.370 125.720 ;
        RECT 47.550 125.620 52.550 125.720 ;
        RECT 53.730 125.620 58.730 125.720 ;
        RECT 59.910 125.620 64.910 125.720 ;
        RECT 66.090 125.620 71.090 125.720 ;
        RECT 28.965 125.420 71.165 125.620 ;
        RECT 30.615 125.220 31.115 125.420 ;
        RECT 31.465 125.220 31.965 125.420 ;
        RECT 38.965 125.070 40.115 125.420 ;
        RECT 43.165 125.220 43.665 125.420 ;
        RECT 44.015 125.220 44.515 125.420 ;
        RECT 51.015 125.120 52.165 125.420 ;
        RECT 55.615 125.170 56.115 125.420 ;
        RECT 56.465 125.170 56.965 125.420 ;
        RECT 63.315 125.120 64.465 125.420 ;
        RECT 68.065 125.220 68.565 125.420 ;
        RECT 68.915 125.220 69.415 125.420 ;
        RECT 0.215 123.395 2.365 124.820 ;
        RECT 97.715 123.395 99.865 125.670 ;
        RECT 0.215 117.705 2.885 123.395 ;
        RECT 12.995 122.870 15.040 123.395 ;
        RECT 28.575 123.220 28.805 123.330 ;
        RECT 34.215 123.270 34.445 123.330 ;
        RECT 34.755 123.270 34.985 123.330 ;
        RECT 34.215 123.220 34.985 123.270 ;
        RECT 40.395 123.270 40.625 123.330 ;
        RECT 40.935 123.270 41.165 123.330 ;
        RECT 46.575 123.270 46.805 123.330 ;
        RECT 47.115 123.270 47.345 123.330 ;
        RECT 40.395 123.220 41.165 123.270 ;
        RECT 46.565 123.220 47.345 123.270 ;
        RECT 52.755 123.270 52.985 123.330 ;
        RECT 53.295 123.270 53.525 123.330 ;
        RECT 58.935 123.270 59.165 123.330 ;
        RECT 59.475 123.270 59.705 123.330 ;
        RECT 52.755 123.220 53.525 123.270 ;
        RECT 58.915 123.220 59.705 123.270 ;
        RECT 65.115 123.270 65.345 123.330 ;
        RECT 65.655 123.270 65.885 123.330 ;
        RECT 65.115 123.220 65.885 123.270 ;
        RECT 71.295 123.220 71.525 123.330 ;
        RECT 28.575 122.970 71.525 123.220 ;
        RECT 28.575 122.870 28.805 122.970 ;
        RECT 34.215 122.920 34.985 122.970 ;
        RECT 34.215 122.870 34.445 122.920 ;
        RECT 34.755 122.870 34.985 122.920 ;
        RECT 40.395 122.920 41.165 122.970 ;
        RECT 46.565 122.920 47.345 122.970 ;
        RECT 40.395 122.870 40.625 122.920 ;
        RECT 40.935 122.870 41.165 122.920 ;
        RECT 46.575 122.870 46.805 122.920 ;
        RECT 47.115 122.870 47.345 122.920 ;
        RECT 52.755 122.920 53.525 122.970 ;
        RECT 58.915 122.920 59.705 122.970 ;
        RECT 52.755 122.870 52.985 122.920 ;
        RECT 53.295 122.870 53.525 122.920 ;
        RECT 58.935 122.870 59.165 122.920 ;
        RECT 59.475 122.870 59.705 122.920 ;
        RECT 65.115 122.920 65.885 122.970 ;
        RECT 65.115 122.870 65.345 122.920 ;
        RECT 65.655 122.870 65.885 122.920 ;
        RECT 71.295 122.870 71.525 122.970 ;
        RECT 86.140 122.870 88.185 123.395 ;
        RECT 12.365 120.670 15.040 122.870 ;
        RECT 29.010 122.670 34.010 122.820 ;
        RECT 35.190 122.670 40.190 122.820 ;
        RECT 41.370 122.670 46.370 122.820 ;
        RECT 47.550 122.670 52.550 122.820 ;
        RECT 53.730 122.670 58.730 122.820 ;
        RECT 59.910 122.670 64.910 122.820 ;
        RECT 66.090 122.670 71.090 122.820 ;
        RECT 28.965 122.470 71.165 122.670 ;
        RECT 30.515 122.170 31.015 122.470 ;
        RECT 31.565 122.170 32.065 122.470 ;
        RECT 38.965 122.220 40.115 122.470 ;
        RECT 43.165 122.320 43.665 122.470 ;
        RECT 44.015 122.320 44.515 122.470 ;
        RECT 51.015 122.220 52.165 122.470 ;
        RECT 55.615 122.320 56.115 122.470 ;
        RECT 56.465 122.320 56.965 122.470 ;
        RECT 63.315 122.220 64.465 122.470 ;
        RECT 68.065 122.320 68.565 122.470 ;
        RECT 68.915 122.320 69.415 122.470 ;
        RECT 85.515 120.670 88.185 122.870 ;
        RECT 12.365 120.630 19.565 120.670 ;
        RECT 80.665 120.630 88.185 120.670 ;
        RECT 12.365 120.520 19.605 120.630 ;
        RECT 25.015 120.570 25.245 120.630 ;
        RECT 25.555 120.570 25.785 120.630 ;
        RECT 25.015 120.520 25.785 120.570 ;
        RECT 31.195 120.570 31.425 120.630 ;
        RECT 31.735 120.570 31.965 120.630 ;
        RECT 37.375 120.570 37.605 120.630 ;
        RECT 37.915 120.570 38.145 120.630 ;
        RECT 31.195 120.520 31.965 120.570 ;
        RECT 37.365 120.520 38.145 120.570 ;
        RECT 43.555 120.570 43.785 120.630 ;
        RECT 44.095 120.570 44.325 120.630 ;
        RECT 43.555 120.520 44.325 120.570 ;
        RECT 49.735 120.570 49.965 120.630 ;
        RECT 50.275 120.570 50.505 120.630 ;
        RECT 55.915 120.570 56.145 120.630 ;
        RECT 56.455 120.570 56.685 120.630 ;
        RECT 49.735 120.520 50.515 120.570 ;
        RECT 55.915 120.520 56.685 120.570 ;
        RECT 62.095 120.570 62.325 120.630 ;
        RECT 62.635 120.570 62.865 120.630 ;
        RECT 68.275 120.570 68.505 120.630 ;
        RECT 68.815 120.570 69.045 120.630 ;
        RECT 62.095 120.520 62.865 120.570 ;
        RECT 68.265 120.520 69.045 120.570 ;
        RECT 74.455 120.570 74.685 120.630 ;
        RECT 74.995 120.570 75.225 120.630 ;
        RECT 74.455 120.520 75.225 120.570 ;
        RECT 80.635 120.520 88.185 120.630 ;
        RECT 12.365 120.320 88.185 120.520 ;
        RECT 12.365 120.170 19.605 120.320 ;
        RECT 25.015 120.220 25.785 120.320 ;
        RECT 25.015 120.170 25.245 120.220 ;
        RECT 25.555 120.170 25.785 120.220 ;
        RECT 31.195 120.220 31.965 120.320 ;
        RECT 37.365 120.220 38.145 120.320 ;
        RECT 31.195 120.170 31.425 120.220 ;
        RECT 31.735 120.170 31.965 120.220 ;
        RECT 37.375 120.170 37.605 120.220 ;
        RECT 37.915 120.170 38.145 120.220 ;
        RECT 43.555 120.220 44.325 120.320 ;
        RECT 43.555 120.170 43.785 120.220 ;
        RECT 44.095 120.170 44.325 120.220 ;
        RECT 49.735 120.220 50.515 120.320 ;
        RECT 55.915 120.220 56.685 120.320 ;
        RECT 49.735 120.170 49.965 120.220 ;
        RECT 50.275 120.170 50.505 120.220 ;
        RECT 55.915 120.170 56.145 120.220 ;
        RECT 56.455 120.170 56.685 120.220 ;
        RECT 62.095 120.220 62.865 120.320 ;
        RECT 68.265 120.220 69.045 120.320 ;
        RECT 62.095 120.170 62.325 120.220 ;
        RECT 62.635 120.170 62.865 120.220 ;
        RECT 68.275 120.170 68.505 120.220 ;
        RECT 68.815 120.170 69.045 120.220 ;
        RECT 74.455 120.220 75.225 120.320 ;
        RECT 74.455 120.170 74.685 120.220 ;
        RECT 74.995 120.170 75.225 120.220 ;
        RECT 80.635 120.170 88.185 120.320 ;
        RECT 12.365 117.970 15.040 120.170 ;
        RECT 12.365 117.930 19.565 117.970 ;
        RECT 12.365 117.820 19.605 117.930 ;
        RECT 25.015 117.920 25.245 117.930 ;
        RECT 25.555 117.920 25.785 117.930 ;
        RECT 25.015 117.820 25.785 117.920 ;
        RECT 31.195 117.870 31.425 117.930 ;
        RECT 31.735 117.870 31.965 117.930 ;
        RECT 37.375 117.870 37.605 117.930 ;
        RECT 37.915 117.870 38.145 117.930 ;
        RECT 31.195 117.820 31.965 117.870 ;
        RECT 37.365 117.820 38.145 117.870 ;
        RECT 43.555 117.870 43.785 117.930 ;
        RECT 44.095 117.870 44.325 117.930 ;
        RECT 43.555 117.820 44.325 117.870 ;
        RECT 49.735 117.870 49.965 117.930 ;
        RECT 50.275 117.870 50.505 117.930 ;
        RECT 55.915 117.870 56.145 117.930 ;
        RECT 56.455 117.870 56.685 117.930 ;
        RECT 49.735 117.820 50.515 117.870 ;
        RECT 55.915 117.820 56.685 117.870 ;
        RECT 62.095 117.870 62.325 117.930 ;
        RECT 62.635 117.870 62.865 117.930 ;
        RECT 68.275 117.870 68.505 117.930 ;
        RECT 68.815 117.870 69.045 117.930 ;
        RECT 62.095 117.820 62.865 117.870 ;
        RECT 68.265 117.820 69.045 117.870 ;
        RECT 74.455 117.870 74.685 117.930 ;
        RECT 74.995 117.870 75.225 117.930 ;
        RECT 74.455 117.820 75.225 117.870 ;
        RECT 80.635 117.920 80.865 117.930 ;
        RECT 85.515 117.920 88.185 120.170 ;
        RECT 80.635 117.820 88.185 117.920 ;
        RECT 12.365 117.705 88.185 117.820 ;
        RECT 97.715 117.705 100.340 123.395 ;
        RECT 0.215 116.045 2.365 117.705 ;
        RECT 12.365 117.620 87.665 117.705 ;
        RECT 12.365 117.470 19.605 117.620 ;
        RECT 25.015 117.570 25.785 117.620 ;
        RECT 25.015 117.470 25.245 117.570 ;
        RECT 25.555 117.470 25.785 117.570 ;
        RECT 31.195 117.520 31.965 117.620 ;
        RECT 37.365 117.520 38.145 117.620 ;
        RECT 31.195 117.470 31.425 117.520 ;
        RECT 31.735 117.470 31.965 117.520 ;
        RECT 37.375 117.470 37.605 117.520 ;
        RECT 37.915 117.470 38.145 117.520 ;
        RECT 43.555 117.520 44.325 117.620 ;
        RECT 43.555 117.470 43.785 117.520 ;
        RECT 44.095 117.470 44.325 117.520 ;
        RECT 49.735 117.520 50.515 117.620 ;
        RECT 55.915 117.520 56.685 117.620 ;
        RECT 49.735 117.470 49.965 117.520 ;
        RECT 50.275 117.470 50.505 117.520 ;
        RECT 55.915 117.470 56.145 117.520 ;
        RECT 56.455 117.470 56.685 117.520 ;
        RECT 62.095 117.520 62.865 117.620 ;
        RECT 68.265 117.520 69.045 117.620 ;
        RECT 62.095 117.470 62.325 117.520 ;
        RECT 62.635 117.470 62.865 117.520 ;
        RECT 68.275 117.470 68.505 117.520 ;
        RECT 68.815 117.470 69.045 117.520 ;
        RECT 74.455 117.520 75.225 117.620 ;
        RECT 74.455 117.470 74.685 117.520 ;
        RECT 74.995 117.470 75.225 117.520 ;
        RECT 80.635 117.470 87.665 117.620 ;
        RECT 12.365 117.420 19.565 117.470 ;
        RECT 80.665 117.420 87.665 117.470 ;
        RECT 12.365 116.045 14.515 117.420 ;
        RECT 85.515 116.045 87.665 117.420 ;
        RECT 97.715 116.045 99.865 117.705 ;
        RECT 0.215 110.520 2.885 116.045 ;
        RECT 0.840 110.355 2.885 110.520 ;
        RECT 12.365 115.270 15.040 116.045 ;
        RECT 85.515 115.270 88.185 116.045 ;
        RECT 12.365 115.120 19.665 115.270 ;
        RECT 80.665 115.230 88.185 115.270 ;
        RECT 25.015 115.170 25.245 115.230 ;
        RECT 25.555 115.170 25.785 115.230 ;
        RECT 25.015 115.120 25.785 115.170 ;
        RECT 31.195 115.170 31.425 115.230 ;
        RECT 31.735 115.170 31.965 115.230 ;
        RECT 37.375 115.170 37.605 115.230 ;
        RECT 37.915 115.170 38.145 115.230 ;
        RECT 31.195 115.120 31.965 115.170 ;
        RECT 37.365 115.120 38.145 115.170 ;
        RECT 43.555 115.170 43.785 115.230 ;
        RECT 44.095 115.170 44.325 115.230 ;
        RECT 43.555 115.120 44.325 115.170 ;
        RECT 49.735 115.170 49.965 115.230 ;
        RECT 50.275 115.170 50.505 115.230 ;
        RECT 55.915 115.170 56.145 115.230 ;
        RECT 56.455 115.170 56.685 115.230 ;
        RECT 49.735 115.120 50.515 115.170 ;
        RECT 55.915 115.120 56.685 115.170 ;
        RECT 62.095 115.170 62.325 115.230 ;
        RECT 62.635 115.170 62.865 115.230 ;
        RECT 68.275 115.170 68.505 115.230 ;
        RECT 68.815 115.170 69.045 115.230 ;
        RECT 62.095 115.120 62.865 115.170 ;
        RECT 68.265 115.120 69.045 115.170 ;
        RECT 74.455 115.170 74.685 115.230 ;
        RECT 74.995 115.170 75.225 115.230 ;
        RECT 74.455 115.120 75.225 115.170 ;
        RECT 80.635 115.120 88.185 115.230 ;
        RECT 12.365 114.920 88.185 115.120 ;
        RECT 12.365 114.720 19.665 114.920 ;
        RECT 25.015 114.820 25.785 114.920 ;
        RECT 25.015 114.770 25.245 114.820 ;
        RECT 25.555 114.770 25.785 114.820 ;
        RECT 31.195 114.820 31.965 114.920 ;
        RECT 37.365 114.820 38.145 114.920 ;
        RECT 31.195 114.770 31.425 114.820 ;
        RECT 31.735 114.770 31.965 114.820 ;
        RECT 37.375 114.770 37.605 114.820 ;
        RECT 37.915 114.770 38.145 114.820 ;
        RECT 43.555 114.820 44.325 114.920 ;
        RECT 43.555 114.770 43.785 114.820 ;
        RECT 44.095 114.770 44.325 114.820 ;
        RECT 49.735 114.820 50.515 114.920 ;
        RECT 55.915 114.820 56.685 114.920 ;
        RECT 49.735 114.770 49.965 114.820 ;
        RECT 50.275 114.770 50.505 114.820 ;
        RECT 55.915 114.770 56.145 114.820 ;
        RECT 56.455 114.770 56.685 114.820 ;
        RECT 62.095 114.820 62.865 114.920 ;
        RECT 68.265 114.820 69.045 114.920 ;
        RECT 62.095 114.770 62.325 114.820 ;
        RECT 62.635 114.770 62.865 114.820 ;
        RECT 68.275 114.770 68.505 114.820 ;
        RECT 68.815 114.770 69.045 114.820 ;
        RECT 74.455 114.820 75.225 114.920 ;
        RECT 74.455 114.770 74.685 114.820 ;
        RECT 74.995 114.770 75.225 114.820 ;
        RECT 80.635 114.770 88.185 114.920 ;
        RECT 12.365 112.570 15.040 114.720 ;
        RECT 85.515 112.570 88.185 114.770 ;
        RECT 12.365 112.420 19.615 112.570 ;
        RECT 80.665 112.530 88.185 112.570 ;
        RECT 25.015 112.470 25.245 112.530 ;
        RECT 25.555 112.470 25.785 112.530 ;
        RECT 25.015 112.420 25.785 112.470 ;
        RECT 31.195 112.470 31.425 112.530 ;
        RECT 31.735 112.470 31.965 112.530 ;
        RECT 37.375 112.470 37.605 112.530 ;
        RECT 37.915 112.470 38.145 112.530 ;
        RECT 31.195 112.420 31.965 112.470 ;
        RECT 37.365 112.420 38.145 112.470 ;
        RECT 43.555 112.470 43.785 112.530 ;
        RECT 44.095 112.470 44.325 112.530 ;
        RECT 43.555 112.420 44.325 112.470 ;
        RECT 49.735 112.470 49.965 112.530 ;
        RECT 50.275 112.470 50.505 112.530 ;
        RECT 55.915 112.470 56.145 112.530 ;
        RECT 56.455 112.470 56.685 112.530 ;
        RECT 49.735 112.420 50.515 112.470 ;
        RECT 55.915 112.420 56.685 112.470 ;
        RECT 62.095 112.470 62.325 112.530 ;
        RECT 62.635 112.470 62.865 112.530 ;
        RECT 68.275 112.470 68.505 112.530 ;
        RECT 68.815 112.470 69.045 112.530 ;
        RECT 62.095 112.420 62.865 112.470 ;
        RECT 68.265 112.420 69.045 112.470 ;
        RECT 74.455 112.470 74.685 112.530 ;
        RECT 74.995 112.470 75.225 112.530 ;
        RECT 74.455 112.420 75.225 112.470 ;
        RECT 80.635 112.420 88.185 112.530 ;
        RECT 12.365 112.220 88.185 112.420 ;
        RECT 12.365 112.020 19.615 112.220 ;
        RECT 25.015 112.120 25.785 112.220 ;
        RECT 25.015 112.070 25.245 112.120 ;
        RECT 25.555 112.070 25.785 112.120 ;
        RECT 31.195 112.120 31.965 112.220 ;
        RECT 37.365 112.120 38.145 112.220 ;
        RECT 31.195 112.070 31.425 112.120 ;
        RECT 31.735 112.070 31.965 112.120 ;
        RECT 37.375 112.070 37.605 112.120 ;
        RECT 37.915 112.070 38.145 112.120 ;
        RECT 43.555 112.120 44.325 112.220 ;
        RECT 43.555 112.070 43.785 112.120 ;
        RECT 44.095 112.070 44.325 112.120 ;
        RECT 49.735 112.120 50.515 112.220 ;
        RECT 55.915 112.120 56.685 112.220 ;
        RECT 49.735 112.070 49.965 112.120 ;
        RECT 50.275 112.070 50.505 112.120 ;
        RECT 55.915 112.070 56.145 112.120 ;
        RECT 56.455 112.070 56.685 112.120 ;
        RECT 62.095 112.120 62.865 112.220 ;
        RECT 68.265 112.120 69.045 112.220 ;
        RECT 62.095 112.070 62.325 112.120 ;
        RECT 62.635 112.070 62.865 112.120 ;
        RECT 68.275 112.070 68.505 112.120 ;
        RECT 68.815 112.070 69.045 112.120 ;
        RECT 74.455 112.120 75.225 112.220 ;
        RECT 74.455 112.070 74.685 112.120 ;
        RECT 74.995 112.070 75.225 112.120 ;
        RECT 80.635 112.070 88.185 112.220 ;
        RECT 12.365 110.470 15.040 112.020 ;
        RECT 85.515 110.470 88.185 112.070 ;
        RECT 12.995 110.355 15.040 110.470 ;
        RECT 86.140 110.355 88.185 110.470 ;
        RECT 97.715 110.370 100.340 116.045 ;
        RECT 98.295 110.355 100.340 110.370 ;
        RECT 31.215 108.970 31.965 109.220 ;
        RECT 37.815 109.170 38.315 109.220 ;
        RECT 37.365 108.970 38.315 109.170 ;
        RECT 38.965 108.970 40.115 109.270 ;
        RECT 49.915 109.170 50.415 109.320 ;
        RECT 43.565 108.970 44.315 109.170 ;
        RECT 49.765 108.970 50.515 109.170 ;
        RECT 51.015 108.970 52.165 109.320 ;
        RECT 55.915 108.970 56.665 109.170 ;
        RECT 62.065 108.970 62.865 109.270 ;
        RECT 63.315 108.970 64.465 109.320 ;
        RECT 68.265 108.970 69.015 109.170 ;
        RECT 29.415 108.770 71.065 108.970 ;
        RECT 29.465 108.680 34.465 108.770 ;
        RECT 35.555 108.680 40.555 108.770 ;
        RECT 41.645 108.680 46.645 108.770 ;
        RECT 47.735 108.680 52.735 108.770 ;
        RECT 53.825 108.680 58.825 108.770 ;
        RECT 59.915 108.680 64.915 108.770 ;
        RECT 66.005 108.680 71.005 108.770 ;
        RECT 29.465 108.020 34.465 108.120 ;
        RECT 35.555 108.020 40.555 108.120 ;
        RECT 41.645 108.020 46.645 108.120 ;
        RECT 47.735 108.020 52.735 108.120 ;
        RECT 53.825 108.020 58.825 108.120 ;
        RECT 59.915 108.020 64.915 108.120 ;
        RECT 66.005 108.020 71.005 108.120 ;
        RECT 29.415 107.820 71.065 108.020 ;
        RECT 30.915 107.470 32.165 107.820 ;
        RECT 43.865 107.570 44.365 107.820 ;
        RECT 55.965 107.570 57.215 107.820 ;
        RECT 30.965 106.720 32.115 107.470 ;
        RECT 30.915 106.470 32.165 106.720 ;
        RECT 37.815 106.470 38.315 106.720 ;
        RECT 49.915 106.470 50.415 106.820 ;
        RECT 56.015 106.670 57.165 107.570 ;
        RECT 68.265 107.520 68.765 107.820 ;
        RECT 55.965 106.470 57.215 106.670 ;
        RECT 62.065 106.470 62.565 106.770 ;
        RECT 29.415 106.270 71.065 106.470 ;
        RECT 29.465 106.180 34.465 106.270 ;
        RECT 35.555 106.180 40.555 106.270 ;
        RECT 41.645 106.180 46.645 106.270 ;
        RECT 47.735 106.180 52.735 106.270 ;
        RECT 53.825 106.180 58.825 106.270 ;
        RECT 59.915 106.180 64.915 106.270 ;
        RECT 66.005 106.180 71.005 106.270 ;
        RECT 29.465 105.520 34.465 105.620 ;
        RECT 35.555 105.520 40.555 105.620 ;
        RECT 41.645 105.520 46.645 105.620 ;
        RECT 47.735 105.520 52.735 105.620 ;
        RECT 53.825 105.520 58.825 105.620 ;
        RECT 59.915 105.520 64.915 105.620 ;
        RECT 66.005 105.520 71.005 105.620 ;
        RECT 29.415 105.320 71.065 105.520 ;
        RECT 31.615 105.070 32.115 105.320 ;
        RECT 32.565 105.020 33.065 105.320 ;
        RECT 33.315 105.020 33.815 105.320 ;
        RECT 37.365 105.220 38.115 105.320 ;
        RECT 43.565 105.170 44.365 105.320 ;
        RECT 43.865 105.070 44.365 105.170 ;
        RECT 45.015 105.120 45.515 105.320 ;
        RECT 45.765 105.120 46.265 105.320 ;
        RECT 49.765 105.170 50.515 105.320 ;
        RECT 56.065 105.020 56.565 105.320 ;
        RECT 57.415 105.120 57.915 105.320 ;
        RECT 58.115 105.120 58.615 105.320 ;
        RECT 62.115 105.170 62.865 105.320 ;
        RECT 68.265 105.170 69.015 105.320 ;
        RECT 68.265 105.020 68.765 105.170 ;
        RECT 31.875 103.470 32.105 103.630 ;
        RECT 37.425 103.470 37.655 103.630 ;
        RECT 37.965 103.470 38.195 103.630 ;
        RECT 43.515 103.470 43.745 103.630 ;
        RECT 44.055 103.470 44.285 103.630 ;
        RECT 49.605 103.470 49.835 103.630 ;
        RECT 50.145 103.470 50.375 103.630 ;
        RECT 55.695 103.470 55.925 103.630 ;
        RECT 56.235 103.470 56.465 103.630 ;
        RECT 61.785 103.470 62.015 103.630 ;
        RECT 62.325 103.470 62.555 103.630 ;
        RECT 67.875 103.470 68.105 103.630 ;
        RECT 31.815 102.870 68.105 103.470 ;
        RECT 31.875 102.670 32.105 102.870 ;
        RECT 37.425 102.670 37.655 102.870 ;
        RECT 37.965 102.670 38.195 102.870 ;
        RECT 43.515 102.670 43.745 102.870 ;
        RECT 44.055 102.670 44.285 102.870 ;
        RECT 49.605 102.670 49.835 102.870 ;
        RECT 50.145 102.670 50.375 102.870 ;
        RECT 55.695 102.670 55.925 102.870 ;
        RECT 56.235 102.670 56.465 102.870 ;
        RECT 61.785 102.670 62.015 102.870 ;
        RECT 62.325 102.670 62.555 102.870 ;
        RECT 67.875 102.670 68.105 102.870 ;
        RECT 31.875 100.370 32.105 100.530 ;
        RECT 37.425 100.370 37.655 100.530 ;
        RECT 37.965 100.370 38.195 100.530 ;
        RECT 43.515 100.370 43.745 100.530 ;
        RECT 44.055 100.370 44.285 100.530 ;
        RECT 49.605 100.370 49.835 100.530 ;
        RECT 50.145 100.370 50.375 100.530 ;
        RECT 55.695 100.370 55.925 100.530 ;
        RECT 56.235 100.370 56.465 100.530 ;
        RECT 61.785 100.370 62.015 100.530 ;
        RECT 62.325 100.370 62.555 100.530 ;
        RECT 67.875 100.370 68.105 100.530 ;
        RECT 31.875 100.320 68.115 100.370 ;
        RECT 31.715 99.820 68.115 100.320 ;
        RECT 31.875 99.770 68.115 99.820 ;
        RECT 31.875 99.570 32.105 99.770 ;
        RECT 37.425 99.570 37.655 99.770 ;
        RECT 37.965 99.570 38.195 99.770 ;
        RECT 43.515 99.570 43.745 99.770 ;
        RECT 44.055 99.570 44.285 99.770 ;
        RECT 49.605 99.570 49.835 99.770 ;
        RECT 50.145 99.570 50.375 99.770 ;
        RECT 55.695 99.570 55.925 99.770 ;
        RECT 56.235 99.570 56.465 99.770 ;
        RECT 61.785 99.570 62.015 99.770 ;
        RECT 62.325 99.570 62.555 99.770 ;
        RECT 67.875 99.570 68.105 99.770 ;
        RECT 29.075 97.370 29.305 97.530 ;
        RECT 34.625 97.370 34.855 97.530 ;
        RECT 35.165 97.370 35.395 97.530 ;
        RECT 40.715 97.370 40.945 97.530 ;
        RECT 41.255 97.370 41.485 97.530 ;
        RECT 46.805 97.370 47.035 97.530 ;
        RECT 47.345 97.370 47.575 97.530 ;
        RECT 52.895 97.370 53.125 97.530 ;
        RECT 53.435 97.370 53.665 97.530 ;
        RECT 58.985 97.370 59.215 97.530 ;
        RECT 59.525 97.370 59.755 97.530 ;
        RECT 65.075 97.370 65.305 97.530 ;
        RECT 65.615 97.370 65.845 97.530 ;
        RECT 71.165 97.370 71.395 97.530 ;
        RECT 29.015 96.770 71.415 97.370 ;
        RECT 29.075 96.570 29.305 96.770 ;
        RECT 34.625 96.570 34.855 96.770 ;
        RECT 35.165 96.570 35.395 96.770 ;
        RECT 40.715 96.570 40.945 96.770 ;
        RECT 41.255 96.570 41.485 96.770 ;
        RECT 46.805 96.570 47.035 96.770 ;
        RECT 47.345 96.570 47.575 96.770 ;
        RECT 52.895 96.570 53.125 96.770 ;
        RECT 53.435 96.570 53.665 96.770 ;
        RECT 58.985 96.570 59.215 96.770 ;
        RECT 59.525 96.570 59.755 96.770 ;
        RECT 65.075 96.570 65.305 96.770 ;
        RECT 65.615 96.570 65.845 96.770 ;
        RECT 71.165 96.570 71.395 96.770 ;
        RECT 29.465 96.370 34.465 96.520 ;
        RECT 35.555 96.370 40.555 96.520 ;
        RECT 41.645 96.370 46.645 96.520 ;
        RECT 47.735 96.370 52.735 96.520 ;
        RECT 53.825 96.370 58.825 96.520 ;
        RECT 59.915 96.370 64.915 96.520 ;
        RECT 66.005 96.370 71.005 96.520 ;
        RECT 29.415 96.170 71.015 96.370 ;
        RECT 30.915 96.070 31.465 96.170 ;
        RECT 31.615 96.070 32.165 96.170 ;
        RECT 55.965 96.070 56.515 96.170 ;
        RECT 56.665 96.070 57.215 96.170 ;
        RECT 29.075 94.370 29.305 94.530 ;
        RECT 34.625 94.370 34.855 94.530 ;
        RECT 35.165 94.370 35.395 94.530 ;
        RECT 40.715 94.370 40.945 94.530 ;
        RECT 41.255 94.370 41.485 94.530 ;
        RECT 46.805 94.370 47.035 94.530 ;
        RECT 47.345 94.370 47.575 94.530 ;
        RECT 52.895 94.370 53.125 94.530 ;
        RECT 53.435 94.370 53.665 94.530 ;
        RECT 58.985 94.370 59.215 94.530 ;
        RECT 59.525 94.370 59.755 94.530 ;
        RECT 65.075 94.370 65.305 94.530 ;
        RECT 65.615 94.370 65.845 94.530 ;
        RECT 71.165 94.370 71.395 94.530 ;
        RECT 29.075 93.770 71.415 94.370 ;
        RECT 29.075 93.570 29.305 93.770 ;
        RECT 34.625 93.570 34.855 93.770 ;
        RECT 35.165 93.570 35.395 93.770 ;
        RECT 40.715 93.570 40.945 93.770 ;
        RECT 41.255 93.570 41.485 93.770 ;
        RECT 46.805 93.570 47.035 93.770 ;
        RECT 47.345 93.570 47.575 93.770 ;
        RECT 52.895 93.570 53.125 93.770 ;
        RECT 53.435 93.570 53.665 93.770 ;
        RECT 58.985 93.570 59.215 93.770 ;
        RECT 59.525 93.570 59.755 93.770 ;
        RECT 65.075 93.570 65.305 93.770 ;
        RECT 65.615 93.570 65.845 93.770 ;
        RECT 71.165 93.570 71.395 93.770 ;
        RECT 29.465 93.370 34.465 93.520 ;
        RECT 35.555 93.370 40.555 93.520 ;
        RECT 41.645 93.370 46.645 93.520 ;
        RECT 47.735 93.370 52.735 93.520 ;
        RECT 53.825 93.370 58.825 93.520 ;
        RECT 59.915 93.370 64.915 93.520 ;
        RECT 66.005 93.370 71.005 93.520 ;
        RECT 29.415 93.170 71.015 93.370 ;
        RECT 30.915 92.970 31.465 93.170 ;
        RECT 31.615 92.970 32.165 93.170 ;
        RECT 55.965 93.070 56.515 93.170 ;
        RECT 56.665 93.070 57.215 93.170 ;
        RECT 31.800 89.400 32.030 89.660 ;
        RECT 37.440 89.400 37.670 89.660 ;
        RECT 37.980 89.400 38.210 89.660 ;
        RECT 43.620 89.400 43.850 89.660 ;
        RECT 44.160 89.400 44.390 89.660 ;
        RECT 49.800 89.400 50.030 89.660 ;
        RECT 50.340 89.400 50.570 89.660 ;
        RECT 55.980 89.400 56.210 89.660 ;
        RECT 56.520 89.400 56.750 89.660 ;
        RECT 62.160 89.400 62.390 89.660 ;
        RECT 62.700 89.400 62.930 89.660 ;
        RECT 68.340 89.400 68.570 89.660 ;
        RECT 31.800 88.700 68.570 89.400 ;
        RECT 31.800 88.340 68.540 88.700 ;
        RECT 31.800 86.450 32.030 86.710 ;
        RECT 37.440 86.450 37.670 86.710 ;
        RECT 37.980 86.450 38.210 86.710 ;
        RECT 43.620 86.450 43.850 86.710 ;
        RECT 44.160 86.450 44.390 86.710 ;
        RECT 49.800 86.450 50.030 86.710 ;
        RECT 50.340 86.450 50.570 86.710 ;
        RECT 55.980 86.450 56.210 86.710 ;
        RECT 56.520 86.450 56.750 86.710 ;
        RECT 62.160 86.450 62.390 86.710 ;
        RECT 62.700 86.450 62.930 86.710 ;
        RECT 68.340 86.450 68.570 86.710 ;
        RECT 31.790 86.000 68.570 86.450 ;
        RECT 31.800 85.750 32.030 86.000 ;
        RECT 37.440 85.750 37.670 86.000 ;
        RECT 37.980 85.750 38.210 86.000 ;
        RECT 43.620 85.750 43.850 86.000 ;
        RECT 44.160 85.750 44.390 86.000 ;
        RECT 49.800 85.750 50.030 86.000 ;
        RECT 50.340 85.750 50.570 86.000 ;
        RECT 55.980 85.750 56.210 86.000 ;
        RECT 56.520 85.750 56.750 86.000 ;
        RECT 62.160 85.750 62.390 86.000 ;
        RECT 62.700 85.750 62.930 86.000 ;
        RECT 68.340 85.750 68.570 86.000 ;
        RECT 32.190 85.600 37.235 85.700 ;
        RECT 38.415 85.600 43.415 85.700 ;
        RECT 44.595 85.600 49.595 85.700 ;
        RECT 50.775 85.600 55.775 85.700 ;
        RECT 56.955 85.600 61.955 85.700 ;
        RECT 63.135 85.600 68.160 85.700 ;
        RECT 32.190 85.200 68.160 85.600 ;
        RECT 49.170 83.150 51.070 83.190 ;
        RECT 45.590 82.760 54.690 83.150 ;
        RECT 45.590 82.400 54.700 82.760 ;
        RECT 45.650 82.000 54.700 82.400 ;
        RECT 45.650 81.800 45.880 82.000 ;
        RECT 47.440 81.800 48.240 82.000 ;
        RECT 49.790 81.800 50.565 82.000 ;
        RECT 52.130 81.800 52.915 82.000 ;
        RECT 54.470 81.800 54.700 82.000 ;
        RECT 57.390 80.200 59.140 80.300 ;
        RECT 41.490 79.300 59.140 80.200 ;
        RECT 41.490 79.150 43.140 79.300 ;
        RECT 46.750 79.175 46.980 79.300 ;
        RECT 49.800 79.175 50.030 79.300 ;
        RECT 50.340 79.175 50.570 79.300 ;
        RECT 53.390 79.175 53.620 79.300 ;
        RECT 47.140 79.025 49.640 79.125 ;
        RECT 50.730 79.025 53.230 79.125 ;
        RECT 47.115 78.950 53.290 79.025 ;
        RECT 47.090 78.600 53.340 78.950 ;
        RECT 32.440 77.290 67.890 77.525 ;
        RECT 32.440 77.150 67.915 77.290 ;
        RECT 32.465 77.060 37.465 77.150 ;
        RECT 38.555 77.060 43.555 77.150 ;
        RECT 44.645 77.060 49.645 77.150 ;
        RECT 50.735 77.060 55.735 77.150 ;
        RECT 56.825 77.060 61.825 77.150 ;
        RECT 62.915 77.060 67.915 77.150 ;
        RECT 32.075 76.775 32.305 77.010 ;
        RECT 37.625 76.775 37.855 77.010 ;
        RECT 38.165 76.775 38.395 77.010 ;
        RECT 43.715 76.775 43.945 77.010 ;
        RECT 44.255 76.775 44.485 77.010 ;
        RECT 49.805 76.775 50.035 77.010 ;
        RECT 50.345 76.775 50.575 77.010 ;
        RECT 55.895 76.775 56.125 77.010 ;
        RECT 56.435 76.775 56.665 77.010 ;
        RECT 61.985 76.775 62.215 77.010 ;
        RECT 62.525 76.775 62.755 77.010 ;
        RECT 68.075 76.775 68.305 77.010 ;
        RECT 32.075 76.350 68.305 76.775 ;
        RECT 32.075 76.050 32.305 76.350 ;
        RECT 37.625 76.050 37.855 76.350 ;
        RECT 38.165 76.050 38.395 76.350 ;
        RECT 43.715 76.050 43.945 76.350 ;
        RECT 44.255 76.050 44.485 76.350 ;
        RECT 49.805 76.050 50.035 76.350 ;
        RECT 50.345 76.050 50.575 76.350 ;
        RECT 55.895 76.050 56.125 76.350 ;
        RECT 56.435 76.050 56.665 76.350 ;
        RECT 61.985 76.050 62.215 76.350 ;
        RECT 62.525 76.050 62.755 76.350 ;
        RECT 68.075 76.050 68.305 76.350 ;
        RECT 32.465 75.900 37.465 76.000 ;
        RECT 38.555 75.900 43.555 76.000 ;
        RECT 44.645 75.900 49.645 76.000 ;
        RECT 50.735 75.900 55.735 76.000 ;
        RECT 56.825 75.900 61.825 76.000 ;
        RECT 62.915 75.900 67.915 76.000 ;
        RECT 32.440 75.770 67.915 75.900 ;
        RECT 32.440 75.525 67.890 75.770 ;
        RECT 39.190 74.050 41.190 75.525 ;
        RECT 46.190 74.050 48.190 75.525 ;
        RECT 52.690 74.050 54.690 75.525 ;
        RECT 59.140 74.050 61.190 75.525 ;
        RECT 35.190 71.050 65.190 74.050 ;
      LAYER via ;
        RECT 32.685 136.640 32.945 136.900 ;
        RECT 33.435 136.640 33.695 136.900 ;
        RECT 34.300 136.865 34.560 137.125 ;
        RECT 34.620 136.865 34.880 137.125 ;
        RECT 40.500 136.865 40.760 137.125 ;
        RECT 40.820 136.865 41.080 137.125 ;
        RECT 45.135 136.640 45.395 136.900 ;
        RECT 45.885 136.640 46.145 136.900 ;
        RECT 46.650 136.865 46.910 137.125 ;
        RECT 46.970 136.865 47.230 137.125 ;
        RECT 52.850 136.865 53.110 137.125 ;
        RECT 53.170 136.865 53.430 137.125 ;
        RECT 57.535 136.640 57.795 136.900 ;
        RECT 58.285 136.640 58.545 136.900 ;
        RECT 59.050 136.865 59.310 137.125 ;
        RECT 59.370 136.865 59.630 137.125 ;
        RECT 65.200 136.865 65.460 137.125 ;
        RECT 65.520 136.865 65.780 137.125 ;
        RECT 30.735 136.290 30.995 136.550 ;
        RECT 31.585 136.290 31.845 136.550 ;
        RECT 43.335 136.290 43.595 136.550 ;
        RECT 44.185 136.290 44.445 136.550 ;
        RECT 55.785 136.290 56.045 136.550 ;
        RECT 56.635 136.290 56.895 136.550 ;
        RECT 68.035 136.290 68.295 136.550 ;
        RECT 68.885 136.290 69.145 136.550 ;
        RECT 32.685 133.940 32.945 134.200 ;
        RECT 33.435 133.940 33.695 134.200 ;
        RECT 34.300 134.165 34.560 134.425 ;
        RECT 34.620 134.165 34.880 134.425 ;
        RECT 40.500 134.165 40.760 134.425 ;
        RECT 40.820 134.165 41.080 134.425 ;
        RECT 45.135 133.940 45.395 134.200 ;
        RECT 45.885 133.940 46.145 134.200 ;
        RECT 46.650 134.165 46.910 134.425 ;
        RECT 46.970 134.165 47.230 134.425 ;
        RECT 52.850 134.165 53.110 134.425 ;
        RECT 53.170 134.165 53.430 134.425 ;
        RECT 57.535 133.940 57.795 134.200 ;
        RECT 58.285 133.940 58.545 134.200 ;
        RECT 59.050 134.165 59.310 134.425 ;
        RECT 59.370 134.165 59.630 134.425 ;
        RECT 65.200 134.165 65.460 134.425 ;
        RECT 65.520 134.165 65.780 134.425 ;
        RECT 30.735 133.590 30.995 133.850 ;
        RECT 31.585 133.590 31.845 133.850 ;
        RECT 43.335 133.590 43.595 133.850 ;
        RECT 44.185 133.590 44.445 133.850 ;
        RECT 55.785 133.590 56.045 133.850 ;
        RECT 56.635 133.590 56.895 133.850 ;
        RECT 68.035 133.540 68.295 133.800 ;
        RECT 68.885 133.540 69.145 133.800 ;
        RECT 32.685 131.240 32.945 131.500 ;
        RECT 33.435 131.240 33.695 131.500 ;
        RECT 34.300 131.465 34.560 131.725 ;
        RECT 34.620 131.465 34.880 131.725 ;
        RECT 40.500 131.465 40.760 131.725 ;
        RECT 40.820 131.465 41.080 131.725 ;
        RECT 45.135 131.240 45.395 131.500 ;
        RECT 45.885 131.240 46.145 131.500 ;
        RECT 46.650 131.465 46.910 131.725 ;
        RECT 46.970 131.465 47.230 131.725 ;
        RECT 52.850 131.465 53.110 131.725 ;
        RECT 53.170 131.465 53.430 131.725 ;
        RECT 57.585 131.240 57.845 131.500 ;
        RECT 58.285 131.240 58.545 131.500 ;
        RECT 59.050 131.465 59.310 131.725 ;
        RECT 59.370 131.465 59.630 131.725 ;
        RECT 65.200 131.465 65.460 131.725 ;
        RECT 65.520 131.465 65.780 131.725 ;
        RECT 30.735 130.890 30.995 131.150 ;
        RECT 31.585 130.890 31.845 131.150 ;
        RECT 43.335 130.890 43.595 131.150 ;
        RECT 44.185 130.890 44.445 131.150 ;
        RECT 55.785 130.840 56.045 131.100 ;
        RECT 56.635 130.840 56.895 131.100 ;
        RECT 68.035 130.890 68.295 131.150 ;
        RECT 68.885 130.890 69.145 131.150 ;
        RECT 34.300 128.765 34.560 129.025 ;
        RECT 34.620 128.765 34.880 129.025 ;
        RECT 40.500 128.765 40.760 129.025 ;
        RECT 40.820 128.765 41.080 129.025 ;
        RECT 46.650 128.765 46.910 129.025 ;
        RECT 46.970 128.765 47.230 129.025 ;
        RECT 52.850 128.765 53.110 129.025 ;
        RECT 53.170 128.765 53.430 129.025 ;
        RECT 59.000 128.765 59.260 129.025 ;
        RECT 59.320 128.765 59.580 129.025 ;
        RECT 65.200 128.765 65.460 129.025 ;
        RECT 65.520 128.765 65.780 129.025 ;
        RECT 30.735 128.190 30.995 128.450 ;
        RECT 31.585 128.190 31.845 128.450 ;
        RECT 39.135 128.240 39.395 128.500 ;
        RECT 39.685 128.240 39.945 128.500 ;
        RECT 43.285 128.190 43.545 128.450 ;
        RECT 44.135 128.190 44.395 128.450 ;
        RECT 51.185 128.240 51.445 128.500 ;
        RECT 51.735 128.240 51.995 128.500 ;
        RECT 55.735 128.190 55.995 128.450 ;
        RECT 56.585 128.190 56.845 128.450 ;
        RECT 63.485 128.190 63.745 128.450 ;
        RECT 64.035 128.190 64.295 128.450 ;
        RECT 68.185 128.190 68.445 128.450 ;
        RECT 69.035 128.190 69.295 128.450 ;
        RECT 34.300 125.865 34.560 126.125 ;
        RECT 34.620 125.865 34.880 126.125 ;
        RECT 40.500 125.865 40.760 126.125 ;
        RECT 40.820 125.865 41.080 126.125 ;
        RECT 46.700 125.865 46.960 126.125 ;
        RECT 47.020 125.865 47.280 126.125 ;
        RECT 52.850 125.865 53.110 126.125 ;
        RECT 53.170 125.865 53.430 126.125 ;
        RECT 59.000 125.865 59.260 126.125 ;
        RECT 59.320 125.865 59.580 126.125 ;
        RECT 65.200 125.865 65.460 126.125 ;
        RECT 65.520 125.865 65.780 126.125 ;
        RECT 30.735 125.290 30.995 125.550 ;
        RECT 31.585 125.290 31.845 125.550 ;
        RECT 39.135 125.190 39.395 125.450 ;
        RECT 39.685 125.190 39.945 125.450 ;
        RECT 43.285 125.290 43.545 125.550 ;
        RECT 44.135 125.290 44.395 125.550 ;
        RECT 51.185 125.290 51.445 125.550 ;
        RECT 51.735 125.290 51.995 125.550 ;
        RECT 55.735 125.240 55.995 125.500 ;
        RECT 56.585 125.240 56.845 125.500 ;
        RECT 63.485 125.290 63.745 125.550 ;
        RECT 64.035 125.290 64.295 125.550 ;
        RECT 68.185 125.290 68.445 125.550 ;
        RECT 69.035 125.290 69.295 125.550 ;
        RECT 0.350 123.580 0.930 124.160 ;
        RECT 1.600 123.580 2.180 124.160 ;
        RECT 97.850 124.430 98.430 125.010 ;
        RECT 99.150 124.430 99.730 125.010 ;
        RECT 34.300 122.965 34.560 123.225 ;
        RECT 34.620 122.965 34.880 123.225 ;
        RECT 40.500 122.965 40.760 123.225 ;
        RECT 40.820 122.965 41.080 123.225 ;
        RECT 46.650 122.965 46.910 123.225 ;
        RECT 46.970 122.965 47.230 123.225 ;
        RECT 52.850 122.965 53.110 123.225 ;
        RECT 53.170 122.965 53.430 123.225 ;
        RECT 59.000 122.965 59.260 123.225 ;
        RECT 59.320 122.965 59.580 123.225 ;
        RECT 65.200 122.965 65.460 123.225 ;
        RECT 65.520 122.965 65.780 123.225 ;
        RECT 30.635 122.240 30.895 122.500 ;
        RECT 31.685 122.240 31.945 122.500 ;
        RECT 43.285 122.390 43.545 122.650 ;
        RECT 44.135 122.390 44.395 122.650 ;
        RECT 51.185 122.390 51.445 122.650 ;
        RECT 51.735 122.390 51.995 122.650 ;
        RECT 55.735 122.390 55.995 122.650 ;
        RECT 56.585 122.390 56.845 122.650 ;
        RECT 63.485 122.390 63.745 122.650 ;
        RECT 64.035 122.390 64.295 122.650 ;
        RECT 68.185 122.390 68.445 122.650 ;
        RECT 69.035 122.390 69.295 122.650 ;
        RECT 25.100 120.265 25.360 120.525 ;
        RECT 25.420 120.265 25.680 120.525 ;
        RECT 31.300 120.265 31.560 120.525 ;
        RECT 31.620 120.265 31.880 120.525 ;
        RECT 37.450 120.265 37.710 120.525 ;
        RECT 37.770 120.265 38.030 120.525 ;
        RECT 43.650 120.265 43.910 120.525 ;
        RECT 43.970 120.265 44.230 120.525 ;
        RECT 49.850 120.265 50.110 120.525 ;
        RECT 50.170 120.265 50.430 120.525 ;
        RECT 56.000 120.265 56.260 120.525 ;
        RECT 56.320 120.265 56.580 120.525 ;
        RECT 62.200 120.265 62.460 120.525 ;
        RECT 62.520 120.265 62.780 120.525 ;
        RECT 68.350 120.265 68.610 120.525 ;
        RECT 68.670 120.265 68.930 120.525 ;
        RECT 74.550 120.265 74.810 120.525 ;
        RECT 74.870 120.265 75.130 120.525 ;
        RECT 25.100 117.615 25.360 117.875 ;
        RECT 25.420 117.615 25.680 117.875 ;
        RECT 31.300 117.565 31.560 117.825 ;
        RECT 31.620 117.565 31.880 117.825 ;
        RECT 37.450 117.565 37.710 117.825 ;
        RECT 37.770 117.565 38.030 117.825 ;
        RECT 43.650 117.565 43.910 117.825 ;
        RECT 43.970 117.565 44.230 117.825 ;
        RECT 49.850 117.565 50.110 117.825 ;
        RECT 50.170 117.565 50.430 117.825 ;
        RECT 56.000 117.565 56.260 117.825 ;
        RECT 56.320 117.565 56.580 117.825 ;
        RECT 62.200 117.565 62.460 117.825 ;
        RECT 62.520 117.565 62.780 117.825 ;
        RECT 68.350 117.565 68.610 117.825 ;
        RECT 68.670 117.565 68.930 117.825 ;
        RECT 74.550 117.565 74.810 117.825 ;
        RECT 74.870 117.565 75.130 117.825 ;
        RECT 25.100 114.865 25.360 115.125 ;
        RECT 25.420 114.865 25.680 115.125 ;
        RECT 31.300 114.865 31.560 115.125 ;
        RECT 31.620 114.865 31.880 115.125 ;
        RECT 37.450 114.865 37.710 115.125 ;
        RECT 37.770 114.865 38.030 115.125 ;
        RECT 43.650 114.865 43.910 115.125 ;
        RECT 43.970 114.865 44.230 115.125 ;
        RECT 49.850 114.865 50.110 115.125 ;
        RECT 50.170 114.865 50.430 115.125 ;
        RECT 56.000 114.865 56.260 115.125 ;
        RECT 56.320 114.865 56.580 115.125 ;
        RECT 62.200 114.865 62.460 115.125 ;
        RECT 62.520 114.865 62.780 115.125 ;
        RECT 68.350 114.865 68.610 115.125 ;
        RECT 68.670 114.865 68.930 115.125 ;
        RECT 74.550 114.865 74.810 115.125 ;
        RECT 74.870 114.865 75.130 115.125 ;
        RECT 25.100 112.165 25.360 112.425 ;
        RECT 25.420 112.165 25.680 112.425 ;
        RECT 31.300 112.165 31.560 112.425 ;
        RECT 31.620 112.165 31.880 112.425 ;
        RECT 37.450 112.165 37.710 112.425 ;
        RECT 37.770 112.165 38.030 112.425 ;
        RECT 43.650 112.165 43.910 112.425 ;
        RECT 43.970 112.165 44.230 112.425 ;
        RECT 49.850 112.165 50.110 112.425 ;
        RECT 50.170 112.165 50.430 112.425 ;
        RECT 56.000 112.165 56.260 112.425 ;
        RECT 56.320 112.165 56.580 112.425 ;
        RECT 62.200 112.165 62.460 112.425 ;
        RECT 62.520 112.165 62.780 112.425 ;
        RECT 68.350 112.165 68.610 112.425 ;
        RECT 68.670 112.165 68.930 112.425 ;
        RECT 74.550 112.165 74.810 112.425 ;
        RECT 74.870 112.165 75.130 112.425 ;
        RECT 31.300 108.915 31.560 109.175 ;
        RECT 31.620 108.915 31.880 109.175 ;
        RECT 37.450 108.865 37.710 109.125 ;
        RECT 37.770 108.865 38.030 109.125 ;
        RECT 39.135 108.890 39.395 109.150 ;
        RECT 39.685 108.890 39.945 109.150 ;
        RECT 43.650 108.865 43.910 109.125 ;
        RECT 43.970 108.865 44.230 109.125 ;
        RECT 49.850 108.865 50.110 109.125 ;
        RECT 50.170 108.865 50.430 109.125 ;
        RECT 51.185 108.890 51.445 109.150 ;
        RECT 51.735 108.890 51.995 109.150 ;
        RECT 56.000 108.865 56.260 109.125 ;
        RECT 56.320 108.865 56.580 109.125 ;
        RECT 62.200 108.965 62.460 109.225 ;
        RECT 62.520 108.965 62.780 109.225 ;
        RECT 63.485 108.940 63.745 109.200 ;
        RECT 64.035 108.940 64.295 109.200 ;
        RECT 68.350 108.865 68.610 109.125 ;
        RECT 68.670 108.865 68.930 109.125 ;
        RECT 31.060 107.540 31.320 107.800 ;
        RECT 31.760 107.540 32.020 107.800 ;
        RECT 56.110 107.640 56.370 107.900 ;
        RECT 56.810 107.640 57.070 107.900 ;
        RECT 31.060 106.390 31.320 106.650 ;
        RECT 31.760 106.390 32.020 106.650 ;
        RECT 56.110 106.340 56.370 106.600 ;
        RECT 56.810 106.340 57.070 106.600 ;
        RECT 32.685 105.090 32.945 105.350 ;
        RECT 33.435 105.090 33.695 105.350 ;
        RECT 45.135 105.190 45.395 105.450 ;
        RECT 45.885 105.190 46.145 105.450 ;
        RECT 57.535 105.190 57.795 105.450 ;
        RECT 58.235 105.190 58.495 105.450 ;
        RECT 40.835 103.040 41.095 103.300 ;
        RECT 52.885 103.040 53.145 103.300 ;
        RECT 37.810 99.940 38.070 100.200 ;
        RECT 38.410 99.940 38.670 100.200 ;
        RECT 40.835 99.940 41.095 100.200 ;
        RECT 50.060 99.940 50.320 100.200 ;
        RECT 50.660 99.940 50.920 100.200 ;
        RECT 52.885 99.940 53.145 100.200 ;
        RECT 62.210 99.940 62.470 100.200 ;
        RECT 62.810 99.940 63.070 100.200 ;
        RECT 37.810 96.940 38.070 97.200 ;
        RECT 38.410 96.940 38.670 97.200 ;
        RECT 50.060 96.940 50.320 97.200 ;
        RECT 50.660 96.940 50.920 97.200 ;
        RECT 62.210 96.940 62.470 97.200 ;
        RECT 62.810 96.940 63.070 97.200 ;
        RECT 31.060 96.140 31.320 96.400 ;
        RECT 31.760 96.140 32.020 96.400 ;
        RECT 56.110 96.140 56.370 96.400 ;
        RECT 56.810 96.140 57.070 96.400 ;
        RECT 37.810 93.940 38.070 94.200 ;
        RECT 38.410 93.940 38.670 94.200 ;
        RECT 49.360 93.935 49.620 94.195 ;
        RECT 50.060 93.940 50.320 94.200 ;
        RECT 50.660 93.940 50.920 94.200 ;
        RECT 62.210 93.940 62.470 94.200 ;
        RECT 62.810 93.940 63.070 94.200 ;
        RECT 31.060 93.040 31.320 93.300 ;
        RECT 31.760 93.040 32.020 93.300 ;
        RECT 56.110 93.140 56.370 93.400 ;
        RECT 56.810 93.140 57.070 93.400 ;
        RECT 41.635 89.045 41.895 89.305 ;
        RECT 42.735 89.045 42.995 89.305 ;
        RECT 57.535 89.045 57.795 89.305 ;
        RECT 58.735 89.045 58.995 89.305 ;
        RECT 41.635 86.095 41.895 86.355 ;
        RECT 42.735 86.095 42.995 86.355 ;
        RECT 57.535 86.095 57.795 86.355 ;
        RECT 58.735 86.095 58.995 86.355 ;
        RECT 47.435 85.295 47.695 85.555 ;
        RECT 47.985 85.295 48.245 85.555 ;
        RECT 52.135 85.295 52.395 85.555 ;
        RECT 52.685 85.295 52.945 85.555 ;
        RECT 49.240 82.910 49.500 83.170 ;
        RECT 49.740 82.910 50.000 83.170 ;
        RECT 50.240 82.910 50.500 83.170 ;
        RECT 50.740 82.910 51.000 83.170 ;
        RECT 47.435 82.445 47.695 82.705 ;
        RECT 47.985 82.445 48.245 82.705 ;
        RECT 52.135 82.495 52.395 82.755 ;
        RECT 52.685 82.495 52.945 82.755 ;
        RECT 41.635 79.795 41.895 80.055 ;
        RECT 42.685 79.795 42.945 80.055 ;
        RECT 57.535 79.895 57.795 80.155 ;
        RECT 58.735 79.895 58.995 80.155 ;
        RECT 41.635 79.345 41.895 79.605 ;
        RECT 42.685 79.345 42.945 79.605 ;
        RECT 57.535 79.445 57.795 79.705 ;
        RECT 58.735 79.445 58.995 79.705 ;
        RECT 47.435 78.695 47.695 78.955 ;
        RECT 47.985 78.695 48.245 78.955 ;
        RECT 52.135 78.695 52.395 78.955 ;
        RECT 52.685 78.695 52.945 78.955 ;
        RECT 41.635 77.195 41.895 77.455 ;
        RECT 42.735 77.195 42.995 77.455 ;
        RECT 57.535 77.195 57.795 77.455 ;
        RECT 58.735 77.195 58.995 77.455 ;
        RECT 47.435 76.445 47.695 76.705 ;
        RECT 47.985 76.445 48.245 76.705 ;
        RECT 52.135 76.445 52.395 76.705 ;
        RECT 52.685 76.445 52.945 76.705 ;
      LAYER met2 ;
        RECT 30.565 130.720 32.015 137.220 ;
        RECT 32.615 136.520 33.015 137.020 ;
        RECT 33.365 136.520 33.765 137.020 ;
        RECT 32.615 133.820 33.015 134.320 ;
        RECT 33.365 133.820 33.765 134.320 ;
        RECT 32.615 131.120 33.015 131.620 ;
        RECT 33.365 131.120 33.765 131.620 ;
        RECT 0.315 123.470 0.965 124.270 ;
        RECT 1.565 123.470 2.215 124.270 ;
        RECT 30.565 122.170 32.015 128.670 ;
        RECT 34.215 122.720 34.965 137.420 ;
        RECT 39.065 128.120 39.465 128.620 ;
        RECT 39.615 128.120 40.015 128.620 ;
        RECT 39.065 125.070 39.465 125.570 ;
        RECT 39.615 125.070 40.015 125.570 ;
        RECT 38.965 122.320 40.115 122.770 ;
        RECT 40.415 122.520 41.165 137.470 ;
        RECT 43.165 130.670 44.615 137.620 ;
        RECT 45.065 136.520 45.465 137.020 ;
        RECT 45.815 136.520 46.215 137.020 ;
        RECT 45.065 133.820 45.465 134.320 ;
        RECT 45.815 133.820 46.215 134.320 ;
        RECT 45.065 131.120 45.465 131.620 ;
        RECT 45.815 131.120 46.215 131.620 ;
        RECT 30.565 122.120 30.965 122.170 ;
        RECT 31.615 122.120 32.015 122.170 ;
        RECT 43.075 122.030 44.735 128.770 ;
        RECT 46.565 122.770 47.315 137.420 ;
        RECT 51.115 128.120 51.515 128.620 ;
        RECT 51.665 128.120 52.065 128.620 ;
        RECT 51.115 125.170 51.515 125.670 ;
        RECT 51.665 125.170 52.065 125.670 ;
        RECT 52.765 122.770 53.515 137.420 ;
        RECT 55.615 130.670 57.065 137.620 ;
        RECT 57.465 136.520 57.865 137.020 ;
        RECT 58.215 136.520 58.615 137.020 ;
        RECT 58.965 135.720 59.715 137.370 ;
        RECT 57.465 133.820 57.865 134.320 ;
        RECT 58.215 133.820 58.615 134.320 ;
        RECT 57.515 131.120 57.915 131.620 ;
        RECT 58.215 131.120 58.615 131.620 ;
        RECT 58.915 131.220 59.715 135.720 ;
        RECT 51.115 122.270 51.515 122.770 ;
        RECT 51.665 122.270 52.065 122.770 ;
        RECT 55.565 122.220 57.015 128.720 ;
        RECT 58.915 122.720 59.665 131.220 ;
        RECT 63.415 128.070 63.815 128.570 ;
        RECT 63.965 128.070 64.365 128.570 ;
        RECT 63.415 125.170 63.815 125.670 ;
        RECT 63.965 125.170 64.365 125.670 ;
        RECT 65.115 122.770 65.865 137.320 ;
        RECT 67.865 130.770 69.315 137.970 ;
        RECT 63.415 122.270 63.815 122.770 ;
        RECT 63.965 122.270 64.365 122.770 ;
        RECT 68.015 122.220 69.465 128.970 ;
        RECT 97.815 124.320 98.465 125.120 ;
        RECT 99.115 124.320 99.765 125.120 ;
        RECT 25.015 111.920 25.765 120.720 ;
        RECT 31.215 108.820 31.965 120.770 ;
        RECT 37.365 108.570 38.115 120.720 ;
        RECT 39.065 108.770 39.465 109.270 ;
        RECT 39.615 108.770 40.015 109.270 ;
        RECT 43.565 108.370 44.315 120.720 ;
        RECT 49.765 108.470 50.515 120.670 ;
        RECT 51.115 108.770 51.515 109.270 ;
        RECT 51.665 108.770 52.065 109.270 ;
        RECT 55.915 108.770 56.665 120.720 ;
        RECT 62.115 108.620 62.865 120.820 ;
        RECT 63.415 108.820 63.815 109.320 ;
        RECT 63.965 108.820 64.365 109.320 ;
        RECT 68.265 108.620 69.015 120.770 ;
        RECT 74.465 111.970 75.215 120.770 ;
        RECT 56.015 107.970 56.465 108.020 ;
        RECT 56.715 107.970 57.165 108.020 ;
        RECT 30.965 107.820 31.415 107.920 ;
        RECT 31.665 107.820 32.115 107.920 ;
        RECT 30.965 92.920 32.115 107.820 ;
        RECT 32.515 105.020 33.865 105.470 ;
        RECT 45.065 105.070 45.465 105.570 ;
        RECT 45.815 105.070 46.215 105.570 ;
        RECT 32.615 104.970 33.015 105.020 ;
        RECT 33.365 104.970 33.765 105.020 ;
        RECT 37.715 93.820 38.765 100.370 ;
        RECT 40.765 99.820 41.165 103.520 ;
        RECT 49.965 94.540 51.015 100.370 ;
        RECT 52.815 99.820 53.215 103.520 ;
        RECT 41.490 77.100 43.140 89.350 ;
        RECT 47.290 76.050 48.390 85.650 ;
        RECT 49.120 82.790 51.120 94.540 ;
        RECT 56.015 93.020 57.165 107.970 ;
        RECT 57.465 105.070 57.865 105.570 ;
        RECT 58.165 105.070 58.565 105.570 ;
        RECT 62.115 93.820 63.165 100.370 ;
        RECT 51.990 76.100 53.090 85.700 ;
        RECT 57.390 77.000 59.140 89.400 ;
      LAYER via2 ;
        RECT 32.675 136.630 32.955 136.910 ;
        RECT 33.425 136.630 33.705 136.910 ;
        RECT 32.675 133.930 32.955 134.210 ;
        RECT 33.425 133.930 33.705 134.210 ;
        RECT 32.675 131.230 32.955 131.510 ;
        RECT 33.425 131.230 33.705 131.510 ;
        RECT 0.500 123.930 0.780 124.210 ;
        RECT 0.500 123.530 0.780 123.810 ;
        RECT 1.750 123.930 2.030 124.210 ;
        RECT 1.750 123.530 2.030 123.810 ;
        RECT 39.125 128.230 39.405 128.510 ;
        RECT 39.675 128.230 39.955 128.510 ;
        RECT 39.125 125.180 39.405 125.460 ;
        RECT 39.675 125.180 39.955 125.460 ;
        RECT 45.125 136.630 45.405 136.910 ;
        RECT 45.875 136.630 46.155 136.910 ;
        RECT 45.125 133.930 45.405 134.210 ;
        RECT 45.875 133.930 46.155 134.210 ;
        RECT 45.125 131.230 45.405 131.510 ;
        RECT 45.875 131.230 46.155 131.510 ;
        RECT 51.175 128.230 51.455 128.510 ;
        RECT 51.725 128.230 52.005 128.510 ;
        RECT 51.175 125.280 51.455 125.560 ;
        RECT 51.725 125.280 52.005 125.560 ;
        RECT 57.525 136.630 57.805 136.910 ;
        RECT 58.275 136.630 58.555 136.910 ;
        RECT 57.525 133.930 57.805 134.210 ;
        RECT 58.275 133.930 58.555 134.210 ;
        RECT 57.575 131.230 57.855 131.510 ;
        RECT 58.275 131.230 58.555 131.510 ;
        RECT 51.175 122.380 51.455 122.660 ;
        RECT 51.725 122.380 52.005 122.660 ;
        RECT 63.475 128.180 63.755 128.460 ;
        RECT 64.025 128.180 64.305 128.460 ;
        RECT 63.475 125.280 63.755 125.560 ;
        RECT 64.025 125.280 64.305 125.560 ;
        RECT 63.475 122.380 63.755 122.660 ;
        RECT 64.025 122.380 64.305 122.660 ;
        RECT 98.000 124.780 98.280 125.060 ;
        RECT 98.000 124.380 98.280 124.660 ;
        RECT 99.300 124.780 99.580 125.060 ;
        RECT 99.300 124.380 99.580 124.660 ;
        RECT 39.125 108.880 39.405 109.160 ;
        RECT 39.675 108.880 39.955 109.160 ;
        RECT 51.175 108.880 51.455 109.160 ;
        RECT 51.725 108.880 52.005 109.160 ;
        RECT 63.475 108.930 63.755 109.210 ;
        RECT 64.025 108.930 64.305 109.210 ;
        RECT 32.675 105.080 32.955 105.360 ;
        RECT 33.425 105.080 33.705 105.360 ;
        RECT 45.125 105.180 45.405 105.460 ;
        RECT 45.875 105.180 46.155 105.460 ;
        RECT 57.525 105.180 57.805 105.460 ;
        RECT 58.225 105.180 58.505 105.460 ;
      LAYER met3 ;
        RECT 0.215 123.420 2.415 158.770 ;
        RECT 13.015 140.770 30.015 158.265 ;
        RECT 32.015 140.770 49.015 158.265 ;
        RECT 51.015 140.770 68.015 158.265 ;
        RECT 70.015 140.770 87.015 158.265 ;
        RECT 32.515 136.470 33.865 137.070 ;
        RECT 44.965 136.470 46.315 137.020 ;
        RECT 57.365 136.470 58.715 137.070 ;
        RECT 32.515 133.770 33.865 134.370 ;
        RECT 44.965 133.770 46.315 134.320 ;
        RECT 57.365 133.770 58.715 134.370 ;
        RECT 32.515 131.070 33.865 131.720 ;
        RECT 44.965 131.070 46.315 131.620 ;
        RECT 57.365 131.070 58.715 131.720 ;
        RECT 38.965 128.020 40.115 128.670 ;
        RECT 51.015 128.120 52.165 128.670 ;
        RECT 63.315 128.020 64.465 128.570 ;
        RECT 38.965 125.070 40.115 125.570 ;
        RECT 51.015 125.120 52.165 125.670 ;
        RECT 63.315 125.120 64.465 125.670 ;
        RECT 97.715 124.320 99.865 158.820 ;
        RECT 38.965 122.220 40.115 122.820 ;
        RECT 51.015 122.220 52.165 122.770 ;
        RECT 63.315 122.220 64.465 122.770 ;
        RECT 38.965 108.770 40.115 109.270 ;
        RECT 51.015 108.770 52.165 109.320 ;
        RECT 63.315 108.820 64.465 109.320 ;
        RECT 32.515 104.870 33.865 105.520 ;
        RECT 44.965 105.020 46.315 105.570 ;
        RECT 57.365 105.020 58.715 105.570 ;
      LAYER via3 ;
        RECT 0.455 158.035 0.775 158.355 ;
        RECT 1.755 158.035 2.075 158.355 ;
        RECT 13.155 157.845 13.475 158.165 ;
        RECT 13.555 157.845 13.875 158.165 ;
        RECT 13.955 157.845 14.275 158.165 ;
        RECT 14.355 157.845 14.675 158.165 ;
        RECT 14.755 157.845 15.075 158.165 ;
        RECT 15.155 157.845 15.475 158.165 ;
        RECT 15.555 157.845 15.875 158.165 ;
        RECT 15.955 157.845 16.275 158.165 ;
        RECT 16.355 157.845 16.675 158.165 ;
        RECT 16.755 157.845 17.075 158.165 ;
        RECT 17.155 157.845 17.475 158.165 ;
        RECT 17.555 157.845 17.875 158.165 ;
        RECT 17.955 157.845 18.275 158.165 ;
        RECT 18.355 157.845 18.675 158.165 ;
        RECT 18.755 157.845 19.075 158.165 ;
        RECT 19.155 157.845 19.475 158.165 ;
        RECT 19.555 157.845 19.875 158.165 ;
        RECT 19.955 157.845 20.275 158.165 ;
        RECT 20.355 157.845 20.675 158.165 ;
        RECT 20.755 157.845 21.075 158.165 ;
        RECT 21.155 157.845 21.475 158.165 ;
        RECT 21.555 157.845 21.875 158.165 ;
        RECT 21.955 157.845 22.275 158.165 ;
        RECT 22.355 157.845 22.675 158.165 ;
        RECT 22.755 157.845 23.075 158.165 ;
        RECT 23.155 157.845 23.475 158.165 ;
        RECT 23.555 157.845 23.875 158.165 ;
        RECT 23.955 157.845 24.275 158.165 ;
        RECT 24.355 157.845 24.675 158.165 ;
        RECT 24.755 157.845 25.075 158.165 ;
        RECT 25.155 157.845 25.475 158.165 ;
        RECT 25.555 157.845 25.875 158.165 ;
        RECT 25.955 157.845 26.275 158.165 ;
        RECT 26.355 157.845 26.675 158.165 ;
        RECT 26.755 157.845 27.075 158.165 ;
        RECT 27.155 157.845 27.475 158.165 ;
        RECT 27.555 157.845 27.875 158.165 ;
        RECT 27.955 157.845 28.275 158.165 ;
        RECT 28.355 157.845 28.675 158.165 ;
        RECT 28.755 157.845 29.075 158.165 ;
        RECT 29.155 157.845 29.475 158.165 ;
        RECT 29.555 157.845 29.875 158.165 ;
        RECT 32.155 157.845 32.475 158.165 ;
        RECT 32.555 157.845 32.875 158.165 ;
        RECT 32.955 157.845 33.275 158.165 ;
        RECT 33.355 157.845 33.675 158.165 ;
        RECT 33.755 157.845 34.075 158.165 ;
        RECT 34.155 157.845 34.475 158.165 ;
        RECT 34.555 157.845 34.875 158.165 ;
        RECT 34.955 157.845 35.275 158.165 ;
        RECT 35.355 157.845 35.675 158.165 ;
        RECT 35.755 157.845 36.075 158.165 ;
        RECT 36.155 157.845 36.475 158.165 ;
        RECT 36.555 157.845 36.875 158.165 ;
        RECT 36.955 157.845 37.275 158.165 ;
        RECT 37.355 157.845 37.675 158.165 ;
        RECT 37.755 157.845 38.075 158.165 ;
        RECT 38.155 157.845 38.475 158.165 ;
        RECT 38.555 157.845 38.875 158.165 ;
        RECT 38.955 157.845 39.275 158.165 ;
        RECT 39.355 157.845 39.675 158.165 ;
        RECT 39.755 157.845 40.075 158.165 ;
        RECT 40.155 157.845 40.475 158.165 ;
        RECT 40.555 157.845 40.875 158.165 ;
        RECT 40.955 157.845 41.275 158.165 ;
        RECT 41.355 157.845 41.675 158.165 ;
        RECT 41.755 157.845 42.075 158.165 ;
        RECT 42.155 157.845 42.475 158.165 ;
        RECT 42.555 157.845 42.875 158.165 ;
        RECT 42.955 157.845 43.275 158.165 ;
        RECT 43.355 157.845 43.675 158.165 ;
        RECT 43.755 157.845 44.075 158.165 ;
        RECT 44.155 157.845 44.475 158.165 ;
        RECT 44.555 157.845 44.875 158.165 ;
        RECT 44.955 157.845 45.275 158.165 ;
        RECT 45.355 157.845 45.675 158.165 ;
        RECT 45.755 157.845 46.075 158.165 ;
        RECT 46.155 157.845 46.475 158.165 ;
        RECT 46.555 157.845 46.875 158.165 ;
        RECT 46.955 157.845 47.275 158.165 ;
        RECT 47.355 157.845 47.675 158.165 ;
        RECT 47.755 157.845 48.075 158.165 ;
        RECT 48.155 157.845 48.475 158.165 ;
        RECT 48.555 157.845 48.875 158.165 ;
        RECT 51.155 157.845 51.475 158.165 ;
        RECT 51.555 157.845 51.875 158.165 ;
        RECT 51.955 157.845 52.275 158.165 ;
        RECT 52.355 157.845 52.675 158.165 ;
        RECT 52.755 157.845 53.075 158.165 ;
        RECT 53.155 157.845 53.475 158.165 ;
        RECT 53.555 157.845 53.875 158.165 ;
        RECT 53.955 157.845 54.275 158.165 ;
        RECT 54.355 157.845 54.675 158.165 ;
        RECT 54.755 157.845 55.075 158.165 ;
        RECT 55.155 157.845 55.475 158.165 ;
        RECT 55.555 157.845 55.875 158.165 ;
        RECT 55.955 157.845 56.275 158.165 ;
        RECT 56.355 157.845 56.675 158.165 ;
        RECT 56.755 157.845 57.075 158.165 ;
        RECT 57.155 157.845 57.475 158.165 ;
        RECT 57.555 157.845 57.875 158.165 ;
        RECT 57.955 157.845 58.275 158.165 ;
        RECT 58.355 157.845 58.675 158.165 ;
        RECT 58.755 157.845 59.075 158.165 ;
        RECT 59.155 157.845 59.475 158.165 ;
        RECT 59.555 157.845 59.875 158.165 ;
        RECT 59.955 157.845 60.275 158.165 ;
        RECT 60.355 157.845 60.675 158.165 ;
        RECT 60.755 157.845 61.075 158.165 ;
        RECT 61.155 157.845 61.475 158.165 ;
        RECT 61.555 157.845 61.875 158.165 ;
        RECT 61.955 157.845 62.275 158.165 ;
        RECT 62.355 157.845 62.675 158.165 ;
        RECT 62.755 157.845 63.075 158.165 ;
        RECT 63.155 157.845 63.475 158.165 ;
        RECT 63.555 157.845 63.875 158.165 ;
        RECT 63.955 157.845 64.275 158.165 ;
        RECT 64.355 157.845 64.675 158.165 ;
        RECT 64.755 157.845 65.075 158.165 ;
        RECT 65.155 157.845 65.475 158.165 ;
        RECT 65.555 157.845 65.875 158.165 ;
        RECT 65.955 157.845 66.275 158.165 ;
        RECT 66.355 157.845 66.675 158.165 ;
        RECT 66.755 157.845 67.075 158.165 ;
        RECT 67.155 157.845 67.475 158.165 ;
        RECT 67.555 157.845 67.875 158.165 ;
        RECT 70.155 157.845 70.475 158.165 ;
        RECT 70.555 157.845 70.875 158.165 ;
        RECT 70.955 157.845 71.275 158.165 ;
        RECT 71.355 157.845 71.675 158.165 ;
        RECT 71.755 157.845 72.075 158.165 ;
        RECT 72.155 157.845 72.475 158.165 ;
        RECT 72.555 157.845 72.875 158.165 ;
        RECT 72.955 157.845 73.275 158.165 ;
        RECT 73.355 157.845 73.675 158.165 ;
        RECT 73.755 157.845 74.075 158.165 ;
        RECT 74.155 157.845 74.475 158.165 ;
        RECT 74.555 157.845 74.875 158.165 ;
        RECT 74.955 157.845 75.275 158.165 ;
        RECT 75.355 157.845 75.675 158.165 ;
        RECT 75.755 157.845 76.075 158.165 ;
        RECT 76.155 157.845 76.475 158.165 ;
        RECT 76.555 157.845 76.875 158.165 ;
        RECT 76.955 157.845 77.275 158.165 ;
        RECT 77.355 157.845 77.675 158.165 ;
        RECT 77.755 157.845 78.075 158.165 ;
        RECT 78.155 157.845 78.475 158.165 ;
        RECT 78.555 157.845 78.875 158.165 ;
        RECT 78.955 157.845 79.275 158.165 ;
        RECT 79.355 157.845 79.675 158.165 ;
        RECT 79.755 157.845 80.075 158.165 ;
        RECT 80.155 157.845 80.475 158.165 ;
        RECT 80.555 157.845 80.875 158.165 ;
        RECT 80.955 157.845 81.275 158.165 ;
        RECT 81.355 157.845 81.675 158.165 ;
        RECT 81.755 157.845 82.075 158.165 ;
        RECT 82.155 157.845 82.475 158.165 ;
        RECT 82.555 157.845 82.875 158.165 ;
        RECT 82.955 157.845 83.275 158.165 ;
        RECT 83.355 157.845 83.675 158.165 ;
        RECT 83.755 157.845 84.075 158.165 ;
        RECT 84.155 157.845 84.475 158.165 ;
        RECT 84.555 157.845 84.875 158.165 ;
        RECT 84.955 157.845 85.275 158.165 ;
        RECT 85.355 157.845 85.675 158.165 ;
        RECT 85.755 157.845 86.075 158.165 ;
        RECT 86.155 157.845 86.475 158.165 ;
        RECT 86.555 157.845 86.875 158.165 ;
        RECT 97.930 158.035 98.250 158.355 ;
        RECT 99.230 158.035 99.550 158.355 ;
        RECT 32.655 136.610 32.975 136.930 ;
        RECT 33.405 136.610 33.725 136.930 ;
        RECT 45.105 136.610 45.425 136.930 ;
        RECT 45.855 136.610 46.175 136.930 ;
        RECT 57.505 136.610 57.825 136.930 ;
        RECT 58.255 136.610 58.575 136.930 ;
        RECT 32.655 133.910 32.975 134.230 ;
        RECT 33.405 133.910 33.725 134.230 ;
        RECT 45.105 133.910 45.425 134.230 ;
        RECT 45.855 133.910 46.175 134.230 ;
        RECT 57.505 133.910 57.825 134.230 ;
        RECT 58.255 133.910 58.575 134.230 ;
        RECT 32.655 131.210 32.975 131.530 ;
        RECT 33.405 131.210 33.725 131.530 ;
        RECT 45.105 131.210 45.425 131.530 ;
        RECT 45.855 131.210 46.175 131.530 ;
        RECT 57.555 131.210 57.875 131.530 ;
        RECT 58.255 131.210 58.575 131.530 ;
        RECT 39.105 128.210 39.425 128.530 ;
        RECT 39.655 128.210 39.975 128.530 ;
        RECT 51.155 128.210 51.475 128.530 ;
        RECT 51.705 128.210 52.025 128.530 ;
        RECT 63.455 128.160 63.775 128.480 ;
        RECT 64.005 128.160 64.325 128.480 ;
        RECT 39.105 125.160 39.425 125.480 ;
        RECT 39.655 125.160 39.975 125.480 ;
        RECT 51.155 125.260 51.475 125.580 ;
        RECT 51.705 125.260 52.025 125.580 ;
        RECT 63.455 125.260 63.775 125.580 ;
        RECT 64.005 125.260 64.325 125.580 ;
        RECT 39.105 122.360 39.425 122.680 ;
        RECT 39.655 122.360 39.975 122.680 ;
        RECT 51.155 122.360 51.475 122.680 ;
        RECT 51.705 122.360 52.025 122.680 ;
        RECT 63.455 122.360 63.775 122.680 ;
        RECT 64.005 122.360 64.325 122.680 ;
        RECT 39.105 108.860 39.425 109.180 ;
        RECT 39.655 108.860 39.975 109.180 ;
        RECT 51.155 108.860 51.475 109.180 ;
        RECT 51.705 108.860 52.025 109.180 ;
        RECT 63.455 108.910 63.775 109.230 ;
        RECT 64.005 108.910 64.325 109.230 ;
        RECT 32.655 105.060 32.975 105.380 ;
        RECT 33.405 105.060 33.725 105.380 ;
        RECT 45.105 105.160 45.425 105.480 ;
        RECT 45.855 105.160 46.175 105.480 ;
        RECT 57.505 105.160 57.825 105.480 ;
        RECT 58.205 105.160 58.525 105.480 ;
      LAYER met4 ;
        RECT 0.165 157.620 99.865 158.820 ;
        RECT 32.515 104.870 33.865 137.620 ;
        RECT 38.965 108.720 40.115 128.670 ;
        RECT 44.965 105.020 46.315 137.870 ;
        RECT 51.015 108.720 52.165 128.670 ;
        RECT 57.365 105.020 58.715 137.920 ;
        RECT 63.315 108.770 64.465 128.720 ;
  END
END MULT_Amp
MACRO MULT_AMPLIFIER
  CLASS BLOCK ;
  FOREIGN MULT_AMPLIFIER ;
  ORIGIN -2326.970 -3148.500 ;
  SIZE 597.030 BY 375.500 ;
  PIN io_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 17.500000 ;
    PORT
      LAYER li1 ;
        RECT 2710.175 3420.110 2710.345 3420.610 ;
        RECT 2715.725 3420.110 2715.895 3420.610 ;
        RECT 2716.265 3420.110 2716.435 3420.610 ;
        RECT 2721.815 3420.110 2721.985 3420.610 ;
        RECT 2722.355 3420.110 2722.525 3420.610 ;
        RECT 2727.905 3420.110 2728.075 3420.610 ;
        RECT 2728.445 3420.110 2728.615 3420.610 ;
        RECT 2733.995 3420.110 2734.165 3420.610 ;
        RECT 2734.535 3420.110 2734.705 3420.610 ;
        RECT 2740.085 3420.110 2740.255 3420.610 ;
        RECT 2740.625 3420.110 2740.795 3420.610 ;
        RECT 2746.175 3420.110 2746.345 3420.610 ;
        RECT 2746.715 3420.110 2746.885 3420.610 ;
        RECT 2752.265 3420.110 2752.435 3420.610 ;
      LAYER mcon ;
        RECT 2710.175 3420.275 2710.345 3420.445 ;
        RECT 2715.725 3420.275 2715.895 3420.445 ;
        RECT 2716.265 3420.275 2716.435 3420.445 ;
        RECT 2721.815 3420.275 2721.985 3420.445 ;
        RECT 2722.355 3420.275 2722.525 3420.445 ;
        RECT 2727.905 3420.275 2728.075 3420.445 ;
        RECT 2728.445 3420.275 2728.615 3420.445 ;
        RECT 2733.995 3420.275 2734.165 3420.445 ;
        RECT 2734.535 3420.275 2734.705 3420.445 ;
        RECT 2740.085 3420.275 2740.255 3420.445 ;
        RECT 2740.625 3420.275 2740.795 3420.445 ;
        RECT 2746.175 3420.275 2746.345 3420.445 ;
        RECT 2746.715 3420.275 2746.885 3420.445 ;
        RECT 2752.265 3420.275 2752.435 3420.445 ;
      LAYER met1 ;
        RECT 2752.300 3420.590 2810.000 3420.700 ;
        RECT 2710.145 3420.480 2710.375 3420.590 ;
        RECT 2715.695 3420.480 2715.925 3420.590 ;
        RECT 2716.235 3420.480 2716.465 3420.590 ;
        RECT 2721.785 3420.530 2722.015 3420.590 ;
        RECT 2722.325 3420.530 2722.555 3420.590 ;
        RECT 2721.785 3420.480 2722.555 3420.530 ;
        RECT 2727.875 3420.530 2728.105 3420.590 ;
        RECT 2728.415 3420.530 2728.645 3420.590 ;
        RECT 2727.875 3420.480 2728.645 3420.530 ;
        RECT 2733.965 3420.530 2734.195 3420.590 ;
        RECT 2734.505 3420.530 2734.735 3420.590 ;
        RECT 2733.965 3420.480 2734.735 3420.530 ;
        RECT 2740.055 3420.530 2740.285 3420.590 ;
        RECT 2740.595 3420.530 2740.825 3420.590 ;
        RECT 2746.145 3420.530 2746.375 3420.590 ;
        RECT 2746.685 3420.530 2746.915 3420.590 ;
        RECT 2740.055 3420.480 2740.835 3420.530 ;
        RECT 2746.135 3420.480 2746.915 3420.530 ;
        RECT 2752.235 3420.480 2810.000 3420.590 ;
        RECT 2710.145 3420.280 2810.000 3420.480 ;
        RECT 2710.145 3420.130 2710.375 3420.280 ;
        RECT 2715.695 3420.130 2715.925 3420.280 ;
        RECT 2716.235 3420.130 2716.465 3420.280 ;
        RECT 2721.785 3420.180 2722.555 3420.280 ;
        RECT 2721.785 3420.130 2722.015 3420.180 ;
        RECT 2722.325 3420.130 2722.555 3420.180 ;
        RECT 2727.875 3420.180 2728.645 3420.280 ;
        RECT 2727.875 3420.130 2728.105 3420.180 ;
        RECT 2728.415 3420.130 2728.645 3420.180 ;
        RECT 2733.965 3420.180 2734.735 3420.280 ;
        RECT 2733.965 3420.130 2734.195 3420.180 ;
        RECT 2734.505 3420.130 2734.735 3420.180 ;
        RECT 2740.055 3420.180 2740.835 3420.280 ;
        RECT 2746.135 3420.180 2746.915 3420.280 ;
        RECT 2740.055 3420.130 2740.285 3420.180 ;
        RECT 2740.595 3420.130 2740.825 3420.180 ;
        RECT 2746.145 3420.130 2746.375 3420.180 ;
        RECT 2746.685 3420.130 2746.915 3420.180 ;
        RECT 2752.235 3420.130 2810.000 3420.280 ;
        RECT 2752.300 3420.000 2810.000 3420.130 ;
        RECT 2753.200 3418.000 2810.000 3420.000 ;
        RECT 2800.600 3389.500 2810.000 3418.000 ;
      LAYER via ;
        RECT 2805.000 3418.500 2806.500 3420.000 ;
        RECT 2808.000 3418.500 2809.500 3420.000 ;
        RECT 2805.000 3416.000 2806.500 3417.500 ;
        RECT 2808.000 3416.000 2809.500 3417.500 ;
        RECT 2805.000 3413.500 2806.500 3415.000 ;
        RECT 2808.000 3413.500 2809.500 3415.000 ;
        RECT 2805.000 3411.000 2806.500 3412.500 ;
        RECT 2808.000 3411.000 2809.500 3412.500 ;
        RECT 2805.000 3408.500 2806.500 3410.000 ;
        RECT 2808.000 3408.500 2809.500 3410.000 ;
        RECT 2805.000 3406.000 2806.500 3407.500 ;
        RECT 2808.000 3406.000 2809.500 3407.500 ;
        RECT 2805.000 3403.500 2806.500 3405.000 ;
        RECT 2808.000 3403.500 2809.500 3405.000 ;
        RECT 2805.000 3401.000 2806.500 3402.500 ;
        RECT 2808.000 3401.000 2809.500 3402.500 ;
        RECT 2805.000 3398.500 2806.500 3400.000 ;
        RECT 2808.000 3398.500 2809.500 3400.000 ;
        RECT 2805.000 3396.000 2806.500 3397.500 ;
        RECT 2808.000 3396.000 2809.500 3397.500 ;
        RECT 2805.000 3393.500 2806.500 3395.000 ;
        RECT 2808.000 3393.500 2809.500 3395.000 ;
        RECT 2805.000 3391.000 2806.500 3392.500 ;
        RECT 2808.000 3391.000 2809.500 3392.500 ;
      LAYER met2 ;
        RECT 2805.000 3418.450 2806.500 3420.050 ;
        RECT 2808.000 3418.450 2809.500 3420.050 ;
        RECT 2805.000 3415.950 2806.500 3417.550 ;
        RECT 2808.000 3415.950 2809.500 3417.550 ;
        RECT 2805.000 3413.450 2806.500 3415.050 ;
        RECT 2808.000 3413.450 2809.500 3415.050 ;
        RECT 2805.000 3410.950 2806.500 3412.550 ;
        RECT 2808.000 3410.950 2809.500 3412.550 ;
        RECT 2805.000 3408.450 2806.500 3410.050 ;
        RECT 2808.000 3408.450 2809.500 3410.050 ;
        RECT 2805.000 3405.950 2806.500 3407.550 ;
        RECT 2808.000 3405.950 2809.500 3407.550 ;
        RECT 2805.000 3403.450 2806.500 3405.050 ;
        RECT 2808.000 3403.450 2809.500 3405.050 ;
        RECT 2805.000 3400.950 2806.500 3402.550 ;
        RECT 2808.000 3400.950 2809.500 3402.550 ;
        RECT 2805.000 3398.450 2806.500 3400.050 ;
        RECT 2808.000 3398.450 2809.500 3400.050 ;
        RECT 2805.000 3395.950 2806.500 3397.550 ;
        RECT 2808.000 3395.950 2809.500 3397.550 ;
        RECT 2805.000 3393.450 2806.500 3395.050 ;
        RECT 2808.000 3393.450 2809.500 3395.050 ;
        RECT 2805.000 3390.950 2806.500 3392.550 ;
        RECT 2808.000 3390.950 2809.500 3392.550 ;
      LAYER via2 ;
        RECT 2805.000 3418.500 2806.500 3420.000 ;
        RECT 2808.000 3418.500 2809.500 3420.000 ;
        RECT 2805.000 3416.000 2806.500 3417.500 ;
        RECT 2808.000 3416.000 2809.500 3417.500 ;
        RECT 2805.000 3413.500 2806.500 3415.000 ;
        RECT 2808.000 3413.500 2809.500 3415.000 ;
        RECT 2805.000 3411.000 2806.500 3412.500 ;
        RECT 2808.000 3411.000 2809.500 3412.500 ;
        RECT 2805.000 3408.500 2806.500 3410.000 ;
        RECT 2808.000 3408.500 2809.500 3410.000 ;
        RECT 2805.000 3406.000 2806.500 3407.500 ;
        RECT 2808.000 3406.000 2809.500 3407.500 ;
        RECT 2805.000 3403.500 2806.500 3405.000 ;
        RECT 2808.000 3403.500 2809.500 3405.000 ;
        RECT 2805.000 3401.000 2806.500 3402.500 ;
        RECT 2808.000 3401.000 2809.500 3402.500 ;
        RECT 2805.000 3398.500 2806.500 3400.000 ;
        RECT 2808.000 3398.500 2809.500 3400.000 ;
        RECT 2805.000 3396.000 2806.500 3397.500 ;
        RECT 2808.000 3396.000 2809.500 3397.500 ;
        RECT 2805.000 3393.500 2806.500 3395.000 ;
        RECT 2808.000 3393.500 2809.500 3395.000 ;
        RECT 2805.000 3391.000 2806.500 3392.500 ;
        RECT 2808.000 3391.000 2809.500 3392.500 ;
      LAYER met3 ;
        RECT 2804.500 3415.500 2810.000 3420.700 ;
        RECT 2804.500 3414.920 2920.000 3415.500 ;
        RECT 2804.500 3389.920 2924.000 3414.920 ;
        RECT 2804.500 3389.500 2920.000 3389.920 ;
    END
  END io_analog[0]
  PIN io_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 17.500000 ;
    PORT
      LAYER li1 ;
        RECT 2710.175 3422.610 2710.345 3423.110 ;
        RECT 2715.725 3422.610 2715.895 3423.110 ;
        RECT 2716.265 3422.610 2716.435 3423.110 ;
        RECT 2721.815 3422.610 2721.985 3423.110 ;
        RECT 2722.355 3422.610 2722.525 3423.110 ;
        RECT 2727.905 3422.610 2728.075 3423.110 ;
        RECT 2728.445 3422.610 2728.615 3423.110 ;
        RECT 2733.995 3422.610 2734.165 3423.110 ;
        RECT 2734.535 3422.610 2734.705 3423.110 ;
        RECT 2740.085 3422.610 2740.255 3423.110 ;
        RECT 2740.625 3422.610 2740.795 3423.110 ;
        RECT 2746.175 3422.610 2746.345 3423.110 ;
        RECT 2746.715 3422.610 2746.885 3423.110 ;
        RECT 2752.265 3422.610 2752.435 3423.110 ;
      LAYER mcon ;
        RECT 2710.175 3422.775 2710.345 3422.945 ;
        RECT 2715.725 3422.775 2715.895 3422.945 ;
        RECT 2716.265 3422.775 2716.435 3422.945 ;
        RECT 2721.815 3422.775 2721.985 3422.945 ;
        RECT 2722.355 3422.775 2722.525 3422.945 ;
        RECT 2727.905 3422.775 2728.075 3422.945 ;
        RECT 2728.445 3422.775 2728.615 3422.945 ;
        RECT 2733.995 3422.775 2734.165 3422.945 ;
        RECT 2734.535 3422.775 2734.705 3422.945 ;
        RECT 2740.085 3422.775 2740.255 3422.945 ;
        RECT 2740.625 3422.775 2740.795 3422.945 ;
        RECT 2746.175 3422.775 2746.345 3422.945 ;
        RECT 2746.715 3422.775 2746.885 3422.945 ;
        RECT 2752.265 3422.775 2752.435 3422.945 ;
      LAYER met1 ;
        RECT 2801.100 3428.300 2858.300 3435.500 ;
        RECT 2801.100 3423.500 2805.400 3428.300 ;
        RECT 2752.500 3423.200 2805.400 3423.500 ;
        RECT 2752.300 3423.090 2805.400 3423.200 ;
        RECT 2710.145 3422.980 2710.375 3423.090 ;
        RECT 2715.695 3422.980 2715.925 3423.090 ;
        RECT 2716.235 3422.980 2716.465 3423.090 ;
        RECT 2721.785 3423.030 2722.015 3423.090 ;
        RECT 2722.325 3423.030 2722.555 3423.090 ;
        RECT 2721.785 3422.980 2722.555 3423.030 ;
        RECT 2727.875 3423.030 2728.105 3423.090 ;
        RECT 2728.415 3423.030 2728.645 3423.090 ;
        RECT 2727.875 3422.980 2728.645 3423.030 ;
        RECT 2733.965 3423.030 2734.195 3423.090 ;
        RECT 2734.505 3423.030 2734.735 3423.090 ;
        RECT 2733.965 3422.980 2734.735 3423.030 ;
        RECT 2740.055 3423.030 2740.285 3423.090 ;
        RECT 2740.595 3423.030 2740.825 3423.090 ;
        RECT 2746.145 3423.030 2746.375 3423.090 ;
        RECT 2746.685 3423.030 2746.915 3423.090 ;
        RECT 2740.055 3422.980 2740.835 3423.030 ;
        RECT 2746.135 3422.980 2746.915 3423.030 ;
        RECT 2752.235 3422.980 2805.400 3423.090 ;
        RECT 2710.135 3422.780 2805.400 3422.980 ;
        RECT 2710.145 3422.630 2710.375 3422.780 ;
        RECT 2715.695 3422.630 2715.925 3422.780 ;
        RECT 2716.235 3422.630 2716.465 3422.780 ;
        RECT 2721.785 3422.680 2722.555 3422.780 ;
        RECT 2721.785 3422.630 2722.015 3422.680 ;
        RECT 2722.325 3422.630 2722.555 3422.680 ;
        RECT 2727.875 3422.680 2728.645 3422.780 ;
        RECT 2727.875 3422.630 2728.105 3422.680 ;
        RECT 2728.415 3422.630 2728.645 3422.680 ;
        RECT 2733.965 3422.680 2734.735 3422.780 ;
        RECT 2733.965 3422.630 2734.195 3422.680 ;
        RECT 2734.505 3422.630 2734.735 3422.680 ;
        RECT 2740.055 3422.680 2740.835 3422.780 ;
        RECT 2746.135 3422.680 2746.915 3422.780 ;
        RECT 2740.055 3422.630 2740.285 3422.680 ;
        RECT 2740.595 3422.630 2740.825 3422.680 ;
        RECT 2746.145 3422.630 2746.375 3422.680 ;
        RECT 2746.685 3422.630 2746.915 3422.680 ;
        RECT 2752.235 3422.630 2805.400 3422.780 ;
        RECT 2752.300 3422.500 2805.400 3422.630 ;
        RECT 2752.500 3421.500 2805.400 3422.500 ;
      LAYER via ;
        RECT 2832.500 3433.000 2834.500 3435.000 ;
        RECT 2836.500 3433.000 2838.500 3435.000 ;
        RECT 2840.500 3433.000 2842.500 3435.000 ;
        RECT 2844.500 3433.000 2846.500 3435.000 ;
        RECT 2848.500 3433.000 2850.500 3435.000 ;
        RECT 2852.500 3433.000 2854.500 3435.000 ;
        RECT 2832.500 3429.000 2834.500 3431.000 ;
        RECT 2836.500 3429.000 2838.500 3431.000 ;
        RECT 2840.500 3429.000 2842.500 3431.000 ;
        RECT 2844.500 3429.000 2846.500 3431.000 ;
        RECT 2848.500 3429.000 2850.500 3431.000 ;
        RECT 2852.500 3429.000 2854.500 3431.000 ;
      LAYER met2 ;
        RECT 2832.500 3432.950 2834.500 3435.050 ;
        RECT 2836.500 3432.950 2838.500 3435.050 ;
        RECT 2840.500 3432.950 2842.500 3435.050 ;
        RECT 2844.500 3432.950 2846.500 3435.050 ;
        RECT 2848.500 3432.950 2850.500 3435.050 ;
        RECT 2852.500 3432.950 2854.500 3435.050 ;
        RECT 2832.500 3428.950 2834.500 3431.050 ;
        RECT 2836.500 3428.950 2838.500 3431.050 ;
        RECT 2840.500 3428.950 2842.500 3431.050 ;
        RECT 2844.500 3428.950 2846.500 3431.050 ;
        RECT 2848.500 3428.950 2850.500 3431.050 ;
        RECT 2852.500 3428.950 2854.500 3431.050 ;
      LAYER via2 ;
        RECT 2832.500 3433.000 2834.500 3435.000 ;
        RECT 2836.500 3433.000 2838.500 3435.000 ;
        RECT 2840.500 3433.000 2842.500 3435.000 ;
        RECT 2844.500 3433.000 2846.500 3435.000 ;
        RECT 2848.500 3433.000 2850.500 3435.000 ;
        RECT 2852.500 3433.000 2854.500 3435.000 ;
        RECT 2832.500 3429.000 2834.500 3431.000 ;
        RECT 2836.500 3429.000 2838.500 3431.000 ;
        RECT 2840.500 3429.000 2842.500 3431.000 ;
        RECT 2844.500 3429.000 2846.500 3431.000 ;
        RECT 2848.500 3429.000 2850.500 3431.000 ;
        RECT 2852.500 3429.000 2854.500 3431.000 ;
      LAYER met3 ;
        RECT 2832.970 3519.800 2857.970 3524.000 ;
        RECT 2831.500 3428.300 2858.300 3519.800 ;
    END
  END io_analog[1]
  PIN io_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 75.400002 ;
    PORT
      LAYER li1 ;
        RECT 2700.860 3434.380 2705.900 3434.550 ;
        RECT 2707.040 3434.380 2712.080 3434.550 ;
        RECT 2713.220 3434.380 2718.260 3434.550 ;
        RECT 2719.400 3434.380 2724.440 3434.550 ;
        RECT 2725.580 3434.380 2730.620 3434.550 ;
        RECT 2731.760 3434.380 2736.800 3434.550 ;
        RECT 2737.940 3434.380 2742.980 3434.550 ;
        RECT 2744.120 3434.380 2749.160 3434.550 ;
        RECT 2750.300 3434.380 2755.340 3434.550 ;
        RECT 2756.480 3434.380 2761.520 3434.550 ;
        RECT 2700.860 3431.680 2705.900 3431.850 ;
        RECT 2707.040 3431.680 2712.080 3431.850 ;
        RECT 2713.220 3431.680 2718.260 3431.850 ;
        RECT 2719.400 3431.680 2724.440 3431.850 ;
        RECT 2725.580 3431.680 2730.620 3431.850 ;
        RECT 2731.760 3431.680 2736.800 3431.850 ;
        RECT 2737.940 3431.680 2742.980 3431.850 ;
        RECT 2744.120 3431.680 2749.160 3431.850 ;
        RECT 2750.300 3431.680 2755.340 3431.850 ;
        RECT 2756.480 3431.680 2761.520 3431.850 ;
        RECT 2700.860 3428.980 2705.900 3429.150 ;
        RECT 2707.040 3428.980 2712.080 3429.150 ;
        RECT 2713.220 3428.980 2718.260 3429.150 ;
        RECT 2719.400 3428.980 2724.440 3429.150 ;
        RECT 2725.580 3428.980 2730.620 3429.150 ;
        RECT 2731.760 3428.980 2736.800 3429.150 ;
        RECT 2737.940 3428.980 2742.980 3429.150 ;
        RECT 2744.120 3428.980 2749.160 3429.150 ;
        RECT 2750.300 3428.980 2755.340 3429.150 ;
        RECT 2756.480 3428.980 2761.520 3429.150 ;
        RECT 2700.860 3426.280 2705.900 3426.450 ;
        RECT 2707.040 3426.280 2712.080 3426.450 ;
        RECT 2713.220 3426.280 2718.260 3426.450 ;
        RECT 2719.400 3426.280 2724.440 3426.450 ;
        RECT 2725.580 3426.280 2730.620 3426.450 ;
        RECT 2731.760 3426.280 2736.800 3426.450 ;
        RECT 2737.940 3426.280 2742.980 3426.450 ;
        RECT 2744.120 3426.280 2749.160 3426.450 ;
        RECT 2750.300 3426.280 2755.340 3426.450 ;
        RECT 2756.480 3426.280 2761.520 3426.450 ;
        RECT 2713.315 3418.170 2718.355 3418.340 ;
        RECT 2719.405 3418.170 2724.445 3418.340 ;
        RECT 2725.495 3418.170 2730.535 3418.340 ;
        RECT 2731.585 3418.170 2736.625 3418.340 ;
        RECT 2737.675 3418.170 2742.715 3418.340 ;
        RECT 2743.765 3418.170 2748.805 3418.340 ;
        RECT 2713.315 3415.070 2718.355 3415.240 ;
        RECT 2719.405 3415.070 2724.445 3415.240 ;
        RECT 2725.495 3415.070 2730.535 3415.240 ;
        RECT 2731.585 3415.070 2736.625 3415.240 ;
        RECT 2737.675 3415.070 2742.715 3415.240 ;
        RECT 2743.765 3415.070 2748.805 3415.240 ;
      LAYER mcon ;
        RECT 2700.955 3434.380 2701.125 3434.550 ;
        RECT 2701.315 3434.380 2701.485 3434.550 ;
        RECT 2701.675 3434.380 2701.845 3434.550 ;
        RECT 2702.035 3434.380 2702.205 3434.550 ;
        RECT 2702.395 3434.380 2702.565 3434.550 ;
        RECT 2702.755 3434.380 2702.925 3434.550 ;
        RECT 2703.115 3434.380 2703.285 3434.550 ;
        RECT 2703.475 3434.380 2703.645 3434.550 ;
        RECT 2703.835 3434.380 2704.005 3434.550 ;
        RECT 2704.195 3434.380 2704.365 3434.550 ;
        RECT 2704.555 3434.380 2704.725 3434.550 ;
        RECT 2704.915 3434.380 2705.085 3434.550 ;
        RECT 2705.275 3434.380 2705.445 3434.550 ;
        RECT 2705.635 3434.380 2705.805 3434.550 ;
        RECT 2707.135 3434.380 2707.305 3434.550 ;
        RECT 2707.495 3434.380 2707.665 3434.550 ;
        RECT 2707.855 3434.380 2708.025 3434.550 ;
        RECT 2708.215 3434.380 2708.385 3434.550 ;
        RECT 2708.575 3434.380 2708.745 3434.550 ;
        RECT 2708.935 3434.380 2709.105 3434.550 ;
        RECT 2709.295 3434.380 2709.465 3434.550 ;
        RECT 2709.655 3434.380 2709.825 3434.550 ;
        RECT 2710.015 3434.380 2710.185 3434.550 ;
        RECT 2710.375 3434.380 2710.545 3434.550 ;
        RECT 2710.735 3434.380 2710.905 3434.550 ;
        RECT 2711.095 3434.380 2711.265 3434.550 ;
        RECT 2711.455 3434.380 2711.625 3434.550 ;
        RECT 2711.815 3434.380 2711.985 3434.550 ;
        RECT 2713.315 3434.380 2713.485 3434.550 ;
        RECT 2713.675 3434.380 2713.845 3434.550 ;
        RECT 2714.035 3434.380 2714.205 3434.550 ;
        RECT 2714.395 3434.380 2714.565 3434.550 ;
        RECT 2714.755 3434.380 2714.925 3434.550 ;
        RECT 2715.115 3434.380 2715.285 3434.550 ;
        RECT 2715.475 3434.380 2715.645 3434.550 ;
        RECT 2715.835 3434.380 2716.005 3434.550 ;
        RECT 2716.195 3434.380 2716.365 3434.550 ;
        RECT 2716.555 3434.380 2716.725 3434.550 ;
        RECT 2716.915 3434.380 2717.085 3434.550 ;
        RECT 2717.275 3434.380 2717.445 3434.550 ;
        RECT 2717.635 3434.380 2717.805 3434.550 ;
        RECT 2717.995 3434.380 2718.165 3434.550 ;
        RECT 2719.495 3434.380 2719.665 3434.550 ;
        RECT 2719.855 3434.380 2720.025 3434.550 ;
        RECT 2720.215 3434.380 2720.385 3434.550 ;
        RECT 2720.575 3434.380 2720.745 3434.550 ;
        RECT 2720.935 3434.380 2721.105 3434.550 ;
        RECT 2721.295 3434.380 2721.465 3434.550 ;
        RECT 2721.655 3434.380 2721.825 3434.550 ;
        RECT 2722.015 3434.380 2722.185 3434.550 ;
        RECT 2722.375 3434.380 2722.545 3434.550 ;
        RECT 2722.735 3434.380 2722.905 3434.550 ;
        RECT 2723.095 3434.380 2723.265 3434.550 ;
        RECT 2723.455 3434.380 2723.625 3434.550 ;
        RECT 2723.815 3434.380 2723.985 3434.550 ;
        RECT 2724.175 3434.380 2724.345 3434.550 ;
        RECT 2725.675 3434.380 2725.845 3434.550 ;
        RECT 2726.035 3434.380 2726.205 3434.550 ;
        RECT 2726.395 3434.380 2726.565 3434.550 ;
        RECT 2726.755 3434.380 2726.925 3434.550 ;
        RECT 2727.115 3434.380 2727.285 3434.550 ;
        RECT 2727.475 3434.380 2727.645 3434.550 ;
        RECT 2727.835 3434.380 2728.005 3434.550 ;
        RECT 2728.195 3434.380 2728.365 3434.550 ;
        RECT 2728.555 3434.380 2728.725 3434.550 ;
        RECT 2728.915 3434.380 2729.085 3434.550 ;
        RECT 2729.275 3434.380 2729.445 3434.550 ;
        RECT 2729.635 3434.380 2729.805 3434.550 ;
        RECT 2729.995 3434.380 2730.165 3434.550 ;
        RECT 2730.355 3434.380 2730.525 3434.550 ;
        RECT 2731.855 3434.380 2732.025 3434.550 ;
        RECT 2732.215 3434.380 2732.385 3434.550 ;
        RECT 2732.575 3434.380 2732.745 3434.550 ;
        RECT 2732.935 3434.380 2733.105 3434.550 ;
        RECT 2733.295 3434.380 2733.465 3434.550 ;
        RECT 2733.655 3434.380 2733.825 3434.550 ;
        RECT 2734.015 3434.380 2734.185 3434.550 ;
        RECT 2734.375 3434.380 2734.545 3434.550 ;
        RECT 2734.735 3434.380 2734.905 3434.550 ;
        RECT 2735.095 3434.380 2735.265 3434.550 ;
        RECT 2735.455 3434.380 2735.625 3434.550 ;
        RECT 2735.815 3434.380 2735.985 3434.550 ;
        RECT 2736.175 3434.380 2736.345 3434.550 ;
        RECT 2736.535 3434.380 2736.705 3434.550 ;
        RECT 2738.035 3434.380 2738.205 3434.550 ;
        RECT 2738.395 3434.380 2738.565 3434.550 ;
        RECT 2738.755 3434.380 2738.925 3434.550 ;
        RECT 2739.115 3434.380 2739.285 3434.550 ;
        RECT 2739.475 3434.380 2739.645 3434.550 ;
        RECT 2739.835 3434.380 2740.005 3434.550 ;
        RECT 2740.195 3434.380 2740.365 3434.550 ;
        RECT 2740.555 3434.380 2740.725 3434.550 ;
        RECT 2740.915 3434.380 2741.085 3434.550 ;
        RECT 2741.275 3434.380 2741.445 3434.550 ;
        RECT 2741.635 3434.380 2741.805 3434.550 ;
        RECT 2741.995 3434.380 2742.165 3434.550 ;
        RECT 2742.355 3434.380 2742.525 3434.550 ;
        RECT 2742.715 3434.380 2742.885 3434.550 ;
        RECT 2744.215 3434.380 2744.385 3434.550 ;
        RECT 2744.575 3434.380 2744.745 3434.550 ;
        RECT 2744.935 3434.380 2745.105 3434.550 ;
        RECT 2745.295 3434.380 2745.465 3434.550 ;
        RECT 2745.655 3434.380 2745.825 3434.550 ;
        RECT 2746.015 3434.380 2746.185 3434.550 ;
        RECT 2746.375 3434.380 2746.545 3434.550 ;
        RECT 2746.735 3434.380 2746.905 3434.550 ;
        RECT 2747.095 3434.380 2747.265 3434.550 ;
        RECT 2747.455 3434.380 2747.625 3434.550 ;
        RECT 2747.815 3434.380 2747.985 3434.550 ;
        RECT 2748.175 3434.380 2748.345 3434.550 ;
        RECT 2748.535 3434.380 2748.705 3434.550 ;
        RECT 2748.895 3434.380 2749.065 3434.550 ;
        RECT 2750.395 3434.380 2750.565 3434.550 ;
        RECT 2750.755 3434.380 2750.925 3434.550 ;
        RECT 2751.115 3434.380 2751.285 3434.550 ;
        RECT 2751.475 3434.380 2751.645 3434.550 ;
        RECT 2751.835 3434.380 2752.005 3434.550 ;
        RECT 2752.195 3434.380 2752.365 3434.550 ;
        RECT 2752.555 3434.380 2752.725 3434.550 ;
        RECT 2752.915 3434.380 2753.085 3434.550 ;
        RECT 2753.275 3434.380 2753.445 3434.550 ;
        RECT 2753.635 3434.380 2753.805 3434.550 ;
        RECT 2753.995 3434.380 2754.165 3434.550 ;
        RECT 2754.355 3434.380 2754.525 3434.550 ;
        RECT 2754.715 3434.380 2754.885 3434.550 ;
        RECT 2755.075 3434.380 2755.245 3434.550 ;
        RECT 2756.575 3434.380 2756.745 3434.550 ;
        RECT 2756.935 3434.380 2757.105 3434.550 ;
        RECT 2757.295 3434.380 2757.465 3434.550 ;
        RECT 2757.655 3434.380 2757.825 3434.550 ;
        RECT 2758.015 3434.380 2758.185 3434.550 ;
        RECT 2758.375 3434.380 2758.545 3434.550 ;
        RECT 2758.735 3434.380 2758.905 3434.550 ;
        RECT 2759.095 3434.380 2759.265 3434.550 ;
        RECT 2759.455 3434.380 2759.625 3434.550 ;
        RECT 2759.815 3434.380 2759.985 3434.550 ;
        RECT 2760.175 3434.380 2760.345 3434.550 ;
        RECT 2760.535 3434.380 2760.705 3434.550 ;
        RECT 2760.895 3434.380 2761.065 3434.550 ;
        RECT 2761.255 3434.380 2761.425 3434.550 ;
        RECT 2700.955 3431.680 2701.125 3431.850 ;
        RECT 2701.315 3431.680 2701.485 3431.850 ;
        RECT 2701.675 3431.680 2701.845 3431.850 ;
        RECT 2702.035 3431.680 2702.205 3431.850 ;
        RECT 2702.395 3431.680 2702.565 3431.850 ;
        RECT 2702.755 3431.680 2702.925 3431.850 ;
        RECT 2703.115 3431.680 2703.285 3431.850 ;
        RECT 2703.475 3431.680 2703.645 3431.850 ;
        RECT 2703.835 3431.680 2704.005 3431.850 ;
        RECT 2704.195 3431.680 2704.365 3431.850 ;
        RECT 2704.555 3431.680 2704.725 3431.850 ;
        RECT 2704.915 3431.680 2705.085 3431.850 ;
        RECT 2705.275 3431.680 2705.445 3431.850 ;
        RECT 2705.635 3431.680 2705.805 3431.850 ;
        RECT 2707.135 3431.680 2707.305 3431.850 ;
        RECT 2707.495 3431.680 2707.665 3431.850 ;
        RECT 2707.855 3431.680 2708.025 3431.850 ;
        RECT 2708.215 3431.680 2708.385 3431.850 ;
        RECT 2708.575 3431.680 2708.745 3431.850 ;
        RECT 2708.935 3431.680 2709.105 3431.850 ;
        RECT 2709.295 3431.680 2709.465 3431.850 ;
        RECT 2709.655 3431.680 2709.825 3431.850 ;
        RECT 2710.015 3431.680 2710.185 3431.850 ;
        RECT 2710.375 3431.680 2710.545 3431.850 ;
        RECT 2710.735 3431.680 2710.905 3431.850 ;
        RECT 2711.095 3431.680 2711.265 3431.850 ;
        RECT 2711.455 3431.680 2711.625 3431.850 ;
        RECT 2711.815 3431.680 2711.985 3431.850 ;
        RECT 2713.315 3431.680 2713.485 3431.850 ;
        RECT 2713.675 3431.680 2713.845 3431.850 ;
        RECT 2714.035 3431.680 2714.205 3431.850 ;
        RECT 2714.395 3431.680 2714.565 3431.850 ;
        RECT 2714.755 3431.680 2714.925 3431.850 ;
        RECT 2715.115 3431.680 2715.285 3431.850 ;
        RECT 2715.475 3431.680 2715.645 3431.850 ;
        RECT 2715.835 3431.680 2716.005 3431.850 ;
        RECT 2716.195 3431.680 2716.365 3431.850 ;
        RECT 2716.555 3431.680 2716.725 3431.850 ;
        RECT 2716.915 3431.680 2717.085 3431.850 ;
        RECT 2717.275 3431.680 2717.445 3431.850 ;
        RECT 2717.635 3431.680 2717.805 3431.850 ;
        RECT 2717.995 3431.680 2718.165 3431.850 ;
        RECT 2719.495 3431.680 2719.665 3431.850 ;
        RECT 2719.855 3431.680 2720.025 3431.850 ;
        RECT 2720.215 3431.680 2720.385 3431.850 ;
        RECT 2720.575 3431.680 2720.745 3431.850 ;
        RECT 2720.935 3431.680 2721.105 3431.850 ;
        RECT 2721.295 3431.680 2721.465 3431.850 ;
        RECT 2721.655 3431.680 2721.825 3431.850 ;
        RECT 2722.015 3431.680 2722.185 3431.850 ;
        RECT 2722.375 3431.680 2722.545 3431.850 ;
        RECT 2722.735 3431.680 2722.905 3431.850 ;
        RECT 2723.095 3431.680 2723.265 3431.850 ;
        RECT 2723.455 3431.680 2723.625 3431.850 ;
        RECT 2723.815 3431.680 2723.985 3431.850 ;
        RECT 2724.175 3431.680 2724.345 3431.850 ;
        RECT 2725.675 3431.680 2725.845 3431.850 ;
        RECT 2726.035 3431.680 2726.205 3431.850 ;
        RECT 2726.395 3431.680 2726.565 3431.850 ;
        RECT 2726.755 3431.680 2726.925 3431.850 ;
        RECT 2727.115 3431.680 2727.285 3431.850 ;
        RECT 2727.475 3431.680 2727.645 3431.850 ;
        RECT 2727.835 3431.680 2728.005 3431.850 ;
        RECT 2728.195 3431.680 2728.365 3431.850 ;
        RECT 2728.555 3431.680 2728.725 3431.850 ;
        RECT 2728.915 3431.680 2729.085 3431.850 ;
        RECT 2729.275 3431.680 2729.445 3431.850 ;
        RECT 2729.635 3431.680 2729.805 3431.850 ;
        RECT 2729.995 3431.680 2730.165 3431.850 ;
        RECT 2730.355 3431.680 2730.525 3431.850 ;
        RECT 2731.855 3431.680 2732.025 3431.850 ;
        RECT 2732.215 3431.680 2732.385 3431.850 ;
        RECT 2732.575 3431.680 2732.745 3431.850 ;
        RECT 2732.935 3431.680 2733.105 3431.850 ;
        RECT 2733.295 3431.680 2733.465 3431.850 ;
        RECT 2733.655 3431.680 2733.825 3431.850 ;
        RECT 2734.015 3431.680 2734.185 3431.850 ;
        RECT 2734.375 3431.680 2734.545 3431.850 ;
        RECT 2734.735 3431.680 2734.905 3431.850 ;
        RECT 2735.095 3431.680 2735.265 3431.850 ;
        RECT 2735.455 3431.680 2735.625 3431.850 ;
        RECT 2735.815 3431.680 2735.985 3431.850 ;
        RECT 2736.175 3431.680 2736.345 3431.850 ;
        RECT 2736.535 3431.680 2736.705 3431.850 ;
        RECT 2738.035 3431.680 2738.205 3431.850 ;
        RECT 2738.395 3431.680 2738.565 3431.850 ;
        RECT 2738.755 3431.680 2738.925 3431.850 ;
        RECT 2739.115 3431.680 2739.285 3431.850 ;
        RECT 2739.475 3431.680 2739.645 3431.850 ;
        RECT 2739.835 3431.680 2740.005 3431.850 ;
        RECT 2740.195 3431.680 2740.365 3431.850 ;
        RECT 2740.555 3431.680 2740.725 3431.850 ;
        RECT 2740.915 3431.680 2741.085 3431.850 ;
        RECT 2741.275 3431.680 2741.445 3431.850 ;
        RECT 2741.635 3431.680 2741.805 3431.850 ;
        RECT 2741.995 3431.680 2742.165 3431.850 ;
        RECT 2742.355 3431.680 2742.525 3431.850 ;
        RECT 2742.715 3431.680 2742.885 3431.850 ;
        RECT 2744.215 3431.680 2744.385 3431.850 ;
        RECT 2744.575 3431.680 2744.745 3431.850 ;
        RECT 2744.935 3431.680 2745.105 3431.850 ;
        RECT 2745.295 3431.680 2745.465 3431.850 ;
        RECT 2745.655 3431.680 2745.825 3431.850 ;
        RECT 2746.015 3431.680 2746.185 3431.850 ;
        RECT 2746.375 3431.680 2746.545 3431.850 ;
        RECT 2746.735 3431.680 2746.905 3431.850 ;
        RECT 2747.095 3431.680 2747.265 3431.850 ;
        RECT 2747.455 3431.680 2747.625 3431.850 ;
        RECT 2747.815 3431.680 2747.985 3431.850 ;
        RECT 2748.175 3431.680 2748.345 3431.850 ;
        RECT 2748.535 3431.680 2748.705 3431.850 ;
        RECT 2748.895 3431.680 2749.065 3431.850 ;
        RECT 2750.395 3431.680 2750.565 3431.850 ;
        RECT 2750.755 3431.680 2750.925 3431.850 ;
        RECT 2751.115 3431.680 2751.285 3431.850 ;
        RECT 2751.475 3431.680 2751.645 3431.850 ;
        RECT 2751.835 3431.680 2752.005 3431.850 ;
        RECT 2752.195 3431.680 2752.365 3431.850 ;
        RECT 2752.555 3431.680 2752.725 3431.850 ;
        RECT 2752.915 3431.680 2753.085 3431.850 ;
        RECT 2753.275 3431.680 2753.445 3431.850 ;
        RECT 2753.635 3431.680 2753.805 3431.850 ;
        RECT 2753.995 3431.680 2754.165 3431.850 ;
        RECT 2754.355 3431.680 2754.525 3431.850 ;
        RECT 2754.715 3431.680 2754.885 3431.850 ;
        RECT 2755.075 3431.680 2755.245 3431.850 ;
        RECT 2756.575 3431.680 2756.745 3431.850 ;
        RECT 2756.935 3431.680 2757.105 3431.850 ;
        RECT 2757.295 3431.680 2757.465 3431.850 ;
        RECT 2757.655 3431.680 2757.825 3431.850 ;
        RECT 2758.015 3431.680 2758.185 3431.850 ;
        RECT 2758.375 3431.680 2758.545 3431.850 ;
        RECT 2758.735 3431.680 2758.905 3431.850 ;
        RECT 2759.095 3431.680 2759.265 3431.850 ;
        RECT 2759.455 3431.680 2759.625 3431.850 ;
        RECT 2759.815 3431.680 2759.985 3431.850 ;
        RECT 2760.175 3431.680 2760.345 3431.850 ;
        RECT 2760.535 3431.680 2760.705 3431.850 ;
        RECT 2760.895 3431.680 2761.065 3431.850 ;
        RECT 2761.255 3431.680 2761.425 3431.850 ;
        RECT 2700.955 3428.980 2701.125 3429.150 ;
        RECT 2701.315 3428.980 2701.485 3429.150 ;
        RECT 2701.675 3428.980 2701.845 3429.150 ;
        RECT 2702.035 3428.980 2702.205 3429.150 ;
        RECT 2702.395 3428.980 2702.565 3429.150 ;
        RECT 2702.755 3428.980 2702.925 3429.150 ;
        RECT 2703.115 3428.980 2703.285 3429.150 ;
        RECT 2703.475 3428.980 2703.645 3429.150 ;
        RECT 2703.835 3428.980 2704.005 3429.150 ;
        RECT 2704.195 3428.980 2704.365 3429.150 ;
        RECT 2704.555 3428.980 2704.725 3429.150 ;
        RECT 2704.915 3428.980 2705.085 3429.150 ;
        RECT 2705.275 3428.980 2705.445 3429.150 ;
        RECT 2705.635 3428.980 2705.805 3429.150 ;
        RECT 2707.135 3428.980 2707.305 3429.150 ;
        RECT 2707.495 3428.980 2707.665 3429.150 ;
        RECT 2707.855 3428.980 2708.025 3429.150 ;
        RECT 2708.215 3428.980 2708.385 3429.150 ;
        RECT 2708.575 3428.980 2708.745 3429.150 ;
        RECT 2708.935 3428.980 2709.105 3429.150 ;
        RECT 2709.295 3428.980 2709.465 3429.150 ;
        RECT 2709.655 3428.980 2709.825 3429.150 ;
        RECT 2710.015 3428.980 2710.185 3429.150 ;
        RECT 2710.375 3428.980 2710.545 3429.150 ;
        RECT 2710.735 3428.980 2710.905 3429.150 ;
        RECT 2711.095 3428.980 2711.265 3429.150 ;
        RECT 2711.455 3428.980 2711.625 3429.150 ;
        RECT 2711.815 3428.980 2711.985 3429.150 ;
        RECT 2713.315 3428.980 2713.485 3429.150 ;
        RECT 2713.675 3428.980 2713.845 3429.150 ;
        RECT 2714.035 3428.980 2714.205 3429.150 ;
        RECT 2714.395 3428.980 2714.565 3429.150 ;
        RECT 2714.755 3428.980 2714.925 3429.150 ;
        RECT 2715.115 3428.980 2715.285 3429.150 ;
        RECT 2715.475 3428.980 2715.645 3429.150 ;
        RECT 2715.835 3428.980 2716.005 3429.150 ;
        RECT 2716.195 3428.980 2716.365 3429.150 ;
        RECT 2716.555 3428.980 2716.725 3429.150 ;
        RECT 2716.915 3428.980 2717.085 3429.150 ;
        RECT 2717.275 3428.980 2717.445 3429.150 ;
        RECT 2717.635 3428.980 2717.805 3429.150 ;
        RECT 2717.995 3428.980 2718.165 3429.150 ;
        RECT 2719.495 3428.980 2719.665 3429.150 ;
        RECT 2719.855 3428.980 2720.025 3429.150 ;
        RECT 2720.215 3428.980 2720.385 3429.150 ;
        RECT 2720.575 3428.980 2720.745 3429.150 ;
        RECT 2720.935 3428.980 2721.105 3429.150 ;
        RECT 2721.295 3428.980 2721.465 3429.150 ;
        RECT 2721.655 3428.980 2721.825 3429.150 ;
        RECT 2722.015 3428.980 2722.185 3429.150 ;
        RECT 2722.375 3428.980 2722.545 3429.150 ;
        RECT 2722.735 3428.980 2722.905 3429.150 ;
        RECT 2723.095 3428.980 2723.265 3429.150 ;
        RECT 2723.455 3428.980 2723.625 3429.150 ;
        RECT 2723.815 3428.980 2723.985 3429.150 ;
        RECT 2724.175 3428.980 2724.345 3429.150 ;
        RECT 2725.675 3428.980 2725.845 3429.150 ;
        RECT 2726.035 3428.980 2726.205 3429.150 ;
        RECT 2726.395 3428.980 2726.565 3429.150 ;
        RECT 2726.755 3428.980 2726.925 3429.150 ;
        RECT 2727.115 3428.980 2727.285 3429.150 ;
        RECT 2727.475 3428.980 2727.645 3429.150 ;
        RECT 2727.835 3428.980 2728.005 3429.150 ;
        RECT 2728.195 3428.980 2728.365 3429.150 ;
        RECT 2728.555 3428.980 2728.725 3429.150 ;
        RECT 2728.915 3428.980 2729.085 3429.150 ;
        RECT 2729.275 3428.980 2729.445 3429.150 ;
        RECT 2729.635 3428.980 2729.805 3429.150 ;
        RECT 2729.995 3428.980 2730.165 3429.150 ;
        RECT 2730.355 3428.980 2730.525 3429.150 ;
        RECT 2731.855 3428.980 2732.025 3429.150 ;
        RECT 2732.215 3428.980 2732.385 3429.150 ;
        RECT 2732.575 3428.980 2732.745 3429.150 ;
        RECT 2732.935 3428.980 2733.105 3429.150 ;
        RECT 2733.295 3428.980 2733.465 3429.150 ;
        RECT 2733.655 3428.980 2733.825 3429.150 ;
        RECT 2734.015 3428.980 2734.185 3429.150 ;
        RECT 2734.375 3428.980 2734.545 3429.150 ;
        RECT 2734.735 3428.980 2734.905 3429.150 ;
        RECT 2735.095 3428.980 2735.265 3429.150 ;
        RECT 2735.455 3428.980 2735.625 3429.150 ;
        RECT 2735.815 3428.980 2735.985 3429.150 ;
        RECT 2736.175 3428.980 2736.345 3429.150 ;
        RECT 2736.535 3428.980 2736.705 3429.150 ;
        RECT 2738.035 3428.980 2738.205 3429.150 ;
        RECT 2738.395 3428.980 2738.565 3429.150 ;
        RECT 2738.755 3428.980 2738.925 3429.150 ;
        RECT 2739.115 3428.980 2739.285 3429.150 ;
        RECT 2739.475 3428.980 2739.645 3429.150 ;
        RECT 2739.835 3428.980 2740.005 3429.150 ;
        RECT 2740.195 3428.980 2740.365 3429.150 ;
        RECT 2740.555 3428.980 2740.725 3429.150 ;
        RECT 2740.915 3428.980 2741.085 3429.150 ;
        RECT 2741.275 3428.980 2741.445 3429.150 ;
        RECT 2741.635 3428.980 2741.805 3429.150 ;
        RECT 2741.995 3428.980 2742.165 3429.150 ;
        RECT 2742.355 3428.980 2742.525 3429.150 ;
        RECT 2742.715 3428.980 2742.885 3429.150 ;
        RECT 2744.215 3428.980 2744.385 3429.150 ;
        RECT 2744.575 3428.980 2744.745 3429.150 ;
        RECT 2744.935 3428.980 2745.105 3429.150 ;
        RECT 2745.295 3428.980 2745.465 3429.150 ;
        RECT 2745.655 3428.980 2745.825 3429.150 ;
        RECT 2746.015 3428.980 2746.185 3429.150 ;
        RECT 2746.375 3428.980 2746.545 3429.150 ;
        RECT 2746.735 3428.980 2746.905 3429.150 ;
        RECT 2747.095 3428.980 2747.265 3429.150 ;
        RECT 2747.455 3428.980 2747.625 3429.150 ;
        RECT 2747.815 3428.980 2747.985 3429.150 ;
        RECT 2748.175 3428.980 2748.345 3429.150 ;
        RECT 2748.535 3428.980 2748.705 3429.150 ;
        RECT 2748.895 3428.980 2749.065 3429.150 ;
        RECT 2750.395 3428.980 2750.565 3429.150 ;
        RECT 2750.755 3428.980 2750.925 3429.150 ;
        RECT 2751.115 3428.980 2751.285 3429.150 ;
        RECT 2751.475 3428.980 2751.645 3429.150 ;
        RECT 2751.835 3428.980 2752.005 3429.150 ;
        RECT 2752.195 3428.980 2752.365 3429.150 ;
        RECT 2752.555 3428.980 2752.725 3429.150 ;
        RECT 2752.915 3428.980 2753.085 3429.150 ;
        RECT 2753.275 3428.980 2753.445 3429.150 ;
        RECT 2753.635 3428.980 2753.805 3429.150 ;
        RECT 2753.995 3428.980 2754.165 3429.150 ;
        RECT 2754.355 3428.980 2754.525 3429.150 ;
        RECT 2754.715 3428.980 2754.885 3429.150 ;
        RECT 2755.075 3428.980 2755.245 3429.150 ;
        RECT 2756.575 3428.980 2756.745 3429.150 ;
        RECT 2756.935 3428.980 2757.105 3429.150 ;
        RECT 2757.295 3428.980 2757.465 3429.150 ;
        RECT 2757.655 3428.980 2757.825 3429.150 ;
        RECT 2758.015 3428.980 2758.185 3429.150 ;
        RECT 2758.375 3428.980 2758.545 3429.150 ;
        RECT 2758.735 3428.980 2758.905 3429.150 ;
        RECT 2759.095 3428.980 2759.265 3429.150 ;
        RECT 2759.455 3428.980 2759.625 3429.150 ;
        RECT 2759.815 3428.980 2759.985 3429.150 ;
        RECT 2760.175 3428.980 2760.345 3429.150 ;
        RECT 2760.535 3428.980 2760.705 3429.150 ;
        RECT 2760.895 3428.980 2761.065 3429.150 ;
        RECT 2761.255 3428.980 2761.425 3429.150 ;
        RECT 2700.955 3426.280 2701.125 3426.450 ;
        RECT 2701.315 3426.280 2701.485 3426.450 ;
        RECT 2701.675 3426.280 2701.845 3426.450 ;
        RECT 2702.035 3426.280 2702.205 3426.450 ;
        RECT 2702.395 3426.280 2702.565 3426.450 ;
        RECT 2702.755 3426.280 2702.925 3426.450 ;
        RECT 2703.115 3426.280 2703.285 3426.450 ;
        RECT 2703.475 3426.280 2703.645 3426.450 ;
        RECT 2703.835 3426.280 2704.005 3426.450 ;
        RECT 2704.195 3426.280 2704.365 3426.450 ;
        RECT 2704.555 3426.280 2704.725 3426.450 ;
        RECT 2704.915 3426.280 2705.085 3426.450 ;
        RECT 2705.275 3426.280 2705.445 3426.450 ;
        RECT 2705.635 3426.280 2705.805 3426.450 ;
        RECT 2707.135 3426.280 2707.305 3426.450 ;
        RECT 2707.495 3426.280 2707.665 3426.450 ;
        RECT 2707.855 3426.280 2708.025 3426.450 ;
        RECT 2708.215 3426.280 2708.385 3426.450 ;
        RECT 2708.575 3426.280 2708.745 3426.450 ;
        RECT 2708.935 3426.280 2709.105 3426.450 ;
        RECT 2709.295 3426.280 2709.465 3426.450 ;
        RECT 2709.655 3426.280 2709.825 3426.450 ;
        RECT 2710.015 3426.280 2710.185 3426.450 ;
        RECT 2710.375 3426.280 2710.545 3426.450 ;
        RECT 2710.735 3426.280 2710.905 3426.450 ;
        RECT 2711.095 3426.280 2711.265 3426.450 ;
        RECT 2711.455 3426.280 2711.625 3426.450 ;
        RECT 2711.815 3426.280 2711.985 3426.450 ;
        RECT 2713.315 3426.280 2713.485 3426.450 ;
        RECT 2713.675 3426.280 2713.845 3426.450 ;
        RECT 2714.035 3426.280 2714.205 3426.450 ;
        RECT 2714.395 3426.280 2714.565 3426.450 ;
        RECT 2714.755 3426.280 2714.925 3426.450 ;
        RECT 2715.115 3426.280 2715.285 3426.450 ;
        RECT 2715.475 3426.280 2715.645 3426.450 ;
        RECT 2715.835 3426.280 2716.005 3426.450 ;
        RECT 2716.195 3426.280 2716.365 3426.450 ;
        RECT 2716.555 3426.280 2716.725 3426.450 ;
        RECT 2716.915 3426.280 2717.085 3426.450 ;
        RECT 2717.275 3426.280 2717.445 3426.450 ;
        RECT 2717.635 3426.280 2717.805 3426.450 ;
        RECT 2717.995 3426.280 2718.165 3426.450 ;
        RECT 2719.495 3426.280 2719.665 3426.450 ;
        RECT 2719.855 3426.280 2720.025 3426.450 ;
        RECT 2720.215 3426.280 2720.385 3426.450 ;
        RECT 2720.575 3426.280 2720.745 3426.450 ;
        RECT 2720.935 3426.280 2721.105 3426.450 ;
        RECT 2721.295 3426.280 2721.465 3426.450 ;
        RECT 2721.655 3426.280 2721.825 3426.450 ;
        RECT 2722.015 3426.280 2722.185 3426.450 ;
        RECT 2722.375 3426.280 2722.545 3426.450 ;
        RECT 2722.735 3426.280 2722.905 3426.450 ;
        RECT 2723.095 3426.280 2723.265 3426.450 ;
        RECT 2723.455 3426.280 2723.625 3426.450 ;
        RECT 2723.815 3426.280 2723.985 3426.450 ;
        RECT 2724.175 3426.280 2724.345 3426.450 ;
        RECT 2725.675 3426.280 2725.845 3426.450 ;
        RECT 2726.035 3426.280 2726.205 3426.450 ;
        RECT 2726.395 3426.280 2726.565 3426.450 ;
        RECT 2726.755 3426.280 2726.925 3426.450 ;
        RECT 2727.115 3426.280 2727.285 3426.450 ;
        RECT 2727.475 3426.280 2727.645 3426.450 ;
        RECT 2727.835 3426.280 2728.005 3426.450 ;
        RECT 2728.195 3426.280 2728.365 3426.450 ;
        RECT 2728.555 3426.280 2728.725 3426.450 ;
        RECT 2728.915 3426.280 2729.085 3426.450 ;
        RECT 2729.275 3426.280 2729.445 3426.450 ;
        RECT 2729.635 3426.280 2729.805 3426.450 ;
        RECT 2729.995 3426.280 2730.165 3426.450 ;
        RECT 2730.355 3426.280 2730.525 3426.450 ;
        RECT 2731.855 3426.280 2732.025 3426.450 ;
        RECT 2732.215 3426.280 2732.385 3426.450 ;
        RECT 2732.575 3426.280 2732.745 3426.450 ;
        RECT 2732.935 3426.280 2733.105 3426.450 ;
        RECT 2733.295 3426.280 2733.465 3426.450 ;
        RECT 2733.655 3426.280 2733.825 3426.450 ;
        RECT 2734.015 3426.280 2734.185 3426.450 ;
        RECT 2734.375 3426.280 2734.545 3426.450 ;
        RECT 2734.735 3426.280 2734.905 3426.450 ;
        RECT 2735.095 3426.280 2735.265 3426.450 ;
        RECT 2735.455 3426.280 2735.625 3426.450 ;
        RECT 2735.815 3426.280 2735.985 3426.450 ;
        RECT 2736.175 3426.280 2736.345 3426.450 ;
        RECT 2736.535 3426.280 2736.705 3426.450 ;
        RECT 2738.035 3426.280 2738.205 3426.450 ;
        RECT 2738.395 3426.280 2738.565 3426.450 ;
        RECT 2738.755 3426.280 2738.925 3426.450 ;
        RECT 2739.115 3426.280 2739.285 3426.450 ;
        RECT 2739.475 3426.280 2739.645 3426.450 ;
        RECT 2739.835 3426.280 2740.005 3426.450 ;
        RECT 2740.195 3426.280 2740.365 3426.450 ;
        RECT 2740.555 3426.280 2740.725 3426.450 ;
        RECT 2740.915 3426.280 2741.085 3426.450 ;
        RECT 2741.275 3426.280 2741.445 3426.450 ;
        RECT 2741.635 3426.280 2741.805 3426.450 ;
        RECT 2741.995 3426.280 2742.165 3426.450 ;
        RECT 2742.355 3426.280 2742.525 3426.450 ;
        RECT 2742.715 3426.280 2742.885 3426.450 ;
        RECT 2744.215 3426.280 2744.385 3426.450 ;
        RECT 2744.575 3426.280 2744.745 3426.450 ;
        RECT 2744.935 3426.280 2745.105 3426.450 ;
        RECT 2745.295 3426.280 2745.465 3426.450 ;
        RECT 2745.655 3426.280 2745.825 3426.450 ;
        RECT 2746.015 3426.280 2746.185 3426.450 ;
        RECT 2746.375 3426.280 2746.545 3426.450 ;
        RECT 2746.735 3426.280 2746.905 3426.450 ;
        RECT 2747.095 3426.280 2747.265 3426.450 ;
        RECT 2747.455 3426.280 2747.625 3426.450 ;
        RECT 2747.815 3426.280 2747.985 3426.450 ;
        RECT 2748.175 3426.280 2748.345 3426.450 ;
        RECT 2748.535 3426.280 2748.705 3426.450 ;
        RECT 2748.895 3426.280 2749.065 3426.450 ;
        RECT 2750.395 3426.280 2750.565 3426.450 ;
        RECT 2750.755 3426.280 2750.925 3426.450 ;
        RECT 2751.115 3426.280 2751.285 3426.450 ;
        RECT 2751.475 3426.280 2751.645 3426.450 ;
        RECT 2751.835 3426.280 2752.005 3426.450 ;
        RECT 2752.195 3426.280 2752.365 3426.450 ;
        RECT 2752.555 3426.280 2752.725 3426.450 ;
        RECT 2752.915 3426.280 2753.085 3426.450 ;
        RECT 2753.275 3426.280 2753.445 3426.450 ;
        RECT 2753.635 3426.280 2753.805 3426.450 ;
        RECT 2753.995 3426.280 2754.165 3426.450 ;
        RECT 2754.355 3426.280 2754.525 3426.450 ;
        RECT 2754.715 3426.280 2754.885 3426.450 ;
        RECT 2755.075 3426.280 2755.245 3426.450 ;
        RECT 2756.575 3426.280 2756.745 3426.450 ;
        RECT 2756.935 3426.280 2757.105 3426.450 ;
        RECT 2757.295 3426.280 2757.465 3426.450 ;
        RECT 2757.655 3426.280 2757.825 3426.450 ;
        RECT 2758.015 3426.280 2758.185 3426.450 ;
        RECT 2758.375 3426.280 2758.545 3426.450 ;
        RECT 2758.735 3426.280 2758.905 3426.450 ;
        RECT 2759.095 3426.280 2759.265 3426.450 ;
        RECT 2759.455 3426.280 2759.625 3426.450 ;
        RECT 2759.815 3426.280 2759.985 3426.450 ;
        RECT 2760.175 3426.280 2760.345 3426.450 ;
        RECT 2760.535 3426.280 2760.705 3426.450 ;
        RECT 2760.895 3426.280 2761.065 3426.450 ;
        RECT 2761.255 3426.280 2761.425 3426.450 ;
        RECT 2713.410 3418.170 2713.580 3418.340 ;
        RECT 2713.770 3418.170 2713.940 3418.340 ;
        RECT 2714.130 3418.170 2714.300 3418.340 ;
        RECT 2714.490 3418.170 2714.660 3418.340 ;
        RECT 2714.850 3418.170 2715.020 3418.340 ;
        RECT 2715.210 3418.170 2715.380 3418.340 ;
        RECT 2715.570 3418.170 2715.740 3418.340 ;
        RECT 2715.930 3418.170 2716.100 3418.340 ;
        RECT 2716.290 3418.170 2716.460 3418.340 ;
        RECT 2716.650 3418.170 2716.820 3418.340 ;
        RECT 2717.010 3418.170 2717.180 3418.340 ;
        RECT 2717.370 3418.170 2717.540 3418.340 ;
        RECT 2717.730 3418.170 2717.900 3418.340 ;
        RECT 2718.090 3418.170 2718.260 3418.340 ;
        RECT 2719.500 3418.170 2719.670 3418.340 ;
        RECT 2719.860 3418.170 2720.030 3418.340 ;
        RECT 2720.220 3418.170 2720.390 3418.340 ;
        RECT 2720.580 3418.170 2720.750 3418.340 ;
        RECT 2720.940 3418.170 2721.110 3418.340 ;
        RECT 2721.300 3418.170 2721.470 3418.340 ;
        RECT 2721.660 3418.170 2721.830 3418.340 ;
        RECT 2722.020 3418.170 2722.190 3418.340 ;
        RECT 2722.380 3418.170 2722.550 3418.340 ;
        RECT 2722.740 3418.170 2722.910 3418.340 ;
        RECT 2723.100 3418.170 2723.270 3418.340 ;
        RECT 2723.460 3418.170 2723.630 3418.340 ;
        RECT 2723.820 3418.170 2723.990 3418.340 ;
        RECT 2724.180 3418.170 2724.350 3418.340 ;
        RECT 2725.590 3418.170 2725.760 3418.340 ;
        RECT 2725.950 3418.170 2726.120 3418.340 ;
        RECT 2726.310 3418.170 2726.480 3418.340 ;
        RECT 2726.670 3418.170 2726.840 3418.340 ;
        RECT 2727.030 3418.170 2727.200 3418.340 ;
        RECT 2727.390 3418.170 2727.560 3418.340 ;
        RECT 2727.750 3418.170 2727.920 3418.340 ;
        RECT 2728.110 3418.170 2728.280 3418.340 ;
        RECT 2728.470 3418.170 2728.640 3418.340 ;
        RECT 2728.830 3418.170 2729.000 3418.340 ;
        RECT 2729.190 3418.170 2729.360 3418.340 ;
        RECT 2729.550 3418.170 2729.720 3418.340 ;
        RECT 2729.910 3418.170 2730.080 3418.340 ;
        RECT 2730.270 3418.170 2730.440 3418.340 ;
        RECT 2731.680 3418.170 2731.850 3418.340 ;
        RECT 2732.040 3418.170 2732.210 3418.340 ;
        RECT 2732.400 3418.170 2732.570 3418.340 ;
        RECT 2732.760 3418.170 2732.930 3418.340 ;
        RECT 2733.120 3418.170 2733.290 3418.340 ;
        RECT 2733.480 3418.170 2733.650 3418.340 ;
        RECT 2733.840 3418.170 2734.010 3418.340 ;
        RECT 2734.200 3418.170 2734.370 3418.340 ;
        RECT 2734.560 3418.170 2734.730 3418.340 ;
        RECT 2734.920 3418.170 2735.090 3418.340 ;
        RECT 2735.280 3418.170 2735.450 3418.340 ;
        RECT 2735.640 3418.170 2735.810 3418.340 ;
        RECT 2736.000 3418.170 2736.170 3418.340 ;
        RECT 2736.360 3418.170 2736.530 3418.340 ;
        RECT 2737.770 3418.170 2737.940 3418.340 ;
        RECT 2738.130 3418.170 2738.300 3418.340 ;
        RECT 2738.490 3418.170 2738.660 3418.340 ;
        RECT 2738.850 3418.170 2739.020 3418.340 ;
        RECT 2739.210 3418.170 2739.380 3418.340 ;
        RECT 2739.570 3418.170 2739.740 3418.340 ;
        RECT 2739.930 3418.170 2740.100 3418.340 ;
        RECT 2740.290 3418.170 2740.460 3418.340 ;
        RECT 2740.650 3418.170 2740.820 3418.340 ;
        RECT 2741.010 3418.170 2741.180 3418.340 ;
        RECT 2741.370 3418.170 2741.540 3418.340 ;
        RECT 2741.730 3418.170 2741.900 3418.340 ;
        RECT 2742.090 3418.170 2742.260 3418.340 ;
        RECT 2742.450 3418.170 2742.620 3418.340 ;
        RECT 2743.860 3418.170 2744.030 3418.340 ;
        RECT 2744.220 3418.170 2744.390 3418.340 ;
        RECT 2744.580 3418.170 2744.750 3418.340 ;
        RECT 2744.940 3418.170 2745.110 3418.340 ;
        RECT 2745.300 3418.170 2745.470 3418.340 ;
        RECT 2745.660 3418.170 2745.830 3418.340 ;
        RECT 2746.020 3418.170 2746.190 3418.340 ;
        RECT 2746.380 3418.170 2746.550 3418.340 ;
        RECT 2746.740 3418.170 2746.910 3418.340 ;
        RECT 2747.100 3418.170 2747.270 3418.340 ;
        RECT 2747.460 3418.170 2747.630 3418.340 ;
        RECT 2747.820 3418.170 2747.990 3418.340 ;
        RECT 2748.180 3418.170 2748.350 3418.340 ;
        RECT 2748.540 3418.170 2748.710 3418.340 ;
        RECT 2713.410 3415.070 2713.580 3415.240 ;
        RECT 2713.770 3415.070 2713.940 3415.240 ;
        RECT 2714.130 3415.070 2714.300 3415.240 ;
        RECT 2714.490 3415.070 2714.660 3415.240 ;
        RECT 2714.850 3415.070 2715.020 3415.240 ;
        RECT 2715.210 3415.070 2715.380 3415.240 ;
        RECT 2715.570 3415.070 2715.740 3415.240 ;
        RECT 2715.930 3415.070 2716.100 3415.240 ;
        RECT 2716.290 3415.070 2716.460 3415.240 ;
        RECT 2716.650 3415.070 2716.820 3415.240 ;
        RECT 2717.010 3415.070 2717.180 3415.240 ;
        RECT 2717.370 3415.070 2717.540 3415.240 ;
        RECT 2717.730 3415.070 2717.900 3415.240 ;
        RECT 2718.090 3415.070 2718.260 3415.240 ;
        RECT 2719.500 3415.070 2719.670 3415.240 ;
        RECT 2719.860 3415.070 2720.030 3415.240 ;
        RECT 2720.220 3415.070 2720.390 3415.240 ;
        RECT 2720.580 3415.070 2720.750 3415.240 ;
        RECT 2720.940 3415.070 2721.110 3415.240 ;
        RECT 2721.300 3415.070 2721.470 3415.240 ;
        RECT 2721.660 3415.070 2721.830 3415.240 ;
        RECT 2722.020 3415.070 2722.190 3415.240 ;
        RECT 2722.380 3415.070 2722.550 3415.240 ;
        RECT 2722.740 3415.070 2722.910 3415.240 ;
        RECT 2723.100 3415.070 2723.270 3415.240 ;
        RECT 2723.460 3415.070 2723.630 3415.240 ;
        RECT 2723.820 3415.070 2723.990 3415.240 ;
        RECT 2724.180 3415.070 2724.350 3415.240 ;
        RECT 2725.590 3415.070 2725.760 3415.240 ;
        RECT 2725.950 3415.070 2726.120 3415.240 ;
        RECT 2726.310 3415.070 2726.480 3415.240 ;
        RECT 2726.670 3415.070 2726.840 3415.240 ;
        RECT 2727.030 3415.070 2727.200 3415.240 ;
        RECT 2727.390 3415.070 2727.560 3415.240 ;
        RECT 2727.750 3415.070 2727.920 3415.240 ;
        RECT 2728.110 3415.070 2728.280 3415.240 ;
        RECT 2728.470 3415.070 2728.640 3415.240 ;
        RECT 2728.830 3415.070 2729.000 3415.240 ;
        RECT 2729.190 3415.070 2729.360 3415.240 ;
        RECT 2729.550 3415.070 2729.720 3415.240 ;
        RECT 2729.910 3415.070 2730.080 3415.240 ;
        RECT 2730.270 3415.070 2730.440 3415.240 ;
        RECT 2731.680 3415.070 2731.850 3415.240 ;
        RECT 2732.040 3415.070 2732.210 3415.240 ;
        RECT 2732.400 3415.070 2732.570 3415.240 ;
        RECT 2732.760 3415.070 2732.930 3415.240 ;
        RECT 2733.120 3415.070 2733.290 3415.240 ;
        RECT 2733.480 3415.070 2733.650 3415.240 ;
        RECT 2733.840 3415.070 2734.010 3415.240 ;
        RECT 2734.200 3415.070 2734.370 3415.240 ;
        RECT 2734.560 3415.070 2734.730 3415.240 ;
        RECT 2734.920 3415.070 2735.090 3415.240 ;
        RECT 2735.280 3415.070 2735.450 3415.240 ;
        RECT 2735.640 3415.070 2735.810 3415.240 ;
        RECT 2736.000 3415.070 2736.170 3415.240 ;
        RECT 2736.360 3415.070 2736.530 3415.240 ;
        RECT 2737.770 3415.070 2737.940 3415.240 ;
        RECT 2738.130 3415.070 2738.300 3415.240 ;
        RECT 2738.490 3415.070 2738.660 3415.240 ;
        RECT 2738.850 3415.070 2739.020 3415.240 ;
        RECT 2739.210 3415.070 2739.380 3415.240 ;
        RECT 2739.570 3415.070 2739.740 3415.240 ;
        RECT 2739.930 3415.070 2740.100 3415.240 ;
        RECT 2740.290 3415.070 2740.460 3415.240 ;
        RECT 2740.650 3415.070 2740.820 3415.240 ;
        RECT 2741.010 3415.070 2741.180 3415.240 ;
        RECT 2741.370 3415.070 2741.540 3415.240 ;
        RECT 2741.730 3415.070 2741.900 3415.240 ;
        RECT 2742.090 3415.070 2742.260 3415.240 ;
        RECT 2742.450 3415.070 2742.620 3415.240 ;
        RECT 2743.860 3415.070 2744.030 3415.240 ;
        RECT 2744.220 3415.070 2744.390 3415.240 ;
        RECT 2744.580 3415.070 2744.750 3415.240 ;
        RECT 2744.940 3415.070 2745.110 3415.240 ;
        RECT 2745.300 3415.070 2745.470 3415.240 ;
        RECT 2745.660 3415.070 2745.830 3415.240 ;
        RECT 2746.020 3415.070 2746.190 3415.240 ;
        RECT 2746.380 3415.070 2746.550 3415.240 ;
        RECT 2746.740 3415.070 2746.910 3415.240 ;
        RECT 2747.100 3415.070 2747.270 3415.240 ;
        RECT 2747.460 3415.070 2747.630 3415.240 ;
        RECT 2747.820 3415.070 2747.990 3415.240 ;
        RECT 2748.180 3415.070 2748.350 3415.240 ;
        RECT 2748.540 3415.070 2748.710 3415.240 ;
      LAYER met1 ;
        RECT 2700.880 3434.480 2705.880 3434.580 ;
        RECT 2707.060 3434.480 2712.060 3434.580 ;
        RECT 2713.240 3434.480 2718.240 3434.580 ;
        RECT 2719.420 3434.480 2724.420 3434.580 ;
        RECT 2725.600 3434.480 2730.600 3434.580 ;
        RECT 2731.780 3434.480 2736.780 3434.580 ;
        RECT 2737.960 3434.480 2742.960 3434.580 ;
        RECT 2744.140 3434.480 2749.140 3434.580 ;
        RECT 2750.320 3434.480 2755.320 3434.580 ;
        RECT 2756.500 3434.480 2761.500 3434.580 ;
        RECT 2700.835 3434.230 2761.585 3434.480 ;
        RECT 2702.435 3434.030 2702.935 3434.230 ;
        RECT 2703.485 3434.030 2703.985 3434.230 ;
        RECT 2714.835 3434.030 2715.335 3434.230 ;
        RECT 2715.935 3434.030 2716.435 3434.230 ;
        RECT 2727.485 3434.030 2727.985 3434.230 ;
        RECT 2728.385 3434.030 2728.885 3434.230 ;
        RECT 2739.785 3433.980 2740.285 3434.230 ;
        RECT 2740.685 3433.980 2741.185 3434.230 ;
        RECT 2752.185 3433.980 2752.685 3434.230 ;
        RECT 2753.035 3433.980 2753.535 3434.230 ;
        RECT 2700.880 3431.780 2705.880 3431.880 ;
        RECT 2707.060 3431.780 2712.060 3431.880 ;
        RECT 2713.240 3431.780 2718.240 3431.880 ;
        RECT 2719.420 3431.780 2724.420 3431.880 ;
        RECT 2725.600 3431.780 2730.600 3431.880 ;
        RECT 2731.780 3431.780 2736.780 3431.880 ;
        RECT 2737.960 3431.780 2742.960 3431.880 ;
        RECT 2744.140 3431.780 2749.140 3431.880 ;
        RECT 2750.320 3431.780 2755.320 3431.880 ;
        RECT 2756.500 3431.780 2761.500 3431.880 ;
        RECT 2700.835 3431.530 2761.585 3431.780 ;
        RECT 2702.435 3431.330 2702.935 3431.530 ;
        RECT 2703.485 3431.330 2703.985 3431.530 ;
        RECT 2714.835 3431.330 2715.335 3431.530 ;
        RECT 2715.935 3431.330 2716.435 3431.530 ;
        RECT 2727.485 3431.330 2727.985 3431.530 ;
        RECT 2728.435 3431.330 2728.935 3431.530 ;
        RECT 2739.785 3431.280 2740.285 3431.530 ;
        RECT 2740.685 3431.280 2741.185 3431.530 ;
        RECT 2752.185 3431.280 2752.685 3431.530 ;
        RECT 2753.035 3431.280 2753.535 3431.530 ;
        RECT 2700.880 3429.080 2705.880 3429.180 ;
        RECT 2707.060 3429.080 2712.060 3429.180 ;
        RECT 2713.240 3429.080 2718.240 3429.180 ;
        RECT 2719.420 3429.080 2724.420 3429.180 ;
        RECT 2725.600 3429.080 2730.600 3429.180 ;
        RECT 2731.780 3429.080 2736.780 3429.180 ;
        RECT 2737.960 3429.080 2742.960 3429.180 ;
        RECT 2744.140 3429.080 2749.140 3429.180 ;
        RECT 2750.320 3429.080 2755.320 3429.180 ;
        RECT 2756.500 3429.080 2761.500 3429.180 ;
        RECT 2700.835 3428.830 2761.585 3429.080 ;
        RECT 2702.435 3428.630 2702.935 3428.830 ;
        RECT 2703.485 3428.630 2703.985 3428.830 ;
        RECT 2714.785 3428.630 2715.285 3428.830 ;
        RECT 2715.985 3428.630 2716.485 3428.830 ;
        RECT 2727.485 3428.630 2727.985 3428.830 ;
        RECT 2728.385 3428.630 2728.885 3428.830 ;
        RECT 2739.835 3428.580 2740.335 3428.830 ;
        RECT 2740.685 3428.580 2741.185 3428.830 ;
        RECT 2752.185 3428.580 2752.685 3428.830 ;
        RECT 2753.035 3428.580 2753.535 3428.830 ;
        RECT 2700.880 3426.380 2705.880 3426.480 ;
        RECT 2707.060 3426.380 2712.060 3426.480 ;
        RECT 2713.240 3426.380 2718.240 3426.480 ;
        RECT 2719.420 3426.380 2724.420 3426.480 ;
        RECT 2725.600 3426.380 2730.600 3426.480 ;
        RECT 2731.780 3426.380 2736.780 3426.480 ;
        RECT 2737.960 3426.380 2742.960 3426.480 ;
        RECT 2744.140 3426.380 2749.140 3426.480 ;
        RECT 2750.320 3426.380 2755.320 3426.480 ;
        RECT 2756.500 3426.380 2761.500 3426.480 ;
        RECT 2700.835 3426.130 2761.585 3426.380 ;
        RECT 2702.435 3425.930 2702.935 3426.130 ;
        RECT 2703.485 3425.930 2703.985 3426.130 ;
        RECT 2714.785 3425.880 2715.285 3426.130 ;
        RECT 2715.985 3425.880 2716.485 3426.130 ;
        RECT 2727.485 3425.930 2727.985 3426.130 ;
        RECT 2728.435 3425.930 2728.935 3426.130 ;
        RECT 2739.785 3425.880 2740.285 3426.130 ;
        RECT 2740.735 3425.880 2741.235 3426.130 ;
        RECT 2752.185 3425.830 2752.685 3426.130 ;
        RECT 2753.035 3425.830 2753.535 3426.130 ;
        RECT 2715.485 3418.730 2717.035 3418.880 ;
        RECT 2714.885 3418.430 2717.035 3418.730 ;
        RECT 2727.935 3418.430 2728.435 3418.580 ;
        RECT 2740.185 3418.430 2741.285 3418.730 ;
        RECT 2746.185 3418.430 2746.685 3418.630 ;
        RECT 2713.285 3418.230 2748.885 3418.430 ;
        RECT 2713.335 3418.140 2718.335 3418.230 ;
        RECT 2719.425 3418.140 2724.425 3418.230 ;
        RECT 2725.515 3418.140 2730.515 3418.230 ;
        RECT 2731.605 3418.140 2736.605 3418.230 ;
        RECT 2737.695 3418.140 2742.695 3418.230 ;
        RECT 2743.785 3418.140 2748.785 3418.230 ;
        RECT 2727.935 3415.330 2728.435 3415.480 ;
        RECT 2746.185 3415.330 2746.685 3415.530 ;
        RECT 2713.285 3415.130 2748.885 3415.330 ;
        RECT 2713.335 3415.040 2718.335 3415.130 ;
        RECT 2719.425 3415.040 2724.425 3415.130 ;
        RECT 2725.515 3415.040 2730.515 3415.130 ;
        RECT 2731.605 3415.040 2736.605 3415.130 ;
        RECT 2737.695 3415.040 2742.695 3415.130 ;
        RECT 2743.785 3415.040 2748.785 3415.130 ;
      LAYER via ;
        RECT 2702.555 3434.100 2702.815 3434.360 ;
        RECT 2703.605 3434.100 2703.865 3434.360 ;
        RECT 2714.955 3434.100 2715.215 3434.360 ;
        RECT 2716.055 3434.100 2716.315 3434.360 ;
        RECT 2727.605 3434.100 2727.865 3434.360 ;
        RECT 2728.505 3434.100 2728.765 3434.360 ;
        RECT 2739.905 3434.050 2740.165 3434.310 ;
        RECT 2740.805 3434.050 2741.065 3434.310 ;
        RECT 2752.305 3434.050 2752.565 3434.310 ;
        RECT 2753.155 3434.050 2753.415 3434.310 ;
        RECT 2702.555 3431.400 2702.815 3431.660 ;
        RECT 2703.605 3431.400 2703.865 3431.660 ;
        RECT 2714.955 3431.400 2715.215 3431.660 ;
        RECT 2716.055 3431.400 2716.315 3431.660 ;
        RECT 2727.605 3431.400 2727.865 3431.660 ;
        RECT 2728.555 3431.400 2728.815 3431.660 ;
        RECT 2739.905 3431.350 2740.165 3431.610 ;
        RECT 2740.805 3431.350 2741.065 3431.610 ;
        RECT 2752.305 3431.350 2752.565 3431.610 ;
        RECT 2753.155 3431.350 2753.415 3431.610 ;
        RECT 2702.555 3428.700 2702.815 3428.960 ;
        RECT 2703.605 3428.700 2703.865 3428.960 ;
        RECT 2714.905 3428.700 2715.165 3428.960 ;
        RECT 2716.105 3428.700 2716.365 3428.960 ;
        RECT 2727.605 3428.700 2727.865 3428.960 ;
        RECT 2728.505 3428.700 2728.765 3428.960 ;
        RECT 2739.955 3428.650 2740.215 3428.910 ;
        RECT 2740.805 3428.650 2741.065 3428.910 ;
        RECT 2752.305 3428.650 2752.565 3428.910 ;
        RECT 2753.155 3428.650 2753.415 3428.910 ;
        RECT 2702.555 3426.000 2702.815 3426.260 ;
        RECT 2703.605 3426.000 2703.865 3426.260 ;
        RECT 2714.905 3425.950 2715.165 3426.210 ;
        RECT 2716.105 3425.950 2716.365 3426.210 ;
        RECT 2727.605 3426.000 2727.865 3426.260 ;
        RECT 2728.555 3426.000 2728.815 3426.260 ;
        RECT 2739.905 3425.950 2740.165 3426.210 ;
        RECT 2740.855 3425.950 2741.115 3426.210 ;
        RECT 2752.305 3425.900 2752.565 3426.160 ;
        RECT 2753.155 3425.900 2753.415 3426.160 ;
        RECT 2716.005 3418.400 2716.265 3418.660 ;
        RECT 2716.555 3418.400 2716.815 3418.660 ;
        RECT 2728.055 3418.250 2728.315 3418.510 ;
        RECT 2740.305 3418.350 2740.565 3418.610 ;
        RECT 2740.905 3418.350 2741.165 3418.610 ;
        RECT 2746.305 3418.300 2746.565 3418.560 ;
        RECT 2728.055 3415.150 2728.315 3415.410 ;
        RECT 2746.305 3415.200 2746.565 3415.460 ;
      LAYER met2 ;
        RECT 2702.485 3425.880 2703.935 3436.680 ;
        RECT 2714.835 3426.680 2716.435 3434.580 ;
        RECT 2714.835 3425.380 2716.885 3426.680 ;
        RECT 2715.935 3418.880 2716.885 3425.380 ;
        RECT 2715.485 3418.230 2717.035 3418.880 ;
        RECT 2727.485 3418.330 2728.935 3434.880 ;
        RECT 2739.785 3426.780 2741.235 3434.880 ;
        RECT 2739.785 3425.780 2741.285 3426.780 ;
        RECT 2752.135 3425.780 2753.585 3436.230 ;
        RECT 2727.985 3415.030 2728.385 3418.330 ;
        RECT 2740.185 3418.230 2741.285 3425.780 ;
        RECT 2745.985 3418.430 2747.435 3418.680 ;
        RECT 2746.235 3415.080 2746.635 3418.430 ;
      LAYER via2 ;
        RECT 2702.670 3435.865 2702.950 3436.145 ;
        RECT 2703.470 3435.865 2703.750 3436.145 ;
        RECT 2752.295 3435.690 2752.575 3435.970 ;
        RECT 2753.145 3435.690 2753.425 3435.970 ;
      LAYER met3 ;
        RECT 2326.970 3511.500 2351.970 3524.000 ;
        RECT 2327.000 3465.500 2352.000 3511.500 ;
        RECT 2327.000 3435.000 2672.500 3465.500 ;
        RECT 2702.485 3435.680 2703.935 3436.380 ;
        RECT 2752.135 3435.590 2753.595 3436.080 ;
      LAYER via3 ;
        RECT 2669.000 3463.500 2670.000 3464.500 ;
        RECT 2671.000 3463.500 2672.000 3464.500 ;
        RECT 2669.000 3462.000 2670.000 3463.000 ;
        RECT 2671.000 3462.000 2672.000 3463.000 ;
        RECT 2669.000 3460.500 2670.000 3461.500 ;
        RECT 2671.000 3460.500 2672.000 3461.500 ;
        RECT 2669.000 3459.000 2670.000 3460.000 ;
        RECT 2671.000 3459.000 2672.000 3460.000 ;
        RECT 2669.000 3457.500 2670.000 3458.500 ;
        RECT 2671.000 3457.500 2672.000 3458.500 ;
        RECT 2669.000 3456.000 2670.000 3457.000 ;
        RECT 2671.000 3456.000 2672.000 3457.000 ;
        RECT 2669.000 3454.500 2670.000 3455.500 ;
        RECT 2671.000 3454.500 2672.000 3455.500 ;
        RECT 2669.000 3453.000 2670.000 3454.000 ;
        RECT 2671.000 3453.000 2672.000 3454.000 ;
        RECT 2669.000 3451.500 2670.000 3452.500 ;
        RECT 2671.000 3451.500 2672.000 3452.500 ;
        RECT 2669.000 3450.000 2670.000 3451.000 ;
        RECT 2671.000 3450.000 2672.000 3451.000 ;
        RECT 2669.000 3448.500 2670.000 3449.500 ;
        RECT 2671.000 3448.500 2672.000 3449.500 ;
        RECT 2669.000 3447.000 2670.000 3448.000 ;
        RECT 2671.000 3447.000 2672.000 3448.000 ;
        RECT 2669.000 3445.500 2670.000 3446.500 ;
        RECT 2671.000 3445.500 2672.000 3446.500 ;
        RECT 2669.000 3444.000 2670.000 3445.000 ;
        RECT 2671.000 3444.000 2672.000 3445.000 ;
        RECT 2669.000 3442.500 2670.000 3443.500 ;
        RECT 2671.000 3442.500 2672.000 3443.500 ;
        RECT 2669.000 3441.000 2670.000 3442.000 ;
        RECT 2671.000 3441.000 2672.000 3442.000 ;
        RECT 2669.000 3439.500 2670.000 3440.500 ;
        RECT 2671.000 3439.500 2672.000 3440.500 ;
        RECT 2669.000 3438.000 2670.000 3439.000 ;
        RECT 2671.000 3438.000 2672.000 3439.000 ;
        RECT 2669.000 3436.500 2670.000 3437.500 ;
        RECT 2671.000 3436.500 2672.000 3437.500 ;
        RECT 2702.650 3435.845 2702.970 3436.165 ;
        RECT 2703.450 3435.845 2703.770 3436.165 ;
        RECT 2752.275 3435.670 2752.595 3435.990 ;
        RECT 2753.125 3435.670 2753.445 3435.990 ;
      LAYER met4 ;
        RECT 2694.780 3465.780 2710.390 3471.535 ;
        RECT 2713.780 3465.780 2729.390 3471.535 ;
        RECT 2732.780 3465.780 2748.390 3471.535 ;
        RECT 2751.780 3465.780 2767.390 3471.535 ;
        RECT 2668.500 3451.700 2672.500 3465.500 ;
        RECT 2694.780 3463.980 2767.390 3465.780 ;
        RECT 2694.780 3455.925 2710.390 3463.980 ;
        RECT 2711.485 3454.880 2712.335 3463.980 ;
        RECT 2713.780 3455.925 2729.390 3463.980 ;
        RECT 2732.780 3455.925 2748.390 3463.980 ;
        RECT 2702.485 3453.930 2712.335 3454.880 ;
        RECT 2749.685 3454.980 2750.485 3463.980 ;
        RECT 2751.780 3455.925 2767.390 3463.980 ;
        RECT 2749.685 3454.330 2753.585 3454.980 ;
        RECT 2702.485 3451.700 2703.935 3453.930 ;
        RECT 2668.500 3444.800 2703.935 3451.700 ;
        RECT 2668.500 3435.000 2672.500 3444.800 ;
        RECT 2702.485 3434.630 2703.935 3444.800 ;
        RECT 2752.135 3433.580 2753.585 3454.330 ;
    END
  END io_analog[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 343.985596 ;
    PORT
      LAYER nwell ;
        RECT 2699.685 3425.530 2762.785 3452.730 ;
        RECT 2710.410 3399.215 2751.460 3405.420 ;
        RECT 2712.210 3399.210 2750.300 3399.215 ;
      LAYER li1 ;
        RECT 2718.085 3452.510 2718.535 3452.830 ;
        RECT 2718.935 3452.510 2719.385 3452.830 ;
        RECT 2730.535 3452.510 2730.985 3452.830 ;
        RECT 2731.385 3452.510 2731.835 3452.830 ;
        RECT 2742.835 3452.510 2743.235 3452.880 ;
        RECT 2743.685 3452.510 2744.085 3452.880 ;
        RECT 2709.165 3452.340 2753.075 3452.510 ;
        RECT 2709.165 3450.580 2709.335 3452.340 ;
        RECT 2710.060 3451.770 2715.100 3451.940 ;
        RECT 2716.240 3451.770 2721.280 3451.940 ;
        RECT 2722.420 3451.770 2727.460 3451.940 ;
        RECT 2728.600 3451.770 2733.640 3451.940 ;
        RECT 2734.780 3451.770 2739.820 3451.940 ;
        RECT 2740.960 3451.770 2746.000 3451.940 ;
        RECT 2747.140 3451.770 2752.180 3451.940 ;
        RECT 2752.905 3450.580 2753.075 3452.340 ;
        RECT 2709.165 3450.410 2753.075 3450.580 ;
        RECT 2709.165 3449.640 2753.075 3449.810 ;
        RECT 2709.165 3447.880 2709.335 3449.640 ;
        RECT 2710.060 3449.070 2715.100 3449.240 ;
        RECT 2716.240 3449.070 2721.280 3449.240 ;
        RECT 2722.420 3449.070 2727.460 3449.240 ;
        RECT 2728.600 3449.070 2733.640 3449.240 ;
        RECT 2734.780 3449.070 2739.820 3449.240 ;
        RECT 2740.960 3449.070 2746.000 3449.240 ;
        RECT 2747.140 3449.070 2752.180 3449.240 ;
        RECT 2752.905 3447.880 2753.075 3449.640 ;
        RECT 2709.165 3447.710 2753.075 3447.880 ;
        RECT 2718.085 3447.110 2719.385 3447.710 ;
        RECT 2730.435 3447.110 2731.885 3447.710 ;
        RECT 2742.735 3447.110 2744.185 3447.710 ;
        RECT 2709.165 3446.940 2753.075 3447.110 ;
        RECT 2709.165 3445.180 2709.335 3446.940 ;
        RECT 2710.060 3446.370 2715.100 3446.540 ;
        RECT 2716.240 3446.370 2721.280 3446.540 ;
        RECT 2722.420 3446.370 2727.460 3446.540 ;
        RECT 2728.600 3446.370 2733.640 3446.540 ;
        RECT 2734.780 3446.370 2739.820 3446.540 ;
        RECT 2740.960 3446.370 2746.000 3446.540 ;
        RECT 2747.140 3446.370 2752.180 3446.540 ;
        RECT 2752.905 3445.180 2753.075 3446.940 ;
        RECT 2709.165 3445.010 2753.075 3445.180 ;
        RECT 2718.035 3444.410 2719.485 3445.010 ;
        RECT 2730.435 3444.410 2731.885 3445.010 ;
        RECT 2742.735 3444.410 2744.185 3445.010 ;
        RECT 2709.165 3444.240 2753.075 3444.410 ;
        RECT 2709.165 3442.480 2709.335 3444.240 ;
        RECT 2710.060 3443.670 2715.100 3443.840 ;
        RECT 2716.240 3443.670 2721.280 3443.840 ;
        RECT 2722.420 3443.670 2727.460 3443.840 ;
        RECT 2728.600 3443.670 2733.640 3443.840 ;
        RECT 2734.780 3443.670 2739.820 3443.840 ;
        RECT 2740.960 3443.670 2746.000 3443.840 ;
        RECT 2747.140 3443.670 2752.180 3443.840 ;
        RECT 2752.905 3442.480 2753.075 3444.240 ;
        RECT 2709.165 3442.310 2753.075 3442.480 ;
        RECT 2709.165 3441.340 2753.075 3441.510 ;
        RECT 2709.165 3439.580 2709.335 3441.340 ;
        RECT 2710.060 3440.770 2715.100 3440.940 ;
        RECT 2716.240 3440.770 2721.280 3440.940 ;
        RECT 2722.420 3440.770 2727.460 3440.940 ;
        RECT 2728.600 3440.770 2733.640 3440.940 ;
        RECT 2734.780 3440.770 2739.820 3440.940 ;
        RECT 2740.960 3440.770 2746.000 3440.940 ;
        RECT 2747.140 3440.770 2752.180 3440.940 ;
        RECT 2752.905 3439.580 2753.075 3441.340 ;
        RECT 2709.165 3439.410 2753.075 3439.580 ;
        RECT 2718.035 3438.610 2719.485 3439.410 ;
        RECT 2730.435 3438.610 2731.885 3439.410 ;
        RECT 2742.735 3438.610 2744.185 3439.410 ;
        RECT 2709.165 3438.440 2753.075 3438.610 ;
        RECT 2709.165 3436.680 2709.335 3438.440 ;
        RECT 2710.060 3437.870 2715.100 3438.040 ;
        RECT 2716.240 3437.870 2721.280 3438.040 ;
        RECT 2722.420 3437.870 2727.460 3438.040 ;
        RECT 2728.600 3437.870 2733.640 3438.040 ;
        RECT 2734.780 3437.870 2739.820 3438.040 ;
        RECT 2740.960 3437.870 2746.000 3438.040 ;
        RECT 2747.140 3437.870 2752.180 3438.040 ;
        RECT 2752.905 3436.680 2753.075 3438.440 ;
        RECT 2709.165 3436.510 2753.075 3436.680 ;
        RECT 2699.965 3435.740 2762.415 3435.910 ;
        RECT 2699.965 3433.980 2700.135 3435.740 ;
        RECT 2700.860 3435.170 2705.900 3435.340 ;
        RECT 2707.040 3435.170 2712.080 3435.340 ;
        RECT 2713.220 3435.170 2718.260 3435.340 ;
        RECT 2719.400 3435.170 2724.440 3435.340 ;
        RECT 2725.580 3435.170 2730.620 3435.340 ;
        RECT 2731.760 3435.170 2736.800 3435.340 ;
        RECT 2737.940 3435.170 2742.980 3435.340 ;
        RECT 2744.120 3435.170 2749.160 3435.340 ;
        RECT 2750.300 3435.170 2755.340 3435.340 ;
        RECT 2756.480 3435.170 2761.520 3435.340 ;
        RECT 2762.245 3433.980 2762.415 3435.740 ;
        RECT 2699.965 3433.810 2762.415 3433.980 ;
        RECT 2708.735 3433.210 2710.285 3433.810 ;
        RECT 2721.385 3433.210 2722.835 3433.810 ;
        RECT 2733.735 3433.210 2735.185 3433.810 ;
        RECT 2745.985 3433.210 2747.435 3433.810 ;
        RECT 2758.485 3433.210 2759.935 3433.810 ;
        RECT 2699.965 3433.040 2762.415 3433.210 ;
        RECT 2699.965 3431.280 2700.135 3433.040 ;
        RECT 2700.860 3432.470 2705.900 3432.640 ;
        RECT 2707.040 3432.470 2712.080 3432.640 ;
        RECT 2713.220 3432.470 2718.260 3432.640 ;
        RECT 2719.400 3432.470 2724.440 3432.640 ;
        RECT 2725.580 3432.470 2730.620 3432.640 ;
        RECT 2731.760 3432.470 2736.800 3432.640 ;
        RECT 2737.940 3432.470 2742.980 3432.640 ;
        RECT 2744.120 3432.470 2749.160 3432.640 ;
        RECT 2750.300 3432.470 2755.340 3432.640 ;
        RECT 2756.480 3432.470 2761.520 3432.640 ;
        RECT 2762.245 3431.280 2762.415 3433.040 ;
        RECT 2699.965 3431.110 2762.415 3431.280 ;
        RECT 2699.965 3430.340 2762.415 3430.510 ;
        RECT 2699.965 3428.580 2700.135 3430.340 ;
        RECT 2700.860 3429.770 2705.900 3429.940 ;
        RECT 2707.040 3429.770 2712.080 3429.940 ;
        RECT 2713.220 3429.770 2718.260 3429.940 ;
        RECT 2719.400 3429.770 2724.440 3429.940 ;
        RECT 2725.580 3429.770 2730.620 3429.940 ;
        RECT 2731.760 3429.770 2736.800 3429.940 ;
        RECT 2737.940 3429.770 2742.980 3429.940 ;
        RECT 2744.120 3429.770 2749.160 3429.940 ;
        RECT 2750.300 3429.770 2755.340 3429.940 ;
        RECT 2756.480 3429.770 2761.520 3429.940 ;
        RECT 2762.245 3428.580 2762.415 3430.340 ;
        RECT 2699.965 3428.410 2762.415 3428.580 ;
        RECT 2708.735 3427.810 2710.285 3428.410 ;
        RECT 2721.385 3427.810 2722.835 3428.410 ;
        RECT 2733.735 3427.810 2735.185 3428.410 ;
        RECT 2745.985 3427.810 2747.435 3428.410 ;
        RECT 2758.485 3427.810 2759.935 3428.410 ;
        RECT 2699.965 3427.640 2762.415 3427.810 ;
        RECT 2699.965 3425.880 2700.135 3427.640 ;
        RECT 2700.860 3427.070 2705.900 3427.240 ;
        RECT 2707.040 3427.070 2712.080 3427.240 ;
        RECT 2713.220 3427.070 2718.260 3427.240 ;
        RECT 2719.400 3427.070 2724.440 3427.240 ;
        RECT 2725.580 3427.070 2730.620 3427.240 ;
        RECT 2731.760 3427.070 2736.800 3427.240 ;
        RECT 2737.940 3427.070 2742.980 3427.240 ;
        RECT 2744.120 3427.070 2749.160 3427.240 ;
        RECT 2750.300 3427.070 2755.340 3427.240 ;
        RECT 2756.480 3427.070 2761.520 3427.240 ;
        RECT 2762.245 3425.880 2762.415 3427.640 ;
        RECT 2699.965 3425.710 2762.415 3425.880 ;
        RECT 2715.160 3404.940 2715.960 3405.410 ;
        RECT 2720.460 3404.940 2721.260 3405.410 ;
        RECT 2727.760 3404.940 2728.560 3405.410 ;
        RECT 2733.860 3404.940 2734.660 3405.410 ;
        RECT 2741.260 3404.940 2742.060 3405.410 ;
        RECT 2746.260 3404.940 2747.060 3405.410 ;
        RECT 2712.390 3404.770 2750.120 3404.940 ;
        RECT 2712.390 3402.510 2712.560 3404.770 ;
        RECT 2715.160 3404.610 2715.960 3404.770 ;
        RECT 2720.460 3404.610 2721.260 3404.770 ;
        RECT 2727.760 3404.610 2728.560 3404.770 ;
        RECT 2733.860 3404.610 2734.660 3404.770 ;
        RECT 2741.260 3404.610 2742.060 3404.770 ;
        RECT 2746.260 3404.610 2747.060 3404.770 ;
        RECT 2713.285 3404.200 2718.325 3404.370 ;
        RECT 2719.465 3404.200 2724.505 3404.370 ;
        RECT 2725.645 3404.200 2730.685 3404.370 ;
        RECT 2731.825 3404.200 2736.865 3404.370 ;
        RECT 2738.005 3404.200 2743.045 3404.370 ;
        RECT 2744.185 3404.200 2749.225 3404.370 ;
        RECT 2749.950 3402.510 2750.120 3404.770 ;
        RECT 2712.390 3402.340 2750.120 3402.510 ;
        RECT 2715.160 3401.990 2715.960 3402.340 ;
        RECT 2720.460 3401.990 2721.260 3402.340 ;
        RECT 2727.760 3401.990 2728.560 3402.340 ;
        RECT 2733.860 3401.990 2734.660 3402.340 ;
        RECT 2741.260 3401.990 2742.060 3402.340 ;
        RECT 2746.260 3401.990 2747.060 3402.340 ;
        RECT 2712.390 3401.820 2750.120 3401.990 ;
        RECT 2712.390 3399.560 2712.560 3401.820 ;
        RECT 2715.160 3401.710 2715.960 3401.820 ;
        RECT 2720.460 3401.710 2721.260 3401.820 ;
        RECT 2727.760 3401.710 2728.560 3401.820 ;
        RECT 2733.860 3401.710 2734.660 3401.820 ;
        RECT 2741.260 3401.710 2742.060 3401.820 ;
        RECT 2746.260 3401.710 2747.060 3401.820 ;
        RECT 2713.285 3401.250 2718.325 3401.420 ;
        RECT 2719.465 3401.250 2724.505 3401.420 ;
        RECT 2725.645 3401.250 2730.685 3401.420 ;
        RECT 2731.825 3401.250 2736.865 3401.420 ;
        RECT 2738.005 3401.250 2743.045 3401.420 ;
        RECT 2744.185 3401.250 2749.225 3401.420 ;
        RECT 2749.950 3399.560 2750.120 3401.820 ;
        RECT 2712.390 3399.390 2750.120 3399.560 ;
      LAYER mcon ;
        RECT 2718.225 3452.570 2718.395 3452.740 ;
        RECT 2719.075 3452.570 2719.245 3452.740 ;
        RECT 2730.675 3452.570 2730.845 3452.740 ;
        RECT 2731.525 3452.570 2731.695 3452.740 ;
        RECT 2742.950 3452.595 2743.120 3452.765 ;
        RECT 2743.800 3452.595 2743.970 3452.765 ;
        RECT 2710.155 3451.770 2710.325 3451.940 ;
        RECT 2710.515 3451.770 2710.685 3451.940 ;
        RECT 2710.875 3451.770 2711.045 3451.940 ;
        RECT 2711.235 3451.770 2711.405 3451.940 ;
        RECT 2711.595 3451.770 2711.765 3451.940 ;
        RECT 2711.955 3451.770 2712.125 3451.940 ;
        RECT 2712.315 3451.770 2712.485 3451.940 ;
        RECT 2712.675 3451.770 2712.845 3451.940 ;
        RECT 2713.035 3451.770 2713.205 3451.940 ;
        RECT 2713.395 3451.770 2713.565 3451.940 ;
        RECT 2713.755 3451.770 2713.925 3451.940 ;
        RECT 2714.115 3451.770 2714.285 3451.940 ;
        RECT 2714.475 3451.770 2714.645 3451.940 ;
        RECT 2714.835 3451.770 2715.005 3451.940 ;
        RECT 2716.335 3451.770 2716.505 3451.940 ;
        RECT 2716.695 3451.770 2716.865 3451.940 ;
        RECT 2717.055 3451.770 2717.225 3451.940 ;
        RECT 2717.415 3451.770 2717.585 3451.940 ;
        RECT 2717.775 3451.770 2717.945 3451.940 ;
        RECT 2718.135 3451.770 2718.305 3451.940 ;
        RECT 2718.495 3451.770 2718.665 3451.940 ;
        RECT 2718.855 3451.770 2719.025 3451.940 ;
        RECT 2719.215 3451.770 2719.385 3451.940 ;
        RECT 2719.575 3451.770 2719.745 3451.940 ;
        RECT 2719.935 3451.770 2720.105 3451.940 ;
        RECT 2720.295 3451.770 2720.465 3451.940 ;
        RECT 2720.655 3451.770 2720.825 3451.940 ;
        RECT 2721.015 3451.770 2721.185 3451.940 ;
        RECT 2722.515 3451.770 2722.685 3451.940 ;
        RECT 2722.875 3451.770 2723.045 3451.940 ;
        RECT 2723.235 3451.770 2723.405 3451.940 ;
        RECT 2723.595 3451.770 2723.765 3451.940 ;
        RECT 2723.955 3451.770 2724.125 3451.940 ;
        RECT 2724.315 3451.770 2724.485 3451.940 ;
        RECT 2724.675 3451.770 2724.845 3451.940 ;
        RECT 2725.035 3451.770 2725.205 3451.940 ;
        RECT 2725.395 3451.770 2725.565 3451.940 ;
        RECT 2725.755 3451.770 2725.925 3451.940 ;
        RECT 2726.115 3451.770 2726.285 3451.940 ;
        RECT 2726.475 3451.770 2726.645 3451.940 ;
        RECT 2726.835 3451.770 2727.005 3451.940 ;
        RECT 2727.195 3451.770 2727.365 3451.940 ;
        RECT 2728.695 3451.770 2728.865 3451.940 ;
        RECT 2729.055 3451.770 2729.225 3451.940 ;
        RECT 2729.415 3451.770 2729.585 3451.940 ;
        RECT 2729.775 3451.770 2729.945 3451.940 ;
        RECT 2730.135 3451.770 2730.305 3451.940 ;
        RECT 2730.495 3451.770 2730.665 3451.940 ;
        RECT 2730.855 3451.770 2731.025 3451.940 ;
        RECT 2731.215 3451.770 2731.385 3451.940 ;
        RECT 2731.575 3451.770 2731.745 3451.940 ;
        RECT 2731.935 3451.770 2732.105 3451.940 ;
        RECT 2732.295 3451.770 2732.465 3451.940 ;
        RECT 2732.655 3451.770 2732.825 3451.940 ;
        RECT 2733.015 3451.770 2733.185 3451.940 ;
        RECT 2733.375 3451.770 2733.545 3451.940 ;
        RECT 2734.875 3451.770 2735.045 3451.940 ;
        RECT 2735.235 3451.770 2735.405 3451.940 ;
        RECT 2735.595 3451.770 2735.765 3451.940 ;
        RECT 2735.955 3451.770 2736.125 3451.940 ;
        RECT 2736.315 3451.770 2736.485 3451.940 ;
        RECT 2736.675 3451.770 2736.845 3451.940 ;
        RECT 2737.035 3451.770 2737.205 3451.940 ;
        RECT 2737.395 3451.770 2737.565 3451.940 ;
        RECT 2737.755 3451.770 2737.925 3451.940 ;
        RECT 2738.115 3451.770 2738.285 3451.940 ;
        RECT 2738.475 3451.770 2738.645 3451.940 ;
        RECT 2738.835 3451.770 2739.005 3451.940 ;
        RECT 2739.195 3451.770 2739.365 3451.940 ;
        RECT 2739.555 3451.770 2739.725 3451.940 ;
        RECT 2741.055 3451.770 2741.225 3451.940 ;
        RECT 2741.415 3451.770 2741.585 3451.940 ;
        RECT 2741.775 3451.770 2741.945 3451.940 ;
        RECT 2742.135 3451.770 2742.305 3451.940 ;
        RECT 2742.495 3451.770 2742.665 3451.940 ;
        RECT 2742.855 3451.770 2743.025 3451.940 ;
        RECT 2743.215 3451.770 2743.385 3451.940 ;
        RECT 2743.575 3451.770 2743.745 3451.940 ;
        RECT 2743.935 3451.770 2744.105 3451.940 ;
        RECT 2744.295 3451.770 2744.465 3451.940 ;
        RECT 2744.655 3451.770 2744.825 3451.940 ;
        RECT 2745.015 3451.770 2745.185 3451.940 ;
        RECT 2745.375 3451.770 2745.545 3451.940 ;
        RECT 2745.735 3451.770 2745.905 3451.940 ;
        RECT 2747.235 3451.770 2747.405 3451.940 ;
        RECT 2747.595 3451.770 2747.765 3451.940 ;
        RECT 2747.955 3451.770 2748.125 3451.940 ;
        RECT 2748.315 3451.770 2748.485 3451.940 ;
        RECT 2748.675 3451.770 2748.845 3451.940 ;
        RECT 2749.035 3451.770 2749.205 3451.940 ;
        RECT 2749.395 3451.770 2749.565 3451.940 ;
        RECT 2749.755 3451.770 2749.925 3451.940 ;
        RECT 2750.115 3451.770 2750.285 3451.940 ;
        RECT 2750.475 3451.770 2750.645 3451.940 ;
        RECT 2750.835 3451.770 2751.005 3451.940 ;
        RECT 2751.195 3451.770 2751.365 3451.940 ;
        RECT 2751.555 3451.770 2751.725 3451.940 ;
        RECT 2751.915 3451.770 2752.085 3451.940 ;
        RECT 2710.155 3449.070 2710.325 3449.240 ;
        RECT 2710.515 3449.070 2710.685 3449.240 ;
        RECT 2710.875 3449.070 2711.045 3449.240 ;
        RECT 2711.235 3449.070 2711.405 3449.240 ;
        RECT 2711.595 3449.070 2711.765 3449.240 ;
        RECT 2711.955 3449.070 2712.125 3449.240 ;
        RECT 2712.315 3449.070 2712.485 3449.240 ;
        RECT 2712.675 3449.070 2712.845 3449.240 ;
        RECT 2713.035 3449.070 2713.205 3449.240 ;
        RECT 2713.395 3449.070 2713.565 3449.240 ;
        RECT 2713.755 3449.070 2713.925 3449.240 ;
        RECT 2714.115 3449.070 2714.285 3449.240 ;
        RECT 2714.475 3449.070 2714.645 3449.240 ;
        RECT 2714.835 3449.070 2715.005 3449.240 ;
        RECT 2716.335 3449.070 2716.505 3449.240 ;
        RECT 2716.695 3449.070 2716.865 3449.240 ;
        RECT 2717.055 3449.070 2717.225 3449.240 ;
        RECT 2717.415 3449.070 2717.585 3449.240 ;
        RECT 2717.775 3449.070 2717.945 3449.240 ;
        RECT 2718.135 3449.070 2718.305 3449.240 ;
        RECT 2718.495 3449.070 2718.665 3449.240 ;
        RECT 2718.855 3449.070 2719.025 3449.240 ;
        RECT 2719.215 3449.070 2719.385 3449.240 ;
        RECT 2719.575 3449.070 2719.745 3449.240 ;
        RECT 2719.935 3449.070 2720.105 3449.240 ;
        RECT 2720.295 3449.070 2720.465 3449.240 ;
        RECT 2720.655 3449.070 2720.825 3449.240 ;
        RECT 2721.015 3449.070 2721.185 3449.240 ;
        RECT 2722.515 3449.070 2722.685 3449.240 ;
        RECT 2722.875 3449.070 2723.045 3449.240 ;
        RECT 2723.235 3449.070 2723.405 3449.240 ;
        RECT 2723.595 3449.070 2723.765 3449.240 ;
        RECT 2723.955 3449.070 2724.125 3449.240 ;
        RECT 2724.315 3449.070 2724.485 3449.240 ;
        RECT 2724.675 3449.070 2724.845 3449.240 ;
        RECT 2725.035 3449.070 2725.205 3449.240 ;
        RECT 2725.395 3449.070 2725.565 3449.240 ;
        RECT 2725.755 3449.070 2725.925 3449.240 ;
        RECT 2726.115 3449.070 2726.285 3449.240 ;
        RECT 2726.475 3449.070 2726.645 3449.240 ;
        RECT 2726.835 3449.070 2727.005 3449.240 ;
        RECT 2727.195 3449.070 2727.365 3449.240 ;
        RECT 2728.695 3449.070 2728.865 3449.240 ;
        RECT 2729.055 3449.070 2729.225 3449.240 ;
        RECT 2729.415 3449.070 2729.585 3449.240 ;
        RECT 2729.775 3449.070 2729.945 3449.240 ;
        RECT 2730.135 3449.070 2730.305 3449.240 ;
        RECT 2730.495 3449.070 2730.665 3449.240 ;
        RECT 2730.855 3449.070 2731.025 3449.240 ;
        RECT 2731.215 3449.070 2731.385 3449.240 ;
        RECT 2731.575 3449.070 2731.745 3449.240 ;
        RECT 2731.935 3449.070 2732.105 3449.240 ;
        RECT 2732.295 3449.070 2732.465 3449.240 ;
        RECT 2732.655 3449.070 2732.825 3449.240 ;
        RECT 2733.015 3449.070 2733.185 3449.240 ;
        RECT 2733.375 3449.070 2733.545 3449.240 ;
        RECT 2734.875 3449.070 2735.045 3449.240 ;
        RECT 2735.235 3449.070 2735.405 3449.240 ;
        RECT 2735.595 3449.070 2735.765 3449.240 ;
        RECT 2735.955 3449.070 2736.125 3449.240 ;
        RECT 2736.315 3449.070 2736.485 3449.240 ;
        RECT 2736.675 3449.070 2736.845 3449.240 ;
        RECT 2737.035 3449.070 2737.205 3449.240 ;
        RECT 2737.395 3449.070 2737.565 3449.240 ;
        RECT 2737.755 3449.070 2737.925 3449.240 ;
        RECT 2738.115 3449.070 2738.285 3449.240 ;
        RECT 2738.475 3449.070 2738.645 3449.240 ;
        RECT 2738.835 3449.070 2739.005 3449.240 ;
        RECT 2739.195 3449.070 2739.365 3449.240 ;
        RECT 2739.555 3449.070 2739.725 3449.240 ;
        RECT 2741.055 3449.070 2741.225 3449.240 ;
        RECT 2741.415 3449.070 2741.585 3449.240 ;
        RECT 2741.775 3449.070 2741.945 3449.240 ;
        RECT 2742.135 3449.070 2742.305 3449.240 ;
        RECT 2742.495 3449.070 2742.665 3449.240 ;
        RECT 2742.855 3449.070 2743.025 3449.240 ;
        RECT 2743.215 3449.070 2743.385 3449.240 ;
        RECT 2743.575 3449.070 2743.745 3449.240 ;
        RECT 2743.935 3449.070 2744.105 3449.240 ;
        RECT 2744.295 3449.070 2744.465 3449.240 ;
        RECT 2744.655 3449.070 2744.825 3449.240 ;
        RECT 2745.015 3449.070 2745.185 3449.240 ;
        RECT 2745.375 3449.070 2745.545 3449.240 ;
        RECT 2745.735 3449.070 2745.905 3449.240 ;
        RECT 2747.235 3449.070 2747.405 3449.240 ;
        RECT 2747.595 3449.070 2747.765 3449.240 ;
        RECT 2747.955 3449.070 2748.125 3449.240 ;
        RECT 2748.315 3449.070 2748.485 3449.240 ;
        RECT 2748.675 3449.070 2748.845 3449.240 ;
        RECT 2749.035 3449.070 2749.205 3449.240 ;
        RECT 2749.395 3449.070 2749.565 3449.240 ;
        RECT 2749.755 3449.070 2749.925 3449.240 ;
        RECT 2750.115 3449.070 2750.285 3449.240 ;
        RECT 2750.475 3449.070 2750.645 3449.240 ;
        RECT 2750.835 3449.070 2751.005 3449.240 ;
        RECT 2751.195 3449.070 2751.365 3449.240 ;
        RECT 2751.555 3449.070 2751.725 3449.240 ;
        RECT 2751.915 3449.070 2752.085 3449.240 ;
        RECT 2718.275 3447.320 2718.445 3447.490 ;
        RECT 2718.975 3447.320 2719.145 3447.490 ;
        RECT 2730.675 3447.320 2730.845 3447.490 ;
        RECT 2731.475 3447.370 2731.645 3447.540 ;
        RECT 2742.950 3447.370 2743.120 3447.540 ;
        RECT 2743.800 3447.370 2743.970 3447.540 ;
        RECT 2710.155 3446.370 2710.325 3446.540 ;
        RECT 2710.515 3446.370 2710.685 3446.540 ;
        RECT 2710.875 3446.370 2711.045 3446.540 ;
        RECT 2711.235 3446.370 2711.405 3446.540 ;
        RECT 2711.595 3446.370 2711.765 3446.540 ;
        RECT 2711.955 3446.370 2712.125 3446.540 ;
        RECT 2712.315 3446.370 2712.485 3446.540 ;
        RECT 2712.675 3446.370 2712.845 3446.540 ;
        RECT 2713.035 3446.370 2713.205 3446.540 ;
        RECT 2713.395 3446.370 2713.565 3446.540 ;
        RECT 2713.755 3446.370 2713.925 3446.540 ;
        RECT 2714.115 3446.370 2714.285 3446.540 ;
        RECT 2714.475 3446.370 2714.645 3446.540 ;
        RECT 2714.835 3446.370 2715.005 3446.540 ;
        RECT 2716.335 3446.370 2716.505 3446.540 ;
        RECT 2716.695 3446.370 2716.865 3446.540 ;
        RECT 2717.055 3446.370 2717.225 3446.540 ;
        RECT 2717.415 3446.370 2717.585 3446.540 ;
        RECT 2717.775 3446.370 2717.945 3446.540 ;
        RECT 2718.135 3446.370 2718.305 3446.540 ;
        RECT 2718.495 3446.370 2718.665 3446.540 ;
        RECT 2718.855 3446.370 2719.025 3446.540 ;
        RECT 2719.215 3446.370 2719.385 3446.540 ;
        RECT 2719.575 3446.370 2719.745 3446.540 ;
        RECT 2719.935 3446.370 2720.105 3446.540 ;
        RECT 2720.295 3446.370 2720.465 3446.540 ;
        RECT 2720.655 3446.370 2720.825 3446.540 ;
        RECT 2721.015 3446.370 2721.185 3446.540 ;
        RECT 2722.515 3446.370 2722.685 3446.540 ;
        RECT 2722.875 3446.370 2723.045 3446.540 ;
        RECT 2723.235 3446.370 2723.405 3446.540 ;
        RECT 2723.595 3446.370 2723.765 3446.540 ;
        RECT 2723.955 3446.370 2724.125 3446.540 ;
        RECT 2724.315 3446.370 2724.485 3446.540 ;
        RECT 2724.675 3446.370 2724.845 3446.540 ;
        RECT 2725.035 3446.370 2725.205 3446.540 ;
        RECT 2725.395 3446.370 2725.565 3446.540 ;
        RECT 2725.755 3446.370 2725.925 3446.540 ;
        RECT 2726.115 3446.370 2726.285 3446.540 ;
        RECT 2726.475 3446.370 2726.645 3446.540 ;
        RECT 2726.835 3446.370 2727.005 3446.540 ;
        RECT 2727.195 3446.370 2727.365 3446.540 ;
        RECT 2728.695 3446.370 2728.865 3446.540 ;
        RECT 2729.055 3446.370 2729.225 3446.540 ;
        RECT 2729.415 3446.370 2729.585 3446.540 ;
        RECT 2729.775 3446.370 2729.945 3446.540 ;
        RECT 2730.135 3446.370 2730.305 3446.540 ;
        RECT 2730.495 3446.370 2730.665 3446.540 ;
        RECT 2730.855 3446.370 2731.025 3446.540 ;
        RECT 2731.215 3446.370 2731.385 3446.540 ;
        RECT 2731.575 3446.370 2731.745 3446.540 ;
        RECT 2731.935 3446.370 2732.105 3446.540 ;
        RECT 2732.295 3446.370 2732.465 3446.540 ;
        RECT 2732.655 3446.370 2732.825 3446.540 ;
        RECT 2733.015 3446.370 2733.185 3446.540 ;
        RECT 2733.375 3446.370 2733.545 3446.540 ;
        RECT 2734.875 3446.370 2735.045 3446.540 ;
        RECT 2735.235 3446.370 2735.405 3446.540 ;
        RECT 2735.595 3446.370 2735.765 3446.540 ;
        RECT 2735.955 3446.370 2736.125 3446.540 ;
        RECT 2736.315 3446.370 2736.485 3446.540 ;
        RECT 2736.675 3446.370 2736.845 3446.540 ;
        RECT 2737.035 3446.370 2737.205 3446.540 ;
        RECT 2737.395 3446.370 2737.565 3446.540 ;
        RECT 2737.755 3446.370 2737.925 3446.540 ;
        RECT 2738.115 3446.370 2738.285 3446.540 ;
        RECT 2738.475 3446.370 2738.645 3446.540 ;
        RECT 2738.835 3446.370 2739.005 3446.540 ;
        RECT 2739.195 3446.370 2739.365 3446.540 ;
        RECT 2739.555 3446.370 2739.725 3446.540 ;
        RECT 2741.055 3446.370 2741.225 3446.540 ;
        RECT 2741.415 3446.370 2741.585 3446.540 ;
        RECT 2741.775 3446.370 2741.945 3446.540 ;
        RECT 2742.135 3446.370 2742.305 3446.540 ;
        RECT 2742.495 3446.370 2742.665 3446.540 ;
        RECT 2742.855 3446.370 2743.025 3446.540 ;
        RECT 2743.215 3446.370 2743.385 3446.540 ;
        RECT 2743.575 3446.370 2743.745 3446.540 ;
        RECT 2743.935 3446.370 2744.105 3446.540 ;
        RECT 2744.295 3446.370 2744.465 3446.540 ;
        RECT 2744.655 3446.370 2744.825 3446.540 ;
        RECT 2745.015 3446.370 2745.185 3446.540 ;
        RECT 2745.375 3446.370 2745.545 3446.540 ;
        RECT 2745.735 3446.370 2745.905 3446.540 ;
        RECT 2747.235 3446.370 2747.405 3446.540 ;
        RECT 2747.595 3446.370 2747.765 3446.540 ;
        RECT 2747.955 3446.370 2748.125 3446.540 ;
        RECT 2748.315 3446.370 2748.485 3446.540 ;
        RECT 2748.675 3446.370 2748.845 3446.540 ;
        RECT 2749.035 3446.370 2749.205 3446.540 ;
        RECT 2749.395 3446.370 2749.565 3446.540 ;
        RECT 2749.755 3446.370 2749.925 3446.540 ;
        RECT 2750.115 3446.370 2750.285 3446.540 ;
        RECT 2750.475 3446.370 2750.645 3446.540 ;
        RECT 2750.835 3446.370 2751.005 3446.540 ;
        RECT 2751.195 3446.370 2751.365 3446.540 ;
        RECT 2751.555 3446.370 2751.725 3446.540 ;
        RECT 2751.915 3446.370 2752.085 3446.540 ;
        RECT 2718.250 3444.645 2718.420 3444.815 ;
        RECT 2719.100 3444.645 2719.270 3444.815 ;
        RECT 2730.650 3444.645 2730.820 3444.815 ;
        RECT 2731.500 3444.645 2731.670 3444.815 ;
        RECT 2742.950 3444.645 2743.120 3444.815 ;
        RECT 2743.800 3444.645 2743.970 3444.815 ;
        RECT 2710.155 3443.670 2710.325 3443.840 ;
        RECT 2710.515 3443.670 2710.685 3443.840 ;
        RECT 2710.875 3443.670 2711.045 3443.840 ;
        RECT 2711.235 3443.670 2711.405 3443.840 ;
        RECT 2711.595 3443.670 2711.765 3443.840 ;
        RECT 2711.955 3443.670 2712.125 3443.840 ;
        RECT 2712.315 3443.670 2712.485 3443.840 ;
        RECT 2712.675 3443.670 2712.845 3443.840 ;
        RECT 2713.035 3443.670 2713.205 3443.840 ;
        RECT 2713.395 3443.670 2713.565 3443.840 ;
        RECT 2713.755 3443.670 2713.925 3443.840 ;
        RECT 2714.115 3443.670 2714.285 3443.840 ;
        RECT 2714.475 3443.670 2714.645 3443.840 ;
        RECT 2714.835 3443.670 2715.005 3443.840 ;
        RECT 2716.335 3443.670 2716.505 3443.840 ;
        RECT 2716.695 3443.670 2716.865 3443.840 ;
        RECT 2717.055 3443.670 2717.225 3443.840 ;
        RECT 2717.415 3443.670 2717.585 3443.840 ;
        RECT 2717.775 3443.670 2717.945 3443.840 ;
        RECT 2718.135 3443.670 2718.305 3443.840 ;
        RECT 2718.495 3443.670 2718.665 3443.840 ;
        RECT 2718.855 3443.670 2719.025 3443.840 ;
        RECT 2719.215 3443.670 2719.385 3443.840 ;
        RECT 2719.575 3443.670 2719.745 3443.840 ;
        RECT 2719.935 3443.670 2720.105 3443.840 ;
        RECT 2720.295 3443.670 2720.465 3443.840 ;
        RECT 2720.655 3443.670 2720.825 3443.840 ;
        RECT 2721.015 3443.670 2721.185 3443.840 ;
        RECT 2722.515 3443.670 2722.685 3443.840 ;
        RECT 2722.875 3443.670 2723.045 3443.840 ;
        RECT 2723.235 3443.670 2723.405 3443.840 ;
        RECT 2723.595 3443.670 2723.765 3443.840 ;
        RECT 2723.955 3443.670 2724.125 3443.840 ;
        RECT 2724.315 3443.670 2724.485 3443.840 ;
        RECT 2724.675 3443.670 2724.845 3443.840 ;
        RECT 2725.035 3443.670 2725.205 3443.840 ;
        RECT 2725.395 3443.670 2725.565 3443.840 ;
        RECT 2725.755 3443.670 2725.925 3443.840 ;
        RECT 2726.115 3443.670 2726.285 3443.840 ;
        RECT 2726.475 3443.670 2726.645 3443.840 ;
        RECT 2726.835 3443.670 2727.005 3443.840 ;
        RECT 2727.195 3443.670 2727.365 3443.840 ;
        RECT 2728.695 3443.670 2728.865 3443.840 ;
        RECT 2729.055 3443.670 2729.225 3443.840 ;
        RECT 2729.415 3443.670 2729.585 3443.840 ;
        RECT 2729.775 3443.670 2729.945 3443.840 ;
        RECT 2730.135 3443.670 2730.305 3443.840 ;
        RECT 2730.495 3443.670 2730.665 3443.840 ;
        RECT 2730.855 3443.670 2731.025 3443.840 ;
        RECT 2731.215 3443.670 2731.385 3443.840 ;
        RECT 2731.575 3443.670 2731.745 3443.840 ;
        RECT 2731.935 3443.670 2732.105 3443.840 ;
        RECT 2732.295 3443.670 2732.465 3443.840 ;
        RECT 2732.655 3443.670 2732.825 3443.840 ;
        RECT 2733.015 3443.670 2733.185 3443.840 ;
        RECT 2733.375 3443.670 2733.545 3443.840 ;
        RECT 2734.875 3443.670 2735.045 3443.840 ;
        RECT 2735.235 3443.670 2735.405 3443.840 ;
        RECT 2735.595 3443.670 2735.765 3443.840 ;
        RECT 2735.955 3443.670 2736.125 3443.840 ;
        RECT 2736.315 3443.670 2736.485 3443.840 ;
        RECT 2736.675 3443.670 2736.845 3443.840 ;
        RECT 2737.035 3443.670 2737.205 3443.840 ;
        RECT 2737.395 3443.670 2737.565 3443.840 ;
        RECT 2737.755 3443.670 2737.925 3443.840 ;
        RECT 2738.115 3443.670 2738.285 3443.840 ;
        RECT 2738.475 3443.670 2738.645 3443.840 ;
        RECT 2738.835 3443.670 2739.005 3443.840 ;
        RECT 2739.195 3443.670 2739.365 3443.840 ;
        RECT 2739.555 3443.670 2739.725 3443.840 ;
        RECT 2741.055 3443.670 2741.225 3443.840 ;
        RECT 2741.415 3443.670 2741.585 3443.840 ;
        RECT 2741.775 3443.670 2741.945 3443.840 ;
        RECT 2742.135 3443.670 2742.305 3443.840 ;
        RECT 2742.495 3443.670 2742.665 3443.840 ;
        RECT 2742.855 3443.670 2743.025 3443.840 ;
        RECT 2743.215 3443.670 2743.385 3443.840 ;
        RECT 2743.575 3443.670 2743.745 3443.840 ;
        RECT 2743.935 3443.670 2744.105 3443.840 ;
        RECT 2744.295 3443.670 2744.465 3443.840 ;
        RECT 2744.655 3443.670 2744.825 3443.840 ;
        RECT 2745.015 3443.670 2745.185 3443.840 ;
        RECT 2745.375 3443.670 2745.545 3443.840 ;
        RECT 2745.735 3443.670 2745.905 3443.840 ;
        RECT 2747.235 3443.670 2747.405 3443.840 ;
        RECT 2747.595 3443.670 2747.765 3443.840 ;
        RECT 2747.955 3443.670 2748.125 3443.840 ;
        RECT 2748.315 3443.670 2748.485 3443.840 ;
        RECT 2748.675 3443.670 2748.845 3443.840 ;
        RECT 2749.035 3443.670 2749.205 3443.840 ;
        RECT 2749.395 3443.670 2749.565 3443.840 ;
        RECT 2749.755 3443.670 2749.925 3443.840 ;
        RECT 2750.115 3443.670 2750.285 3443.840 ;
        RECT 2750.475 3443.670 2750.645 3443.840 ;
        RECT 2750.835 3443.670 2751.005 3443.840 ;
        RECT 2751.195 3443.670 2751.365 3443.840 ;
        RECT 2751.555 3443.670 2751.725 3443.840 ;
        RECT 2751.915 3443.670 2752.085 3443.840 ;
        RECT 2710.155 3440.770 2710.325 3440.940 ;
        RECT 2710.515 3440.770 2710.685 3440.940 ;
        RECT 2710.875 3440.770 2711.045 3440.940 ;
        RECT 2711.235 3440.770 2711.405 3440.940 ;
        RECT 2711.595 3440.770 2711.765 3440.940 ;
        RECT 2711.955 3440.770 2712.125 3440.940 ;
        RECT 2712.315 3440.770 2712.485 3440.940 ;
        RECT 2712.675 3440.770 2712.845 3440.940 ;
        RECT 2713.035 3440.770 2713.205 3440.940 ;
        RECT 2713.395 3440.770 2713.565 3440.940 ;
        RECT 2713.755 3440.770 2713.925 3440.940 ;
        RECT 2714.115 3440.770 2714.285 3440.940 ;
        RECT 2714.475 3440.770 2714.645 3440.940 ;
        RECT 2714.835 3440.770 2715.005 3440.940 ;
        RECT 2716.335 3440.770 2716.505 3440.940 ;
        RECT 2716.695 3440.770 2716.865 3440.940 ;
        RECT 2717.055 3440.770 2717.225 3440.940 ;
        RECT 2717.415 3440.770 2717.585 3440.940 ;
        RECT 2717.775 3440.770 2717.945 3440.940 ;
        RECT 2718.135 3440.770 2718.305 3440.940 ;
        RECT 2718.495 3440.770 2718.665 3440.940 ;
        RECT 2718.855 3440.770 2719.025 3440.940 ;
        RECT 2719.215 3440.770 2719.385 3440.940 ;
        RECT 2719.575 3440.770 2719.745 3440.940 ;
        RECT 2719.935 3440.770 2720.105 3440.940 ;
        RECT 2720.295 3440.770 2720.465 3440.940 ;
        RECT 2720.655 3440.770 2720.825 3440.940 ;
        RECT 2721.015 3440.770 2721.185 3440.940 ;
        RECT 2722.515 3440.770 2722.685 3440.940 ;
        RECT 2722.875 3440.770 2723.045 3440.940 ;
        RECT 2723.235 3440.770 2723.405 3440.940 ;
        RECT 2723.595 3440.770 2723.765 3440.940 ;
        RECT 2723.955 3440.770 2724.125 3440.940 ;
        RECT 2724.315 3440.770 2724.485 3440.940 ;
        RECT 2724.675 3440.770 2724.845 3440.940 ;
        RECT 2725.035 3440.770 2725.205 3440.940 ;
        RECT 2725.395 3440.770 2725.565 3440.940 ;
        RECT 2725.755 3440.770 2725.925 3440.940 ;
        RECT 2726.115 3440.770 2726.285 3440.940 ;
        RECT 2726.475 3440.770 2726.645 3440.940 ;
        RECT 2726.835 3440.770 2727.005 3440.940 ;
        RECT 2727.195 3440.770 2727.365 3440.940 ;
        RECT 2728.695 3440.770 2728.865 3440.940 ;
        RECT 2729.055 3440.770 2729.225 3440.940 ;
        RECT 2729.415 3440.770 2729.585 3440.940 ;
        RECT 2729.775 3440.770 2729.945 3440.940 ;
        RECT 2730.135 3440.770 2730.305 3440.940 ;
        RECT 2730.495 3440.770 2730.665 3440.940 ;
        RECT 2730.855 3440.770 2731.025 3440.940 ;
        RECT 2731.215 3440.770 2731.385 3440.940 ;
        RECT 2731.575 3440.770 2731.745 3440.940 ;
        RECT 2731.935 3440.770 2732.105 3440.940 ;
        RECT 2732.295 3440.770 2732.465 3440.940 ;
        RECT 2732.655 3440.770 2732.825 3440.940 ;
        RECT 2733.015 3440.770 2733.185 3440.940 ;
        RECT 2733.375 3440.770 2733.545 3440.940 ;
        RECT 2734.875 3440.770 2735.045 3440.940 ;
        RECT 2735.235 3440.770 2735.405 3440.940 ;
        RECT 2735.595 3440.770 2735.765 3440.940 ;
        RECT 2735.955 3440.770 2736.125 3440.940 ;
        RECT 2736.315 3440.770 2736.485 3440.940 ;
        RECT 2736.675 3440.770 2736.845 3440.940 ;
        RECT 2737.035 3440.770 2737.205 3440.940 ;
        RECT 2737.395 3440.770 2737.565 3440.940 ;
        RECT 2737.755 3440.770 2737.925 3440.940 ;
        RECT 2738.115 3440.770 2738.285 3440.940 ;
        RECT 2738.475 3440.770 2738.645 3440.940 ;
        RECT 2738.835 3440.770 2739.005 3440.940 ;
        RECT 2739.195 3440.770 2739.365 3440.940 ;
        RECT 2739.555 3440.770 2739.725 3440.940 ;
        RECT 2741.055 3440.770 2741.225 3440.940 ;
        RECT 2741.415 3440.770 2741.585 3440.940 ;
        RECT 2741.775 3440.770 2741.945 3440.940 ;
        RECT 2742.135 3440.770 2742.305 3440.940 ;
        RECT 2742.495 3440.770 2742.665 3440.940 ;
        RECT 2742.855 3440.770 2743.025 3440.940 ;
        RECT 2743.215 3440.770 2743.385 3440.940 ;
        RECT 2743.575 3440.770 2743.745 3440.940 ;
        RECT 2743.935 3440.770 2744.105 3440.940 ;
        RECT 2744.295 3440.770 2744.465 3440.940 ;
        RECT 2744.655 3440.770 2744.825 3440.940 ;
        RECT 2745.015 3440.770 2745.185 3440.940 ;
        RECT 2745.375 3440.770 2745.545 3440.940 ;
        RECT 2745.735 3440.770 2745.905 3440.940 ;
        RECT 2747.235 3440.770 2747.405 3440.940 ;
        RECT 2747.595 3440.770 2747.765 3440.940 ;
        RECT 2747.955 3440.770 2748.125 3440.940 ;
        RECT 2748.315 3440.770 2748.485 3440.940 ;
        RECT 2748.675 3440.770 2748.845 3440.940 ;
        RECT 2749.035 3440.770 2749.205 3440.940 ;
        RECT 2749.395 3440.770 2749.565 3440.940 ;
        RECT 2749.755 3440.770 2749.925 3440.940 ;
        RECT 2750.115 3440.770 2750.285 3440.940 ;
        RECT 2750.475 3440.770 2750.645 3440.940 ;
        RECT 2750.835 3440.770 2751.005 3440.940 ;
        RECT 2751.195 3440.770 2751.365 3440.940 ;
        RECT 2751.555 3440.770 2751.725 3440.940 ;
        RECT 2751.915 3440.770 2752.085 3440.940 ;
        RECT 2718.275 3438.845 2718.445 3439.015 ;
        RECT 2719.075 3438.845 2719.245 3439.015 ;
        RECT 2730.650 3438.820 2730.820 3438.990 ;
        RECT 2731.500 3438.820 2731.670 3438.990 ;
        RECT 2742.950 3438.820 2743.120 3438.990 ;
        RECT 2743.800 3438.820 2743.970 3438.990 ;
        RECT 2710.155 3437.870 2710.325 3438.040 ;
        RECT 2710.515 3437.870 2710.685 3438.040 ;
        RECT 2710.875 3437.870 2711.045 3438.040 ;
        RECT 2711.235 3437.870 2711.405 3438.040 ;
        RECT 2711.595 3437.870 2711.765 3438.040 ;
        RECT 2711.955 3437.870 2712.125 3438.040 ;
        RECT 2712.315 3437.870 2712.485 3438.040 ;
        RECT 2712.675 3437.870 2712.845 3438.040 ;
        RECT 2713.035 3437.870 2713.205 3438.040 ;
        RECT 2713.395 3437.870 2713.565 3438.040 ;
        RECT 2713.755 3437.870 2713.925 3438.040 ;
        RECT 2714.115 3437.870 2714.285 3438.040 ;
        RECT 2714.475 3437.870 2714.645 3438.040 ;
        RECT 2714.835 3437.870 2715.005 3438.040 ;
        RECT 2716.335 3437.870 2716.505 3438.040 ;
        RECT 2716.695 3437.870 2716.865 3438.040 ;
        RECT 2717.055 3437.870 2717.225 3438.040 ;
        RECT 2717.415 3437.870 2717.585 3438.040 ;
        RECT 2717.775 3437.870 2717.945 3438.040 ;
        RECT 2718.135 3437.870 2718.305 3438.040 ;
        RECT 2718.495 3437.870 2718.665 3438.040 ;
        RECT 2718.855 3437.870 2719.025 3438.040 ;
        RECT 2719.215 3437.870 2719.385 3438.040 ;
        RECT 2719.575 3437.870 2719.745 3438.040 ;
        RECT 2719.935 3437.870 2720.105 3438.040 ;
        RECT 2720.295 3437.870 2720.465 3438.040 ;
        RECT 2720.655 3437.870 2720.825 3438.040 ;
        RECT 2721.015 3437.870 2721.185 3438.040 ;
        RECT 2722.515 3437.870 2722.685 3438.040 ;
        RECT 2722.875 3437.870 2723.045 3438.040 ;
        RECT 2723.235 3437.870 2723.405 3438.040 ;
        RECT 2723.595 3437.870 2723.765 3438.040 ;
        RECT 2723.955 3437.870 2724.125 3438.040 ;
        RECT 2724.315 3437.870 2724.485 3438.040 ;
        RECT 2724.675 3437.870 2724.845 3438.040 ;
        RECT 2725.035 3437.870 2725.205 3438.040 ;
        RECT 2725.395 3437.870 2725.565 3438.040 ;
        RECT 2725.755 3437.870 2725.925 3438.040 ;
        RECT 2726.115 3437.870 2726.285 3438.040 ;
        RECT 2726.475 3437.870 2726.645 3438.040 ;
        RECT 2726.835 3437.870 2727.005 3438.040 ;
        RECT 2727.195 3437.870 2727.365 3438.040 ;
        RECT 2728.695 3437.870 2728.865 3438.040 ;
        RECT 2729.055 3437.870 2729.225 3438.040 ;
        RECT 2729.415 3437.870 2729.585 3438.040 ;
        RECT 2729.775 3437.870 2729.945 3438.040 ;
        RECT 2730.135 3437.870 2730.305 3438.040 ;
        RECT 2730.495 3437.870 2730.665 3438.040 ;
        RECT 2730.855 3437.870 2731.025 3438.040 ;
        RECT 2731.215 3437.870 2731.385 3438.040 ;
        RECT 2731.575 3437.870 2731.745 3438.040 ;
        RECT 2731.935 3437.870 2732.105 3438.040 ;
        RECT 2732.295 3437.870 2732.465 3438.040 ;
        RECT 2732.655 3437.870 2732.825 3438.040 ;
        RECT 2733.015 3437.870 2733.185 3438.040 ;
        RECT 2733.375 3437.870 2733.545 3438.040 ;
        RECT 2734.875 3437.870 2735.045 3438.040 ;
        RECT 2735.235 3437.870 2735.405 3438.040 ;
        RECT 2735.595 3437.870 2735.765 3438.040 ;
        RECT 2735.955 3437.870 2736.125 3438.040 ;
        RECT 2736.315 3437.870 2736.485 3438.040 ;
        RECT 2736.675 3437.870 2736.845 3438.040 ;
        RECT 2737.035 3437.870 2737.205 3438.040 ;
        RECT 2737.395 3437.870 2737.565 3438.040 ;
        RECT 2737.755 3437.870 2737.925 3438.040 ;
        RECT 2738.115 3437.870 2738.285 3438.040 ;
        RECT 2738.475 3437.870 2738.645 3438.040 ;
        RECT 2738.835 3437.870 2739.005 3438.040 ;
        RECT 2739.195 3437.870 2739.365 3438.040 ;
        RECT 2739.555 3437.870 2739.725 3438.040 ;
        RECT 2741.055 3437.870 2741.225 3438.040 ;
        RECT 2741.415 3437.870 2741.585 3438.040 ;
        RECT 2741.775 3437.870 2741.945 3438.040 ;
        RECT 2742.135 3437.870 2742.305 3438.040 ;
        RECT 2742.495 3437.870 2742.665 3438.040 ;
        RECT 2742.855 3437.870 2743.025 3438.040 ;
        RECT 2743.215 3437.870 2743.385 3438.040 ;
        RECT 2743.575 3437.870 2743.745 3438.040 ;
        RECT 2743.935 3437.870 2744.105 3438.040 ;
        RECT 2744.295 3437.870 2744.465 3438.040 ;
        RECT 2744.655 3437.870 2744.825 3438.040 ;
        RECT 2745.015 3437.870 2745.185 3438.040 ;
        RECT 2745.375 3437.870 2745.545 3438.040 ;
        RECT 2745.735 3437.870 2745.905 3438.040 ;
        RECT 2747.235 3437.870 2747.405 3438.040 ;
        RECT 2747.595 3437.870 2747.765 3438.040 ;
        RECT 2747.955 3437.870 2748.125 3438.040 ;
        RECT 2748.315 3437.870 2748.485 3438.040 ;
        RECT 2748.675 3437.870 2748.845 3438.040 ;
        RECT 2749.035 3437.870 2749.205 3438.040 ;
        RECT 2749.395 3437.870 2749.565 3438.040 ;
        RECT 2749.755 3437.870 2749.925 3438.040 ;
        RECT 2750.115 3437.870 2750.285 3438.040 ;
        RECT 2750.475 3437.870 2750.645 3438.040 ;
        RECT 2750.835 3437.870 2751.005 3438.040 ;
        RECT 2751.195 3437.870 2751.365 3438.040 ;
        RECT 2751.555 3437.870 2751.725 3438.040 ;
        RECT 2751.915 3437.870 2752.085 3438.040 ;
        RECT 2700.955 3435.170 2701.125 3435.340 ;
        RECT 2701.315 3435.170 2701.485 3435.340 ;
        RECT 2701.675 3435.170 2701.845 3435.340 ;
        RECT 2702.035 3435.170 2702.205 3435.340 ;
        RECT 2702.395 3435.170 2702.565 3435.340 ;
        RECT 2702.755 3435.170 2702.925 3435.340 ;
        RECT 2703.115 3435.170 2703.285 3435.340 ;
        RECT 2703.475 3435.170 2703.645 3435.340 ;
        RECT 2703.835 3435.170 2704.005 3435.340 ;
        RECT 2704.195 3435.170 2704.365 3435.340 ;
        RECT 2704.555 3435.170 2704.725 3435.340 ;
        RECT 2704.915 3435.170 2705.085 3435.340 ;
        RECT 2705.275 3435.170 2705.445 3435.340 ;
        RECT 2705.635 3435.170 2705.805 3435.340 ;
        RECT 2707.135 3435.170 2707.305 3435.340 ;
        RECT 2707.495 3435.170 2707.665 3435.340 ;
        RECT 2707.855 3435.170 2708.025 3435.340 ;
        RECT 2708.215 3435.170 2708.385 3435.340 ;
        RECT 2708.575 3435.170 2708.745 3435.340 ;
        RECT 2708.935 3435.170 2709.105 3435.340 ;
        RECT 2709.295 3435.170 2709.465 3435.340 ;
        RECT 2709.655 3435.170 2709.825 3435.340 ;
        RECT 2710.015 3435.170 2710.185 3435.340 ;
        RECT 2710.375 3435.170 2710.545 3435.340 ;
        RECT 2710.735 3435.170 2710.905 3435.340 ;
        RECT 2711.095 3435.170 2711.265 3435.340 ;
        RECT 2711.455 3435.170 2711.625 3435.340 ;
        RECT 2711.815 3435.170 2711.985 3435.340 ;
        RECT 2713.315 3435.170 2713.485 3435.340 ;
        RECT 2713.675 3435.170 2713.845 3435.340 ;
        RECT 2714.035 3435.170 2714.205 3435.340 ;
        RECT 2714.395 3435.170 2714.565 3435.340 ;
        RECT 2714.755 3435.170 2714.925 3435.340 ;
        RECT 2715.115 3435.170 2715.285 3435.340 ;
        RECT 2715.475 3435.170 2715.645 3435.340 ;
        RECT 2715.835 3435.170 2716.005 3435.340 ;
        RECT 2716.195 3435.170 2716.365 3435.340 ;
        RECT 2716.555 3435.170 2716.725 3435.340 ;
        RECT 2716.915 3435.170 2717.085 3435.340 ;
        RECT 2717.275 3435.170 2717.445 3435.340 ;
        RECT 2717.635 3435.170 2717.805 3435.340 ;
        RECT 2717.995 3435.170 2718.165 3435.340 ;
        RECT 2719.495 3435.170 2719.665 3435.340 ;
        RECT 2719.855 3435.170 2720.025 3435.340 ;
        RECT 2720.215 3435.170 2720.385 3435.340 ;
        RECT 2720.575 3435.170 2720.745 3435.340 ;
        RECT 2720.935 3435.170 2721.105 3435.340 ;
        RECT 2721.295 3435.170 2721.465 3435.340 ;
        RECT 2721.655 3435.170 2721.825 3435.340 ;
        RECT 2722.015 3435.170 2722.185 3435.340 ;
        RECT 2722.375 3435.170 2722.545 3435.340 ;
        RECT 2722.735 3435.170 2722.905 3435.340 ;
        RECT 2723.095 3435.170 2723.265 3435.340 ;
        RECT 2723.455 3435.170 2723.625 3435.340 ;
        RECT 2723.815 3435.170 2723.985 3435.340 ;
        RECT 2724.175 3435.170 2724.345 3435.340 ;
        RECT 2725.675 3435.170 2725.845 3435.340 ;
        RECT 2726.035 3435.170 2726.205 3435.340 ;
        RECT 2726.395 3435.170 2726.565 3435.340 ;
        RECT 2726.755 3435.170 2726.925 3435.340 ;
        RECT 2727.115 3435.170 2727.285 3435.340 ;
        RECT 2727.475 3435.170 2727.645 3435.340 ;
        RECT 2727.835 3435.170 2728.005 3435.340 ;
        RECT 2728.195 3435.170 2728.365 3435.340 ;
        RECT 2728.555 3435.170 2728.725 3435.340 ;
        RECT 2728.915 3435.170 2729.085 3435.340 ;
        RECT 2729.275 3435.170 2729.445 3435.340 ;
        RECT 2729.635 3435.170 2729.805 3435.340 ;
        RECT 2729.995 3435.170 2730.165 3435.340 ;
        RECT 2730.355 3435.170 2730.525 3435.340 ;
        RECT 2731.855 3435.170 2732.025 3435.340 ;
        RECT 2732.215 3435.170 2732.385 3435.340 ;
        RECT 2732.575 3435.170 2732.745 3435.340 ;
        RECT 2732.935 3435.170 2733.105 3435.340 ;
        RECT 2733.295 3435.170 2733.465 3435.340 ;
        RECT 2733.655 3435.170 2733.825 3435.340 ;
        RECT 2734.015 3435.170 2734.185 3435.340 ;
        RECT 2734.375 3435.170 2734.545 3435.340 ;
        RECT 2734.735 3435.170 2734.905 3435.340 ;
        RECT 2735.095 3435.170 2735.265 3435.340 ;
        RECT 2735.455 3435.170 2735.625 3435.340 ;
        RECT 2735.815 3435.170 2735.985 3435.340 ;
        RECT 2736.175 3435.170 2736.345 3435.340 ;
        RECT 2736.535 3435.170 2736.705 3435.340 ;
        RECT 2738.035 3435.170 2738.205 3435.340 ;
        RECT 2738.395 3435.170 2738.565 3435.340 ;
        RECT 2738.755 3435.170 2738.925 3435.340 ;
        RECT 2739.115 3435.170 2739.285 3435.340 ;
        RECT 2739.475 3435.170 2739.645 3435.340 ;
        RECT 2739.835 3435.170 2740.005 3435.340 ;
        RECT 2740.195 3435.170 2740.365 3435.340 ;
        RECT 2740.555 3435.170 2740.725 3435.340 ;
        RECT 2740.915 3435.170 2741.085 3435.340 ;
        RECT 2741.275 3435.170 2741.445 3435.340 ;
        RECT 2741.635 3435.170 2741.805 3435.340 ;
        RECT 2741.995 3435.170 2742.165 3435.340 ;
        RECT 2742.355 3435.170 2742.525 3435.340 ;
        RECT 2742.715 3435.170 2742.885 3435.340 ;
        RECT 2744.215 3435.170 2744.385 3435.340 ;
        RECT 2744.575 3435.170 2744.745 3435.340 ;
        RECT 2744.935 3435.170 2745.105 3435.340 ;
        RECT 2745.295 3435.170 2745.465 3435.340 ;
        RECT 2745.655 3435.170 2745.825 3435.340 ;
        RECT 2746.015 3435.170 2746.185 3435.340 ;
        RECT 2746.375 3435.170 2746.545 3435.340 ;
        RECT 2746.735 3435.170 2746.905 3435.340 ;
        RECT 2747.095 3435.170 2747.265 3435.340 ;
        RECT 2747.455 3435.170 2747.625 3435.340 ;
        RECT 2747.815 3435.170 2747.985 3435.340 ;
        RECT 2748.175 3435.170 2748.345 3435.340 ;
        RECT 2748.535 3435.170 2748.705 3435.340 ;
        RECT 2748.895 3435.170 2749.065 3435.340 ;
        RECT 2750.395 3435.170 2750.565 3435.340 ;
        RECT 2750.755 3435.170 2750.925 3435.340 ;
        RECT 2751.115 3435.170 2751.285 3435.340 ;
        RECT 2751.475 3435.170 2751.645 3435.340 ;
        RECT 2751.835 3435.170 2752.005 3435.340 ;
        RECT 2752.195 3435.170 2752.365 3435.340 ;
        RECT 2752.555 3435.170 2752.725 3435.340 ;
        RECT 2752.915 3435.170 2753.085 3435.340 ;
        RECT 2753.275 3435.170 2753.445 3435.340 ;
        RECT 2753.635 3435.170 2753.805 3435.340 ;
        RECT 2753.995 3435.170 2754.165 3435.340 ;
        RECT 2754.355 3435.170 2754.525 3435.340 ;
        RECT 2754.715 3435.170 2754.885 3435.340 ;
        RECT 2755.075 3435.170 2755.245 3435.340 ;
        RECT 2756.575 3435.170 2756.745 3435.340 ;
        RECT 2756.935 3435.170 2757.105 3435.340 ;
        RECT 2757.295 3435.170 2757.465 3435.340 ;
        RECT 2757.655 3435.170 2757.825 3435.340 ;
        RECT 2758.015 3435.170 2758.185 3435.340 ;
        RECT 2758.375 3435.170 2758.545 3435.340 ;
        RECT 2758.735 3435.170 2758.905 3435.340 ;
        RECT 2759.095 3435.170 2759.265 3435.340 ;
        RECT 2759.455 3435.170 2759.625 3435.340 ;
        RECT 2759.815 3435.170 2759.985 3435.340 ;
        RECT 2760.175 3435.170 2760.345 3435.340 ;
        RECT 2760.535 3435.170 2760.705 3435.340 ;
        RECT 2760.895 3435.170 2761.065 3435.340 ;
        RECT 2761.255 3435.170 2761.425 3435.340 ;
        RECT 2708.975 3433.445 2709.145 3433.615 ;
        RECT 2709.875 3433.445 2710.045 3433.615 ;
        RECT 2721.625 3433.445 2721.795 3433.615 ;
        RECT 2722.425 3433.445 2722.595 3433.615 ;
        RECT 2733.975 3433.445 2734.145 3433.615 ;
        RECT 2734.775 3433.445 2734.945 3433.615 ;
        RECT 2746.225 3433.445 2746.395 3433.615 ;
        RECT 2747.025 3433.445 2747.195 3433.615 ;
        RECT 2758.725 3433.445 2758.895 3433.615 ;
        RECT 2759.525 3433.445 2759.695 3433.615 ;
        RECT 2700.955 3432.470 2701.125 3432.640 ;
        RECT 2701.315 3432.470 2701.485 3432.640 ;
        RECT 2701.675 3432.470 2701.845 3432.640 ;
        RECT 2702.035 3432.470 2702.205 3432.640 ;
        RECT 2702.395 3432.470 2702.565 3432.640 ;
        RECT 2702.755 3432.470 2702.925 3432.640 ;
        RECT 2703.115 3432.470 2703.285 3432.640 ;
        RECT 2703.475 3432.470 2703.645 3432.640 ;
        RECT 2703.835 3432.470 2704.005 3432.640 ;
        RECT 2704.195 3432.470 2704.365 3432.640 ;
        RECT 2704.555 3432.470 2704.725 3432.640 ;
        RECT 2704.915 3432.470 2705.085 3432.640 ;
        RECT 2705.275 3432.470 2705.445 3432.640 ;
        RECT 2705.635 3432.470 2705.805 3432.640 ;
        RECT 2707.135 3432.470 2707.305 3432.640 ;
        RECT 2707.495 3432.470 2707.665 3432.640 ;
        RECT 2707.855 3432.470 2708.025 3432.640 ;
        RECT 2708.215 3432.470 2708.385 3432.640 ;
        RECT 2708.575 3432.470 2708.745 3432.640 ;
        RECT 2708.935 3432.470 2709.105 3432.640 ;
        RECT 2709.295 3432.470 2709.465 3432.640 ;
        RECT 2709.655 3432.470 2709.825 3432.640 ;
        RECT 2710.015 3432.470 2710.185 3432.640 ;
        RECT 2710.375 3432.470 2710.545 3432.640 ;
        RECT 2710.735 3432.470 2710.905 3432.640 ;
        RECT 2711.095 3432.470 2711.265 3432.640 ;
        RECT 2711.455 3432.470 2711.625 3432.640 ;
        RECT 2711.815 3432.470 2711.985 3432.640 ;
        RECT 2713.315 3432.470 2713.485 3432.640 ;
        RECT 2713.675 3432.470 2713.845 3432.640 ;
        RECT 2714.035 3432.470 2714.205 3432.640 ;
        RECT 2714.395 3432.470 2714.565 3432.640 ;
        RECT 2714.755 3432.470 2714.925 3432.640 ;
        RECT 2715.115 3432.470 2715.285 3432.640 ;
        RECT 2715.475 3432.470 2715.645 3432.640 ;
        RECT 2715.835 3432.470 2716.005 3432.640 ;
        RECT 2716.195 3432.470 2716.365 3432.640 ;
        RECT 2716.555 3432.470 2716.725 3432.640 ;
        RECT 2716.915 3432.470 2717.085 3432.640 ;
        RECT 2717.275 3432.470 2717.445 3432.640 ;
        RECT 2717.635 3432.470 2717.805 3432.640 ;
        RECT 2717.995 3432.470 2718.165 3432.640 ;
        RECT 2719.495 3432.470 2719.665 3432.640 ;
        RECT 2719.855 3432.470 2720.025 3432.640 ;
        RECT 2720.215 3432.470 2720.385 3432.640 ;
        RECT 2720.575 3432.470 2720.745 3432.640 ;
        RECT 2720.935 3432.470 2721.105 3432.640 ;
        RECT 2721.295 3432.470 2721.465 3432.640 ;
        RECT 2721.655 3432.470 2721.825 3432.640 ;
        RECT 2722.015 3432.470 2722.185 3432.640 ;
        RECT 2722.375 3432.470 2722.545 3432.640 ;
        RECT 2722.735 3432.470 2722.905 3432.640 ;
        RECT 2723.095 3432.470 2723.265 3432.640 ;
        RECT 2723.455 3432.470 2723.625 3432.640 ;
        RECT 2723.815 3432.470 2723.985 3432.640 ;
        RECT 2724.175 3432.470 2724.345 3432.640 ;
        RECT 2725.675 3432.470 2725.845 3432.640 ;
        RECT 2726.035 3432.470 2726.205 3432.640 ;
        RECT 2726.395 3432.470 2726.565 3432.640 ;
        RECT 2726.755 3432.470 2726.925 3432.640 ;
        RECT 2727.115 3432.470 2727.285 3432.640 ;
        RECT 2727.475 3432.470 2727.645 3432.640 ;
        RECT 2727.835 3432.470 2728.005 3432.640 ;
        RECT 2728.195 3432.470 2728.365 3432.640 ;
        RECT 2728.555 3432.470 2728.725 3432.640 ;
        RECT 2728.915 3432.470 2729.085 3432.640 ;
        RECT 2729.275 3432.470 2729.445 3432.640 ;
        RECT 2729.635 3432.470 2729.805 3432.640 ;
        RECT 2729.995 3432.470 2730.165 3432.640 ;
        RECT 2730.355 3432.470 2730.525 3432.640 ;
        RECT 2731.855 3432.470 2732.025 3432.640 ;
        RECT 2732.215 3432.470 2732.385 3432.640 ;
        RECT 2732.575 3432.470 2732.745 3432.640 ;
        RECT 2732.935 3432.470 2733.105 3432.640 ;
        RECT 2733.295 3432.470 2733.465 3432.640 ;
        RECT 2733.655 3432.470 2733.825 3432.640 ;
        RECT 2734.015 3432.470 2734.185 3432.640 ;
        RECT 2734.375 3432.470 2734.545 3432.640 ;
        RECT 2734.735 3432.470 2734.905 3432.640 ;
        RECT 2735.095 3432.470 2735.265 3432.640 ;
        RECT 2735.455 3432.470 2735.625 3432.640 ;
        RECT 2735.815 3432.470 2735.985 3432.640 ;
        RECT 2736.175 3432.470 2736.345 3432.640 ;
        RECT 2736.535 3432.470 2736.705 3432.640 ;
        RECT 2738.035 3432.470 2738.205 3432.640 ;
        RECT 2738.395 3432.470 2738.565 3432.640 ;
        RECT 2738.755 3432.470 2738.925 3432.640 ;
        RECT 2739.115 3432.470 2739.285 3432.640 ;
        RECT 2739.475 3432.470 2739.645 3432.640 ;
        RECT 2739.835 3432.470 2740.005 3432.640 ;
        RECT 2740.195 3432.470 2740.365 3432.640 ;
        RECT 2740.555 3432.470 2740.725 3432.640 ;
        RECT 2740.915 3432.470 2741.085 3432.640 ;
        RECT 2741.275 3432.470 2741.445 3432.640 ;
        RECT 2741.635 3432.470 2741.805 3432.640 ;
        RECT 2741.995 3432.470 2742.165 3432.640 ;
        RECT 2742.355 3432.470 2742.525 3432.640 ;
        RECT 2742.715 3432.470 2742.885 3432.640 ;
        RECT 2744.215 3432.470 2744.385 3432.640 ;
        RECT 2744.575 3432.470 2744.745 3432.640 ;
        RECT 2744.935 3432.470 2745.105 3432.640 ;
        RECT 2745.295 3432.470 2745.465 3432.640 ;
        RECT 2745.655 3432.470 2745.825 3432.640 ;
        RECT 2746.015 3432.470 2746.185 3432.640 ;
        RECT 2746.375 3432.470 2746.545 3432.640 ;
        RECT 2746.735 3432.470 2746.905 3432.640 ;
        RECT 2747.095 3432.470 2747.265 3432.640 ;
        RECT 2747.455 3432.470 2747.625 3432.640 ;
        RECT 2747.815 3432.470 2747.985 3432.640 ;
        RECT 2748.175 3432.470 2748.345 3432.640 ;
        RECT 2748.535 3432.470 2748.705 3432.640 ;
        RECT 2748.895 3432.470 2749.065 3432.640 ;
        RECT 2750.395 3432.470 2750.565 3432.640 ;
        RECT 2750.755 3432.470 2750.925 3432.640 ;
        RECT 2751.115 3432.470 2751.285 3432.640 ;
        RECT 2751.475 3432.470 2751.645 3432.640 ;
        RECT 2751.835 3432.470 2752.005 3432.640 ;
        RECT 2752.195 3432.470 2752.365 3432.640 ;
        RECT 2752.555 3432.470 2752.725 3432.640 ;
        RECT 2752.915 3432.470 2753.085 3432.640 ;
        RECT 2753.275 3432.470 2753.445 3432.640 ;
        RECT 2753.635 3432.470 2753.805 3432.640 ;
        RECT 2753.995 3432.470 2754.165 3432.640 ;
        RECT 2754.355 3432.470 2754.525 3432.640 ;
        RECT 2754.715 3432.470 2754.885 3432.640 ;
        RECT 2755.075 3432.470 2755.245 3432.640 ;
        RECT 2756.575 3432.470 2756.745 3432.640 ;
        RECT 2756.935 3432.470 2757.105 3432.640 ;
        RECT 2757.295 3432.470 2757.465 3432.640 ;
        RECT 2757.655 3432.470 2757.825 3432.640 ;
        RECT 2758.015 3432.470 2758.185 3432.640 ;
        RECT 2758.375 3432.470 2758.545 3432.640 ;
        RECT 2758.735 3432.470 2758.905 3432.640 ;
        RECT 2759.095 3432.470 2759.265 3432.640 ;
        RECT 2759.455 3432.470 2759.625 3432.640 ;
        RECT 2759.815 3432.470 2759.985 3432.640 ;
        RECT 2760.175 3432.470 2760.345 3432.640 ;
        RECT 2760.535 3432.470 2760.705 3432.640 ;
        RECT 2760.895 3432.470 2761.065 3432.640 ;
        RECT 2761.255 3432.470 2761.425 3432.640 ;
        RECT 2700.955 3429.770 2701.125 3429.940 ;
        RECT 2701.315 3429.770 2701.485 3429.940 ;
        RECT 2701.675 3429.770 2701.845 3429.940 ;
        RECT 2702.035 3429.770 2702.205 3429.940 ;
        RECT 2702.395 3429.770 2702.565 3429.940 ;
        RECT 2702.755 3429.770 2702.925 3429.940 ;
        RECT 2703.115 3429.770 2703.285 3429.940 ;
        RECT 2703.475 3429.770 2703.645 3429.940 ;
        RECT 2703.835 3429.770 2704.005 3429.940 ;
        RECT 2704.195 3429.770 2704.365 3429.940 ;
        RECT 2704.555 3429.770 2704.725 3429.940 ;
        RECT 2704.915 3429.770 2705.085 3429.940 ;
        RECT 2705.275 3429.770 2705.445 3429.940 ;
        RECT 2705.635 3429.770 2705.805 3429.940 ;
        RECT 2707.135 3429.770 2707.305 3429.940 ;
        RECT 2707.495 3429.770 2707.665 3429.940 ;
        RECT 2707.855 3429.770 2708.025 3429.940 ;
        RECT 2708.215 3429.770 2708.385 3429.940 ;
        RECT 2708.575 3429.770 2708.745 3429.940 ;
        RECT 2708.935 3429.770 2709.105 3429.940 ;
        RECT 2709.295 3429.770 2709.465 3429.940 ;
        RECT 2709.655 3429.770 2709.825 3429.940 ;
        RECT 2710.015 3429.770 2710.185 3429.940 ;
        RECT 2710.375 3429.770 2710.545 3429.940 ;
        RECT 2710.735 3429.770 2710.905 3429.940 ;
        RECT 2711.095 3429.770 2711.265 3429.940 ;
        RECT 2711.455 3429.770 2711.625 3429.940 ;
        RECT 2711.815 3429.770 2711.985 3429.940 ;
        RECT 2713.315 3429.770 2713.485 3429.940 ;
        RECT 2713.675 3429.770 2713.845 3429.940 ;
        RECT 2714.035 3429.770 2714.205 3429.940 ;
        RECT 2714.395 3429.770 2714.565 3429.940 ;
        RECT 2714.755 3429.770 2714.925 3429.940 ;
        RECT 2715.115 3429.770 2715.285 3429.940 ;
        RECT 2715.475 3429.770 2715.645 3429.940 ;
        RECT 2715.835 3429.770 2716.005 3429.940 ;
        RECT 2716.195 3429.770 2716.365 3429.940 ;
        RECT 2716.555 3429.770 2716.725 3429.940 ;
        RECT 2716.915 3429.770 2717.085 3429.940 ;
        RECT 2717.275 3429.770 2717.445 3429.940 ;
        RECT 2717.635 3429.770 2717.805 3429.940 ;
        RECT 2717.995 3429.770 2718.165 3429.940 ;
        RECT 2719.495 3429.770 2719.665 3429.940 ;
        RECT 2719.855 3429.770 2720.025 3429.940 ;
        RECT 2720.215 3429.770 2720.385 3429.940 ;
        RECT 2720.575 3429.770 2720.745 3429.940 ;
        RECT 2720.935 3429.770 2721.105 3429.940 ;
        RECT 2721.295 3429.770 2721.465 3429.940 ;
        RECT 2721.655 3429.770 2721.825 3429.940 ;
        RECT 2722.015 3429.770 2722.185 3429.940 ;
        RECT 2722.375 3429.770 2722.545 3429.940 ;
        RECT 2722.735 3429.770 2722.905 3429.940 ;
        RECT 2723.095 3429.770 2723.265 3429.940 ;
        RECT 2723.455 3429.770 2723.625 3429.940 ;
        RECT 2723.815 3429.770 2723.985 3429.940 ;
        RECT 2724.175 3429.770 2724.345 3429.940 ;
        RECT 2725.675 3429.770 2725.845 3429.940 ;
        RECT 2726.035 3429.770 2726.205 3429.940 ;
        RECT 2726.395 3429.770 2726.565 3429.940 ;
        RECT 2726.755 3429.770 2726.925 3429.940 ;
        RECT 2727.115 3429.770 2727.285 3429.940 ;
        RECT 2727.475 3429.770 2727.645 3429.940 ;
        RECT 2727.835 3429.770 2728.005 3429.940 ;
        RECT 2728.195 3429.770 2728.365 3429.940 ;
        RECT 2728.555 3429.770 2728.725 3429.940 ;
        RECT 2728.915 3429.770 2729.085 3429.940 ;
        RECT 2729.275 3429.770 2729.445 3429.940 ;
        RECT 2729.635 3429.770 2729.805 3429.940 ;
        RECT 2729.995 3429.770 2730.165 3429.940 ;
        RECT 2730.355 3429.770 2730.525 3429.940 ;
        RECT 2731.855 3429.770 2732.025 3429.940 ;
        RECT 2732.215 3429.770 2732.385 3429.940 ;
        RECT 2732.575 3429.770 2732.745 3429.940 ;
        RECT 2732.935 3429.770 2733.105 3429.940 ;
        RECT 2733.295 3429.770 2733.465 3429.940 ;
        RECT 2733.655 3429.770 2733.825 3429.940 ;
        RECT 2734.015 3429.770 2734.185 3429.940 ;
        RECT 2734.375 3429.770 2734.545 3429.940 ;
        RECT 2734.735 3429.770 2734.905 3429.940 ;
        RECT 2735.095 3429.770 2735.265 3429.940 ;
        RECT 2735.455 3429.770 2735.625 3429.940 ;
        RECT 2735.815 3429.770 2735.985 3429.940 ;
        RECT 2736.175 3429.770 2736.345 3429.940 ;
        RECT 2736.535 3429.770 2736.705 3429.940 ;
        RECT 2738.035 3429.770 2738.205 3429.940 ;
        RECT 2738.395 3429.770 2738.565 3429.940 ;
        RECT 2738.755 3429.770 2738.925 3429.940 ;
        RECT 2739.115 3429.770 2739.285 3429.940 ;
        RECT 2739.475 3429.770 2739.645 3429.940 ;
        RECT 2739.835 3429.770 2740.005 3429.940 ;
        RECT 2740.195 3429.770 2740.365 3429.940 ;
        RECT 2740.555 3429.770 2740.725 3429.940 ;
        RECT 2740.915 3429.770 2741.085 3429.940 ;
        RECT 2741.275 3429.770 2741.445 3429.940 ;
        RECT 2741.635 3429.770 2741.805 3429.940 ;
        RECT 2741.995 3429.770 2742.165 3429.940 ;
        RECT 2742.355 3429.770 2742.525 3429.940 ;
        RECT 2742.715 3429.770 2742.885 3429.940 ;
        RECT 2744.215 3429.770 2744.385 3429.940 ;
        RECT 2744.575 3429.770 2744.745 3429.940 ;
        RECT 2744.935 3429.770 2745.105 3429.940 ;
        RECT 2745.295 3429.770 2745.465 3429.940 ;
        RECT 2745.655 3429.770 2745.825 3429.940 ;
        RECT 2746.015 3429.770 2746.185 3429.940 ;
        RECT 2746.375 3429.770 2746.545 3429.940 ;
        RECT 2746.735 3429.770 2746.905 3429.940 ;
        RECT 2747.095 3429.770 2747.265 3429.940 ;
        RECT 2747.455 3429.770 2747.625 3429.940 ;
        RECT 2747.815 3429.770 2747.985 3429.940 ;
        RECT 2748.175 3429.770 2748.345 3429.940 ;
        RECT 2748.535 3429.770 2748.705 3429.940 ;
        RECT 2748.895 3429.770 2749.065 3429.940 ;
        RECT 2750.395 3429.770 2750.565 3429.940 ;
        RECT 2750.755 3429.770 2750.925 3429.940 ;
        RECT 2751.115 3429.770 2751.285 3429.940 ;
        RECT 2751.475 3429.770 2751.645 3429.940 ;
        RECT 2751.835 3429.770 2752.005 3429.940 ;
        RECT 2752.195 3429.770 2752.365 3429.940 ;
        RECT 2752.555 3429.770 2752.725 3429.940 ;
        RECT 2752.915 3429.770 2753.085 3429.940 ;
        RECT 2753.275 3429.770 2753.445 3429.940 ;
        RECT 2753.635 3429.770 2753.805 3429.940 ;
        RECT 2753.995 3429.770 2754.165 3429.940 ;
        RECT 2754.355 3429.770 2754.525 3429.940 ;
        RECT 2754.715 3429.770 2754.885 3429.940 ;
        RECT 2755.075 3429.770 2755.245 3429.940 ;
        RECT 2756.575 3429.770 2756.745 3429.940 ;
        RECT 2756.935 3429.770 2757.105 3429.940 ;
        RECT 2757.295 3429.770 2757.465 3429.940 ;
        RECT 2757.655 3429.770 2757.825 3429.940 ;
        RECT 2758.015 3429.770 2758.185 3429.940 ;
        RECT 2758.375 3429.770 2758.545 3429.940 ;
        RECT 2758.735 3429.770 2758.905 3429.940 ;
        RECT 2759.095 3429.770 2759.265 3429.940 ;
        RECT 2759.455 3429.770 2759.625 3429.940 ;
        RECT 2759.815 3429.770 2759.985 3429.940 ;
        RECT 2760.175 3429.770 2760.345 3429.940 ;
        RECT 2760.535 3429.770 2760.705 3429.940 ;
        RECT 2760.895 3429.770 2761.065 3429.940 ;
        RECT 2761.255 3429.770 2761.425 3429.940 ;
        RECT 2708.975 3428.045 2709.145 3428.215 ;
        RECT 2709.875 3428.095 2710.045 3428.265 ;
        RECT 2721.625 3428.045 2721.795 3428.215 ;
        RECT 2722.425 3428.045 2722.595 3428.215 ;
        RECT 2733.975 3428.045 2734.145 3428.215 ;
        RECT 2734.775 3428.045 2734.945 3428.215 ;
        RECT 2746.225 3428.045 2746.395 3428.215 ;
        RECT 2747.025 3428.045 2747.195 3428.215 ;
        RECT 2758.725 3428.045 2758.895 3428.215 ;
        RECT 2759.525 3428.045 2759.695 3428.215 ;
        RECT 2700.955 3427.070 2701.125 3427.240 ;
        RECT 2701.315 3427.070 2701.485 3427.240 ;
        RECT 2701.675 3427.070 2701.845 3427.240 ;
        RECT 2702.035 3427.070 2702.205 3427.240 ;
        RECT 2702.395 3427.070 2702.565 3427.240 ;
        RECT 2702.755 3427.070 2702.925 3427.240 ;
        RECT 2703.115 3427.070 2703.285 3427.240 ;
        RECT 2703.475 3427.070 2703.645 3427.240 ;
        RECT 2703.835 3427.070 2704.005 3427.240 ;
        RECT 2704.195 3427.070 2704.365 3427.240 ;
        RECT 2704.555 3427.070 2704.725 3427.240 ;
        RECT 2704.915 3427.070 2705.085 3427.240 ;
        RECT 2705.275 3427.070 2705.445 3427.240 ;
        RECT 2705.635 3427.070 2705.805 3427.240 ;
        RECT 2707.135 3427.070 2707.305 3427.240 ;
        RECT 2707.495 3427.070 2707.665 3427.240 ;
        RECT 2707.855 3427.070 2708.025 3427.240 ;
        RECT 2708.215 3427.070 2708.385 3427.240 ;
        RECT 2708.575 3427.070 2708.745 3427.240 ;
        RECT 2708.935 3427.070 2709.105 3427.240 ;
        RECT 2709.295 3427.070 2709.465 3427.240 ;
        RECT 2709.655 3427.070 2709.825 3427.240 ;
        RECT 2710.015 3427.070 2710.185 3427.240 ;
        RECT 2710.375 3427.070 2710.545 3427.240 ;
        RECT 2710.735 3427.070 2710.905 3427.240 ;
        RECT 2711.095 3427.070 2711.265 3427.240 ;
        RECT 2711.455 3427.070 2711.625 3427.240 ;
        RECT 2711.815 3427.070 2711.985 3427.240 ;
        RECT 2713.315 3427.070 2713.485 3427.240 ;
        RECT 2713.675 3427.070 2713.845 3427.240 ;
        RECT 2714.035 3427.070 2714.205 3427.240 ;
        RECT 2714.395 3427.070 2714.565 3427.240 ;
        RECT 2714.755 3427.070 2714.925 3427.240 ;
        RECT 2715.115 3427.070 2715.285 3427.240 ;
        RECT 2715.475 3427.070 2715.645 3427.240 ;
        RECT 2715.835 3427.070 2716.005 3427.240 ;
        RECT 2716.195 3427.070 2716.365 3427.240 ;
        RECT 2716.555 3427.070 2716.725 3427.240 ;
        RECT 2716.915 3427.070 2717.085 3427.240 ;
        RECT 2717.275 3427.070 2717.445 3427.240 ;
        RECT 2717.635 3427.070 2717.805 3427.240 ;
        RECT 2717.995 3427.070 2718.165 3427.240 ;
        RECT 2719.495 3427.070 2719.665 3427.240 ;
        RECT 2719.855 3427.070 2720.025 3427.240 ;
        RECT 2720.215 3427.070 2720.385 3427.240 ;
        RECT 2720.575 3427.070 2720.745 3427.240 ;
        RECT 2720.935 3427.070 2721.105 3427.240 ;
        RECT 2721.295 3427.070 2721.465 3427.240 ;
        RECT 2721.655 3427.070 2721.825 3427.240 ;
        RECT 2722.015 3427.070 2722.185 3427.240 ;
        RECT 2722.375 3427.070 2722.545 3427.240 ;
        RECT 2722.735 3427.070 2722.905 3427.240 ;
        RECT 2723.095 3427.070 2723.265 3427.240 ;
        RECT 2723.455 3427.070 2723.625 3427.240 ;
        RECT 2723.815 3427.070 2723.985 3427.240 ;
        RECT 2724.175 3427.070 2724.345 3427.240 ;
        RECT 2725.675 3427.070 2725.845 3427.240 ;
        RECT 2726.035 3427.070 2726.205 3427.240 ;
        RECT 2726.395 3427.070 2726.565 3427.240 ;
        RECT 2726.755 3427.070 2726.925 3427.240 ;
        RECT 2727.115 3427.070 2727.285 3427.240 ;
        RECT 2727.475 3427.070 2727.645 3427.240 ;
        RECT 2727.835 3427.070 2728.005 3427.240 ;
        RECT 2728.195 3427.070 2728.365 3427.240 ;
        RECT 2728.555 3427.070 2728.725 3427.240 ;
        RECT 2728.915 3427.070 2729.085 3427.240 ;
        RECT 2729.275 3427.070 2729.445 3427.240 ;
        RECT 2729.635 3427.070 2729.805 3427.240 ;
        RECT 2729.995 3427.070 2730.165 3427.240 ;
        RECT 2730.355 3427.070 2730.525 3427.240 ;
        RECT 2731.855 3427.070 2732.025 3427.240 ;
        RECT 2732.215 3427.070 2732.385 3427.240 ;
        RECT 2732.575 3427.070 2732.745 3427.240 ;
        RECT 2732.935 3427.070 2733.105 3427.240 ;
        RECT 2733.295 3427.070 2733.465 3427.240 ;
        RECT 2733.655 3427.070 2733.825 3427.240 ;
        RECT 2734.015 3427.070 2734.185 3427.240 ;
        RECT 2734.375 3427.070 2734.545 3427.240 ;
        RECT 2734.735 3427.070 2734.905 3427.240 ;
        RECT 2735.095 3427.070 2735.265 3427.240 ;
        RECT 2735.455 3427.070 2735.625 3427.240 ;
        RECT 2735.815 3427.070 2735.985 3427.240 ;
        RECT 2736.175 3427.070 2736.345 3427.240 ;
        RECT 2736.535 3427.070 2736.705 3427.240 ;
        RECT 2738.035 3427.070 2738.205 3427.240 ;
        RECT 2738.395 3427.070 2738.565 3427.240 ;
        RECT 2738.755 3427.070 2738.925 3427.240 ;
        RECT 2739.115 3427.070 2739.285 3427.240 ;
        RECT 2739.475 3427.070 2739.645 3427.240 ;
        RECT 2739.835 3427.070 2740.005 3427.240 ;
        RECT 2740.195 3427.070 2740.365 3427.240 ;
        RECT 2740.555 3427.070 2740.725 3427.240 ;
        RECT 2740.915 3427.070 2741.085 3427.240 ;
        RECT 2741.275 3427.070 2741.445 3427.240 ;
        RECT 2741.635 3427.070 2741.805 3427.240 ;
        RECT 2741.995 3427.070 2742.165 3427.240 ;
        RECT 2742.355 3427.070 2742.525 3427.240 ;
        RECT 2742.715 3427.070 2742.885 3427.240 ;
        RECT 2744.215 3427.070 2744.385 3427.240 ;
        RECT 2744.575 3427.070 2744.745 3427.240 ;
        RECT 2744.935 3427.070 2745.105 3427.240 ;
        RECT 2745.295 3427.070 2745.465 3427.240 ;
        RECT 2745.655 3427.070 2745.825 3427.240 ;
        RECT 2746.015 3427.070 2746.185 3427.240 ;
        RECT 2746.375 3427.070 2746.545 3427.240 ;
        RECT 2746.735 3427.070 2746.905 3427.240 ;
        RECT 2747.095 3427.070 2747.265 3427.240 ;
        RECT 2747.455 3427.070 2747.625 3427.240 ;
        RECT 2747.815 3427.070 2747.985 3427.240 ;
        RECT 2748.175 3427.070 2748.345 3427.240 ;
        RECT 2748.535 3427.070 2748.705 3427.240 ;
        RECT 2748.895 3427.070 2749.065 3427.240 ;
        RECT 2750.395 3427.070 2750.565 3427.240 ;
        RECT 2750.755 3427.070 2750.925 3427.240 ;
        RECT 2751.115 3427.070 2751.285 3427.240 ;
        RECT 2751.475 3427.070 2751.645 3427.240 ;
        RECT 2751.835 3427.070 2752.005 3427.240 ;
        RECT 2752.195 3427.070 2752.365 3427.240 ;
        RECT 2752.555 3427.070 2752.725 3427.240 ;
        RECT 2752.915 3427.070 2753.085 3427.240 ;
        RECT 2753.275 3427.070 2753.445 3427.240 ;
        RECT 2753.635 3427.070 2753.805 3427.240 ;
        RECT 2753.995 3427.070 2754.165 3427.240 ;
        RECT 2754.355 3427.070 2754.525 3427.240 ;
        RECT 2754.715 3427.070 2754.885 3427.240 ;
        RECT 2755.075 3427.070 2755.245 3427.240 ;
        RECT 2756.575 3427.070 2756.745 3427.240 ;
        RECT 2756.935 3427.070 2757.105 3427.240 ;
        RECT 2757.295 3427.070 2757.465 3427.240 ;
        RECT 2757.655 3427.070 2757.825 3427.240 ;
        RECT 2758.015 3427.070 2758.185 3427.240 ;
        RECT 2758.375 3427.070 2758.545 3427.240 ;
        RECT 2758.735 3427.070 2758.905 3427.240 ;
        RECT 2759.095 3427.070 2759.265 3427.240 ;
        RECT 2759.455 3427.070 2759.625 3427.240 ;
        RECT 2759.815 3427.070 2759.985 3427.240 ;
        RECT 2760.175 3427.070 2760.345 3427.240 ;
        RECT 2760.535 3427.070 2760.705 3427.240 ;
        RECT 2760.895 3427.070 2761.065 3427.240 ;
        RECT 2761.255 3427.070 2761.425 3427.240 ;
        RECT 2715.295 3404.745 2715.825 3405.275 ;
        RECT 2720.595 3404.745 2721.125 3405.275 ;
        RECT 2727.895 3404.745 2728.425 3405.275 ;
        RECT 2733.995 3404.745 2734.525 3405.275 ;
        RECT 2741.395 3404.745 2741.925 3405.275 ;
        RECT 2746.395 3404.745 2746.925 3405.275 ;
        RECT 2713.380 3404.200 2713.550 3404.370 ;
        RECT 2713.740 3404.200 2713.910 3404.370 ;
        RECT 2714.100 3404.200 2714.270 3404.370 ;
        RECT 2714.460 3404.200 2714.630 3404.370 ;
        RECT 2714.820 3404.200 2714.990 3404.370 ;
        RECT 2715.180 3404.200 2715.350 3404.370 ;
        RECT 2715.540 3404.200 2715.710 3404.370 ;
        RECT 2715.900 3404.200 2716.070 3404.370 ;
        RECT 2716.260 3404.200 2716.430 3404.370 ;
        RECT 2716.620 3404.200 2716.790 3404.370 ;
        RECT 2716.980 3404.200 2717.150 3404.370 ;
        RECT 2717.340 3404.200 2717.510 3404.370 ;
        RECT 2717.700 3404.200 2717.870 3404.370 ;
        RECT 2718.060 3404.200 2718.230 3404.370 ;
        RECT 2719.560 3404.200 2719.730 3404.370 ;
        RECT 2719.920 3404.200 2720.090 3404.370 ;
        RECT 2720.280 3404.200 2720.450 3404.370 ;
        RECT 2720.640 3404.200 2720.810 3404.370 ;
        RECT 2721.000 3404.200 2721.170 3404.370 ;
        RECT 2721.360 3404.200 2721.530 3404.370 ;
        RECT 2721.720 3404.200 2721.890 3404.370 ;
        RECT 2722.080 3404.200 2722.250 3404.370 ;
        RECT 2722.440 3404.200 2722.610 3404.370 ;
        RECT 2722.800 3404.200 2722.970 3404.370 ;
        RECT 2723.160 3404.200 2723.330 3404.370 ;
        RECT 2723.520 3404.200 2723.690 3404.370 ;
        RECT 2723.880 3404.200 2724.050 3404.370 ;
        RECT 2724.240 3404.200 2724.410 3404.370 ;
        RECT 2725.740 3404.200 2725.910 3404.370 ;
        RECT 2726.100 3404.200 2726.270 3404.370 ;
        RECT 2726.460 3404.200 2726.630 3404.370 ;
        RECT 2726.820 3404.200 2726.990 3404.370 ;
        RECT 2727.180 3404.200 2727.350 3404.370 ;
        RECT 2727.540 3404.200 2727.710 3404.370 ;
        RECT 2727.900 3404.200 2728.070 3404.370 ;
        RECT 2728.260 3404.200 2728.430 3404.370 ;
        RECT 2728.620 3404.200 2728.790 3404.370 ;
        RECT 2728.980 3404.200 2729.150 3404.370 ;
        RECT 2729.340 3404.200 2729.510 3404.370 ;
        RECT 2729.700 3404.200 2729.870 3404.370 ;
        RECT 2730.060 3404.200 2730.230 3404.370 ;
        RECT 2730.420 3404.200 2730.590 3404.370 ;
        RECT 2731.920 3404.200 2732.090 3404.370 ;
        RECT 2732.280 3404.200 2732.450 3404.370 ;
        RECT 2732.640 3404.200 2732.810 3404.370 ;
        RECT 2733.000 3404.200 2733.170 3404.370 ;
        RECT 2733.360 3404.200 2733.530 3404.370 ;
        RECT 2733.720 3404.200 2733.890 3404.370 ;
        RECT 2734.080 3404.200 2734.250 3404.370 ;
        RECT 2734.440 3404.200 2734.610 3404.370 ;
        RECT 2734.800 3404.200 2734.970 3404.370 ;
        RECT 2735.160 3404.200 2735.330 3404.370 ;
        RECT 2735.520 3404.200 2735.690 3404.370 ;
        RECT 2735.880 3404.200 2736.050 3404.370 ;
        RECT 2736.240 3404.200 2736.410 3404.370 ;
        RECT 2736.600 3404.200 2736.770 3404.370 ;
        RECT 2738.100 3404.200 2738.270 3404.370 ;
        RECT 2738.460 3404.200 2738.630 3404.370 ;
        RECT 2738.820 3404.200 2738.990 3404.370 ;
        RECT 2739.180 3404.200 2739.350 3404.370 ;
        RECT 2739.540 3404.200 2739.710 3404.370 ;
        RECT 2739.900 3404.200 2740.070 3404.370 ;
        RECT 2740.260 3404.200 2740.430 3404.370 ;
        RECT 2740.620 3404.200 2740.790 3404.370 ;
        RECT 2740.980 3404.200 2741.150 3404.370 ;
        RECT 2741.340 3404.200 2741.510 3404.370 ;
        RECT 2741.700 3404.200 2741.870 3404.370 ;
        RECT 2742.060 3404.200 2742.230 3404.370 ;
        RECT 2742.420 3404.200 2742.590 3404.370 ;
        RECT 2742.780 3404.200 2742.950 3404.370 ;
        RECT 2744.280 3404.200 2744.450 3404.370 ;
        RECT 2744.640 3404.200 2744.810 3404.370 ;
        RECT 2745.000 3404.200 2745.170 3404.370 ;
        RECT 2745.360 3404.200 2745.530 3404.370 ;
        RECT 2745.720 3404.200 2745.890 3404.370 ;
        RECT 2746.080 3404.200 2746.250 3404.370 ;
        RECT 2746.440 3404.200 2746.610 3404.370 ;
        RECT 2746.800 3404.200 2746.970 3404.370 ;
        RECT 2747.160 3404.200 2747.330 3404.370 ;
        RECT 2747.520 3404.200 2747.690 3404.370 ;
        RECT 2747.880 3404.200 2748.050 3404.370 ;
        RECT 2748.240 3404.200 2748.410 3404.370 ;
        RECT 2748.600 3404.200 2748.770 3404.370 ;
        RECT 2748.960 3404.200 2749.130 3404.370 ;
        RECT 2715.295 3401.845 2715.825 3402.375 ;
        RECT 2720.595 3401.845 2721.125 3402.375 ;
        RECT 2727.895 3401.845 2728.425 3402.375 ;
        RECT 2733.995 3401.845 2734.525 3402.375 ;
        RECT 2741.395 3401.845 2741.925 3402.375 ;
        RECT 2746.395 3401.845 2746.925 3402.375 ;
        RECT 2713.380 3401.250 2713.550 3401.420 ;
        RECT 2713.740 3401.250 2713.910 3401.420 ;
        RECT 2714.100 3401.250 2714.270 3401.420 ;
        RECT 2714.460 3401.250 2714.630 3401.420 ;
        RECT 2714.820 3401.250 2714.990 3401.420 ;
        RECT 2715.180 3401.250 2715.350 3401.420 ;
        RECT 2715.540 3401.250 2715.710 3401.420 ;
        RECT 2715.900 3401.250 2716.070 3401.420 ;
        RECT 2716.260 3401.250 2716.430 3401.420 ;
        RECT 2716.620 3401.250 2716.790 3401.420 ;
        RECT 2716.980 3401.250 2717.150 3401.420 ;
        RECT 2717.340 3401.250 2717.510 3401.420 ;
        RECT 2717.700 3401.250 2717.870 3401.420 ;
        RECT 2718.060 3401.250 2718.230 3401.420 ;
        RECT 2719.560 3401.250 2719.730 3401.420 ;
        RECT 2719.920 3401.250 2720.090 3401.420 ;
        RECT 2720.280 3401.250 2720.450 3401.420 ;
        RECT 2720.640 3401.250 2720.810 3401.420 ;
        RECT 2721.000 3401.250 2721.170 3401.420 ;
        RECT 2721.360 3401.250 2721.530 3401.420 ;
        RECT 2721.720 3401.250 2721.890 3401.420 ;
        RECT 2722.080 3401.250 2722.250 3401.420 ;
        RECT 2722.440 3401.250 2722.610 3401.420 ;
        RECT 2722.800 3401.250 2722.970 3401.420 ;
        RECT 2723.160 3401.250 2723.330 3401.420 ;
        RECT 2723.520 3401.250 2723.690 3401.420 ;
        RECT 2723.880 3401.250 2724.050 3401.420 ;
        RECT 2724.240 3401.250 2724.410 3401.420 ;
        RECT 2725.740 3401.250 2725.910 3401.420 ;
        RECT 2726.100 3401.250 2726.270 3401.420 ;
        RECT 2726.460 3401.250 2726.630 3401.420 ;
        RECT 2726.820 3401.250 2726.990 3401.420 ;
        RECT 2727.180 3401.250 2727.350 3401.420 ;
        RECT 2727.540 3401.250 2727.710 3401.420 ;
        RECT 2727.900 3401.250 2728.070 3401.420 ;
        RECT 2728.260 3401.250 2728.430 3401.420 ;
        RECT 2728.620 3401.250 2728.790 3401.420 ;
        RECT 2728.980 3401.250 2729.150 3401.420 ;
        RECT 2729.340 3401.250 2729.510 3401.420 ;
        RECT 2729.700 3401.250 2729.870 3401.420 ;
        RECT 2730.060 3401.250 2730.230 3401.420 ;
        RECT 2730.420 3401.250 2730.590 3401.420 ;
        RECT 2731.920 3401.250 2732.090 3401.420 ;
        RECT 2732.280 3401.250 2732.450 3401.420 ;
        RECT 2732.640 3401.250 2732.810 3401.420 ;
        RECT 2733.000 3401.250 2733.170 3401.420 ;
        RECT 2733.360 3401.250 2733.530 3401.420 ;
        RECT 2733.720 3401.250 2733.890 3401.420 ;
        RECT 2734.080 3401.250 2734.250 3401.420 ;
        RECT 2734.440 3401.250 2734.610 3401.420 ;
        RECT 2734.800 3401.250 2734.970 3401.420 ;
        RECT 2735.160 3401.250 2735.330 3401.420 ;
        RECT 2735.520 3401.250 2735.690 3401.420 ;
        RECT 2735.880 3401.250 2736.050 3401.420 ;
        RECT 2736.240 3401.250 2736.410 3401.420 ;
        RECT 2736.600 3401.250 2736.770 3401.420 ;
        RECT 2738.100 3401.250 2738.270 3401.420 ;
        RECT 2738.460 3401.250 2738.630 3401.420 ;
        RECT 2738.820 3401.250 2738.990 3401.420 ;
        RECT 2739.180 3401.250 2739.350 3401.420 ;
        RECT 2739.540 3401.250 2739.710 3401.420 ;
        RECT 2739.900 3401.250 2740.070 3401.420 ;
        RECT 2740.260 3401.250 2740.430 3401.420 ;
        RECT 2740.620 3401.250 2740.790 3401.420 ;
        RECT 2740.980 3401.250 2741.150 3401.420 ;
        RECT 2741.340 3401.250 2741.510 3401.420 ;
        RECT 2741.700 3401.250 2741.870 3401.420 ;
        RECT 2742.060 3401.250 2742.230 3401.420 ;
        RECT 2742.420 3401.250 2742.590 3401.420 ;
        RECT 2742.780 3401.250 2742.950 3401.420 ;
        RECT 2744.280 3401.250 2744.450 3401.420 ;
        RECT 2744.640 3401.250 2744.810 3401.420 ;
        RECT 2745.000 3401.250 2745.170 3401.420 ;
        RECT 2745.360 3401.250 2745.530 3401.420 ;
        RECT 2745.720 3401.250 2745.890 3401.420 ;
        RECT 2746.080 3401.250 2746.250 3401.420 ;
        RECT 2746.440 3401.250 2746.610 3401.420 ;
        RECT 2746.800 3401.250 2746.970 3401.420 ;
        RECT 2747.160 3401.250 2747.330 3401.420 ;
        RECT 2747.520 3401.250 2747.690 3401.420 ;
        RECT 2747.880 3401.250 2748.050 3401.420 ;
        RECT 2748.240 3401.250 2748.410 3401.420 ;
        RECT 2748.600 3401.250 2748.770 3401.420 ;
        RECT 2748.960 3401.250 2749.130 3401.420 ;
      LAYER met1 ;
        RECT 2718.025 3452.450 2718.595 3452.860 ;
        RECT 2718.875 3452.450 2719.445 3452.860 ;
        RECT 2730.475 3452.450 2731.045 3452.860 ;
        RECT 2731.325 3452.450 2731.895 3452.860 ;
        RECT 2742.775 3452.450 2743.295 3452.910 ;
        RECT 2743.625 3452.450 2744.145 3452.910 ;
        RECT 2718.035 3452.030 2718.535 3452.280 ;
        RECT 2718.885 3452.030 2719.385 3452.280 ;
        RECT 2730.485 3452.030 2730.985 3452.280 ;
        RECT 2731.335 3452.030 2731.835 3452.280 ;
        RECT 2742.785 3452.030 2743.285 3452.230 ;
        RECT 2743.635 3452.030 2744.135 3452.230 ;
        RECT 2710.035 3451.830 2752.235 3452.030 ;
        RECT 2710.080 3451.740 2715.080 3451.830 ;
        RECT 2716.260 3451.740 2721.260 3451.830 ;
        RECT 2722.440 3451.740 2727.440 3451.830 ;
        RECT 2728.620 3451.740 2733.620 3451.830 ;
        RECT 2734.800 3451.740 2739.800 3451.830 ;
        RECT 2740.980 3451.740 2745.980 3451.830 ;
        RECT 2747.160 3451.740 2752.160 3451.830 ;
        RECT 2718.035 3449.330 2718.535 3449.580 ;
        RECT 2718.885 3449.330 2719.385 3449.580 ;
        RECT 2730.485 3449.330 2730.985 3449.580 ;
        RECT 2731.335 3449.330 2731.835 3449.580 ;
        RECT 2742.785 3449.330 2743.285 3449.530 ;
        RECT 2743.635 3449.330 2744.135 3449.530 ;
        RECT 2710.035 3449.130 2752.235 3449.330 ;
        RECT 2710.080 3449.040 2715.080 3449.130 ;
        RECT 2716.260 3449.040 2721.260 3449.130 ;
        RECT 2722.440 3449.040 2727.440 3449.130 ;
        RECT 2728.620 3449.040 2733.620 3449.130 ;
        RECT 2734.800 3449.040 2739.800 3449.130 ;
        RECT 2740.980 3449.040 2745.980 3449.130 ;
        RECT 2747.160 3449.040 2752.160 3449.130 ;
        RECT 2718.085 3447.610 2719.385 3447.780 ;
        RECT 2718.075 3447.200 2719.385 3447.610 ;
        RECT 2730.475 3447.200 2731.045 3447.610 ;
        RECT 2731.275 3447.250 2731.845 3447.660 ;
        RECT 2742.775 3447.250 2743.295 3447.660 ;
        RECT 2743.625 3447.250 2744.145 3447.660 ;
        RECT 2718.085 3447.030 2719.385 3447.200 ;
        RECT 2718.035 3446.630 2718.535 3446.880 ;
        RECT 2718.885 3446.630 2719.385 3446.880 ;
        RECT 2730.485 3446.630 2730.985 3446.930 ;
        RECT 2731.335 3446.630 2731.835 3446.930 ;
        RECT 2742.785 3446.630 2743.285 3446.830 ;
        RECT 2743.635 3446.630 2744.135 3446.830 ;
        RECT 2710.035 3446.430 2752.235 3446.630 ;
        RECT 2710.080 3446.340 2715.080 3446.430 ;
        RECT 2716.260 3446.340 2721.260 3446.430 ;
        RECT 2722.440 3446.340 2727.440 3446.430 ;
        RECT 2728.620 3446.340 2733.620 3446.430 ;
        RECT 2734.800 3446.340 2739.800 3446.430 ;
        RECT 2740.980 3446.340 2745.980 3446.430 ;
        RECT 2747.160 3446.340 2752.160 3446.430 ;
        RECT 2718.075 3444.500 2718.595 3444.960 ;
        RECT 2718.925 3444.500 2719.445 3444.960 ;
        RECT 2730.475 3444.500 2730.995 3444.960 ;
        RECT 2731.325 3444.500 2731.845 3444.960 ;
        RECT 2742.775 3444.500 2743.295 3444.960 ;
        RECT 2743.625 3444.500 2744.145 3444.960 ;
        RECT 2718.085 3443.980 2718.585 3444.280 ;
        RECT 2718.935 3443.980 2719.435 3444.280 ;
        RECT 2730.485 3443.980 2730.985 3444.330 ;
        RECT 2731.335 3443.980 2731.835 3444.330 ;
        RECT 2742.785 3443.980 2743.285 3444.280 ;
        RECT 2743.635 3443.980 2744.135 3444.280 ;
        RECT 2710.085 3443.870 2752.285 3443.980 ;
        RECT 2710.080 3443.780 2752.285 3443.870 ;
        RECT 2710.080 3443.640 2715.080 3443.780 ;
        RECT 2716.260 3443.640 2721.260 3443.780 ;
        RECT 2722.440 3443.640 2727.440 3443.780 ;
        RECT 2728.620 3443.640 2733.620 3443.780 ;
        RECT 2734.800 3443.640 2739.800 3443.780 ;
        RECT 2740.980 3443.640 2745.980 3443.780 ;
        RECT 2747.160 3443.640 2752.160 3443.780 ;
        RECT 2718.085 3441.080 2718.585 3441.380 ;
        RECT 2718.935 3441.080 2719.435 3441.380 ;
        RECT 2730.485 3441.080 2730.985 3441.430 ;
        RECT 2731.335 3441.080 2731.835 3441.430 ;
        RECT 2742.785 3441.080 2743.285 3441.380 ;
        RECT 2743.635 3441.080 2744.135 3441.380 ;
        RECT 2710.035 3440.880 2752.235 3441.080 ;
        RECT 2710.080 3440.740 2715.080 3440.880 ;
        RECT 2716.260 3440.740 2721.260 3440.880 ;
        RECT 2722.440 3440.740 2727.440 3440.880 ;
        RECT 2728.620 3440.740 2733.620 3440.880 ;
        RECT 2734.800 3440.740 2739.800 3440.880 ;
        RECT 2740.980 3440.740 2745.980 3440.880 ;
        RECT 2747.160 3440.740 2752.160 3440.880 ;
        RECT 2718.075 3438.700 2718.645 3439.160 ;
        RECT 2718.875 3438.700 2719.445 3439.160 ;
        RECT 2730.475 3438.700 2730.995 3439.110 ;
        RECT 2731.325 3438.700 2731.845 3439.110 ;
        RECT 2742.775 3438.700 2743.295 3439.110 ;
        RECT 2743.625 3438.700 2744.145 3439.110 ;
        RECT 2718.085 3438.180 2718.585 3438.480 ;
        RECT 2718.935 3438.180 2719.435 3438.480 ;
        RECT 2730.485 3438.180 2730.985 3438.530 ;
        RECT 2731.335 3438.180 2731.835 3438.530 ;
        RECT 2742.785 3438.180 2743.285 3438.480 ;
        RECT 2743.635 3438.180 2744.135 3438.480 ;
        RECT 2710.035 3437.980 2752.235 3438.180 ;
        RECT 2710.080 3437.840 2715.080 3437.980 ;
        RECT 2716.260 3437.840 2721.260 3437.980 ;
        RECT 2722.440 3437.840 2727.440 3437.980 ;
        RECT 2728.620 3437.840 2733.620 3437.980 ;
        RECT 2734.800 3437.840 2739.800 3437.980 ;
        RECT 2740.980 3437.840 2745.980 3437.980 ;
        RECT 2747.160 3437.840 2752.160 3437.980 ;
        RECT 2708.685 3435.480 2709.185 3435.830 ;
        RECT 2709.835 3435.480 2710.335 3435.830 ;
        RECT 2721.435 3435.480 2721.935 3435.780 ;
        RECT 2722.285 3435.480 2722.785 3435.780 ;
        RECT 2733.735 3435.480 2734.235 3435.780 ;
        RECT 2734.685 3435.480 2735.185 3435.780 ;
        RECT 2745.985 3435.480 2746.485 3435.780 ;
        RECT 2746.935 3435.480 2747.435 3435.780 ;
        RECT 2758.535 3435.480 2759.035 3435.780 ;
        RECT 2759.385 3435.480 2759.885 3435.780 ;
        RECT 2700.835 3435.230 2761.585 3435.480 ;
        RECT 2700.880 3435.140 2705.880 3435.230 ;
        RECT 2707.060 3435.140 2712.060 3435.230 ;
        RECT 2713.240 3435.140 2718.240 3435.230 ;
        RECT 2719.420 3435.140 2724.420 3435.230 ;
        RECT 2725.600 3435.140 2730.600 3435.230 ;
        RECT 2731.780 3435.140 2736.780 3435.230 ;
        RECT 2737.960 3435.140 2742.960 3435.230 ;
        RECT 2744.140 3435.140 2749.140 3435.230 ;
        RECT 2750.320 3435.140 2755.320 3435.230 ;
        RECT 2756.500 3435.140 2761.500 3435.230 ;
        RECT 2708.775 3433.300 2709.345 3433.760 ;
        RECT 2709.675 3433.300 2710.245 3433.760 ;
        RECT 2721.425 3433.300 2721.995 3433.760 ;
        RECT 2722.225 3433.300 2722.795 3433.760 ;
        RECT 2733.775 3433.300 2734.345 3433.760 ;
        RECT 2734.575 3433.300 2735.145 3433.760 ;
        RECT 2746.025 3433.300 2746.595 3433.760 ;
        RECT 2746.825 3433.300 2747.395 3433.760 ;
        RECT 2758.525 3433.300 2759.095 3433.760 ;
        RECT 2759.325 3433.300 2759.895 3433.760 ;
        RECT 2708.685 3432.830 2709.185 3433.130 ;
        RECT 2709.835 3432.830 2710.335 3433.130 ;
        RECT 2721.435 3432.830 2721.935 3433.080 ;
        RECT 2722.285 3432.830 2722.785 3433.130 ;
        RECT 2733.735 3432.830 2734.235 3433.130 ;
        RECT 2734.685 3432.830 2735.185 3433.130 ;
        RECT 2745.985 3432.830 2746.485 3433.080 ;
        RECT 2746.935 3432.830 2747.435 3433.080 ;
        RECT 2758.535 3432.830 2759.035 3433.080 ;
        RECT 2759.385 3432.830 2759.885 3433.080 ;
        RECT 2700.835 3432.580 2761.585 3432.830 ;
        RECT 2700.880 3432.440 2705.880 3432.580 ;
        RECT 2707.060 3432.440 2712.060 3432.580 ;
        RECT 2713.240 3432.440 2718.240 3432.580 ;
        RECT 2719.420 3432.440 2724.420 3432.580 ;
        RECT 2725.600 3432.440 2730.600 3432.580 ;
        RECT 2731.780 3432.440 2736.780 3432.580 ;
        RECT 2737.960 3432.440 2742.960 3432.580 ;
        RECT 2744.140 3432.440 2749.140 3432.580 ;
        RECT 2750.320 3432.440 2755.320 3432.580 ;
        RECT 2756.500 3432.440 2761.500 3432.580 ;
        RECT 2708.685 3430.130 2709.185 3430.430 ;
        RECT 2709.835 3430.130 2710.335 3430.430 ;
        RECT 2721.385 3430.130 2721.885 3430.380 ;
        RECT 2722.235 3430.130 2722.735 3430.380 ;
        RECT 2733.735 3430.130 2734.235 3430.380 ;
        RECT 2734.635 3430.130 2735.135 3430.380 ;
        RECT 2745.985 3430.130 2746.485 3430.380 ;
        RECT 2746.935 3430.130 2747.435 3430.380 ;
        RECT 2758.535 3430.130 2759.035 3430.380 ;
        RECT 2759.385 3430.130 2759.885 3430.380 ;
        RECT 2700.835 3429.880 2761.585 3430.130 ;
        RECT 2700.880 3429.740 2705.880 3429.880 ;
        RECT 2707.060 3429.740 2712.060 3429.880 ;
        RECT 2713.240 3429.740 2718.240 3429.880 ;
        RECT 2719.420 3429.740 2724.420 3429.880 ;
        RECT 2725.600 3429.740 2730.600 3429.880 ;
        RECT 2731.780 3429.740 2736.780 3429.880 ;
        RECT 2737.960 3429.740 2742.960 3429.880 ;
        RECT 2744.140 3429.740 2749.140 3429.880 ;
        RECT 2750.320 3429.740 2755.320 3429.880 ;
        RECT 2756.500 3429.740 2761.500 3429.880 ;
        RECT 2708.775 3427.900 2709.345 3428.360 ;
        RECT 2709.675 3427.950 2710.245 3428.410 ;
        RECT 2721.425 3427.900 2721.995 3428.360 ;
        RECT 2722.225 3427.900 2722.795 3428.360 ;
        RECT 2733.775 3427.900 2734.345 3428.360 ;
        RECT 2734.575 3427.900 2735.145 3428.360 ;
        RECT 2746.025 3427.900 2746.595 3428.360 ;
        RECT 2746.825 3427.900 2747.395 3428.360 ;
        RECT 2758.525 3427.900 2759.095 3428.360 ;
        RECT 2759.325 3427.900 2759.895 3428.360 ;
        RECT 2708.685 3427.430 2709.185 3427.680 ;
        RECT 2709.835 3427.430 2710.335 3427.680 ;
        RECT 2721.335 3427.430 2721.835 3427.730 ;
        RECT 2722.285 3427.430 2722.785 3427.730 ;
        RECT 2733.735 3427.430 2734.235 3427.680 ;
        RECT 2734.685 3427.430 2735.185 3427.680 ;
        RECT 2745.985 3427.430 2746.485 3427.680 ;
        RECT 2746.935 3427.430 2747.435 3427.680 ;
        RECT 2758.535 3427.430 2759.035 3427.630 ;
        RECT 2759.385 3427.430 2759.885 3427.630 ;
        RECT 2700.835 3427.180 2761.585 3427.430 ;
        RECT 2700.880 3427.040 2705.880 3427.180 ;
        RECT 2707.060 3427.040 2712.060 3427.180 ;
        RECT 2713.240 3427.040 2718.240 3427.180 ;
        RECT 2719.420 3427.040 2724.420 3427.180 ;
        RECT 2725.600 3427.040 2730.600 3427.180 ;
        RECT 2731.780 3427.040 2736.780 3427.180 ;
        RECT 2737.960 3427.040 2742.960 3427.180 ;
        RECT 2744.140 3427.040 2749.140 3427.180 ;
        RECT 2750.320 3427.040 2755.320 3427.180 ;
        RECT 2756.500 3427.040 2761.500 3427.180 ;
        RECT 2715.100 3405.410 2716.020 3405.440 ;
        RECT 2720.400 3405.410 2721.320 3405.440 ;
        RECT 2727.700 3405.410 2728.620 3405.440 ;
        RECT 2733.800 3405.410 2734.720 3405.440 ;
        RECT 2741.200 3405.410 2742.120 3405.440 ;
        RECT 2746.200 3405.410 2747.120 3405.440 ;
        RECT 2713.260 3404.310 2749.260 3405.410 ;
        RECT 2713.260 3404.110 2718.360 3404.310 ;
        RECT 2719.460 3404.170 2724.485 3404.310 ;
        RECT 2725.660 3404.170 2730.665 3404.310 ;
        RECT 2731.845 3404.170 2736.860 3404.310 ;
        RECT 2719.460 3404.110 2724.460 3404.170 ;
        RECT 2725.660 3404.110 2730.660 3404.170 ;
        RECT 2731.860 3404.110 2736.860 3404.170 ;
        RECT 2737.960 3404.110 2743.060 3404.310 ;
        RECT 2744.160 3404.110 2749.260 3404.310 ;
        RECT 2715.100 3402.510 2716.020 3402.540 ;
        RECT 2720.400 3402.510 2721.320 3402.540 ;
        RECT 2727.700 3402.510 2728.620 3402.540 ;
        RECT 2733.800 3402.510 2734.720 3402.540 ;
        RECT 2741.200 3402.510 2742.120 3402.540 ;
        RECT 2746.200 3402.510 2747.120 3402.540 ;
        RECT 2713.260 3401.360 2749.260 3402.510 ;
        RECT 2713.260 3401.310 2718.305 3401.360 ;
        RECT 2713.305 3401.220 2718.305 3401.310 ;
        RECT 2719.485 3401.220 2724.485 3401.360 ;
        RECT 2725.665 3401.220 2730.665 3401.360 ;
        RECT 2731.845 3401.220 2736.845 3401.360 ;
        RECT 2738.025 3401.220 2743.025 3401.360 ;
        RECT 2744.205 3401.310 2749.260 3401.360 ;
        RECT 2744.205 3401.220 2749.205 3401.310 ;
      LAYER via ;
        RECT 2718.180 3452.525 2718.440 3452.785 ;
        RECT 2719.030 3452.525 2719.290 3452.785 ;
        RECT 2730.630 3452.525 2730.890 3452.785 ;
        RECT 2731.480 3452.525 2731.740 3452.785 ;
        RECT 2742.905 3452.550 2743.165 3452.810 ;
        RECT 2743.755 3452.550 2744.015 3452.810 ;
        RECT 2718.155 3451.950 2718.415 3452.210 ;
        RECT 2719.005 3451.950 2719.265 3452.210 ;
        RECT 2730.605 3451.950 2730.865 3452.210 ;
        RECT 2731.455 3451.950 2731.715 3452.210 ;
        RECT 2742.905 3451.900 2743.165 3452.160 ;
        RECT 2743.755 3451.900 2744.015 3452.160 ;
        RECT 2718.155 3449.250 2718.415 3449.510 ;
        RECT 2719.005 3449.250 2719.265 3449.510 ;
        RECT 2730.605 3449.250 2730.865 3449.510 ;
        RECT 2731.455 3449.250 2731.715 3449.510 ;
        RECT 2742.905 3449.200 2743.165 3449.460 ;
        RECT 2743.755 3449.200 2744.015 3449.460 ;
        RECT 2718.230 3447.275 2718.490 3447.535 ;
        RECT 2718.930 3447.275 2719.190 3447.535 ;
        RECT 2730.630 3447.275 2730.890 3447.535 ;
        RECT 2731.430 3447.325 2731.690 3447.585 ;
        RECT 2742.905 3447.325 2743.165 3447.585 ;
        RECT 2743.755 3447.325 2744.015 3447.585 ;
        RECT 2718.155 3446.550 2718.415 3446.810 ;
        RECT 2719.005 3446.550 2719.265 3446.810 ;
        RECT 2730.605 3446.600 2730.865 3446.860 ;
        RECT 2731.455 3446.600 2731.715 3446.860 ;
        RECT 2742.905 3446.500 2743.165 3446.760 ;
        RECT 2743.755 3446.500 2744.015 3446.760 ;
        RECT 2718.205 3444.600 2718.465 3444.860 ;
        RECT 2719.055 3444.600 2719.315 3444.860 ;
        RECT 2730.605 3444.600 2730.865 3444.860 ;
        RECT 2731.455 3444.600 2731.715 3444.860 ;
        RECT 2742.905 3444.600 2743.165 3444.860 ;
        RECT 2743.755 3444.600 2744.015 3444.860 ;
        RECT 2718.205 3443.950 2718.465 3444.210 ;
        RECT 2719.055 3443.950 2719.315 3444.210 ;
        RECT 2730.605 3444.000 2730.865 3444.260 ;
        RECT 2731.455 3444.000 2731.715 3444.260 ;
        RECT 2742.905 3443.950 2743.165 3444.210 ;
        RECT 2743.755 3443.950 2744.015 3444.210 ;
        RECT 2718.205 3441.050 2718.465 3441.310 ;
        RECT 2719.055 3441.050 2719.315 3441.310 ;
        RECT 2730.605 3441.100 2730.865 3441.360 ;
        RECT 2731.455 3441.100 2731.715 3441.360 ;
        RECT 2742.905 3441.050 2743.165 3441.310 ;
        RECT 2743.755 3441.050 2744.015 3441.310 ;
        RECT 2718.230 3438.800 2718.490 3439.060 ;
        RECT 2719.030 3438.800 2719.290 3439.060 ;
        RECT 2730.605 3438.775 2730.865 3439.035 ;
        RECT 2731.455 3438.775 2731.715 3439.035 ;
        RECT 2742.905 3438.775 2743.165 3439.035 ;
        RECT 2743.755 3438.775 2744.015 3439.035 ;
        RECT 2718.205 3438.150 2718.465 3438.410 ;
        RECT 2719.055 3438.150 2719.315 3438.410 ;
        RECT 2730.605 3438.200 2730.865 3438.460 ;
        RECT 2731.455 3438.200 2731.715 3438.460 ;
        RECT 2742.905 3438.150 2743.165 3438.410 ;
        RECT 2743.755 3438.150 2744.015 3438.410 ;
        RECT 2708.805 3435.500 2709.065 3435.760 ;
        RECT 2709.955 3435.500 2710.215 3435.760 ;
        RECT 2721.555 3435.450 2721.815 3435.710 ;
        RECT 2722.405 3435.450 2722.665 3435.710 ;
        RECT 2733.855 3435.450 2734.115 3435.710 ;
        RECT 2734.805 3435.450 2735.065 3435.710 ;
        RECT 2746.105 3435.450 2746.365 3435.710 ;
        RECT 2747.055 3435.450 2747.315 3435.710 ;
        RECT 2758.655 3435.450 2758.915 3435.710 ;
        RECT 2759.505 3435.450 2759.765 3435.710 ;
        RECT 2708.930 3433.400 2709.190 3433.660 ;
        RECT 2709.830 3433.400 2710.090 3433.660 ;
        RECT 2721.580 3433.400 2721.840 3433.660 ;
        RECT 2722.380 3433.400 2722.640 3433.660 ;
        RECT 2733.930 3433.400 2734.190 3433.660 ;
        RECT 2734.730 3433.400 2734.990 3433.660 ;
        RECT 2746.180 3433.400 2746.440 3433.660 ;
        RECT 2746.980 3433.400 2747.240 3433.660 ;
        RECT 2758.680 3433.400 2758.940 3433.660 ;
        RECT 2759.480 3433.400 2759.740 3433.660 ;
        RECT 2708.805 3432.800 2709.065 3433.060 ;
        RECT 2709.955 3432.800 2710.215 3433.060 ;
        RECT 2721.555 3432.750 2721.815 3433.010 ;
        RECT 2722.405 3432.800 2722.665 3433.060 ;
        RECT 2733.855 3432.800 2734.115 3433.060 ;
        RECT 2734.805 3432.800 2735.065 3433.060 ;
        RECT 2746.105 3432.750 2746.365 3433.010 ;
        RECT 2747.055 3432.750 2747.315 3433.010 ;
        RECT 2758.655 3432.750 2758.915 3433.010 ;
        RECT 2759.505 3432.750 2759.765 3433.010 ;
        RECT 2708.805 3430.100 2709.065 3430.360 ;
        RECT 2709.955 3430.100 2710.215 3430.360 ;
        RECT 2721.505 3430.050 2721.765 3430.310 ;
        RECT 2722.355 3430.050 2722.615 3430.310 ;
        RECT 2733.855 3430.050 2734.115 3430.310 ;
        RECT 2734.755 3430.050 2735.015 3430.310 ;
        RECT 2746.105 3430.050 2746.365 3430.310 ;
        RECT 2747.055 3430.050 2747.315 3430.310 ;
        RECT 2758.655 3430.050 2758.915 3430.310 ;
        RECT 2759.505 3430.050 2759.765 3430.310 ;
        RECT 2708.930 3428.000 2709.190 3428.260 ;
        RECT 2709.830 3428.050 2710.090 3428.310 ;
        RECT 2721.580 3428.000 2721.840 3428.260 ;
        RECT 2722.380 3428.000 2722.640 3428.260 ;
        RECT 2733.930 3428.000 2734.190 3428.260 ;
        RECT 2734.730 3428.000 2734.990 3428.260 ;
        RECT 2746.180 3428.000 2746.440 3428.260 ;
        RECT 2746.980 3428.000 2747.240 3428.260 ;
        RECT 2758.680 3428.000 2758.940 3428.260 ;
        RECT 2759.480 3428.000 2759.740 3428.260 ;
        RECT 2708.805 3427.350 2709.065 3427.610 ;
        RECT 2709.955 3427.350 2710.215 3427.610 ;
        RECT 2721.455 3427.400 2721.715 3427.660 ;
        RECT 2722.405 3427.400 2722.665 3427.660 ;
        RECT 2733.855 3427.350 2734.115 3427.610 ;
        RECT 2734.805 3427.350 2735.065 3427.610 ;
        RECT 2746.105 3427.350 2746.365 3427.610 ;
        RECT 2747.055 3427.350 2747.315 3427.610 ;
        RECT 2758.655 3427.300 2758.915 3427.560 ;
        RECT 2759.505 3427.300 2759.765 3427.560 ;
        RECT 2715.270 3404.720 2715.850 3405.300 ;
        RECT 2720.570 3404.720 2721.150 3405.300 ;
        RECT 2727.870 3404.720 2728.450 3405.300 ;
        RECT 2733.970 3404.720 2734.550 3405.300 ;
        RECT 2741.370 3404.720 2741.950 3405.300 ;
        RECT 2746.370 3404.720 2746.950 3405.300 ;
        RECT 2715.270 3401.820 2715.850 3402.400 ;
        RECT 2720.570 3401.820 2721.150 3402.400 ;
        RECT 2727.870 3401.820 2728.450 3402.400 ;
        RECT 2733.970 3401.820 2734.550 3402.400 ;
        RECT 2741.370 3401.820 2741.950 3402.400 ;
        RECT 2746.370 3401.820 2746.950 3402.400 ;
      LAYER met2 ;
        RECT 2717.985 3446.430 2719.435 3452.930 ;
        RECT 2730.435 3446.430 2731.885 3452.930 ;
        RECT 2742.735 3445.180 2744.185 3453.080 ;
        RECT 2718.135 3444.480 2718.535 3444.980 ;
        RECT 2718.985 3444.480 2719.385 3444.980 ;
        RECT 2730.535 3444.530 2730.935 3444.980 ;
        RECT 2731.385 3444.530 2731.785 3444.980 ;
        RECT 2742.835 3444.530 2743.235 3444.980 ;
        RECT 2743.685 3444.530 2744.085 3444.980 ;
        RECT 2718.035 3437.980 2719.485 3444.480 ;
        RECT 2730.435 3438.030 2731.885 3444.530 ;
        RECT 2742.735 3438.030 2744.185 3444.530 ;
        RECT 2708.735 3427.230 2710.285 3435.930 ;
        RECT 2721.385 3427.180 2722.835 3435.930 ;
        RECT 2733.735 3427.230 2735.185 3435.980 ;
        RECT 2745.985 3426.030 2747.435 3435.930 ;
        RECT 2758.485 3427.130 2759.935 3435.880 ;
        RECT 2715.160 3404.560 2715.960 3405.460 ;
        RECT 2720.460 3404.560 2721.260 3405.460 ;
        RECT 2727.760 3404.560 2728.560 3405.460 ;
        RECT 2733.860 3404.560 2734.660 3405.460 ;
        RECT 2741.260 3404.560 2742.060 3405.460 ;
        RECT 2746.260 3404.560 2747.060 3405.460 ;
        RECT 2715.160 3401.660 2715.960 3402.560 ;
        RECT 2720.460 3401.660 2721.260 3402.560 ;
        RECT 2727.760 3401.660 2728.560 3402.560 ;
        RECT 2733.860 3401.660 2734.660 3402.560 ;
        RECT 2741.260 3401.660 2742.060 3402.560 ;
        RECT 2746.260 3401.660 2747.060 3402.560 ;
      LAYER via2 ;
        RECT 2718.170 3452.515 2718.450 3452.795 ;
        RECT 2719.020 3452.515 2719.300 3452.795 ;
        RECT 2718.220 3447.265 2718.500 3447.545 ;
        RECT 2718.920 3447.265 2719.200 3447.545 ;
        RECT 2730.620 3452.515 2730.900 3452.795 ;
        RECT 2731.470 3452.515 2731.750 3452.795 ;
        RECT 2730.620 3447.265 2730.900 3447.545 ;
        RECT 2731.420 3447.315 2731.700 3447.595 ;
        RECT 2742.895 3452.540 2743.175 3452.820 ;
        RECT 2743.745 3452.540 2744.025 3452.820 ;
        RECT 2742.895 3447.315 2743.175 3447.595 ;
        RECT 2743.745 3447.315 2744.025 3447.595 ;
        RECT 2718.195 3444.590 2718.475 3444.870 ;
        RECT 2719.045 3444.590 2719.325 3444.870 ;
        RECT 2730.595 3444.590 2730.875 3444.870 ;
        RECT 2731.445 3444.590 2731.725 3444.870 ;
        RECT 2742.895 3444.590 2743.175 3444.870 ;
        RECT 2743.745 3444.590 2744.025 3444.870 ;
        RECT 2718.220 3438.790 2718.500 3439.070 ;
        RECT 2719.020 3438.790 2719.300 3439.070 ;
        RECT 2730.595 3438.765 2730.875 3439.045 ;
        RECT 2731.445 3438.765 2731.725 3439.045 ;
        RECT 2742.895 3438.765 2743.175 3439.045 ;
        RECT 2743.745 3438.765 2744.025 3439.045 ;
        RECT 2708.920 3433.390 2709.200 3433.670 ;
        RECT 2709.820 3433.390 2710.100 3433.670 ;
        RECT 2708.920 3427.990 2709.200 3428.270 ;
        RECT 2709.820 3428.040 2710.100 3428.320 ;
        RECT 2721.570 3433.390 2721.850 3433.670 ;
        RECT 2722.370 3433.390 2722.650 3433.670 ;
        RECT 2721.570 3427.990 2721.850 3428.270 ;
        RECT 2722.370 3427.990 2722.650 3428.270 ;
        RECT 2733.920 3433.390 2734.200 3433.670 ;
        RECT 2734.720 3433.390 2735.000 3433.670 ;
        RECT 2733.920 3427.990 2734.200 3428.270 ;
        RECT 2734.720 3427.990 2735.000 3428.270 ;
        RECT 2746.170 3433.390 2746.450 3433.670 ;
        RECT 2746.970 3433.390 2747.250 3433.670 ;
        RECT 2746.170 3427.990 2746.450 3428.270 ;
        RECT 2746.970 3427.990 2747.250 3428.270 ;
        RECT 2758.670 3433.390 2758.950 3433.670 ;
        RECT 2759.470 3433.390 2759.750 3433.670 ;
        RECT 2758.670 3427.990 2758.950 3428.270 ;
        RECT 2759.470 3427.990 2759.750 3428.270 ;
        RECT 2715.220 3404.670 2715.900 3405.350 ;
        RECT 2720.520 3404.670 2721.200 3405.350 ;
        RECT 2727.820 3404.670 2728.500 3405.350 ;
        RECT 2733.920 3404.670 2734.600 3405.350 ;
        RECT 2741.320 3404.670 2742.000 3405.350 ;
        RECT 2746.320 3404.670 2747.000 3405.350 ;
        RECT 2715.220 3401.770 2715.900 3402.450 ;
        RECT 2720.520 3401.770 2721.200 3402.450 ;
        RECT 2727.820 3401.770 2728.500 3402.450 ;
        RECT 2733.920 3401.770 2734.600 3402.450 ;
        RECT 2741.320 3401.770 2742.000 3402.450 ;
        RECT 2746.320 3401.770 2747.000 3402.450 ;
      LAYER met3 ;
        RECT 2707.835 3452.280 2765.735 3454.080 ;
        RECT 2763.685 3447.930 2765.735 3452.280 ;
        RECT 2706.635 3446.780 2765.735 3447.930 ;
        RECT 2763.685 3444.980 2765.735 3446.780 ;
        RECT 2708.585 3443.880 2765.735 3444.980 ;
        RECT 2763.685 3439.180 2765.735 3443.880 ;
        RECT 2708.185 3438.280 2765.735 3439.180 ;
        RECT 2763.685 3434.630 2765.735 3438.280 ;
        RECT 2697.435 3432.830 2765.735 3434.630 ;
        RECT 2763.685 3428.980 2765.735 3432.830 ;
        RECT 2699.285 3427.280 2765.735 3428.980 ;
        RECT 2714.960 3401.610 2747.260 3407.710 ;
        RECT 2895.000 3223.000 2912.000 3223.500 ;
        RECT 2755.000 3222.920 2912.000 3223.000 ;
        RECT 2755.000 3198.920 2924.000 3222.920 ;
        RECT 2755.000 3172.920 2912.000 3198.920 ;
        RECT 2755.000 3149.000 2924.000 3172.920 ;
        RECT 2755.000 3148.500 2899.000 3149.000 ;
        RECT 2911.700 3148.920 2924.000 3149.000 ;
      LAYER via3 ;
        RECT 2756.000 3433.000 2757.000 3434.000 ;
        RECT 2758.000 3433.000 2759.000 3434.000 ;
        RECT 2760.000 3433.000 2761.000 3434.000 ;
        RECT 2762.000 3433.000 2763.000 3434.000 ;
        RECT 2764.000 3433.000 2765.000 3434.000 ;
        RECT 2756.000 3427.500 2757.000 3428.500 ;
        RECT 2758.000 3427.500 2759.000 3428.500 ;
        RECT 2760.000 3427.500 2761.000 3428.500 ;
        RECT 2762.000 3427.500 2763.000 3428.500 ;
        RECT 2764.095 3427.700 2765.215 3428.420 ;
        RECT 2735.000 3404.000 2736.000 3405.000 ;
        RECT 2737.000 3404.000 2738.000 3405.000 ;
        RECT 2739.000 3404.000 2740.000 3405.000 ;
        RECT 2741.000 3404.000 2742.000 3405.000 ;
        RECT 2743.000 3404.000 2744.000 3405.000 ;
        RECT 2745.000 3404.000 2746.000 3405.000 ;
        RECT 2735.000 3402.500 2736.000 3403.500 ;
        RECT 2737.000 3402.500 2738.000 3403.500 ;
        RECT 2739.000 3402.500 2740.000 3403.500 ;
        RECT 2741.000 3402.500 2742.000 3403.500 ;
        RECT 2743.000 3402.500 2744.000 3403.500 ;
        RECT 2745.455 3403.200 2745.775 3403.520 ;
        RECT 2756.000 3214.000 2760.000 3218.000 ;
        RECT 2765.000 3214.000 2769.000 3218.000 ;
        RECT 2756.000 3206.000 2760.000 3210.000 ;
        RECT 2765.000 3206.000 2769.000 3210.000 ;
        RECT 2756.000 3198.000 2760.000 3202.000 ;
        RECT 2765.000 3198.000 2769.000 3202.000 ;
        RECT 2756.000 3190.000 2760.000 3194.000 ;
        RECT 2765.000 3190.000 2769.000 3194.000 ;
        RECT 2756.000 3182.000 2760.000 3186.000 ;
        RECT 2765.000 3182.000 2769.000 3186.000 ;
        RECT 2756.000 3174.000 2760.000 3178.000 ;
        RECT 2765.000 3174.000 2769.000 3178.000 ;
        RECT 2756.000 3166.000 2760.000 3170.000 ;
        RECT 2765.000 3166.000 2769.000 3170.000 ;
        RECT 2756.000 3158.000 2760.000 3162.000 ;
        RECT 2765.000 3158.000 2769.000 3162.000 ;
        RECT 2756.000 3150.000 2760.000 3154.000 ;
        RECT 2765.000 3150.000 2769.000 3154.000 ;
      LAYER met4 ;
        RECT 2755.000 3405.500 2770.000 3434.500 ;
        RECT 2733.500 3402.000 2770.000 3405.500 ;
        RECT 2755.000 3148.500 2770.000 3402.000 ;
    END
  END vccd1
  PIN vssa1
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 183.797394 ;
    PORT
      LAYER pwell ;
        RECT 2681.070 3438.225 2696.950 3438.655 ;
        RECT 2681.070 3431.795 2681.500 3438.225 ;
        RECT 2696.520 3431.795 2696.950 3438.225 ;
        RECT 2681.070 3431.365 2696.950 3431.795 ;
        RECT 2766.370 3438.225 2782.250 3438.655 ;
        RECT 2766.370 3431.795 2766.800 3438.225 ;
        RECT 2781.820 3431.795 2782.250 3438.225 ;
        RECT 2766.370 3431.365 2782.250 3431.795 ;
        RECT 2681.070 3430.875 2696.950 3431.305 ;
        RECT 2681.070 3424.445 2681.500 3430.875 ;
        RECT 2696.520 3424.445 2696.950 3430.875 ;
        RECT 2681.070 3424.015 2696.950 3424.445 ;
        RECT 2766.370 3430.875 2782.250 3431.305 ;
        RECT 2766.370 3424.445 2766.800 3430.875 ;
        RECT 2781.820 3424.445 2782.250 3430.875 ;
        RECT 2709.535 3421.680 2753.075 3424.040 ;
        RECT 2766.370 3424.015 2782.250 3424.445 ;
        RECT 2709.535 3419.180 2753.075 3421.540 ;
        RECT 2712.335 3416.180 2749.785 3419.040 ;
        RECT 2712.335 3413.080 2749.785 3415.940 ;
        RECT 2709.535 3410.080 2753.075 3412.940 ;
        RECT 2709.535 3407.080 2753.075 3409.940 ;
        RECT 2726.110 3395.310 2736.380 3398.170 ;
        RECT 2727.210 3392.420 2735.300 3395.310 ;
        RECT 2712.535 3389.560 2749.985 3392.420 ;
        RECT 2714.930 3382.460 2715.790 3383.560 ;
        RECT 2746.780 3382.460 2747.640 3383.560 ;
        RECT 2714.930 3367.460 2715.790 3368.560 ;
        RECT 2746.780 3367.460 2747.640 3368.560 ;
        RECT 2714.930 3352.460 2715.790 3353.560 ;
        RECT 2746.780 3352.460 2747.640 3353.560 ;
        RECT 2714.930 3337.460 2715.790 3338.560 ;
        RECT 2746.780 3337.460 2747.640 3338.560 ;
        RECT 2714.930 3322.460 2715.790 3323.560 ;
        RECT 2746.780 3322.460 2747.640 3323.560 ;
      LAYER li1 ;
        RECT 2681.200 3438.355 2696.820 3438.525 ;
        RECT 2681.200 3431.665 2681.370 3438.355 ;
        RECT 2687.135 3431.665 2687.585 3431.730 ;
        RECT 2696.650 3431.665 2696.820 3438.355 ;
        RECT 2681.200 3431.495 2696.820 3431.665 ;
        RECT 2766.500 3438.355 2782.120 3438.525 ;
        RECT 2766.500 3431.665 2766.670 3438.355 ;
        RECT 2781.950 3431.665 2782.120 3438.355 ;
        RECT 2766.500 3431.495 2782.120 3431.665 ;
        RECT 2687.135 3431.175 2687.585 3431.495 ;
        RECT 2773.385 3431.175 2774.085 3431.495 ;
        RECT 2681.200 3431.005 2696.820 3431.175 ;
        RECT 2681.200 3424.315 2681.370 3431.005 ;
        RECT 2696.650 3424.315 2696.820 3431.005 ;
        RECT 2681.200 3424.145 2696.820 3424.315 ;
        RECT 2766.500 3431.005 2782.120 3431.175 ;
        RECT 2766.500 3424.315 2766.670 3431.005 ;
        RECT 2781.950 3424.315 2782.120 3431.005 ;
        RECT 2766.500 3424.145 2782.120 3424.315 ;
        RECT 2687.035 3423.630 2687.485 3424.145 ;
        RECT 2688.085 3423.630 2688.535 3424.145 ;
        RECT 2709.665 3423.740 2752.945 3423.910 ;
        RECT 2773.585 3423.780 2773.935 3424.145 ;
        RECT 2774.385 3423.780 2774.735 3424.145 ;
        RECT 2709.665 3421.980 2709.835 3423.740 ;
        RECT 2752.775 3421.980 2752.945 3423.740 ;
        RECT 2709.665 3421.810 2752.945 3421.980 ;
        RECT 2719.635 3421.410 2720.185 3421.810 ;
        RECT 2723.935 3421.410 2724.485 3421.810 ;
        RECT 2729.985 3421.410 2730.535 3421.810 ;
        RECT 2734.235 3421.410 2734.785 3421.810 ;
        RECT 2742.085 3421.410 2742.635 3421.810 ;
        RECT 2746.485 3421.410 2747.035 3421.810 ;
        RECT 2709.665 3421.240 2752.945 3421.410 ;
        RECT 2709.665 3419.480 2709.835 3421.240 ;
        RECT 2752.775 3419.480 2752.945 3421.240 ;
        RECT 2709.665 3419.310 2752.945 3419.480 ;
        RECT 2712.465 3418.740 2749.655 3418.910 ;
        RECT 2712.465 3416.480 2712.635 3418.740 ;
        RECT 2713.315 3416.880 2718.355 3417.050 ;
        RECT 2719.405 3416.880 2724.445 3417.050 ;
        RECT 2725.495 3416.880 2730.535 3417.050 ;
        RECT 2731.585 3416.880 2736.625 3417.050 ;
        RECT 2737.675 3416.880 2742.715 3417.050 ;
        RECT 2743.765 3416.880 2748.805 3417.050 ;
        RECT 2749.485 3416.480 2749.655 3418.740 ;
        RECT 2712.465 3416.310 2749.655 3416.480 ;
        RECT 2715.935 3415.810 2716.785 3416.310 ;
        RECT 2740.485 3415.810 2741.335 3416.310 ;
        RECT 2712.465 3415.640 2749.655 3415.810 ;
        RECT 2712.465 3413.380 2712.635 3415.640 ;
        RECT 2713.315 3413.780 2718.355 3413.950 ;
        RECT 2719.405 3413.780 2724.445 3413.950 ;
        RECT 2725.495 3413.780 2730.535 3413.950 ;
        RECT 2731.585 3413.780 2736.625 3413.950 ;
        RECT 2737.675 3413.780 2742.715 3413.950 ;
        RECT 2743.765 3413.780 2748.805 3413.950 ;
        RECT 2749.485 3413.380 2749.655 3415.640 ;
        RECT 2712.465 3413.210 2749.655 3413.380 ;
        RECT 2709.665 3412.640 2752.945 3412.810 ;
        RECT 2709.665 3410.380 2709.835 3412.640 ;
        RECT 2710.515 3412.070 2715.555 3412.240 ;
        RECT 2716.605 3412.070 2721.645 3412.240 ;
        RECT 2722.695 3412.070 2727.735 3412.240 ;
        RECT 2728.785 3412.070 2733.825 3412.240 ;
        RECT 2734.875 3412.070 2739.915 3412.240 ;
        RECT 2740.965 3412.070 2746.005 3412.240 ;
        RECT 2747.055 3412.070 2752.095 3412.240 ;
        RECT 2752.775 3410.380 2752.945 3412.640 ;
        RECT 2709.665 3410.210 2752.945 3410.380 ;
        RECT 2715.785 3409.810 2716.385 3410.210 ;
        RECT 2721.885 3409.810 2722.485 3410.210 ;
        RECT 2727.935 3409.810 2728.535 3410.210 ;
        RECT 2734.035 3409.810 2734.635 3410.210 ;
        RECT 2740.185 3409.810 2740.785 3410.210 ;
        RECT 2746.235 3409.810 2746.835 3410.210 ;
        RECT 2709.665 3409.640 2752.945 3409.810 ;
        RECT 2709.665 3407.380 2709.835 3409.640 ;
        RECT 2710.515 3409.070 2715.555 3409.240 ;
        RECT 2716.605 3409.070 2721.645 3409.240 ;
        RECT 2722.695 3409.070 2727.735 3409.240 ;
        RECT 2728.785 3409.070 2733.825 3409.240 ;
        RECT 2734.875 3409.070 2739.915 3409.240 ;
        RECT 2740.965 3409.070 2746.005 3409.240 ;
        RECT 2747.055 3409.070 2752.095 3409.240 ;
        RECT 2752.775 3407.380 2752.945 3409.640 ;
        RECT 2709.665 3407.210 2752.945 3407.380 ;
        RECT 2726.240 3397.870 2736.250 3398.040 ;
        RECT 2726.240 3395.610 2726.410 3397.870 ;
        RECT 2727.090 3396.010 2728.380 3396.180 ;
        RECT 2729.430 3396.010 2730.720 3396.180 ;
        RECT 2731.770 3396.010 2733.060 3396.180 ;
        RECT 2734.110 3396.010 2735.400 3396.180 ;
        RECT 2736.080 3395.610 2736.250 3397.870 ;
        RECT 2726.240 3395.440 2736.250 3395.610 ;
        RECT 2727.060 3394.915 2728.160 3395.440 ;
        RECT 2729.660 3394.915 2730.760 3395.440 ;
        RECT 2731.760 3394.915 2732.860 3395.440 ;
        RECT 2734.510 3394.915 2735.610 3395.440 ;
        RECT 2727.060 3394.860 2735.610 3394.915 ;
        RECT 2727.340 3394.745 2735.170 3394.860 ;
        RECT 2727.340 3392.985 2727.510 3394.745 ;
        RECT 2735.000 3392.985 2735.170 3394.745 ;
        RECT 2715.260 3392.290 2716.160 3392.810 ;
        RECT 2720.960 3392.290 2721.860 3392.810 ;
        RECT 2725.860 3392.290 2726.760 3392.860 ;
        RECT 2727.340 3392.815 2735.170 3392.985 ;
        RECT 2729.710 3392.290 2730.610 3392.815 ;
        RECT 2731.910 3392.290 2732.810 3392.815 ;
        RECT 2735.510 3392.290 2736.410 3392.810 ;
        RECT 2740.860 3392.290 2741.760 3392.860 ;
        RECT 2745.860 3392.290 2746.760 3392.860 ;
        RECT 2712.665 3392.120 2749.855 3392.290 ;
        RECT 2712.665 3389.860 2712.835 3392.120 ;
        RECT 2749.685 3389.860 2749.855 3392.120 ;
        RECT 2712.665 3389.690 2749.855 3389.860 ;
        RECT 2715.060 3382.630 2715.660 3383.390 ;
        RECT 2746.910 3382.630 2747.510 3383.390 ;
        RECT 2715.060 3367.630 2715.660 3368.390 ;
        RECT 2746.910 3367.630 2747.510 3368.390 ;
        RECT 2715.060 3352.630 2715.660 3353.390 ;
        RECT 2746.910 3352.630 2747.510 3353.390 ;
        RECT 2715.060 3337.630 2715.660 3338.390 ;
        RECT 2746.910 3337.630 2747.510 3338.390 ;
        RECT 2715.060 3322.630 2715.660 3323.390 ;
        RECT 2746.910 3322.630 2747.510 3323.390 ;
        RECT 2717.045 3314.710 2722.775 3316.870 ;
        RECT 2724.645 3314.710 2730.375 3316.870 ;
        RECT 2732.195 3314.740 2737.925 3316.900 ;
        RECT 2739.745 3314.740 2745.475 3316.900 ;
      LAYER mcon ;
        RECT 2687.175 3424.050 2687.345 3424.220 ;
        RECT 2687.175 3423.690 2687.345 3423.860 ;
        RECT 2688.225 3424.050 2688.395 3424.220 ;
        RECT 2773.675 3423.920 2773.845 3424.090 ;
        RECT 2688.225 3423.690 2688.395 3423.860 ;
        RECT 2774.475 3423.920 2774.645 3424.090 ;
        RECT 2719.645 3421.340 2720.175 3421.870 ;
        RECT 2723.945 3421.340 2724.475 3421.870 ;
        RECT 2729.995 3421.340 2730.525 3421.870 ;
        RECT 2734.245 3421.340 2734.775 3421.870 ;
        RECT 2742.095 3421.340 2742.625 3421.870 ;
        RECT 2746.495 3421.340 2747.025 3421.870 ;
        RECT 2713.410 3416.880 2713.580 3417.050 ;
        RECT 2713.770 3416.880 2713.940 3417.050 ;
        RECT 2714.130 3416.880 2714.300 3417.050 ;
        RECT 2714.490 3416.880 2714.660 3417.050 ;
        RECT 2714.850 3416.880 2715.020 3417.050 ;
        RECT 2715.210 3416.880 2715.380 3417.050 ;
        RECT 2715.570 3416.880 2715.740 3417.050 ;
        RECT 2715.930 3416.880 2716.100 3417.050 ;
        RECT 2716.290 3416.880 2716.460 3417.050 ;
        RECT 2716.650 3416.880 2716.820 3417.050 ;
        RECT 2717.010 3416.880 2717.180 3417.050 ;
        RECT 2717.370 3416.880 2717.540 3417.050 ;
        RECT 2717.730 3416.880 2717.900 3417.050 ;
        RECT 2718.090 3416.880 2718.260 3417.050 ;
        RECT 2719.500 3416.880 2719.670 3417.050 ;
        RECT 2719.860 3416.880 2720.030 3417.050 ;
        RECT 2720.220 3416.880 2720.390 3417.050 ;
        RECT 2720.580 3416.880 2720.750 3417.050 ;
        RECT 2720.940 3416.880 2721.110 3417.050 ;
        RECT 2721.300 3416.880 2721.470 3417.050 ;
        RECT 2721.660 3416.880 2721.830 3417.050 ;
        RECT 2722.020 3416.880 2722.190 3417.050 ;
        RECT 2722.380 3416.880 2722.550 3417.050 ;
        RECT 2722.740 3416.880 2722.910 3417.050 ;
        RECT 2723.100 3416.880 2723.270 3417.050 ;
        RECT 2723.460 3416.880 2723.630 3417.050 ;
        RECT 2723.820 3416.880 2723.990 3417.050 ;
        RECT 2724.180 3416.880 2724.350 3417.050 ;
        RECT 2725.590 3416.880 2725.760 3417.050 ;
        RECT 2725.950 3416.880 2726.120 3417.050 ;
        RECT 2726.310 3416.880 2726.480 3417.050 ;
        RECT 2726.670 3416.880 2726.840 3417.050 ;
        RECT 2727.030 3416.880 2727.200 3417.050 ;
        RECT 2727.390 3416.880 2727.560 3417.050 ;
        RECT 2727.750 3416.880 2727.920 3417.050 ;
        RECT 2728.110 3416.880 2728.280 3417.050 ;
        RECT 2728.470 3416.880 2728.640 3417.050 ;
        RECT 2728.830 3416.880 2729.000 3417.050 ;
        RECT 2729.190 3416.880 2729.360 3417.050 ;
        RECT 2729.550 3416.880 2729.720 3417.050 ;
        RECT 2729.910 3416.880 2730.080 3417.050 ;
        RECT 2730.270 3416.880 2730.440 3417.050 ;
        RECT 2731.680 3416.880 2731.850 3417.050 ;
        RECT 2732.040 3416.880 2732.210 3417.050 ;
        RECT 2732.400 3416.880 2732.570 3417.050 ;
        RECT 2732.760 3416.880 2732.930 3417.050 ;
        RECT 2733.120 3416.880 2733.290 3417.050 ;
        RECT 2733.480 3416.880 2733.650 3417.050 ;
        RECT 2733.840 3416.880 2734.010 3417.050 ;
        RECT 2734.200 3416.880 2734.370 3417.050 ;
        RECT 2734.560 3416.880 2734.730 3417.050 ;
        RECT 2734.920 3416.880 2735.090 3417.050 ;
        RECT 2735.280 3416.880 2735.450 3417.050 ;
        RECT 2735.640 3416.880 2735.810 3417.050 ;
        RECT 2736.000 3416.880 2736.170 3417.050 ;
        RECT 2736.360 3416.880 2736.530 3417.050 ;
        RECT 2737.770 3416.880 2737.940 3417.050 ;
        RECT 2738.130 3416.880 2738.300 3417.050 ;
        RECT 2738.490 3416.880 2738.660 3417.050 ;
        RECT 2738.850 3416.880 2739.020 3417.050 ;
        RECT 2739.210 3416.880 2739.380 3417.050 ;
        RECT 2739.570 3416.880 2739.740 3417.050 ;
        RECT 2739.930 3416.880 2740.100 3417.050 ;
        RECT 2740.290 3416.880 2740.460 3417.050 ;
        RECT 2740.650 3416.880 2740.820 3417.050 ;
        RECT 2741.010 3416.880 2741.180 3417.050 ;
        RECT 2741.370 3416.880 2741.540 3417.050 ;
        RECT 2741.730 3416.880 2741.900 3417.050 ;
        RECT 2742.090 3416.880 2742.260 3417.050 ;
        RECT 2742.450 3416.880 2742.620 3417.050 ;
        RECT 2743.860 3416.880 2744.030 3417.050 ;
        RECT 2744.220 3416.880 2744.390 3417.050 ;
        RECT 2744.580 3416.880 2744.750 3417.050 ;
        RECT 2744.940 3416.880 2745.110 3417.050 ;
        RECT 2745.300 3416.880 2745.470 3417.050 ;
        RECT 2745.660 3416.880 2745.830 3417.050 ;
        RECT 2746.020 3416.880 2746.190 3417.050 ;
        RECT 2746.380 3416.880 2746.550 3417.050 ;
        RECT 2746.740 3416.880 2746.910 3417.050 ;
        RECT 2747.100 3416.880 2747.270 3417.050 ;
        RECT 2747.460 3416.880 2747.630 3417.050 ;
        RECT 2747.820 3416.880 2747.990 3417.050 ;
        RECT 2748.180 3416.880 2748.350 3417.050 ;
        RECT 2748.540 3416.880 2748.710 3417.050 ;
        RECT 2716.095 3415.970 2716.265 3416.140 ;
        RECT 2716.455 3415.970 2716.625 3416.140 ;
        RECT 2740.645 3415.970 2740.815 3416.140 ;
        RECT 2741.005 3415.970 2741.175 3416.140 ;
        RECT 2713.410 3413.780 2713.580 3413.950 ;
        RECT 2713.770 3413.780 2713.940 3413.950 ;
        RECT 2714.130 3413.780 2714.300 3413.950 ;
        RECT 2714.490 3413.780 2714.660 3413.950 ;
        RECT 2714.850 3413.780 2715.020 3413.950 ;
        RECT 2715.210 3413.780 2715.380 3413.950 ;
        RECT 2715.570 3413.780 2715.740 3413.950 ;
        RECT 2715.930 3413.780 2716.100 3413.950 ;
        RECT 2716.290 3413.780 2716.460 3413.950 ;
        RECT 2716.650 3413.780 2716.820 3413.950 ;
        RECT 2717.010 3413.780 2717.180 3413.950 ;
        RECT 2717.370 3413.780 2717.540 3413.950 ;
        RECT 2717.730 3413.780 2717.900 3413.950 ;
        RECT 2718.090 3413.780 2718.260 3413.950 ;
        RECT 2719.500 3413.780 2719.670 3413.950 ;
        RECT 2719.860 3413.780 2720.030 3413.950 ;
        RECT 2720.220 3413.780 2720.390 3413.950 ;
        RECT 2720.580 3413.780 2720.750 3413.950 ;
        RECT 2720.940 3413.780 2721.110 3413.950 ;
        RECT 2721.300 3413.780 2721.470 3413.950 ;
        RECT 2721.660 3413.780 2721.830 3413.950 ;
        RECT 2722.020 3413.780 2722.190 3413.950 ;
        RECT 2722.380 3413.780 2722.550 3413.950 ;
        RECT 2722.740 3413.780 2722.910 3413.950 ;
        RECT 2723.100 3413.780 2723.270 3413.950 ;
        RECT 2723.460 3413.780 2723.630 3413.950 ;
        RECT 2723.820 3413.780 2723.990 3413.950 ;
        RECT 2724.180 3413.780 2724.350 3413.950 ;
        RECT 2725.590 3413.780 2725.760 3413.950 ;
        RECT 2725.950 3413.780 2726.120 3413.950 ;
        RECT 2726.310 3413.780 2726.480 3413.950 ;
        RECT 2726.670 3413.780 2726.840 3413.950 ;
        RECT 2727.030 3413.780 2727.200 3413.950 ;
        RECT 2727.390 3413.780 2727.560 3413.950 ;
        RECT 2727.750 3413.780 2727.920 3413.950 ;
        RECT 2728.110 3413.780 2728.280 3413.950 ;
        RECT 2728.470 3413.780 2728.640 3413.950 ;
        RECT 2728.830 3413.780 2729.000 3413.950 ;
        RECT 2729.190 3413.780 2729.360 3413.950 ;
        RECT 2729.550 3413.780 2729.720 3413.950 ;
        RECT 2729.910 3413.780 2730.080 3413.950 ;
        RECT 2730.270 3413.780 2730.440 3413.950 ;
        RECT 2731.680 3413.780 2731.850 3413.950 ;
        RECT 2732.040 3413.780 2732.210 3413.950 ;
        RECT 2732.400 3413.780 2732.570 3413.950 ;
        RECT 2732.760 3413.780 2732.930 3413.950 ;
        RECT 2733.120 3413.780 2733.290 3413.950 ;
        RECT 2733.480 3413.780 2733.650 3413.950 ;
        RECT 2733.840 3413.780 2734.010 3413.950 ;
        RECT 2734.200 3413.780 2734.370 3413.950 ;
        RECT 2734.560 3413.780 2734.730 3413.950 ;
        RECT 2734.920 3413.780 2735.090 3413.950 ;
        RECT 2735.280 3413.780 2735.450 3413.950 ;
        RECT 2735.640 3413.780 2735.810 3413.950 ;
        RECT 2736.000 3413.780 2736.170 3413.950 ;
        RECT 2736.360 3413.780 2736.530 3413.950 ;
        RECT 2737.770 3413.780 2737.940 3413.950 ;
        RECT 2738.130 3413.780 2738.300 3413.950 ;
        RECT 2738.490 3413.780 2738.660 3413.950 ;
        RECT 2738.850 3413.780 2739.020 3413.950 ;
        RECT 2739.210 3413.780 2739.380 3413.950 ;
        RECT 2739.570 3413.780 2739.740 3413.950 ;
        RECT 2739.930 3413.780 2740.100 3413.950 ;
        RECT 2740.290 3413.780 2740.460 3413.950 ;
        RECT 2740.650 3413.780 2740.820 3413.950 ;
        RECT 2741.010 3413.780 2741.180 3413.950 ;
        RECT 2741.370 3413.780 2741.540 3413.950 ;
        RECT 2741.730 3413.780 2741.900 3413.950 ;
        RECT 2742.090 3413.780 2742.260 3413.950 ;
        RECT 2742.450 3413.780 2742.620 3413.950 ;
        RECT 2743.860 3413.780 2744.030 3413.950 ;
        RECT 2744.220 3413.780 2744.390 3413.950 ;
        RECT 2744.580 3413.780 2744.750 3413.950 ;
        RECT 2744.940 3413.780 2745.110 3413.950 ;
        RECT 2745.300 3413.780 2745.470 3413.950 ;
        RECT 2745.660 3413.780 2745.830 3413.950 ;
        RECT 2746.020 3413.780 2746.190 3413.950 ;
        RECT 2746.380 3413.780 2746.550 3413.950 ;
        RECT 2746.740 3413.780 2746.910 3413.950 ;
        RECT 2747.100 3413.780 2747.270 3413.950 ;
        RECT 2747.460 3413.780 2747.630 3413.950 ;
        RECT 2747.820 3413.780 2747.990 3413.950 ;
        RECT 2748.180 3413.780 2748.350 3413.950 ;
        RECT 2748.540 3413.780 2748.710 3413.950 ;
        RECT 2710.610 3412.070 2710.780 3412.240 ;
        RECT 2710.970 3412.070 2711.140 3412.240 ;
        RECT 2711.330 3412.070 2711.500 3412.240 ;
        RECT 2711.690 3412.070 2711.860 3412.240 ;
        RECT 2712.050 3412.070 2712.220 3412.240 ;
        RECT 2712.410 3412.070 2712.580 3412.240 ;
        RECT 2712.770 3412.070 2712.940 3412.240 ;
        RECT 2713.130 3412.070 2713.300 3412.240 ;
        RECT 2713.490 3412.070 2713.660 3412.240 ;
        RECT 2713.850 3412.070 2714.020 3412.240 ;
        RECT 2714.210 3412.070 2714.380 3412.240 ;
        RECT 2714.570 3412.070 2714.740 3412.240 ;
        RECT 2714.930 3412.070 2715.100 3412.240 ;
        RECT 2715.290 3412.070 2715.460 3412.240 ;
        RECT 2716.700 3412.070 2716.870 3412.240 ;
        RECT 2717.060 3412.070 2717.230 3412.240 ;
        RECT 2717.420 3412.070 2717.590 3412.240 ;
        RECT 2717.780 3412.070 2717.950 3412.240 ;
        RECT 2718.140 3412.070 2718.310 3412.240 ;
        RECT 2718.500 3412.070 2718.670 3412.240 ;
        RECT 2718.860 3412.070 2719.030 3412.240 ;
        RECT 2719.220 3412.070 2719.390 3412.240 ;
        RECT 2719.580 3412.070 2719.750 3412.240 ;
        RECT 2719.940 3412.070 2720.110 3412.240 ;
        RECT 2720.300 3412.070 2720.470 3412.240 ;
        RECT 2720.660 3412.070 2720.830 3412.240 ;
        RECT 2721.020 3412.070 2721.190 3412.240 ;
        RECT 2721.380 3412.070 2721.550 3412.240 ;
        RECT 2722.790 3412.070 2722.960 3412.240 ;
        RECT 2723.150 3412.070 2723.320 3412.240 ;
        RECT 2723.510 3412.070 2723.680 3412.240 ;
        RECT 2723.870 3412.070 2724.040 3412.240 ;
        RECT 2724.230 3412.070 2724.400 3412.240 ;
        RECT 2724.590 3412.070 2724.760 3412.240 ;
        RECT 2724.950 3412.070 2725.120 3412.240 ;
        RECT 2725.310 3412.070 2725.480 3412.240 ;
        RECT 2725.670 3412.070 2725.840 3412.240 ;
        RECT 2726.030 3412.070 2726.200 3412.240 ;
        RECT 2726.390 3412.070 2726.560 3412.240 ;
        RECT 2726.750 3412.070 2726.920 3412.240 ;
        RECT 2727.110 3412.070 2727.280 3412.240 ;
        RECT 2727.470 3412.070 2727.640 3412.240 ;
        RECT 2728.880 3412.070 2729.050 3412.240 ;
        RECT 2729.240 3412.070 2729.410 3412.240 ;
        RECT 2729.600 3412.070 2729.770 3412.240 ;
        RECT 2729.960 3412.070 2730.130 3412.240 ;
        RECT 2730.320 3412.070 2730.490 3412.240 ;
        RECT 2730.680 3412.070 2730.850 3412.240 ;
        RECT 2731.040 3412.070 2731.210 3412.240 ;
        RECT 2731.400 3412.070 2731.570 3412.240 ;
        RECT 2731.760 3412.070 2731.930 3412.240 ;
        RECT 2732.120 3412.070 2732.290 3412.240 ;
        RECT 2732.480 3412.070 2732.650 3412.240 ;
        RECT 2732.840 3412.070 2733.010 3412.240 ;
        RECT 2733.200 3412.070 2733.370 3412.240 ;
        RECT 2733.560 3412.070 2733.730 3412.240 ;
        RECT 2734.970 3412.070 2735.140 3412.240 ;
        RECT 2735.330 3412.070 2735.500 3412.240 ;
        RECT 2735.690 3412.070 2735.860 3412.240 ;
        RECT 2736.050 3412.070 2736.220 3412.240 ;
        RECT 2736.410 3412.070 2736.580 3412.240 ;
        RECT 2736.770 3412.070 2736.940 3412.240 ;
        RECT 2737.130 3412.070 2737.300 3412.240 ;
        RECT 2737.490 3412.070 2737.660 3412.240 ;
        RECT 2737.850 3412.070 2738.020 3412.240 ;
        RECT 2738.210 3412.070 2738.380 3412.240 ;
        RECT 2738.570 3412.070 2738.740 3412.240 ;
        RECT 2738.930 3412.070 2739.100 3412.240 ;
        RECT 2739.290 3412.070 2739.460 3412.240 ;
        RECT 2739.650 3412.070 2739.820 3412.240 ;
        RECT 2741.060 3412.070 2741.230 3412.240 ;
        RECT 2741.420 3412.070 2741.590 3412.240 ;
        RECT 2741.780 3412.070 2741.950 3412.240 ;
        RECT 2742.140 3412.070 2742.310 3412.240 ;
        RECT 2742.500 3412.070 2742.670 3412.240 ;
        RECT 2742.860 3412.070 2743.030 3412.240 ;
        RECT 2743.220 3412.070 2743.390 3412.240 ;
        RECT 2743.580 3412.070 2743.750 3412.240 ;
        RECT 2743.940 3412.070 2744.110 3412.240 ;
        RECT 2744.300 3412.070 2744.470 3412.240 ;
        RECT 2744.660 3412.070 2744.830 3412.240 ;
        RECT 2745.020 3412.070 2745.190 3412.240 ;
        RECT 2745.380 3412.070 2745.550 3412.240 ;
        RECT 2745.740 3412.070 2745.910 3412.240 ;
        RECT 2747.150 3412.070 2747.320 3412.240 ;
        RECT 2747.510 3412.070 2747.680 3412.240 ;
        RECT 2747.870 3412.070 2748.040 3412.240 ;
        RECT 2748.230 3412.070 2748.400 3412.240 ;
        RECT 2748.590 3412.070 2748.760 3412.240 ;
        RECT 2748.950 3412.070 2749.120 3412.240 ;
        RECT 2749.310 3412.070 2749.480 3412.240 ;
        RECT 2749.670 3412.070 2749.840 3412.240 ;
        RECT 2750.030 3412.070 2750.200 3412.240 ;
        RECT 2750.390 3412.070 2750.560 3412.240 ;
        RECT 2750.750 3412.070 2750.920 3412.240 ;
        RECT 2751.110 3412.070 2751.280 3412.240 ;
        RECT 2751.470 3412.070 2751.640 3412.240 ;
        RECT 2751.830 3412.070 2752.000 3412.240 ;
        RECT 2715.820 3409.945 2715.990 3410.115 ;
        RECT 2716.180 3409.945 2716.350 3410.115 ;
        RECT 2721.920 3409.945 2722.090 3410.115 ;
        RECT 2722.280 3409.945 2722.450 3410.115 ;
        RECT 2727.970 3409.945 2728.140 3410.115 ;
        RECT 2728.330 3409.945 2728.500 3410.115 ;
        RECT 2734.070 3409.945 2734.240 3410.115 ;
        RECT 2734.430 3409.945 2734.600 3410.115 ;
        RECT 2740.220 3409.895 2740.390 3410.065 ;
        RECT 2740.580 3409.895 2740.750 3410.065 ;
        RECT 2746.270 3409.945 2746.440 3410.115 ;
        RECT 2746.630 3409.945 2746.800 3410.115 ;
        RECT 2710.610 3409.070 2710.780 3409.240 ;
        RECT 2710.970 3409.070 2711.140 3409.240 ;
        RECT 2711.330 3409.070 2711.500 3409.240 ;
        RECT 2711.690 3409.070 2711.860 3409.240 ;
        RECT 2712.050 3409.070 2712.220 3409.240 ;
        RECT 2712.410 3409.070 2712.580 3409.240 ;
        RECT 2712.770 3409.070 2712.940 3409.240 ;
        RECT 2713.130 3409.070 2713.300 3409.240 ;
        RECT 2713.490 3409.070 2713.660 3409.240 ;
        RECT 2713.850 3409.070 2714.020 3409.240 ;
        RECT 2714.210 3409.070 2714.380 3409.240 ;
        RECT 2714.570 3409.070 2714.740 3409.240 ;
        RECT 2714.930 3409.070 2715.100 3409.240 ;
        RECT 2715.290 3409.070 2715.460 3409.240 ;
        RECT 2716.700 3409.070 2716.870 3409.240 ;
        RECT 2717.060 3409.070 2717.230 3409.240 ;
        RECT 2717.420 3409.070 2717.590 3409.240 ;
        RECT 2717.780 3409.070 2717.950 3409.240 ;
        RECT 2718.140 3409.070 2718.310 3409.240 ;
        RECT 2718.500 3409.070 2718.670 3409.240 ;
        RECT 2718.860 3409.070 2719.030 3409.240 ;
        RECT 2719.220 3409.070 2719.390 3409.240 ;
        RECT 2719.580 3409.070 2719.750 3409.240 ;
        RECT 2719.940 3409.070 2720.110 3409.240 ;
        RECT 2720.300 3409.070 2720.470 3409.240 ;
        RECT 2720.660 3409.070 2720.830 3409.240 ;
        RECT 2721.020 3409.070 2721.190 3409.240 ;
        RECT 2721.380 3409.070 2721.550 3409.240 ;
        RECT 2722.790 3409.070 2722.960 3409.240 ;
        RECT 2723.150 3409.070 2723.320 3409.240 ;
        RECT 2723.510 3409.070 2723.680 3409.240 ;
        RECT 2723.870 3409.070 2724.040 3409.240 ;
        RECT 2724.230 3409.070 2724.400 3409.240 ;
        RECT 2724.590 3409.070 2724.760 3409.240 ;
        RECT 2724.950 3409.070 2725.120 3409.240 ;
        RECT 2725.310 3409.070 2725.480 3409.240 ;
        RECT 2725.670 3409.070 2725.840 3409.240 ;
        RECT 2726.030 3409.070 2726.200 3409.240 ;
        RECT 2726.390 3409.070 2726.560 3409.240 ;
        RECT 2726.750 3409.070 2726.920 3409.240 ;
        RECT 2727.110 3409.070 2727.280 3409.240 ;
        RECT 2727.470 3409.070 2727.640 3409.240 ;
        RECT 2728.880 3409.070 2729.050 3409.240 ;
        RECT 2729.240 3409.070 2729.410 3409.240 ;
        RECT 2729.600 3409.070 2729.770 3409.240 ;
        RECT 2729.960 3409.070 2730.130 3409.240 ;
        RECT 2730.320 3409.070 2730.490 3409.240 ;
        RECT 2730.680 3409.070 2730.850 3409.240 ;
        RECT 2731.040 3409.070 2731.210 3409.240 ;
        RECT 2731.400 3409.070 2731.570 3409.240 ;
        RECT 2731.760 3409.070 2731.930 3409.240 ;
        RECT 2732.120 3409.070 2732.290 3409.240 ;
        RECT 2732.480 3409.070 2732.650 3409.240 ;
        RECT 2732.840 3409.070 2733.010 3409.240 ;
        RECT 2733.200 3409.070 2733.370 3409.240 ;
        RECT 2733.560 3409.070 2733.730 3409.240 ;
        RECT 2734.970 3409.070 2735.140 3409.240 ;
        RECT 2735.330 3409.070 2735.500 3409.240 ;
        RECT 2735.690 3409.070 2735.860 3409.240 ;
        RECT 2736.050 3409.070 2736.220 3409.240 ;
        RECT 2736.410 3409.070 2736.580 3409.240 ;
        RECT 2736.770 3409.070 2736.940 3409.240 ;
        RECT 2737.130 3409.070 2737.300 3409.240 ;
        RECT 2737.490 3409.070 2737.660 3409.240 ;
        RECT 2737.850 3409.070 2738.020 3409.240 ;
        RECT 2738.210 3409.070 2738.380 3409.240 ;
        RECT 2738.570 3409.070 2738.740 3409.240 ;
        RECT 2738.930 3409.070 2739.100 3409.240 ;
        RECT 2739.290 3409.070 2739.460 3409.240 ;
        RECT 2739.650 3409.070 2739.820 3409.240 ;
        RECT 2741.060 3409.070 2741.230 3409.240 ;
        RECT 2741.420 3409.070 2741.590 3409.240 ;
        RECT 2741.780 3409.070 2741.950 3409.240 ;
        RECT 2742.140 3409.070 2742.310 3409.240 ;
        RECT 2742.500 3409.070 2742.670 3409.240 ;
        RECT 2742.860 3409.070 2743.030 3409.240 ;
        RECT 2743.220 3409.070 2743.390 3409.240 ;
        RECT 2743.580 3409.070 2743.750 3409.240 ;
        RECT 2743.940 3409.070 2744.110 3409.240 ;
        RECT 2744.300 3409.070 2744.470 3409.240 ;
        RECT 2744.660 3409.070 2744.830 3409.240 ;
        RECT 2745.020 3409.070 2745.190 3409.240 ;
        RECT 2745.380 3409.070 2745.550 3409.240 ;
        RECT 2745.740 3409.070 2745.910 3409.240 ;
        RECT 2747.150 3409.070 2747.320 3409.240 ;
        RECT 2747.510 3409.070 2747.680 3409.240 ;
        RECT 2747.870 3409.070 2748.040 3409.240 ;
        RECT 2748.230 3409.070 2748.400 3409.240 ;
        RECT 2748.590 3409.070 2748.760 3409.240 ;
        RECT 2748.950 3409.070 2749.120 3409.240 ;
        RECT 2749.310 3409.070 2749.480 3409.240 ;
        RECT 2749.670 3409.070 2749.840 3409.240 ;
        RECT 2750.030 3409.070 2750.200 3409.240 ;
        RECT 2750.390 3409.070 2750.560 3409.240 ;
        RECT 2750.750 3409.070 2750.920 3409.240 ;
        RECT 2751.110 3409.070 2751.280 3409.240 ;
        RECT 2751.470 3409.070 2751.640 3409.240 ;
        RECT 2751.830 3409.070 2752.000 3409.240 ;
        RECT 2727.290 3396.010 2727.460 3396.180 ;
        RECT 2727.650 3396.010 2727.820 3396.180 ;
        RECT 2728.010 3396.010 2728.180 3396.180 ;
        RECT 2729.630 3396.010 2729.800 3396.180 ;
        RECT 2729.990 3396.010 2730.160 3396.180 ;
        RECT 2730.350 3396.010 2730.520 3396.180 ;
        RECT 2731.970 3396.010 2732.140 3396.180 ;
        RECT 2732.330 3396.010 2732.500 3396.180 ;
        RECT 2732.690 3396.010 2732.860 3396.180 ;
        RECT 2734.310 3396.010 2734.480 3396.180 ;
        RECT 2734.670 3396.010 2734.840 3396.180 ;
        RECT 2735.030 3396.010 2735.200 3396.180 ;
        RECT 2727.165 3394.970 2728.055 3395.500 ;
        RECT 2729.765 3394.970 2730.655 3395.500 ;
        RECT 2731.865 3394.970 2732.755 3395.500 ;
        RECT 2734.615 3394.970 2735.505 3395.500 ;
        RECT 2715.265 3392.220 2716.155 3392.750 ;
        RECT 2720.965 3392.220 2721.855 3392.750 ;
        RECT 2725.865 3392.270 2726.755 3392.800 ;
        RECT 2729.715 3392.270 2730.605 3392.800 ;
        RECT 2731.915 3392.270 2732.805 3392.800 ;
        RECT 2735.515 3392.220 2736.405 3392.750 ;
        RECT 2740.865 3392.270 2741.755 3392.800 ;
        RECT 2745.865 3392.270 2746.755 3392.800 ;
        RECT 2715.095 3382.745 2715.625 3383.275 ;
        RECT 2746.945 3382.745 2747.475 3383.275 ;
        RECT 2715.095 3367.745 2715.625 3368.275 ;
        RECT 2746.945 3367.745 2747.475 3368.275 ;
        RECT 2715.095 3352.745 2715.625 3353.275 ;
        RECT 2746.945 3352.745 2747.475 3353.275 ;
        RECT 2715.095 3337.745 2715.625 3338.275 ;
        RECT 2746.945 3337.745 2747.475 3338.275 ;
        RECT 2715.095 3322.745 2715.625 3323.275 ;
        RECT 2746.945 3322.745 2747.475 3323.275 ;
        RECT 2717.125 3314.805 2722.695 3316.775 ;
        RECT 2724.725 3314.805 2730.295 3316.775 ;
        RECT 2732.275 3314.835 2737.845 3316.805 ;
        RECT 2739.825 3314.835 2745.395 3316.805 ;
      LAYER met1 ;
        RECT 2687.005 3424.280 2687.515 3424.340 ;
        RECT 2688.055 3424.280 2688.565 3424.340 ;
        RECT 2686.985 3423.630 2687.535 3424.280 ;
        RECT 2688.035 3423.630 2688.585 3424.280 ;
        RECT 2773.555 3424.230 2773.965 3424.290 ;
        RECT 2774.355 3424.230 2774.765 3424.290 ;
        RECT 2773.535 3423.780 2773.985 3424.230 ;
        RECT 2774.335 3423.780 2774.785 3424.230 ;
        RECT 2773.555 3423.720 2773.965 3423.780 ;
        RECT 2774.355 3423.720 2774.765 3423.780 ;
        RECT 2687.005 3423.570 2687.515 3423.630 ;
        RECT 2688.055 3423.570 2688.565 3423.630 ;
        RECT 2719.575 3421.300 2720.245 3421.910 ;
        RECT 2723.875 3421.300 2724.545 3421.910 ;
        RECT 2729.925 3421.300 2730.595 3421.910 ;
        RECT 2734.175 3421.300 2734.845 3421.910 ;
        RECT 2742.025 3421.300 2742.695 3421.910 ;
        RECT 2746.425 3421.300 2747.095 3421.910 ;
        RECT 2713.335 3416.930 2718.335 3417.080 ;
        RECT 2719.425 3416.930 2724.425 3417.080 ;
        RECT 2725.515 3416.930 2730.515 3417.080 ;
        RECT 2731.605 3416.930 2736.605 3417.080 ;
        RECT 2737.695 3416.930 2742.695 3417.080 ;
        RECT 2743.785 3416.930 2748.785 3417.080 ;
        RECT 2713.285 3416.730 2748.885 3416.930 ;
        RECT 2715.485 3416.530 2715.985 3416.730 ;
        RECT 2739.935 3416.530 2740.435 3416.730 ;
        RECT 2716.025 3415.800 2716.695 3416.310 ;
        RECT 2740.575 3415.800 2741.245 3416.310 ;
        RECT 2713.335 3413.830 2718.335 3413.980 ;
        RECT 2719.425 3413.830 2724.425 3413.980 ;
        RECT 2725.515 3413.830 2730.515 3413.980 ;
        RECT 2731.605 3413.830 2736.605 3413.980 ;
        RECT 2737.695 3413.830 2742.695 3413.980 ;
        RECT 2743.785 3413.830 2748.785 3413.980 ;
        RECT 2713.285 3413.630 2748.885 3413.830 ;
        RECT 2715.485 3413.430 2715.985 3413.630 ;
        RECT 2739.935 3413.430 2740.435 3413.630 ;
        RECT 2724.885 3412.430 2725.435 3412.580 ;
        RECT 2749.285 3412.430 2749.835 3412.680 ;
        RECT 2710.485 3412.230 2752.085 3412.430 ;
        RECT 2710.535 3412.040 2715.535 3412.230 ;
        RECT 2716.625 3412.040 2721.625 3412.230 ;
        RECT 2722.715 3412.040 2727.715 3412.230 ;
        RECT 2728.805 3412.040 2733.805 3412.230 ;
        RECT 2734.895 3412.040 2739.895 3412.230 ;
        RECT 2740.985 3412.040 2745.985 3412.230 ;
        RECT 2747.075 3412.040 2752.075 3412.230 ;
        RECT 2715.685 3409.430 2716.485 3410.330 ;
        RECT 2721.785 3409.430 2722.585 3410.330 ;
        RECT 2724.885 3409.430 2725.435 3409.580 ;
        RECT 2727.835 3409.430 2728.635 3410.330 ;
        RECT 2733.975 3410.280 2734.695 3410.310 ;
        RECT 2746.175 3410.280 2746.895 3410.310 ;
        RECT 2733.935 3409.430 2734.735 3410.280 ;
        RECT 2740.125 3410.230 2740.845 3410.260 ;
        RECT 2740.085 3409.430 2740.885 3410.230 ;
        RECT 2746.135 3409.430 2746.935 3410.280 ;
        RECT 2749.285 3409.430 2749.835 3409.680 ;
        RECT 2710.485 3409.230 2752.085 3409.430 ;
        RECT 2710.535 3409.040 2715.535 3409.230 ;
        RECT 2716.625 3409.040 2721.625 3409.230 ;
        RECT 2722.715 3409.040 2727.715 3409.230 ;
        RECT 2728.805 3409.040 2733.805 3409.230 ;
        RECT 2734.895 3409.040 2739.895 3409.230 ;
        RECT 2740.985 3409.040 2745.985 3409.230 ;
        RECT 2747.075 3409.040 2752.075 3409.230 ;
        RECT 2727.110 3396.110 2728.360 3396.210 ;
        RECT 2729.450 3396.110 2730.700 3396.210 ;
        RECT 2731.790 3396.110 2733.040 3396.210 ;
        RECT 2734.130 3396.110 2735.380 3396.210 ;
        RECT 2727.060 3395.910 2735.410 3396.110 ;
        RECT 2727.060 3395.640 2735.610 3395.910 ;
        RECT 2727.000 3395.560 2735.670 3395.640 ;
        RECT 2727.000 3394.830 2728.220 3395.560 ;
        RECT 2729.600 3394.830 2730.820 3395.560 ;
        RECT 2731.700 3394.830 2732.920 3395.560 ;
        RECT 2734.450 3394.830 2735.670 3395.560 ;
        RECT 2715.200 3392.130 2716.220 3392.840 ;
        RECT 2720.900 3392.130 2721.920 3392.840 ;
        RECT 2725.800 3392.180 2726.820 3392.890 ;
        RECT 2729.650 3392.180 2730.670 3392.890 ;
        RECT 2731.850 3392.180 2732.870 3392.890 ;
        RECT 2735.450 3392.130 2736.470 3392.840 ;
        RECT 2740.800 3392.180 2741.820 3392.890 ;
        RECT 2745.800 3392.180 2746.820 3392.890 ;
        RECT 2715.000 3382.680 2715.720 3383.340 ;
        RECT 2746.850 3382.680 2747.570 3383.340 ;
        RECT 2715.000 3367.680 2715.720 3368.340 ;
        RECT 2746.850 3367.680 2747.570 3368.340 ;
        RECT 2715.000 3352.680 2715.720 3353.340 ;
        RECT 2746.850 3352.680 2747.570 3353.340 ;
        RECT 2715.000 3337.680 2715.720 3338.340 ;
        RECT 2746.850 3337.680 2747.570 3338.340 ;
        RECT 2715.000 3322.680 2715.720 3323.340 ;
        RECT 2746.850 3322.680 2747.570 3323.340 ;
        RECT 2716.260 3314.510 2746.260 3317.010 ;
      LAYER via ;
        RECT 2687.130 3423.985 2687.390 3424.245 ;
        RECT 2687.130 3423.665 2687.390 3423.925 ;
        RECT 2688.180 3423.985 2688.440 3424.245 ;
        RECT 2688.180 3423.665 2688.440 3423.925 ;
        RECT 2773.630 3423.875 2773.890 3424.135 ;
        RECT 2774.430 3423.875 2774.690 3424.135 ;
        RECT 2719.780 3421.475 2720.040 3421.735 ;
        RECT 2724.080 3421.475 2724.340 3421.735 ;
        RECT 2730.130 3421.475 2730.390 3421.735 ;
        RECT 2734.380 3421.475 2734.640 3421.735 ;
        RECT 2742.230 3421.475 2742.490 3421.735 ;
        RECT 2746.630 3421.475 2746.890 3421.735 ;
        RECT 2715.605 3416.600 2715.865 3416.860 ;
        RECT 2740.055 3416.600 2740.315 3416.860 ;
        RECT 2716.230 3415.925 2716.490 3416.185 ;
        RECT 2740.780 3415.925 2741.040 3416.185 ;
        RECT 2715.605 3413.500 2715.865 3413.760 ;
        RECT 2740.055 3413.500 2740.315 3413.760 ;
        RECT 2725.030 3412.250 2725.290 3412.510 ;
        RECT 2749.430 3412.350 2749.690 3412.610 ;
        RECT 2715.795 3409.900 2716.055 3410.160 ;
        RECT 2716.115 3409.900 2716.375 3410.160 ;
        RECT 2721.895 3409.900 2722.155 3410.160 ;
        RECT 2722.215 3409.900 2722.475 3410.160 ;
        RECT 2727.945 3409.900 2728.205 3410.160 ;
        RECT 2728.265 3409.900 2728.525 3410.160 ;
        RECT 2725.030 3409.250 2725.290 3409.510 ;
        RECT 2734.045 3409.900 2734.305 3410.160 ;
        RECT 2734.365 3409.900 2734.625 3410.160 ;
        RECT 2740.195 3409.850 2740.455 3410.110 ;
        RECT 2740.515 3409.850 2740.775 3410.110 ;
        RECT 2746.245 3409.900 2746.505 3410.160 ;
        RECT 2746.565 3409.900 2746.825 3410.160 ;
        RECT 2749.430 3409.350 2749.690 3409.610 ;
        RECT 2727.160 3394.945 2728.060 3395.525 ;
        RECT 2729.760 3394.945 2730.660 3395.525 ;
        RECT 2731.860 3394.945 2732.760 3395.525 ;
        RECT 2734.610 3394.945 2735.510 3395.525 ;
        RECT 2715.260 3392.195 2716.160 3392.775 ;
        RECT 2720.960 3392.195 2721.860 3392.775 ;
        RECT 2725.860 3392.245 2726.760 3392.825 ;
        RECT 2729.710 3392.245 2730.610 3392.825 ;
        RECT 2731.910 3392.245 2732.810 3392.825 ;
        RECT 2735.510 3392.195 2736.410 3392.775 ;
        RECT 2740.860 3392.245 2741.760 3392.825 ;
        RECT 2745.860 3392.245 2746.760 3392.825 ;
        RECT 2715.070 3382.720 2715.650 3383.300 ;
        RECT 2746.920 3382.720 2747.500 3383.300 ;
        RECT 2715.070 3367.720 2715.650 3368.300 ;
        RECT 2746.920 3367.720 2747.500 3368.300 ;
        RECT 2715.070 3352.720 2715.650 3353.300 ;
        RECT 2746.920 3352.720 2747.500 3353.300 ;
        RECT 2715.070 3337.720 2715.650 3338.300 ;
        RECT 2746.920 3337.720 2747.500 3338.300 ;
        RECT 2715.070 3322.720 2715.650 3323.300 ;
        RECT 2746.920 3322.720 2747.500 3323.300 ;
        RECT 2717.035 3314.705 2722.735 3316.565 ;
        RECT 2724.585 3314.705 2730.285 3316.565 ;
        RECT 2732.185 3314.705 2737.885 3316.565 ;
        RECT 2739.785 3314.755 2745.485 3316.615 ;
      LAYER met2 ;
        RECT 2687.035 3423.580 2687.485 3424.330 ;
        RECT 2688.085 3423.580 2688.535 3424.330 ;
        RECT 2773.585 3423.730 2773.935 3424.280 ;
        RECT 2774.385 3423.730 2774.735 3424.280 ;
        RECT 2719.635 3421.280 2720.185 3421.930 ;
        RECT 2723.935 3421.280 2724.485 3421.930 ;
        RECT 2729.985 3421.280 2730.535 3421.930 ;
        RECT 2734.235 3421.280 2734.785 3421.930 ;
        RECT 2742.085 3421.280 2742.635 3421.930 ;
        RECT 2746.485 3421.280 2747.035 3421.930 ;
        RECT 2715.535 3416.480 2715.935 3417.080 ;
        RECT 2739.985 3416.480 2740.385 3417.080 ;
        RECT 2715.535 3415.630 2716.835 3416.480 ;
        RECT 2739.985 3415.630 2741.335 3416.480 ;
        RECT 2715.535 3413.380 2715.935 3415.630 ;
        RECT 2739.985 3413.380 2740.385 3415.630 ;
        RECT 2715.785 3409.730 2716.385 3410.330 ;
        RECT 2721.885 3409.730 2722.485 3410.330 ;
        RECT 2724.935 3409.130 2725.385 3412.730 ;
        RECT 2727.935 3409.730 2728.535 3410.330 ;
        RECT 2734.035 3409.730 2734.635 3410.330 ;
        RECT 2740.185 3409.680 2740.785 3410.280 ;
        RECT 2746.235 3409.730 2746.835 3410.330 ;
        RECT 2749.335 3409.230 2749.785 3412.830 ;
        RECT 2727.060 3394.810 2728.160 3395.660 ;
        RECT 2729.660 3394.810 2730.760 3395.660 ;
        RECT 2731.760 3394.810 2732.860 3395.660 ;
        RECT 2734.510 3394.810 2735.610 3395.660 ;
        RECT 2715.260 3392.110 2716.160 3392.860 ;
        RECT 2720.960 3392.110 2721.860 3392.860 ;
        RECT 2725.860 3392.160 2726.760 3392.910 ;
        RECT 2729.710 3392.160 2730.610 3392.910 ;
        RECT 2731.910 3392.160 2732.810 3392.910 ;
        RECT 2735.510 3392.110 2736.410 3392.860 ;
        RECT 2740.860 3392.160 2741.760 3392.910 ;
        RECT 2745.860 3392.160 2746.760 3392.910 ;
        RECT 2715.060 3382.660 2715.660 3383.360 ;
        RECT 2746.910 3382.660 2747.510 3383.360 ;
        RECT 2715.060 3367.660 2715.660 3368.360 ;
        RECT 2746.910 3367.660 2747.510 3368.360 ;
        RECT 2715.060 3352.660 2715.660 3353.360 ;
        RECT 2746.910 3352.660 2747.510 3353.360 ;
        RECT 2715.060 3337.660 2715.660 3338.360 ;
        RECT 2746.910 3337.660 2747.510 3338.360 ;
        RECT 2715.060 3322.660 2715.660 3323.360 ;
        RECT 2746.910 3322.660 2747.510 3323.360 ;
        RECT 2716.960 3314.560 2722.810 3316.710 ;
        RECT 2724.510 3314.560 2730.360 3316.710 ;
        RECT 2732.110 3314.560 2737.960 3316.710 ;
        RECT 2739.710 3314.610 2745.560 3316.760 ;
      LAYER via2 ;
        RECT 2687.120 3423.815 2687.400 3424.095 ;
        RECT 2688.170 3423.815 2688.450 3424.095 ;
        RECT 2773.620 3423.865 2773.900 3424.145 ;
        RECT 2774.420 3423.865 2774.700 3424.145 ;
        RECT 2719.770 3421.465 2720.050 3421.745 ;
        RECT 2724.070 3421.465 2724.350 3421.745 ;
        RECT 2730.120 3421.465 2730.400 3421.745 ;
        RECT 2734.370 3421.465 2734.650 3421.745 ;
        RECT 2742.220 3421.465 2742.500 3421.745 ;
        RECT 2746.620 3421.465 2746.900 3421.745 ;
        RECT 2716.220 3415.915 2716.500 3416.195 ;
        RECT 2740.770 3415.915 2741.050 3416.195 ;
        RECT 2715.945 3409.890 2716.225 3410.170 ;
        RECT 2722.045 3409.890 2722.325 3410.170 ;
        RECT 2728.095 3409.890 2728.375 3410.170 ;
        RECT 2734.195 3409.890 2734.475 3410.170 ;
        RECT 2746.395 3409.890 2746.675 3410.170 ;
        RECT 2727.070 3394.895 2728.150 3395.575 ;
        RECT 2729.670 3394.895 2730.750 3395.575 ;
        RECT 2731.770 3394.895 2732.850 3395.575 ;
        RECT 2734.520 3394.895 2735.600 3395.575 ;
        RECT 2715.370 3392.345 2715.650 3392.625 ;
        RECT 2715.770 3392.345 2716.050 3392.625 ;
        RECT 2721.070 3392.345 2721.350 3392.625 ;
        RECT 2721.470 3392.345 2721.750 3392.625 ;
        RECT 2725.970 3392.395 2726.250 3392.675 ;
        RECT 2726.370 3392.395 2726.650 3392.675 ;
        RECT 2729.820 3392.395 2730.100 3392.675 ;
        RECT 2730.220 3392.395 2730.500 3392.675 ;
        RECT 2732.020 3392.395 2732.300 3392.675 ;
        RECT 2732.420 3392.395 2732.700 3392.675 ;
        RECT 2735.620 3392.345 2735.900 3392.625 ;
        RECT 2736.020 3392.345 2736.300 3392.625 ;
        RECT 2740.970 3392.395 2741.250 3392.675 ;
        RECT 2741.370 3392.395 2741.650 3392.675 ;
        RECT 2745.970 3392.395 2746.250 3392.675 ;
        RECT 2746.370 3392.395 2746.650 3392.675 ;
        RECT 2715.220 3382.870 2715.500 3383.150 ;
        RECT 2747.070 3382.870 2747.350 3383.150 ;
        RECT 2715.220 3367.870 2715.500 3368.150 ;
        RECT 2747.070 3367.870 2747.350 3368.150 ;
        RECT 2715.220 3352.870 2715.500 3353.150 ;
        RECT 2747.070 3352.870 2747.350 3353.150 ;
        RECT 2715.220 3337.870 2715.500 3338.150 ;
        RECT 2747.070 3337.870 2747.350 3338.150 ;
        RECT 2715.220 3322.870 2715.500 3323.150 ;
        RECT 2747.070 3322.870 2747.350 3323.150 ;
        RECT 2717.145 3314.695 2722.625 3316.575 ;
        RECT 2724.695 3314.695 2730.175 3316.575 ;
        RECT 2732.295 3314.695 2737.775 3316.575 ;
        RECT 2739.895 3314.745 2745.375 3316.625 ;
      LAYER met3 ;
        RECT 2552.970 3514.500 2576.970 3524.000 ;
        RECT 2602.970 3514.500 2626.970 3524.000 ;
        RECT 2552.500 3496.300 2629.000 3514.500 ;
        RECT 2686.935 3422.630 2688.685 3424.330 ;
        RECT 2684.435 3422.580 2707.785 3422.630 ;
        RECT 2773.535 3422.580 2774.835 3424.280 ;
        RECT 2684.435 3422.500 2780.485 3422.580 ;
        RECT 2578.500 3420.780 2780.485 3422.500 ;
        RECT 2578.500 3417.280 2708.500 3420.780 ;
        RECT 2755.235 3420.730 2780.485 3420.780 ;
        RECT 2755.585 3417.280 2756.685 3420.730 ;
        RECT 2578.500 3414.980 2756.685 3417.280 ;
        RECT 2578.500 3411.380 2708.500 3414.980 ;
        RECT 2755.585 3411.380 2756.685 3414.980 ;
        RECT 2578.500 3410.070 2756.685 3411.380 ;
        RECT 2578.500 3409.080 2758.750 3410.070 ;
        RECT 2578.500 3407.500 2708.500 3409.080 ;
        RECT 2578.500 3395.810 2718.000 3396.500 ;
        RECT 2754.070 3396.200 2758.750 3409.080 ;
        RECT 2754.070 3396.000 2758.800 3396.200 ;
        RECT 2747.500 3395.810 2758.800 3396.000 ;
        RECT 2578.500 3392.600 2758.800 3395.810 ;
        RECT 2578.500 3392.500 2755.500 3392.600 ;
        RECT 2578.500 3392.010 2747.810 3392.500 ;
        RECT 2578.500 3380.000 2718.000 3392.010 ;
        RECT 2714.710 3316.810 2716.310 3380.000 ;
        RECT 2746.210 3316.810 2747.810 3392.010 ;
        RECT 2714.710 3314.410 2747.810 3316.810 ;
      LAYER via3 ;
        RECT 2580.000 3507.000 2583.000 3510.000 ;
        RECT 2585.000 3507.000 2588.000 3510.000 ;
        RECT 2590.000 3507.000 2593.000 3510.000 ;
        RECT 2595.000 3507.000 2598.000 3510.000 ;
        RECT 2600.000 3507.000 2603.000 3510.000 ;
        RECT 2580.000 3503.000 2583.000 3506.000 ;
        RECT 2585.000 3503.000 2588.000 3506.000 ;
        RECT 2590.000 3503.000 2593.000 3506.000 ;
        RECT 2595.000 3503.000 2598.000 3506.000 ;
        RECT 2600.000 3503.000 2603.000 3506.000 ;
        RECT 2580.000 3499.000 2583.000 3502.000 ;
        RECT 2585.000 3499.000 2588.000 3502.000 ;
        RECT 2590.000 3499.000 2593.000 3502.000 ;
        RECT 2595.000 3499.000 2598.000 3502.000 ;
        RECT 2600.000 3499.000 2603.000 3502.000 ;
        RECT 2580.000 3419.000 2583.000 3422.000 ;
        RECT 2585.000 3419.000 2588.000 3422.000 ;
        RECT 2590.000 3419.000 2593.000 3422.000 ;
        RECT 2595.000 3419.000 2598.000 3422.000 ;
        RECT 2600.000 3419.000 2603.000 3422.000 ;
        RECT 2580.000 3414.000 2583.000 3417.000 ;
        RECT 2585.000 3414.000 2588.000 3417.000 ;
        RECT 2590.000 3414.000 2593.000 3417.000 ;
        RECT 2595.000 3414.000 2598.000 3417.000 ;
        RECT 2600.000 3414.000 2603.000 3417.000 ;
        RECT 2580.000 3409.000 2583.000 3412.000 ;
        RECT 2585.000 3409.000 2588.000 3412.000 ;
        RECT 2590.000 3409.000 2593.000 3412.000 ;
        RECT 2595.000 3409.000 2598.000 3412.000 ;
        RECT 2600.000 3409.000 2603.000 3412.000 ;
        RECT 2740.325 3409.820 2740.645 3410.140 ;
        RECT 2580.000 3391.000 2583.000 3394.000 ;
        RECT 2585.000 3391.000 2588.000 3394.000 ;
        RECT 2590.000 3391.000 2593.000 3394.000 ;
        RECT 2595.000 3391.000 2598.000 3394.000 ;
        RECT 2600.000 3391.000 2603.000 3394.000 ;
        RECT 2580.000 3386.000 2583.000 3389.000 ;
        RECT 2585.000 3386.000 2588.000 3389.000 ;
        RECT 2590.000 3386.000 2593.000 3389.000 ;
        RECT 2595.000 3386.000 2598.000 3389.000 ;
        RECT 2600.000 3386.000 2603.000 3389.000 ;
        RECT 2580.000 3381.000 2583.000 3384.000 ;
        RECT 2585.000 3381.000 2588.000 3384.000 ;
        RECT 2590.000 3381.000 2593.000 3384.000 ;
        RECT 2595.000 3381.000 2598.000 3384.000 ;
        RECT 2600.000 3381.000 2603.000 3384.000 ;
      LAYER met4 ;
        RECT 2578.500 3507.000 2604.100 3511.000 ;
        RECT 2578.500 3380.000 2604.000 3507.000 ;
        RECT 2740.180 3409.725 2740.790 3410.235 ;
    END
  END vssa1
  OBS
      LAYER li1 ;
        RECT 2709.675 3451.210 2709.845 3451.710 ;
        RECT 2715.315 3451.210 2715.485 3451.710 ;
        RECT 2715.855 3451.210 2716.025 3451.710 ;
        RECT 2721.495 3451.210 2721.665 3451.710 ;
        RECT 2722.035 3451.210 2722.205 3451.710 ;
        RECT 2727.675 3451.210 2727.845 3451.710 ;
        RECT 2728.215 3451.210 2728.385 3451.710 ;
        RECT 2733.855 3451.210 2734.025 3451.710 ;
        RECT 2734.395 3451.210 2734.565 3451.710 ;
        RECT 2740.035 3451.210 2740.205 3451.710 ;
        RECT 2740.575 3451.210 2740.745 3451.710 ;
        RECT 2746.215 3451.210 2746.385 3451.710 ;
        RECT 2746.755 3451.210 2746.925 3451.710 ;
        RECT 2752.395 3451.210 2752.565 3451.710 ;
        RECT 2710.060 3450.980 2715.100 3451.150 ;
        RECT 2716.240 3450.980 2721.280 3451.150 ;
        RECT 2722.420 3450.980 2727.460 3451.150 ;
        RECT 2728.600 3450.980 2733.640 3451.150 ;
        RECT 2734.780 3450.980 2739.820 3451.150 ;
        RECT 2740.960 3450.980 2746.000 3451.150 ;
        RECT 2747.140 3450.980 2752.180 3451.150 ;
        RECT 2709.675 3448.510 2709.845 3449.010 ;
        RECT 2715.315 3448.510 2715.485 3449.010 ;
        RECT 2715.855 3448.510 2716.025 3449.010 ;
        RECT 2721.495 3448.510 2721.665 3449.010 ;
        RECT 2722.035 3448.510 2722.205 3449.010 ;
        RECT 2727.675 3448.510 2727.845 3449.010 ;
        RECT 2728.215 3448.510 2728.385 3449.010 ;
        RECT 2733.855 3448.510 2734.025 3449.010 ;
        RECT 2734.395 3448.510 2734.565 3449.010 ;
        RECT 2740.035 3448.510 2740.205 3449.010 ;
        RECT 2740.575 3448.510 2740.745 3449.010 ;
        RECT 2746.215 3448.510 2746.385 3449.010 ;
        RECT 2746.755 3448.510 2746.925 3449.010 ;
        RECT 2752.395 3448.510 2752.565 3449.010 ;
        RECT 2710.060 3448.280 2715.100 3448.450 ;
        RECT 2716.240 3448.280 2721.280 3448.450 ;
        RECT 2722.420 3448.280 2727.460 3448.450 ;
        RECT 2728.600 3448.280 2733.640 3448.450 ;
        RECT 2734.780 3448.280 2739.820 3448.450 ;
        RECT 2740.960 3448.280 2746.000 3448.450 ;
        RECT 2747.140 3448.280 2752.180 3448.450 ;
        RECT 2709.675 3445.810 2709.845 3446.310 ;
        RECT 2715.315 3445.810 2715.485 3446.310 ;
        RECT 2715.855 3445.810 2716.025 3446.310 ;
        RECT 2721.495 3445.810 2721.665 3446.310 ;
        RECT 2722.035 3445.810 2722.205 3446.310 ;
        RECT 2727.675 3445.810 2727.845 3446.310 ;
        RECT 2728.215 3445.810 2728.385 3446.310 ;
        RECT 2733.855 3445.810 2734.025 3446.310 ;
        RECT 2734.395 3445.810 2734.565 3446.310 ;
        RECT 2740.035 3445.810 2740.205 3446.310 ;
        RECT 2740.575 3445.810 2740.745 3446.310 ;
        RECT 2746.215 3445.810 2746.385 3446.310 ;
        RECT 2746.755 3445.810 2746.925 3446.310 ;
        RECT 2752.395 3445.810 2752.565 3446.310 ;
        RECT 2710.060 3445.580 2715.100 3445.750 ;
        RECT 2716.240 3445.580 2721.280 3445.750 ;
        RECT 2722.420 3445.580 2727.460 3445.750 ;
        RECT 2728.600 3445.580 2733.640 3445.750 ;
        RECT 2734.780 3445.580 2739.820 3445.750 ;
        RECT 2740.960 3445.580 2746.000 3445.750 ;
        RECT 2747.140 3445.580 2752.180 3445.750 ;
        RECT 2709.675 3443.110 2709.845 3443.610 ;
        RECT 2715.315 3443.110 2715.485 3443.610 ;
        RECT 2715.855 3443.110 2716.025 3443.610 ;
        RECT 2721.495 3443.110 2721.665 3443.610 ;
        RECT 2722.035 3443.110 2722.205 3443.610 ;
        RECT 2727.675 3443.110 2727.845 3443.610 ;
        RECT 2728.215 3443.110 2728.385 3443.610 ;
        RECT 2733.855 3443.110 2734.025 3443.610 ;
        RECT 2734.395 3443.110 2734.565 3443.610 ;
        RECT 2740.035 3443.110 2740.205 3443.610 ;
        RECT 2740.575 3443.110 2740.745 3443.610 ;
        RECT 2746.215 3443.110 2746.385 3443.610 ;
        RECT 2746.755 3443.110 2746.925 3443.610 ;
        RECT 2752.395 3443.110 2752.565 3443.610 ;
        RECT 2710.060 3442.880 2715.100 3443.050 ;
        RECT 2716.240 3442.880 2721.280 3443.050 ;
        RECT 2722.420 3442.880 2727.460 3443.050 ;
        RECT 2728.600 3442.880 2733.640 3443.050 ;
        RECT 2734.780 3442.880 2739.820 3443.050 ;
        RECT 2740.960 3442.880 2746.000 3443.050 ;
        RECT 2747.140 3442.880 2752.180 3443.050 ;
        RECT 2709.675 3440.210 2709.845 3440.710 ;
        RECT 2715.315 3440.210 2715.485 3440.710 ;
        RECT 2715.855 3440.210 2716.025 3440.710 ;
        RECT 2721.495 3440.210 2721.665 3440.710 ;
        RECT 2722.035 3440.210 2722.205 3440.710 ;
        RECT 2727.675 3440.210 2727.845 3440.710 ;
        RECT 2728.215 3440.210 2728.385 3440.710 ;
        RECT 2733.855 3440.210 2734.025 3440.710 ;
        RECT 2734.395 3440.210 2734.565 3440.710 ;
        RECT 2740.035 3440.210 2740.205 3440.710 ;
        RECT 2740.575 3440.210 2740.745 3440.710 ;
        RECT 2746.215 3440.210 2746.385 3440.710 ;
        RECT 2746.755 3440.210 2746.925 3440.710 ;
        RECT 2752.395 3440.210 2752.565 3440.710 ;
        RECT 2710.060 3439.980 2715.100 3440.150 ;
        RECT 2716.240 3439.980 2721.280 3440.150 ;
        RECT 2722.420 3439.980 2727.460 3440.150 ;
        RECT 2728.600 3439.980 2733.640 3440.150 ;
        RECT 2734.780 3439.980 2739.820 3440.150 ;
        RECT 2740.960 3439.980 2746.000 3440.150 ;
        RECT 2747.140 3439.980 2752.180 3440.150 ;
        RECT 2681.850 3432.145 2684.010 3437.875 ;
        RECT 2694.010 3432.145 2696.170 3437.875 ;
        RECT 2709.675 3437.310 2709.845 3437.810 ;
        RECT 2715.315 3437.310 2715.485 3437.810 ;
        RECT 2715.855 3437.310 2716.025 3437.810 ;
        RECT 2721.495 3437.310 2721.665 3437.810 ;
        RECT 2722.035 3437.310 2722.205 3437.810 ;
        RECT 2727.675 3437.310 2727.845 3437.810 ;
        RECT 2728.215 3437.310 2728.385 3437.810 ;
        RECT 2733.855 3437.310 2734.025 3437.810 ;
        RECT 2734.395 3437.310 2734.565 3437.810 ;
        RECT 2740.035 3437.310 2740.205 3437.810 ;
        RECT 2740.575 3437.310 2740.745 3437.810 ;
        RECT 2746.215 3437.310 2746.385 3437.810 ;
        RECT 2746.755 3437.310 2746.925 3437.810 ;
        RECT 2752.395 3437.310 2752.565 3437.810 ;
        RECT 2710.060 3437.080 2715.100 3437.250 ;
        RECT 2716.240 3437.080 2721.280 3437.250 ;
        RECT 2722.420 3437.080 2727.460 3437.250 ;
        RECT 2728.600 3437.080 2733.640 3437.250 ;
        RECT 2734.780 3437.080 2739.820 3437.250 ;
        RECT 2740.960 3437.080 2746.000 3437.250 ;
        RECT 2747.140 3437.080 2752.180 3437.250 ;
        RECT 2700.475 3434.610 2700.645 3435.110 ;
        RECT 2706.115 3434.610 2706.285 3435.110 ;
        RECT 2706.655 3434.610 2706.825 3435.110 ;
        RECT 2712.295 3434.610 2712.465 3435.110 ;
        RECT 2712.835 3434.610 2713.005 3435.110 ;
        RECT 2718.475 3434.610 2718.645 3435.110 ;
        RECT 2719.015 3434.610 2719.185 3435.110 ;
        RECT 2724.655 3434.610 2724.825 3435.110 ;
        RECT 2725.195 3434.610 2725.365 3435.110 ;
        RECT 2730.835 3434.610 2731.005 3435.110 ;
        RECT 2731.375 3434.610 2731.545 3435.110 ;
        RECT 2737.015 3434.610 2737.185 3435.110 ;
        RECT 2737.555 3434.610 2737.725 3435.110 ;
        RECT 2743.195 3434.610 2743.365 3435.110 ;
        RECT 2743.735 3434.610 2743.905 3435.110 ;
        RECT 2749.375 3434.610 2749.545 3435.110 ;
        RECT 2749.915 3434.610 2750.085 3435.110 ;
        RECT 2755.555 3434.610 2755.725 3435.110 ;
        RECT 2756.095 3434.610 2756.265 3435.110 ;
        RECT 2761.735 3434.610 2761.905 3435.110 ;
        RECT 2700.475 3431.910 2700.645 3432.410 ;
        RECT 2706.115 3431.910 2706.285 3432.410 ;
        RECT 2706.655 3431.910 2706.825 3432.410 ;
        RECT 2712.295 3431.910 2712.465 3432.410 ;
        RECT 2712.835 3431.910 2713.005 3432.410 ;
        RECT 2718.475 3431.910 2718.645 3432.410 ;
        RECT 2719.015 3431.910 2719.185 3432.410 ;
        RECT 2724.655 3431.910 2724.825 3432.410 ;
        RECT 2725.195 3431.910 2725.365 3432.410 ;
        RECT 2730.835 3431.910 2731.005 3432.410 ;
        RECT 2731.375 3431.910 2731.545 3432.410 ;
        RECT 2737.015 3431.910 2737.185 3432.410 ;
        RECT 2737.555 3431.910 2737.725 3432.410 ;
        RECT 2743.195 3431.910 2743.365 3432.410 ;
        RECT 2743.735 3431.910 2743.905 3432.410 ;
        RECT 2749.375 3431.910 2749.545 3432.410 ;
        RECT 2749.915 3431.910 2750.085 3432.410 ;
        RECT 2755.555 3431.910 2755.725 3432.410 ;
        RECT 2756.095 3431.910 2756.265 3432.410 ;
        RECT 2761.735 3431.910 2761.905 3432.410 ;
        RECT 2767.150 3432.145 2769.310 3437.875 ;
        RECT 2779.310 3432.145 2781.470 3437.875 ;
        RECT 2681.850 3424.795 2684.010 3430.525 ;
        RECT 2694.010 3424.795 2696.170 3430.525 ;
        RECT 2700.475 3429.210 2700.645 3429.710 ;
        RECT 2706.115 3429.210 2706.285 3429.710 ;
        RECT 2706.655 3429.210 2706.825 3429.710 ;
        RECT 2712.295 3429.210 2712.465 3429.710 ;
        RECT 2712.835 3429.210 2713.005 3429.710 ;
        RECT 2718.475 3429.210 2718.645 3429.710 ;
        RECT 2719.015 3429.210 2719.185 3429.710 ;
        RECT 2724.655 3429.210 2724.825 3429.710 ;
        RECT 2725.195 3429.210 2725.365 3429.710 ;
        RECT 2730.835 3429.210 2731.005 3429.710 ;
        RECT 2731.375 3429.210 2731.545 3429.710 ;
        RECT 2737.015 3429.210 2737.185 3429.710 ;
        RECT 2737.555 3429.210 2737.725 3429.710 ;
        RECT 2743.195 3429.210 2743.365 3429.710 ;
        RECT 2743.735 3429.210 2743.905 3429.710 ;
        RECT 2749.375 3429.210 2749.545 3429.710 ;
        RECT 2749.915 3429.210 2750.085 3429.710 ;
        RECT 2755.555 3429.210 2755.725 3429.710 ;
        RECT 2756.095 3429.210 2756.265 3429.710 ;
        RECT 2761.735 3429.210 2761.905 3429.710 ;
        RECT 2700.475 3426.510 2700.645 3427.010 ;
        RECT 2706.115 3426.510 2706.285 3427.010 ;
        RECT 2706.655 3426.510 2706.825 3427.010 ;
        RECT 2712.295 3426.510 2712.465 3427.010 ;
        RECT 2712.835 3426.510 2713.005 3427.010 ;
        RECT 2718.475 3426.510 2718.645 3427.010 ;
        RECT 2719.015 3426.510 2719.185 3427.010 ;
        RECT 2724.655 3426.510 2724.825 3427.010 ;
        RECT 2725.195 3426.510 2725.365 3427.010 ;
        RECT 2730.835 3426.510 2731.005 3427.010 ;
        RECT 2731.375 3426.510 2731.545 3427.010 ;
        RECT 2737.015 3426.510 2737.185 3427.010 ;
        RECT 2737.555 3426.510 2737.725 3427.010 ;
        RECT 2743.195 3426.510 2743.365 3427.010 ;
        RECT 2743.735 3426.510 2743.905 3427.010 ;
        RECT 2749.375 3426.510 2749.545 3427.010 ;
        RECT 2749.915 3426.510 2750.085 3427.010 ;
        RECT 2755.555 3426.510 2755.725 3427.010 ;
        RECT 2756.095 3426.510 2756.265 3427.010 ;
        RECT 2761.735 3426.510 2761.905 3427.010 ;
        RECT 2767.150 3424.795 2769.310 3430.525 ;
        RECT 2779.310 3424.795 2781.470 3430.525 ;
        RECT 2710.515 3423.170 2715.555 3423.340 ;
        RECT 2716.605 3423.170 2721.645 3423.340 ;
        RECT 2722.695 3423.170 2727.735 3423.340 ;
        RECT 2728.785 3423.170 2733.825 3423.340 ;
        RECT 2734.875 3423.170 2739.915 3423.340 ;
        RECT 2740.965 3423.170 2746.005 3423.340 ;
        RECT 2747.055 3423.170 2752.095 3423.340 ;
        RECT 2710.515 3422.380 2715.555 3422.550 ;
        RECT 2716.605 3422.380 2721.645 3422.550 ;
        RECT 2722.695 3422.380 2727.735 3422.550 ;
        RECT 2728.785 3422.380 2733.825 3422.550 ;
        RECT 2734.875 3422.380 2739.915 3422.550 ;
        RECT 2740.965 3422.380 2746.005 3422.550 ;
        RECT 2747.055 3422.380 2752.095 3422.550 ;
        RECT 2710.515 3420.670 2715.555 3420.840 ;
        RECT 2716.605 3420.670 2721.645 3420.840 ;
        RECT 2722.695 3420.670 2727.735 3420.840 ;
        RECT 2728.785 3420.670 2733.825 3420.840 ;
        RECT 2734.875 3420.670 2739.915 3420.840 ;
        RECT 2740.965 3420.670 2746.005 3420.840 ;
        RECT 2747.055 3420.670 2752.095 3420.840 ;
        RECT 2710.515 3419.880 2715.555 3420.050 ;
        RECT 2716.605 3419.880 2721.645 3420.050 ;
        RECT 2722.695 3419.880 2727.735 3420.050 ;
        RECT 2728.785 3419.880 2733.825 3420.050 ;
        RECT 2734.875 3419.880 2739.915 3420.050 ;
        RECT 2740.965 3419.880 2746.005 3420.050 ;
        RECT 2747.055 3419.880 2752.095 3420.050 ;
        RECT 2712.975 3417.110 2713.145 3418.110 ;
        RECT 2718.525 3417.110 2718.695 3418.110 ;
        RECT 2719.065 3417.110 2719.235 3418.110 ;
        RECT 2724.615 3417.110 2724.785 3418.110 ;
        RECT 2725.155 3417.110 2725.325 3418.110 ;
        RECT 2730.705 3417.110 2730.875 3418.110 ;
        RECT 2731.245 3417.110 2731.415 3418.110 ;
        RECT 2736.795 3417.110 2736.965 3418.110 ;
        RECT 2737.335 3417.110 2737.505 3418.110 ;
        RECT 2742.885 3417.110 2743.055 3418.110 ;
        RECT 2743.425 3417.110 2743.595 3418.110 ;
        RECT 2748.975 3417.110 2749.145 3418.110 ;
        RECT 2712.975 3414.010 2713.145 3415.010 ;
        RECT 2718.525 3414.010 2718.695 3415.010 ;
        RECT 2719.065 3414.010 2719.235 3415.010 ;
        RECT 2724.615 3414.010 2724.785 3415.010 ;
        RECT 2725.155 3414.010 2725.325 3415.010 ;
        RECT 2730.705 3414.010 2730.875 3415.010 ;
        RECT 2731.245 3414.010 2731.415 3415.010 ;
        RECT 2736.795 3414.010 2736.965 3415.010 ;
        RECT 2737.335 3414.010 2737.505 3415.010 ;
        RECT 2742.885 3414.010 2743.055 3415.010 ;
        RECT 2743.425 3414.010 2743.595 3415.010 ;
        RECT 2748.975 3414.010 2749.145 3415.010 ;
        RECT 2710.175 3411.010 2710.345 3412.010 ;
        RECT 2715.725 3411.010 2715.895 3412.010 ;
        RECT 2716.265 3411.010 2716.435 3412.010 ;
        RECT 2721.815 3411.010 2721.985 3412.010 ;
        RECT 2722.355 3411.010 2722.525 3412.010 ;
        RECT 2727.905 3411.010 2728.075 3412.010 ;
        RECT 2728.445 3411.010 2728.615 3412.010 ;
        RECT 2733.995 3411.010 2734.165 3412.010 ;
        RECT 2734.535 3411.010 2734.705 3412.010 ;
        RECT 2740.085 3411.010 2740.255 3412.010 ;
        RECT 2740.625 3411.010 2740.795 3412.010 ;
        RECT 2746.175 3411.010 2746.345 3412.010 ;
        RECT 2746.715 3411.010 2746.885 3412.010 ;
        RECT 2752.265 3411.010 2752.435 3412.010 ;
        RECT 2710.515 3410.780 2715.555 3410.950 ;
        RECT 2716.605 3410.780 2721.645 3410.950 ;
        RECT 2722.695 3410.780 2727.735 3410.950 ;
        RECT 2728.785 3410.780 2733.825 3410.950 ;
        RECT 2734.875 3410.780 2739.915 3410.950 ;
        RECT 2740.965 3410.780 2746.005 3410.950 ;
        RECT 2747.055 3410.780 2752.095 3410.950 ;
        RECT 2710.175 3408.010 2710.345 3409.010 ;
        RECT 2715.725 3408.010 2715.895 3409.010 ;
        RECT 2716.265 3408.010 2716.435 3409.010 ;
        RECT 2721.815 3408.010 2721.985 3409.010 ;
        RECT 2722.355 3408.010 2722.525 3409.010 ;
        RECT 2727.905 3408.010 2728.075 3409.010 ;
        RECT 2728.445 3408.010 2728.615 3409.010 ;
        RECT 2733.995 3408.010 2734.165 3409.010 ;
        RECT 2734.535 3408.010 2734.705 3409.010 ;
        RECT 2740.085 3408.010 2740.255 3409.010 ;
        RECT 2740.625 3408.010 2740.795 3409.010 ;
        RECT 2746.175 3408.010 2746.345 3409.010 ;
        RECT 2746.715 3408.010 2746.885 3409.010 ;
        RECT 2752.265 3408.010 2752.435 3409.010 ;
        RECT 2710.515 3407.780 2715.555 3407.950 ;
        RECT 2716.605 3407.780 2721.645 3407.950 ;
        RECT 2722.695 3407.780 2727.735 3407.950 ;
        RECT 2728.785 3407.780 2733.825 3407.950 ;
        RECT 2734.875 3407.780 2739.915 3407.950 ;
        RECT 2740.965 3407.780 2746.005 3407.950 ;
        RECT 2747.055 3407.780 2752.095 3407.950 ;
        RECT 2712.900 3403.140 2713.070 3404.140 ;
        RECT 2718.540 3403.140 2718.710 3404.140 ;
        RECT 2719.080 3403.140 2719.250 3404.140 ;
        RECT 2724.720 3403.140 2724.890 3404.140 ;
        RECT 2725.260 3403.140 2725.430 3404.140 ;
        RECT 2730.900 3403.140 2731.070 3404.140 ;
        RECT 2731.440 3403.140 2731.610 3404.140 ;
        RECT 2737.080 3403.140 2737.250 3404.140 ;
        RECT 2737.620 3403.140 2737.790 3404.140 ;
        RECT 2743.260 3403.140 2743.430 3404.140 ;
        RECT 2743.800 3403.140 2743.970 3404.140 ;
        RECT 2749.440 3403.140 2749.610 3404.140 ;
        RECT 2713.285 3402.910 2718.325 3403.080 ;
        RECT 2719.465 3402.910 2724.505 3403.080 ;
        RECT 2725.645 3402.910 2730.685 3403.080 ;
        RECT 2731.825 3402.910 2736.865 3403.080 ;
        RECT 2738.005 3402.910 2743.045 3403.080 ;
        RECT 2744.185 3402.910 2749.225 3403.080 ;
        RECT 2712.900 3400.190 2713.070 3401.190 ;
        RECT 2718.540 3400.190 2718.710 3401.190 ;
        RECT 2719.080 3400.190 2719.250 3401.190 ;
        RECT 2724.720 3400.190 2724.890 3401.190 ;
        RECT 2725.260 3400.190 2725.430 3401.190 ;
        RECT 2730.900 3400.190 2731.070 3401.190 ;
        RECT 2731.440 3400.190 2731.610 3401.190 ;
        RECT 2737.080 3400.190 2737.250 3401.190 ;
        RECT 2737.620 3400.190 2737.790 3401.190 ;
        RECT 2743.260 3400.190 2743.430 3401.190 ;
        RECT 2743.800 3400.190 2743.970 3401.190 ;
        RECT 2749.440 3400.190 2749.610 3401.190 ;
        RECT 2713.285 3399.960 2718.325 3400.130 ;
        RECT 2719.465 3399.960 2724.505 3400.130 ;
        RECT 2725.645 3399.960 2730.685 3400.130 ;
        RECT 2731.825 3399.960 2736.865 3400.130 ;
        RECT 2738.005 3399.960 2743.045 3400.130 ;
        RECT 2744.185 3399.960 2749.225 3400.130 ;
        RECT 2727.090 3397.300 2728.380 3397.470 ;
        RECT 2729.430 3397.300 2730.720 3397.470 ;
        RECT 2731.770 3397.300 2733.060 3397.470 ;
        RECT 2734.110 3397.300 2735.400 3397.470 ;
        RECT 2726.750 3396.240 2726.920 3397.240 ;
        RECT 2728.550 3396.240 2728.720 3397.240 ;
        RECT 2729.090 3396.240 2729.260 3397.240 ;
        RECT 2730.890 3396.240 2731.060 3397.240 ;
        RECT 2731.430 3396.240 2731.600 3397.240 ;
        RECT 2733.230 3396.240 2733.400 3397.240 ;
        RECT 2733.770 3396.240 2733.940 3397.240 ;
        RECT 2735.570 3396.240 2735.740 3397.240 ;
        RECT 2728.190 3394.175 2730.730 3394.345 ;
        RECT 2731.780 3394.175 2734.320 3394.345 ;
        RECT 2727.850 3393.615 2728.020 3394.115 ;
        RECT 2730.900 3393.615 2731.070 3394.115 ;
        RECT 2731.440 3393.615 2731.610 3394.115 ;
        RECT 2734.490 3393.615 2734.660 3394.115 ;
        RECT 2728.190 3393.385 2730.730 3393.555 ;
        RECT 2731.780 3393.385 2734.320 3393.555 ;
        RECT 2713.515 3391.550 2718.555 3391.720 ;
        RECT 2719.605 3391.550 2724.645 3391.720 ;
        RECT 2725.695 3391.550 2730.735 3391.720 ;
        RECT 2731.785 3391.550 2736.825 3391.720 ;
        RECT 2737.875 3391.550 2742.915 3391.720 ;
        RECT 2743.965 3391.550 2749.005 3391.720 ;
        RECT 2713.175 3390.490 2713.345 3391.490 ;
        RECT 2718.725 3390.490 2718.895 3391.490 ;
        RECT 2719.265 3390.490 2719.435 3391.490 ;
        RECT 2724.815 3390.490 2724.985 3391.490 ;
        RECT 2725.355 3390.490 2725.525 3391.490 ;
        RECT 2730.905 3390.490 2731.075 3391.490 ;
        RECT 2731.445 3390.490 2731.615 3391.490 ;
        RECT 2736.995 3390.490 2737.165 3391.490 ;
        RECT 2737.535 3390.490 2737.705 3391.490 ;
        RECT 2743.085 3390.490 2743.255 3391.490 ;
        RECT 2743.625 3390.490 2743.795 3391.490 ;
        RECT 2749.175 3390.490 2749.345 3391.490 ;
        RECT 2713.515 3390.260 2718.555 3390.430 ;
        RECT 2719.605 3390.260 2724.645 3390.430 ;
        RECT 2725.695 3390.260 2730.735 3390.430 ;
        RECT 2731.785 3390.260 2736.825 3390.430 ;
        RECT 2737.875 3390.260 2742.915 3390.430 ;
        RECT 2743.965 3390.260 2749.005 3390.430 ;
        RECT 2717.045 3385.870 2722.775 3388.030 ;
        RECT 2724.645 3385.870 2730.375 3388.030 ;
        RECT 2732.195 3385.900 2737.925 3388.060 ;
        RECT 2739.745 3385.900 2745.475 3388.060 ;
      LAYER mcon ;
        RECT 2709.675 3451.375 2709.845 3451.545 ;
        RECT 2715.315 3451.375 2715.485 3451.545 ;
        RECT 2715.855 3451.375 2716.025 3451.545 ;
        RECT 2721.495 3451.375 2721.665 3451.545 ;
        RECT 2722.035 3451.375 2722.205 3451.545 ;
        RECT 2727.675 3451.375 2727.845 3451.545 ;
        RECT 2728.215 3451.375 2728.385 3451.545 ;
        RECT 2733.855 3451.375 2734.025 3451.545 ;
        RECT 2734.395 3451.375 2734.565 3451.545 ;
        RECT 2740.035 3451.375 2740.205 3451.545 ;
        RECT 2740.575 3451.375 2740.745 3451.545 ;
        RECT 2746.215 3451.375 2746.385 3451.545 ;
        RECT 2746.755 3451.375 2746.925 3451.545 ;
        RECT 2752.395 3451.375 2752.565 3451.545 ;
        RECT 2710.155 3450.980 2710.325 3451.150 ;
        RECT 2710.515 3450.980 2710.685 3451.150 ;
        RECT 2710.875 3450.980 2711.045 3451.150 ;
        RECT 2711.235 3450.980 2711.405 3451.150 ;
        RECT 2711.595 3450.980 2711.765 3451.150 ;
        RECT 2711.955 3450.980 2712.125 3451.150 ;
        RECT 2712.315 3450.980 2712.485 3451.150 ;
        RECT 2712.675 3450.980 2712.845 3451.150 ;
        RECT 2713.035 3450.980 2713.205 3451.150 ;
        RECT 2713.395 3450.980 2713.565 3451.150 ;
        RECT 2713.755 3450.980 2713.925 3451.150 ;
        RECT 2714.115 3450.980 2714.285 3451.150 ;
        RECT 2714.475 3450.980 2714.645 3451.150 ;
        RECT 2714.835 3450.980 2715.005 3451.150 ;
        RECT 2716.335 3450.980 2716.505 3451.150 ;
        RECT 2716.695 3450.980 2716.865 3451.150 ;
        RECT 2717.055 3450.980 2717.225 3451.150 ;
        RECT 2717.415 3450.980 2717.585 3451.150 ;
        RECT 2717.775 3450.980 2717.945 3451.150 ;
        RECT 2718.135 3450.980 2718.305 3451.150 ;
        RECT 2718.495 3450.980 2718.665 3451.150 ;
        RECT 2718.855 3450.980 2719.025 3451.150 ;
        RECT 2719.215 3450.980 2719.385 3451.150 ;
        RECT 2719.575 3450.980 2719.745 3451.150 ;
        RECT 2719.935 3450.980 2720.105 3451.150 ;
        RECT 2720.295 3450.980 2720.465 3451.150 ;
        RECT 2720.655 3450.980 2720.825 3451.150 ;
        RECT 2721.015 3450.980 2721.185 3451.150 ;
        RECT 2722.515 3450.980 2722.685 3451.150 ;
        RECT 2722.875 3450.980 2723.045 3451.150 ;
        RECT 2723.235 3450.980 2723.405 3451.150 ;
        RECT 2723.595 3450.980 2723.765 3451.150 ;
        RECT 2723.955 3450.980 2724.125 3451.150 ;
        RECT 2724.315 3450.980 2724.485 3451.150 ;
        RECT 2724.675 3450.980 2724.845 3451.150 ;
        RECT 2725.035 3450.980 2725.205 3451.150 ;
        RECT 2725.395 3450.980 2725.565 3451.150 ;
        RECT 2725.755 3450.980 2725.925 3451.150 ;
        RECT 2726.115 3450.980 2726.285 3451.150 ;
        RECT 2726.475 3450.980 2726.645 3451.150 ;
        RECT 2726.835 3450.980 2727.005 3451.150 ;
        RECT 2727.195 3450.980 2727.365 3451.150 ;
        RECT 2728.695 3450.980 2728.865 3451.150 ;
        RECT 2729.055 3450.980 2729.225 3451.150 ;
        RECT 2729.415 3450.980 2729.585 3451.150 ;
        RECT 2729.775 3450.980 2729.945 3451.150 ;
        RECT 2730.135 3450.980 2730.305 3451.150 ;
        RECT 2730.495 3450.980 2730.665 3451.150 ;
        RECT 2730.855 3450.980 2731.025 3451.150 ;
        RECT 2731.215 3450.980 2731.385 3451.150 ;
        RECT 2731.575 3450.980 2731.745 3451.150 ;
        RECT 2731.935 3450.980 2732.105 3451.150 ;
        RECT 2732.295 3450.980 2732.465 3451.150 ;
        RECT 2732.655 3450.980 2732.825 3451.150 ;
        RECT 2733.015 3450.980 2733.185 3451.150 ;
        RECT 2733.375 3450.980 2733.545 3451.150 ;
        RECT 2734.875 3450.980 2735.045 3451.150 ;
        RECT 2735.235 3450.980 2735.405 3451.150 ;
        RECT 2735.595 3450.980 2735.765 3451.150 ;
        RECT 2735.955 3450.980 2736.125 3451.150 ;
        RECT 2736.315 3450.980 2736.485 3451.150 ;
        RECT 2736.675 3450.980 2736.845 3451.150 ;
        RECT 2737.035 3450.980 2737.205 3451.150 ;
        RECT 2737.395 3450.980 2737.565 3451.150 ;
        RECT 2737.755 3450.980 2737.925 3451.150 ;
        RECT 2738.115 3450.980 2738.285 3451.150 ;
        RECT 2738.475 3450.980 2738.645 3451.150 ;
        RECT 2738.835 3450.980 2739.005 3451.150 ;
        RECT 2739.195 3450.980 2739.365 3451.150 ;
        RECT 2739.555 3450.980 2739.725 3451.150 ;
        RECT 2741.055 3450.980 2741.225 3451.150 ;
        RECT 2741.415 3450.980 2741.585 3451.150 ;
        RECT 2741.775 3450.980 2741.945 3451.150 ;
        RECT 2742.135 3450.980 2742.305 3451.150 ;
        RECT 2742.495 3450.980 2742.665 3451.150 ;
        RECT 2742.855 3450.980 2743.025 3451.150 ;
        RECT 2743.215 3450.980 2743.385 3451.150 ;
        RECT 2743.575 3450.980 2743.745 3451.150 ;
        RECT 2743.935 3450.980 2744.105 3451.150 ;
        RECT 2744.295 3450.980 2744.465 3451.150 ;
        RECT 2744.655 3450.980 2744.825 3451.150 ;
        RECT 2745.015 3450.980 2745.185 3451.150 ;
        RECT 2745.375 3450.980 2745.545 3451.150 ;
        RECT 2745.735 3450.980 2745.905 3451.150 ;
        RECT 2747.235 3450.980 2747.405 3451.150 ;
        RECT 2747.595 3450.980 2747.765 3451.150 ;
        RECT 2747.955 3450.980 2748.125 3451.150 ;
        RECT 2748.315 3450.980 2748.485 3451.150 ;
        RECT 2748.675 3450.980 2748.845 3451.150 ;
        RECT 2749.035 3450.980 2749.205 3451.150 ;
        RECT 2749.395 3450.980 2749.565 3451.150 ;
        RECT 2749.755 3450.980 2749.925 3451.150 ;
        RECT 2750.115 3450.980 2750.285 3451.150 ;
        RECT 2750.475 3450.980 2750.645 3451.150 ;
        RECT 2750.835 3450.980 2751.005 3451.150 ;
        RECT 2751.195 3450.980 2751.365 3451.150 ;
        RECT 2751.555 3450.980 2751.725 3451.150 ;
        RECT 2751.915 3450.980 2752.085 3451.150 ;
        RECT 2709.675 3448.675 2709.845 3448.845 ;
        RECT 2715.315 3448.675 2715.485 3448.845 ;
        RECT 2715.855 3448.675 2716.025 3448.845 ;
        RECT 2721.495 3448.675 2721.665 3448.845 ;
        RECT 2722.035 3448.675 2722.205 3448.845 ;
        RECT 2727.675 3448.675 2727.845 3448.845 ;
        RECT 2728.215 3448.675 2728.385 3448.845 ;
        RECT 2733.855 3448.675 2734.025 3448.845 ;
        RECT 2734.395 3448.675 2734.565 3448.845 ;
        RECT 2740.035 3448.675 2740.205 3448.845 ;
        RECT 2740.575 3448.675 2740.745 3448.845 ;
        RECT 2746.215 3448.675 2746.385 3448.845 ;
        RECT 2746.755 3448.675 2746.925 3448.845 ;
        RECT 2752.395 3448.675 2752.565 3448.845 ;
        RECT 2710.155 3448.280 2710.325 3448.450 ;
        RECT 2710.515 3448.280 2710.685 3448.450 ;
        RECT 2710.875 3448.280 2711.045 3448.450 ;
        RECT 2711.235 3448.280 2711.405 3448.450 ;
        RECT 2711.595 3448.280 2711.765 3448.450 ;
        RECT 2711.955 3448.280 2712.125 3448.450 ;
        RECT 2712.315 3448.280 2712.485 3448.450 ;
        RECT 2712.675 3448.280 2712.845 3448.450 ;
        RECT 2713.035 3448.280 2713.205 3448.450 ;
        RECT 2713.395 3448.280 2713.565 3448.450 ;
        RECT 2713.755 3448.280 2713.925 3448.450 ;
        RECT 2714.115 3448.280 2714.285 3448.450 ;
        RECT 2714.475 3448.280 2714.645 3448.450 ;
        RECT 2714.835 3448.280 2715.005 3448.450 ;
        RECT 2716.335 3448.280 2716.505 3448.450 ;
        RECT 2716.695 3448.280 2716.865 3448.450 ;
        RECT 2717.055 3448.280 2717.225 3448.450 ;
        RECT 2717.415 3448.280 2717.585 3448.450 ;
        RECT 2717.775 3448.280 2717.945 3448.450 ;
        RECT 2718.135 3448.280 2718.305 3448.450 ;
        RECT 2718.495 3448.280 2718.665 3448.450 ;
        RECT 2718.855 3448.280 2719.025 3448.450 ;
        RECT 2719.215 3448.280 2719.385 3448.450 ;
        RECT 2719.575 3448.280 2719.745 3448.450 ;
        RECT 2719.935 3448.280 2720.105 3448.450 ;
        RECT 2720.295 3448.280 2720.465 3448.450 ;
        RECT 2720.655 3448.280 2720.825 3448.450 ;
        RECT 2721.015 3448.280 2721.185 3448.450 ;
        RECT 2722.515 3448.280 2722.685 3448.450 ;
        RECT 2722.875 3448.280 2723.045 3448.450 ;
        RECT 2723.235 3448.280 2723.405 3448.450 ;
        RECT 2723.595 3448.280 2723.765 3448.450 ;
        RECT 2723.955 3448.280 2724.125 3448.450 ;
        RECT 2724.315 3448.280 2724.485 3448.450 ;
        RECT 2724.675 3448.280 2724.845 3448.450 ;
        RECT 2725.035 3448.280 2725.205 3448.450 ;
        RECT 2725.395 3448.280 2725.565 3448.450 ;
        RECT 2725.755 3448.280 2725.925 3448.450 ;
        RECT 2726.115 3448.280 2726.285 3448.450 ;
        RECT 2726.475 3448.280 2726.645 3448.450 ;
        RECT 2726.835 3448.280 2727.005 3448.450 ;
        RECT 2727.195 3448.280 2727.365 3448.450 ;
        RECT 2728.695 3448.280 2728.865 3448.450 ;
        RECT 2729.055 3448.280 2729.225 3448.450 ;
        RECT 2729.415 3448.280 2729.585 3448.450 ;
        RECT 2729.775 3448.280 2729.945 3448.450 ;
        RECT 2730.135 3448.280 2730.305 3448.450 ;
        RECT 2730.495 3448.280 2730.665 3448.450 ;
        RECT 2730.855 3448.280 2731.025 3448.450 ;
        RECT 2731.215 3448.280 2731.385 3448.450 ;
        RECT 2731.575 3448.280 2731.745 3448.450 ;
        RECT 2731.935 3448.280 2732.105 3448.450 ;
        RECT 2732.295 3448.280 2732.465 3448.450 ;
        RECT 2732.655 3448.280 2732.825 3448.450 ;
        RECT 2733.015 3448.280 2733.185 3448.450 ;
        RECT 2733.375 3448.280 2733.545 3448.450 ;
        RECT 2734.875 3448.280 2735.045 3448.450 ;
        RECT 2735.235 3448.280 2735.405 3448.450 ;
        RECT 2735.595 3448.280 2735.765 3448.450 ;
        RECT 2735.955 3448.280 2736.125 3448.450 ;
        RECT 2736.315 3448.280 2736.485 3448.450 ;
        RECT 2736.675 3448.280 2736.845 3448.450 ;
        RECT 2737.035 3448.280 2737.205 3448.450 ;
        RECT 2737.395 3448.280 2737.565 3448.450 ;
        RECT 2737.755 3448.280 2737.925 3448.450 ;
        RECT 2738.115 3448.280 2738.285 3448.450 ;
        RECT 2738.475 3448.280 2738.645 3448.450 ;
        RECT 2738.835 3448.280 2739.005 3448.450 ;
        RECT 2739.195 3448.280 2739.365 3448.450 ;
        RECT 2739.555 3448.280 2739.725 3448.450 ;
        RECT 2741.055 3448.280 2741.225 3448.450 ;
        RECT 2741.415 3448.280 2741.585 3448.450 ;
        RECT 2741.775 3448.280 2741.945 3448.450 ;
        RECT 2742.135 3448.280 2742.305 3448.450 ;
        RECT 2742.495 3448.280 2742.665 3448.450 ;
        RECT 2742.855 3448.280 2743.025 3448.450 ;
        RECT 2743.215 3448.280 2743.385 3448.450 ;
        RECT 2743.575 3448.280 2743.745 3448.450 ;
        RECT 2743.935 3448.280 2744.105 3448.450 ;
        RECT 2744.295 3448.280 2744.465 3448.450 ;
        RECT 2744.655 3448.280 2744.825 3448.450 ;
        RECT 2745.015 3448.280 2745.185 3448.450 ;
        RECT 2745.375 3448.280 2745.545 3448.450 ;
        RECT 2745.735 3448.280 2745.905 3448.450 ;
        RECT 2747.235 3448.280 2747.405 3448.450 ;
        RECT 2747.595 3448.280 2747.765 3448.450 ;
        RECT 2747.955 3448.280 2748.125 3448.450 ;
        RECT 2748.315 3448.280 2748.485 3448.450 ;
        RECT 2748.675 3448.280 2748.845 3448.450 ;
        RECT 2749.035 3448.280 2749.205 3448.450 ;
        RECT 2749.395 3448.280 2749.565 3448.450 ;
        RECT 2749.755 3448.280 2749.925 3448.450 ;
        RECT 2750.115 3448.280 2750.285 3448.450 ;
        RECT 2750.475 3448.280 2750.645 3448.450 ;
        RECT 2750.835 3448.280 2751.005 3448.450 ;
        RECT 2751.195 3448.280 2751.365 3448.450 ;
        RECT 2751.555 3448.280 2751.725 3448.450 ;
        RECT 2751.915 3448.280 2752.085 3448.450 ;
        RECT 2709.675 3445.975 2709.845 3446.145 ;
        RECT 2715.315 3445.975 2715.485 3446.145 ;
        RECT 2715.855 3445.975 2716.025 3446.145 ;
        RECT 2721.495 3445.975 2721.665 3446.145 ;
        RECT 2722.035 3445.975 2722.205 3446.145 ;
        RECT 2727.675 3445.975 2727.845 3446.145 ;
        RECT 2728.215 3445.975 2728.385 3446.145 ;
        RECT 2733.855 3445.975 2734.025 3446.145 ;
        RECT 2734.395 3445.975 2734.565 3446.145 ;
        RECT 2740.035 3445.975 2740.205 3446.145 ;
        RECT 2740.575 3445.975 2740.745 3446.145 ;
        RECT 2746.215 3445.975 2746.385 3446.145 ;
        RECT 2746.755 3445.975 2746.925 3446.145 ;
        RECT 2752.395 3445.975 2752.565 3446.145 ;
        RECT 2710.155 3445.580 2710.325 3445.750 ;
        RECT 2710.515 3445.580 2710.685 3445.750 ;
        RECT 2710.875 3445.580 2711.045 3445.750 ;
        RECT 2711.235 3445.580 2711.405 3445.750 ;
        RECT 2711.595 3445.580 2711.765 3445.750 ;
        RECT 2711.955 3445.580 2712.125 3445.750 ;
        RECT 2712.315 3445.580 2712.485 3445.750 ;
        RECT 2712.675 3445.580 2712.845 3445.750 ;
        RECT 2713.035 3445.580 2713.205 3445.750 ;
        RECT 2713.395 3445.580 2713.565 3445.750 ;
        RECT 2713.755 3445.580 2713.925 3445.750 ;
        RECT 2714.115 3445.580 2714.285 3445.750 ;
        RECT 2714.475 3445.580 2714.645 3445.750 ;
        RECT 2714.835 3445.580 2715.005 3445.750 ;
        RECT 2716.335 3445.580 2716.505 3445.750 ;
        RECT 2716.695 3445.580 2716.865 3445.750 ;
        RECT 2717.055 3445.580 2717.225 3445.750 ;
        RECT 2717.415 3445.580 2717.585 3445.750 ;
        RECT 2717.775 3445.580 2717.945 3445.750 ;
        RECT 2718.135 3445.580 2718.305 3445.750 ;
        RECT 2718.495 3445.580 2718.665 3445.750 ;
        RECT 2718.855 3445.580 2719.025 3445.750 ;
        RECT 2719.215 3445.580 2719.385 3445.750 ;
        RECT 2719.575 3445.580 2719.745 3445.750 ;
        RECT 2719.935 3445.580 2720.105 3445.750 ;
        RECT 2720.295 3445.580 2720.465 3445.750 ;
        RECT 2720.655 3445.580 2720.825 3445.750 ;
        RECT 2721.015 3445.580 2721.185 3445.750 ;
        RECT 2722.515 3445.580 2722.685 3445.750 ;
        RECT 2722.875 3445.580 2723.045 3445.750 ;
        RECT 2723.235 3445.580 2723.405 3445.750 ;
        RECT 2723.595 3445.580 2723.765 3445.750 ;
        RECT 2723.955 3445.580 2724.125 3445.750 ;
        RECT 2724.315 3445.580 2724.485 3445.750 ;
        RECT 2724.675 3445.580 2724.845 3445.750 ;
        RECT 2725.035 3445.580 2725.205 3445.750 ;
        RECT 2725.395 3445.580 2725.565 3445.750 ;
        RECT 2725.755 3445.580 2725.925 3445.750 ;
        RECT 2726.115 3445.580 2726.285 3445.750 ;
        RECT 2726.475 3445.580 2726.645 3445.750 ;
        RECT 2726.835 3445.580 2727.005 3445.750 ;
        RECT 2727.195 3445.580 2727.365 3445.750 ;
        RECT 2728.695 3445.580 2728.865 3445.750 ;
        RECT 2729.055 3445.580 2729.225 3445.750 ;
        RECT 2729.415 3445.580 2729.585 3445.750 ;
        RECT 2729.775 3445.580 2729.945 3445.750 ;
        RECT 2730.135 3445.580 2730.305 3445.750 ;
        RECT 2730.495 3445.580 2730.665 3445.750 ;
        RECT 2730.855 3445.580 2731.025 3445.750 ;
        RECT 2731.215 3445.580 2731.385 3445.750 ;
        RECT 2731.575 3445.580 2731.745 3445.750 ;
        RECT 2731.935 3445.580 2732.105 3445.750 ;
        RECT 2732.295 3445.580 2732.465 3445.750 ;
        RECT 2732.655 3445.580 2732.825 3445.750 ;
        RECT 2733.015 3445.580 2733.185 3445.750 ;
        RECT 2733.375 3445.580 2733.545 3445.750 ;
        RECT 2734.875 3445.580 2735.045 3445.750 ;
        RECT 2735.235 3445.580 2735.405 3445.750 ;
        RECT 2735.595 3445.580 2735.765 3445.750 ;
        RECT 2735.955 3445.580 2736.125 3445.750 ;
        RECT 2736.315 3445.580 2736.485 3445.750 ;
        RECT 2736.675 3445.580 2736.845 3445.750 ;
        RECT 2737.035 3445.580 2737.205 3445.750 ;
        RECT 2737.395 3445.580 2737.565 3445.750 ;
        RECT 2737.755 3445.580 2737.925 3445.750 ;
        RECT 2738.115 3445.580 2738.285 3445.750 ;
        RECT 2738.475 3445.580 2738.645 3445.750 ;
        RECT 2738.835 3445.580 2739.005 3445.750 ;
        RECT 2739.195 3445.580 2739.365 3445.750 ;
        RECT 2739.555 3445.580 2739.725 3445.750 ;
        RECT 2741.055 3445.580 2741.225 3445.750 ;
        RECT 2741.415 3445.580 2741.585 3445.750 ;
        RECT 2741.775 3445.580 2741.945 3445.750 ;
        RECT 2742.135 3445.580 2742.305 3445.750 ;
        RECT 2742.495 3445.580 2742.665 3445.750 ;
        RECT 2742.855 3445.580 2743.025 3445.750 ;
        RECT 2743.215 3445.580 2743.385 3445.750 ;
        RECT 2743.575 3445.580 2743.745 3445.750 ;
        RECT 2743.935 3445.580 2744.105 3445.750 ;
        RECT 2744.295 3445.580 2744.465 3445.750 ;
        RECT 2744.655 3445.580 2744.825 3445.750 ;
        RECT 2745.015 3445.580 2745.185 3445.750 ;
        RECT 2745.375 3445.580 2745.545 3445.750 ;
        RECT 2745.735 3445.580 2745.905 3445.750 ;
        RECT 2747.235 3445.580 2747.405 3445.750 ;
        RECT 2747.595 3445.580 2747.765 3445.750 ;
        RECT 2747.955 3445.580 2748.125 3445.750 ;
        RECT 2748.315 3445.580 2748.485 3445.750 ;
        RECT 2748.675 3445.580 2748.845 3445.750 ;
        RECT 2749.035 3445.580 2749.205 3445.750 ;
        RECT 2749.395 3445.580 2749.565 3445.750 ;
        RECT 2749.755 3445.580 2749.925 3445.750 ;
        RECT 2750.115 3445.580 2750.285 3445.750 ;
        RECT 2750.475 3445.580 2750.645 3445.750 ;
        RECT 2750.835 3445.580 2751.005 3445.750 ;
        RECT 2751.195 3445.580 2751.365 3445.750 ;
        RECT 2751.555 3445.580 2751.725 3445.750 ;
        RECT 2751.915 3445.580 2752.085 3445.750 ;
        RECT 2709.675 3443.275 2709.845 3443.445 ;
        RECT 2715.315 3443.275 2715.485 3443.445 ;
        RECT 2715.855 3443.275 2716.025 3443.445 ;
        RECT 2721.495 3443.275 2721.665 3443.445 ;
        RECT 2722.035 3443.275 2722.205 3443.445 ;
        RECT 2727.675 3443.275 2727.845 3443.445 ;
        RECT 2728.215 3443.275 2728.385 3443.445 ;
        RECT 2733.855 3443.275 2734.025 3443.445 ;
        RECT 2734.395 3443.275 2734.565 3443.445 ;
        RECT 2740.035 3443.275 2740.205 3443.445 ;
        RECT 2740.575 3443.275 2740.745 3443.445 ;
        RECT 2746.215 3443.275 2746.385 3443.445 ;
        RECT 2746.755 3443.275 2746.925 3443.445 ;
        RECT 2752.395 3443.275 2752.565 3443.445 ;
        RECT 2710.155 3442.880 2710.325 3443.050 ;
        RECT 2710.515 3442.880 2710.685 3443.050 ;
        RECT 2710.875 3442.880 2711.045 3443.050 ;
        RECT 2711.235 3442.880 2711.405 3443.050 ;
        RECT 2711.595 3442.880 2711.765 3443.050 ;
        RECT 2711.955 3442.880 2712.125 3443.050 ;
        RECT 2712.315 3442.880 2712.485 3443.050 ;
        RECT 2712.675 3442.880 2712.845 3443.050 ;
        RECT 2713.035 3442.880 2713.205 3443.050 ;
        RECT 2713.395 3442.880 2713.565 3443.050 ;
        RECT 2713.755 3442.880 2713.925 3443.050 ;
        RECT 2714.115 3442.880 2714.285 3443.050 ;
        RECT 2714.475 3442.880 2714.645 3443.050 ;
        RECT 2714.835 3442.880 2715.005 3443.050 ;
        RECT 2716.335 3442.880 2716.505 3443.050 ;
        RECT 2716.695 3442.880 2716.865 3443.050 ;
        RECT 2717.055 3442.880 2717.225 3443.050 ;
        RECT 2717.415 3442.880 2717.585 3443.050 ;
        RECT 2717.775 3442.880 2717.945 3443.050 ;
        RECT 2718.135 3442.880 2718.305 3443.050 ;
        RECT 2718.495 3442.880 2718.665 3443.050 ;
        RECT 2718.855 3442.880 2719.025 3443.050 ;
        RECT 2719.215 3442.880 2719.385 3443.050 ;
        RECT 2719.575 3442.880 2719.745 3443.050 ;
        RECT 2719.935 3442.880 2720.105 3443.050 ;
        RECT 2720.295 3442.880 2720.465 3443.050 ;
        RECT 2720.655 3442.880 2720.825 3443.050 ;
        RECT 2721.015 3442.880 2721.185 3443.050 ;
        RECT 2722.515 3442.880 2722.685 3443.050 ;
        RECT 2722.875 3442.880 2723.045 3443.050 ;
        RECT 2723.235 3442.880 2723.405 3443.050 ;
        RECT 2723.595 3442.880 2723.765 3443.050 ;
        RECT 2723.955 3442.880 2724.125 3443.050 ;
        RECT 2724.315 3442.880 2724.485 3443.050 ;
        RECT 2724.675 3442.880 2724.845 3443.050 ;
        RECT 2725.035 3442.880 2725.205 3443.050 ;
        RECT 2725.395 3442.880 2725.565 3443.050 ;
        RECT 2725.755 3442.880 2725.925 3443.050 ;
        RECT 2726.115 3442.880 2726.285 3443.050 ;
        RECT 2726.475 3442.880 2726.645 3443.050 ;
        RECT 2726.835 3442.880 2727.005 3443.050 ;
        RECT 2727.195 3442.880 2727.365 3443.050 ;
        RECT 2728.695 3442.880 2728.865 3443.050 ;
        RECT 2729.055 3442.880 2729.225 3443.050 ;
        RECT 2729.415 3442.880 2729.585 3443.050 ;
        RECT 2729.775 3442.880 2729.945 3443.050 ;
        RECT 2730.135 3442.880 2730.305 3443.050 ;
        RECT 2730.495 3442.880 2730.665 3443.050 ;
        RECT 2730.855 3442.880 2731.025 3443.050 ;
        RECT 2731.215 3442.880 2731.385 3443.050 ;
        RECT 2731.575 3442.880 2731.745 3443.050 ;
        RECT 2731.935 3442.880 2732.105 3443.050 ;
        RECT 2732.295 3442.880 2732.465 3443.050 ;
        RECT 2732.655 3442.880 2732.825 3443.050 ;
        RECT 2733.015 3442.880 2733.185 3443.050 ;
        RECT 2733.375 3442.880 2733.545 3443.050 ;
        RECT 2734.875 3442.880 2735.045 3443.050 ;
        RECT 2735.235 3442.880 2735.405 3443.050 ;
        RECT 2735.595 3442.880 2735.765 3443.050 ;
        RECT 2735.955 3442.880 2736.125 3443.050 ;
        RECT 2736.315 3442.880 2736.485 3443.050 ;
        RECT 2736.675 3442.880 2736.845 3443.050 ;
        RECT 2737.035 3442.880 2737.205 3443.050 ;
        RECT 2737.395 3442.880 2737.565 3443.050 ;
        RECT 2737.755 3442.880 2737.925 3443.050 ;
        RECT 2738.115 3442.880 2738.285 3443.050 ;
        RECT 2738.475 3442.880 2738.645 3443.050 ;
        RECT 2738.835 3442.880 2739.005 3443.050 ;
        RECT 2739.195 3442.880 2739.365 3443.050 ;
        RECT 2739.555 3442.880 2739.725 3443.050 ;
        RECT 2741.055 3442.880 2741.225 3443.050 ;
        RECT 2741.415 3442.880 2741.585 3443.050 ;
        RECT 2741.775 3442.880 2741.945 3443.050 ;
        RECT 2742.135 3442.880 2742.305 3443.050 ;
        RECT 2742.495 3442.880 2742.665 3443.050 ;
        RECT 2742.855 3442.880 2743.025 3443.050 ;
        RECT 2743.215 3442.880 2743.385 3443.050 ;
        RECT 2743.575 3442.880 2743.745 3443.050 ;
        RECT 2743.935 3442.880 2744.105 3443.050 ;
        RECT 2744.295 3442.880 2744.465 3443.050 ;
        RECT 2744.655 3442.880 2744.825 3443.050 ;
        RECT 2745.015 3442.880 2745.185 3443.050 ;
        RECT 2745.375 3442.880 2745.545 3443.050 ;
        RECT 2745.735 3442.880 2745.905 3443.050 ;
        RECT 2747.235 3442.880 2747.405 3443.050 ;
        RECT 2747.595 3442.880 2747.765 3443.050 ;
        RECT 2747.955 3442.880 2748.125 3443.050 ;
        RECT 2748.315 3442.880 2748.485 3443.050 ;
        RECT 2748.675 3442.880 2748.845 3443.050 ;
        RECT 2749.035 3442.880 2749.205 3443.050 ;
        RECT 2749.395 3442.880 2749.565 3443.050 ;
        RECT 2749.755 3442.880 2749.925 3443.050 ;
        RECT 2750.115 3442.880 2750.285 3443.050 ;
        RECT 2750.475 3442.880 2750.645 3443.050 ;
        RECT 2750.835 3442.880 2751.005 3443.050 ;
        RECT 2751.195 3442.880 2751.365 3443.050 ;
        RECT 2751.555 3442.880 2751.725 3443.050 ;
        RECT 2751.915 3442.880 2752.085 3443.050 ;
        RECT 2709.675 3440.375 2709.845 3440.545 ;
        RECT 2715.315 3440.375 2715.485 3440.545 ;
        RECT 2715.855 3440.375 2716.025 3440.545 ;
        RECT 2721.495 3440.375 2721.665 3440.545 ;
        RECT 2722.035 3440.375 2722.205 3440.545 ;
        RECT 2727.675 3440.375 2727.845 3440.545 ;
        RECT 2728.215 3440.375 2728.385 3440.545 ;
        RECT 2733.855 3440.375 2734.025 3440.545 ;
        RECT 2734.395 3440.375 2734.565 3440.545 ;
        RECT 2740.035 3440.375 2740.205 3440.545 ;
        RECT 2740.575 3440.375 2740.745 3440.545 ;
        RECT 2746.215 3440.375 2746.385 3440.545 ;
        RECT 2746.755 3440.375 2746.925 3440.545 ;
        RECT 2752.395 3440.375 2752.565 3440.545 ;
        RECT 2710.155 3439.980 2710.325 3440.150 ;
        RECT 2710.515 3439.980 2710.685 3440.150 ;
        RECT 2710.875 3439.980 2711.045 3440.150 ;
        RECT 2711.235 3439.980 2711.405 3440.150 ;
        RECT 2711.595 3439.980 2711.765 3440.150 ;
        RECT 2711.955 3439.980 2712.125 3440.150 ;
        RECT 2712.315 3439.980 2712.485 3440.150 ;
        RECT 2712.675 3439.980 2712.845 3440.150 ;
        RECT 2713.035 3439.980 2713.205 3440.150 ;
        RECT 2713.395 3439.980 2713.565 3440.150 ;
        RECT 2713.755 3439.980 2713.925 3440.150 ;
        RECT 2714.115 3439.980 2714.285 3440.150 ;
        RECT 2714.475 3439.980 2714.645 3440.150 ;
        RECT 2714.835 3439.980 2715.005 3440.150 ;
        RECT 2716.335 3439.980 2716.505 3440.150 ;
        RECT 2716.695 3439.980 2716.865 3440.150 ;
        RECT 2717.055 3439.980 2717.225 3440.150 ;
        RECT 2717.415 3439.980 2717.585 3440.150 ;
        RECT 2717.775 3439.980 2717.945 3440.150 ;
        RECT 2718.135 3439.980 2718.305 3440.150 ;
        RECT 2718.495 3439.980 2718.665 3440.150 ;
        RECT 2718.855 3439.980 2719.025 3440.150 ;
        RECT 2719.215 3439.980 2719.385 3440.150 ;
        RECT 2719.575 3439.980 2719.745 3440.150 ;
        RECT 2719.935 3439.980 2720.105 3440.150 ;
        RECT 2720.295 3439.980 2720.465 3440.150 ;
        RECT 2720.655 3439.980 2720.825 3440.150 ;
        RECT 2721.015 3439.980 2721.185 3440.150 ;
        RECT 2722.515 3439.980 2722.685 3440.150 ;
        RECT 2722.875 3439.980 2723.045 3440.150 ;
        RECT 2723.235 3439.980 2723.405 3440.150 ;
        RECT 2723.595 3439.980 2723.765 3440.150 ;
        RECT 2723.955 3439.980 2724.125 3440.150 ;
        RECT 2724.315 3439.980 2724.485 3440.150 ;
        RECT 2724.675 3439.980 2724.845 3440.150 ;
        RECT 2725.035 3439.980 2725.205 3440.150 ;
        RECT 2725.395 3439.980 2725.565 3440.150 ;
        RECT 2725.755 3439.980 2725.925 3440.150 ;
        RECT 2726.115 3439.980 2726.285 3440.150 ;
        RECT 2726.475 3439.980 2726.645 3440.150 ;
        RECT 2726.835 3439.980 2727.005 3440.150 ;
        RECT 2727.195 3439.980 2727.365 3440.150 ;
        RECT 2728.695 3439.980 2728.865 3440.150 ;
        RECT 2729.055 3439.980 2729.225 3440.150 ;
        RECT 2729.415 3439.980 2729.585 3440.150 ;
        RECT 2729.775 3439.980 2729.945 3440.150 ;
        RECT 2730.135 3439.980 2730.305 3440.150 ;
        RECT 2730.495 3439.980 2730.665 3440.150 ;
        RECT 2730.855 3439.980 2731.025 3440.150 ;
        RECT 2731.215 3439.980 2731.385 3440.150 ;
        RECT 2731.575 3439.980 2731.745 3440.150 ;
        RECT 2731.935 3439.980 2732.105 3440.150 ;
        RECT 2732.295 3439.980 2732.465 3440.150 ;
        RECT 2732.655 3439.980 2732.825 3440.150 ;
        RECT 2733.015 3439.980 2733.185 3440.150 ;
        RECT 2733.375 3439.980 2733.545 3440.150 ;
        RECT 2734.875 3439.980 2735.045 3440.150 ;
        RECT 2735.235 3439.980 2735.405 3440.150 ;
        RECT 2735.595 3439.980 2735.765 3440.150 ;
        RECT 2735.955 3439.980 2736.125 3440.150 ;
        RECT 2736.315 3439.980 2736.485 3440.150 ;
        RECT 2736.675 3439.980 2736.845 3440.150 ;
        RECT 2737.035 3439.980 2737.205 3440.150 ;
        RECT 2737.395 3439.980 2737.565 3440.150 ;
        RECT 2737.755 3439.980 2737.925 3440.150 ;
        RECT 2738.115 3439.980 2738.285 3440.150 ;
        RECT 2738.475 3439.980 2738.645 3440.150 ;
        RECT 2738.835 3439.980 2739.005 3440.150 ;
        RECT 2739.195 3439.980 2739.365 3440.150 ;
        RECT 2739.555 3439.980 2739.725 3440.150 ;
        RECT 2741.055 3439.980 2741.225 3440.150 ;
        RECT 2741.415 3439.980 2741.585 3440.150 ;
        RECT 2741.775 3439.980 2741.945 3440.150 ;
        RECT 2742.135 3439.980 2742.305 3440.150 ;
        RECT 2742.495 3439.980 2742.665 3440.150 ;
        RECT 2742.855 3439.980 2743.025 3440.150 ;
        RECT 2743.215 3439.980 2743.385 3440.150 ;
        RECT 2743.575 3439.980 2743.745 3440.150 ;
        RECT 2743.935 3439.980 2744.105 3440.150 ;
        RECT 2744.295 3439.980 2744.465 3440.150 ;
        RECT 2744.655 3439.980 2744.825 3440.150 ;
        RECT 2745.015 3439.980 2745.185 3440.150 ;
        RECT 2745.375 3439.980 2745.545 3440.150 ;
        RECT 2745.735 3439.980 2745.905 3440.150 ;
        RECT 2747.235 3439.980 2747.405 3440.150 ;
        RECT 2747.595 3439.980 2747.765 3440.150 ;
        RECT 2747.955 3439.980 2748.125 3440.150 ;
        RECT 2748.315 3439.980 2748.485 3440.150 ;
        RECT 2748.675 3439.980 2748.845 3440.150 ;
        RECT 2749.035 3439.980 2749.205 3440.150 ;
        RECT 2749.395 3439.980 2749.565 3440.150 ;
        RECT 2749.755 3439.980 2749.925 3440.150 ;
        RECT 2750.115 3439.980 2750.285 3440.150 ;
        RECT 2750.475 3439.980 2750.645 3440.150 ;
        RECT 2750.835 3439.980 2751.005 3440.150 ;
        RECT 2751.195 3439.980 2751.365 3440.150 ;
        RECT 2751.555 3439.980 2751.725 3440.150 ;
        RECT 2751.915 3439.980 2752.085 3440.150 ;
        RECT 2681.945 3432.225 2683.915 3437.795 ;
        RECT 2694.100 3432.225 2696.070 3437.795 ;
        RECT 2709.675 3437.475 2709.845 3437.645 ;
        RECT 2715.315 3437.475 2715.485 3437.645 ;
        RECT 2715.855 3437.475 2716.025 3437.645 ;
        RECT 2721.495 3437.475 2721.665 3437.645 ;
        RECT 2722.035 3437.475 2722.205 3437.645 ;
        RECT 2727.675 3437.475 2727.845 3437.645 ;
        RECT 2728.215 3437.475 2728.385 3437.645 ;
        RECT 2733.855 3437.475 2734.025 3437.645 ;
        RECT 2734.395 3437.475 2734.565 3437.645 ;
        RECT 2740.035 3437.475 2740.205 3437.645 ;
        RECT 2740.575 3437.475 2740.745 3437.645 ;
        RECT 2746.215 3437.475 2746.385 3437.645 ;
        RECT 2746.755 3437.475 2746.925 3437.645 ;
        RECT 2752.395 3437.475 2752.565 3437.645 ;
        RECT 2710.155 3437.080 2710.325 3437.250 ;
        RECT 2710.515 3437.080 2710.685 3437.250 ;
        RECT 2710.875 3437.080 2711.045 3437.250 ;
        RECT 2711.235 3437.080 2711.405 3437.250 ;
        RECT 2711.595 3437.080 2711.765 3437.250 ;
        RECT 2711.955 3437.080 2712.125 3437.250 ;
        RECT 2712.315 3437.080 2712.485 3437.250 ;
        RECT 2712.675 3437.080 2712.845 3437.250 ;
        RECT 2713.035 3437.080 2713.205 3437.250 ;
        RECT 2713.395 3437.080 2713.565 3437.250 ;
        RECT 2713.755 3437.080 2713.925 3437.250 ;
        RECT 2714.115 3437.080 2714.285 3437.250 ;
        RECT 2714.475 3437.080 2714.645 3437.250 ;
        RECT 2714.835 3437.080 2715.005 3437.250 ;
        RECT 2716.335 3437.080 2716.505 3437.250 ;
        RECT 2716.695 3437.080 2716.865 3437.250 ;
        RECT 2717.055 3437.080 2717.225 3437.250 ;
        RECT 2717.415 3437.080 2717.585 3437.250 ;
        RECT 2717.775 3437.080 2717.945 3437.250 ;
        RECT 2718.135 3437.080 2718.305 3437.250 ;
        RECT 2718.495 3437.080 2718.665 3437.250 ;
        RECT 2718.855 3437.080 2719.025 3437.250 ;
        RECT 2719.215 3437.080 2719.385 3437.250 ;
        RECT 2719.575 3437.080 2719.745 3437.250 ;
        RECT 2719.935 3437.080 2720.105 3437.250 ;
        RECT 2720.295 3437.080 2720.465 3437.250 ;
        RECT 2720.655 3437.080 2720.825 3437.250 ;
        RECT 2721.015 3437.080 2721.185 3437.250 ;
        RECT 2722.515 3437.080 2722.685 3437.250 ;
        RECT 2722.875 3437.080 2723.045 3437.250 ;
        RECT 2723.235 3437.080 2723.405 3437.250 ;
        RECT 2723.595 3437.080 2723.765 3437.250 ;
        RECT 2723.955 3437.080 2724.125 3437.250 ;
        RECT 2724.315 3437.080 2724.485 3437.250 ;
        RECT 2724.675 3437.080 2724.845 3437.250 ;
        RECT 2725.035 3437.080 2725.205 3437.250 ;
        RECT 2725.395 3437.080 2725.565 3437.250 ;
        RECT 2725.755 3437.080 2725.925 3437.250 ;
        RECT 2726.115 3437.080 2726.285 3437.250 ;
        RECT 2726.475 3437.080 2726.645 3437.250 ;
        RECT 2726.835 3437.080 2727.005 3437.250 ;
        RECT 2727.195 3437.080 2727.365 3437.250 ;
        RECT 2728.695 3437.080 2728.865 3437.250 ;
        RECT 2729.055 3437.080 2729.225 3437.250 ;
        RECT 2729.415 3437.080 2729.585 3437.250 ;
        RECT 2729.775 3437.080 2729.945 3437.250 ;
        RECT 2730.135 3437.080 2730.305 3437.250 ;
        RECT 2730.495 3437.080 2730.665 3437.250 ;
        RECT 2730.855 3437.080 2731.025 3437.250 ;
        RECT 2731.215 3437.080 2731.385 3437.250 ;
        RECT 2731.575 3437.080 2731.745 3437.250 ;
        RECT 2731.935 3437.080 2732.105 3437.250 ;
        RECT 2732.295 3437.080 2732.465 3437.250 ;
        RECT 2732.655 3437.080 2732.825 3437.250 ;
        RECT 2733.015 3437.080 2733.185 3437.250 ;
        RECT 2733.375 3437.080 2733.545 3437.250 ;
        RECT 2734.875 3437.080 2735.045 3437.250 ;
        RECT 2735.235 3437.080 2735.405 3437.250 ;
        RECT 2735.595 3437.080 2735.765 3437.250 ;
        RECT 2735.955 3437.080 2736.125 3437.250 ;
        RECT 2736.315 3437.080 2736.485 3437.250 ;
        RECT 2736.675 3437.080 2736.845 3437.250 ;
        RECT 2737.035 3437.080 2737.205 3437.250 ;
        RECT 2737.395 3437.080 2737.565 3437.250 ;
        RECT 2737.755 3437.080 2737.925 3437.250 ;
        RECT 2738.115 3437.080 2738.285 3437.250 ;
        RECT 2738.475 3437.080 2738.645 3437.250 ;
        RECT 2738.835 3437.080 2739.005 3437.250 ;
        RECT 2739.195 3437.080 2739.365 3437.250 ;
        RECT 2739.555 3437.080 2739.725 3437.250 ;
        RECT 2741.055 3437.080 2741.225 3437.250 ;
        RECT 2741.415 3437.080 2741.585 3437.250 ;
        RECT 2741.775 3437.080 2741.945 3437.250 ;
        RECT 2742.135 3437.080 2742.305 3437.250 ;
        RECT 2742.495 3437.080 2742.665 3437.250 ;
        RECT 2742.855 3437.080 2743.025 3437.250 ;
        RECT 2743.215 3437.080 2743.385 3437.250 ;
        RECT 2743.575 3437.080 2743.745 3437.250 ;
        RECT 2743.935 3437.080 2744.105 3437.250 ;
        RECT 2744.295 3437.080 2744.465 3437.250 ;
        RECT 2744.655 3437.080 2744.825 3437.250 ;
        RECT 2745.015 3437.080 2745.185 3437.250 ;
        RECT 2745.375 3437.080 2745.545 3437.250 ;
        RECT 2745.735 3437.080 2745.905 3437.250 ;
        RECT 2747.235 3437.080 2747.405 3437.250 ;
        RECT 2747.595 3437.080 2747.765 3437.250 ;
        RECT 2747.955 3437.080 2748.125 3437.250 ;
        RECT 2748.315 3437.080 2748.485 3437.250 ;
        RECT 2748.675 3437.080 2748.845 3437.250 ;
        RECT 2749.035 3437.080 2749.205 3437.250 ;
        RECT 2749.395 3437.080 2749.565 3437.250 ;
        RECT 2749.755 3437.080 2749.925 3437.250 ;
        RECT 2750.115 3437.080 2750.285 3437.250 ;
        RECT 2750.475 3437.080 2750.645 3437.250 ;
        RECT 2750.835 3437.080 2751.005 3437.250 ;
        RECT 2751.195 3437.080 2751.365 3437.250 ;
        RECT 2751.555 3437.080 2751.725 3437.250 ;
        RECT 2751.915 3437.080 2752.085 3437.250 ;
        RECT 2700.475 3434.775 2700.645 3434.945 ;
        RECT 2706.115 3434.775 2706.285 3434.945 ;
        RECT 2706.655 3434.775 2706.825 3434.945 ;
        RECT 2712.295 3434.775 2712.465 3434.945 ;
        RECT 2712.835 3434.775 2713.005 3434.945 ;
        RECT 2718.475 3434.775 2718.645 3434.945 ;
        RECT 2719.015 3434.775 2719.185 3434.945 ;
        RECT 2724.655 3434.775 2724.825 3434.945 ;
        RECT 2725.195 3434.775 2725.365 3434.945 ;
        RECT 2730.835 3434.775 2731.005 3434.945 ;
        RECT 2731.375 3434.775 2731.545 3434.945 ;
        RECT 2737.015 3434.775 2737.185 3434.945 ;
        RECT 2737.555 3434.775 2737.725 3434.945 ;
        RECT 2743.195 3434.775 2743.365 3434.945 ;
        RECT 2743.735 3434.775 2743.905 3434.945 ;
        RECT 2749.375 3434.775 2749.545 3434.945 ;
        RECT 2749.915 3434.775 2750.085 3434.945 ;
        RECT 2755.555 3434.775 2755.725 3434.945 ;
        RECT 2756.095 3434.775 2756.265 3434.945 ;
        RECT 2761.735 3434.775 2761.905 3434.945 ;
        RECT 2700.475 3432.075 2700.645 3432.245 ;
        RECT 2706.115 3432.075 2706.285 3432.245 ;
        RECT 2706.655 3432.075 2706.825 3432.245 ;
        RECT 2712.295 3432.075 2712.465 3432.245 ;
        RECT 2712.835 3432.075 2713.005 3432.245 ;
        RECT 2718.475 3432.075 2718.645 3432.245 ;
        RECT 2719.015 3432.075 2719.185 3432.245 ;
        RECT 2724.655 3432.075 2724.825 3432.245 ;
        RECT 2725.195 3432.075 2725.365 3432.245 ;
        RECT 2730.835 3432.075 2731.005 3432.245 ;
        RECT 2731.375 3432.075 2731.545 3432.245 ;
        RECT 2737.015 3432.075 2737.185 3432.245 ;
        RECT 2737.555 3432.075 2737.725 3432.245 ;
        RECT 2743.195 3432.075 2743.365 3432.245 ;
        RECT 2743.735 3432.075 2743.905 3432.245 ;
        RECT 2749.375 3432.075 2749.545 3432.245 ;
        RECT 2749.915 3432.075 2750.085 3432.245 ;
        RECT 2755.555 3432.075 2755.725 3432.245 ;
        RECT 2756.095 3432.075 2756.265 3432.245 ;
        RECT 2761.735 3432.075 2761.905 3432.245 ;
        RECT 2767.245 3432.225 2769.215 3437.795 ;
        RECT 2779.400 3432.225 2781.370 3437.795 ;
        RECT 2681.945 3424.875 2683.915 3430.445 ;
        RECT 2694.100 3424.875 2696.070 3430.445 ;
        RECT 2700.475 3429.375 2700.645 3429.545 ;
        RECT 2706.115 3429.375 2706.285 3429.545 ;
        RECT 2706.655 3429.375 2706.825 3429.545 ;
        RECT 2712.295 3429.375 2712.465 3429.545 ;
        RECT 2712.835 3429.375 2713.005 3429.545 ;
        RECT 2718.475 3429.375 2718.645 3429.545 ;
        RECT 2719.015 3429.375 2719.185 3429.545 ;
        RECT 2724.655 3429.375 2724.825 3429.545 ;
        RECT 2725.195 3429.375 2725.365 3429.545 ;
        RECT 2730.835 3429.375 2731.005 3429.545 ;
        RECT 2731.375 3429.375 2731.545 3429.545 ;
        RECT 2737.015 3429.375 2737.185 3429.545 ;
        RECT 2737.555 3429.375 2737.725 3429.545 ;
        RECT 2743.195 3429.375 2743.365 3429.545 ;
        RECT 2743.735 3429.375 2743.905 3429.545 ;
        RECT 2749.375 3429.375 2749.545 3429.545 ;
        RECT 2749.915 3429.375 2750.085 3429.545 ;
        RECT 2755.555 3429.375 2755.725 3429.545 ;
        RECT 2756.095 3429.375 2756.265 3429.545 ;
        RECT 2761.735 3429.375 2761.905 3429.545 ;
        RECT 2700.475 3426.675 2700.645 3426.845 ;
        RECT 2706.115 3426.675 2706.285 3426.845 ;
        RECT 2706.655 3426.675 2706.825 3426.845 ;
        RECT 2712.295 3426.675 2712.465 3426.845 ;
        RECT 2712.835 3426.675 2713.005 3426.845 ;
        RECT 2718.475 3426.675 2718.645 3426.845 ;
        RECT 2719.015 3426.675 2719.185 3426.845 ;
        RECT 2724.655 3426.675 2724.825 3426.845 ;
        RECT 2725.195 3426.675 2725.365 3426.845 ;
        RECT 2730.835 3426.675 2731.005 3426.845 ;
        RECT 2731.375 3426.675 2731.545 3426.845 ;
        RECT 2737.015 3426.675 2737.185 3426.845 ;
        RECT 2737.555 3426.675 2737.725 3426.845 ;
        RECT 2743.195 3426.675 2743.365 3426.845 ;
        RECT 2743.735 3426.675 2743.905 3426.845 ;
        RECT 2749.375 3426.675 2749.545 3426.845 ;
        RECT 2749.915 3426.675 2750.085 3426.845 ;
        RECT 2755.555 3426.675 2755.725 3426.845 ;
        RECT 2756.095 3426.675 2756.265 3426.845 ;
        RECT 2761.735 3426.675 2761.905 3426.845 ;
        RECT 2767.245 3424.875 2769.215 3430.445 ;
        RECT 2779.400 3424.875 2781.370 3430.445 ;
        RECT 2710.610 3423.170 2710.780 3423.340 ;
        RECT 2710.970 3423.170 2711.140 3423.340 ;
        RECT 2711.330 3423.170 2711.500 3423.340 ;
        RECT 2711.690 3423.170 2711.860 3423.340 ;
        RECT 2712.050 3423.170 2712.220 3423.340 ;
        RECT 2712.410 3423.170 2712.580 3423.340 ;
        RECT 2712.770 3423.170 2712.940 3423.340 ;
        RECT 2713.130 3423.170 2713.300 3423.340 ;
        RECT 2713.490 3423.170 2713.660 3423.340 ;
        RECT 2713.850 3423.170 2714.020 3423.340 ;
        RECT 2714.210 3423.170 2714.380 3423.340 ;
        RECT 2714.570 3423.170 2714.740 3423.340 ;
        RECT 2714.930 3423.170 2715.100 3423.340 ;
        RECT 2715.290 3423.170 2715.460 3423.340 ;
        RECT 2716.700 3423.170 2716.870 3423.340 ;
        RECT 2717.060 3423.170 2717.230 3423.340 ;
        RECT 2717.420 3423.170 2717.590 3423.340 ;
        RECT 2717.780 3423.170 2717.950 3423.340 ;
        RECT 2718.140 3423.170 2718.310 3423.340 ;
        RECT 2718.500 3423.170 2718.670 3423.340 ;
        RECT 2718.860 3423.170 2719.030 3423.340 ;
        RECT 2719.220 3423.170 2719.390 3423.340 ;
        RECT 2719.580 3423.170 2719.750 3423.340 ;
        RECT 2719.940 3423.170 2720.110 3423.340 ;
        RECT 2720.300 3423.170 2720.470 3423.340 ;
        RECT 2720.660 3423.170 2720.830 3423.340 ;
        RECT 2721.020 3423.170 2721.190 3423.340 ;
        RECT 2721.380 3423.170 2721.550 3423.340 ;
        RECT 2722.790 3423.170 2722.960 3423.340 ;
        RECT 2723.150 3423.170 2723.320 3423.340 ;
        RECT 2723.510 3423.170 2723.680 3423.340 ;
        RECT 2723.870 3423.170 2724.040 3423.340 ;
        RECT 2724.230 3423.170 2724.400 3423.340 ;
        RECT 2724.590 3423.170 2724.760 3423.340 ;
        RECT 2724.950 3423.170 2725.120 3423.340 ;
        RECT 2725.310 3423.170 2725.480 3423.340 ;
        RECT 2725.670 3423.170 2725.840 3423.340 ;
        RECT 2726.030 3423.170 2726.200 3423.340 ;
        RECT 2726.390 3423.170 2726.560 3423.340 ;
        RECT 2726.750 3423.170 2726.920 3423.340 ;
        RECT 2727.110 3423.170 2727.280 3423.340 ;
        RECT 2727.470 3423.170 2727.640 3423.340 ;
        RECT 2728.880 3423.170 2729.050 3423.340 ;
        RECT 2729.240 3423.170 2729.410 3423.340 ;
        RECT 2729.600 3423.170 2729.770 3423.340 ;
        RECT 2729.960 3423.170 2730.130 3423.340 ;
        RECT 2730.320 3423.170 2730.490 3423.340 ;
        RECT 2730.680 3423.170 2730.850 3423.340 ;
        RECT 2731.040 3423.170 2731.210 3423.340 ;
        RECT 2731.400 3423.170 2731.570 3423.340 ;
        RECT 2731.760 3423.170 2731.930 3423.340 ;
        RECT 2732.120 3423.170 2732.290 3423.340 ;
        RECT 2732.480 3423.170 2732.650 3423.340 ;
        RECT 2732.840 3423.170 2733.010 3423.340 ;
        RECT 2733.200 3423.170 2733.370 3423.340 ;
        RECT 2733.560 3423.170 2733.730 3423.340 ;
        RECT 2734.970 3423.170 2735.140 3423.340 ;
        RECT 2735.330 3423.170 2735.500 3423.340 ;
        RECT 2735.690 3423.170 2735.860 3423.340 ;
        RECT 2736.050 3423.170 2736.220 3423.340 ;
        RECT 2736.410 3423.170 2736.580 3423.340 ;
        RECT 2736.770 3423.170 2736.940 3423.340 ;
        RECT 2737.130 3423.170 2737.300 3423.340 ;
        RECT 2737.490 3423.170 2737.660 3423.340 ;
        RECT 2737.850 3423.170 2738.020 3423.340 ;
        RECT 2738.210 3423.170 2738.380 3423.340 ;
        RECT 2738.570 3423.170 2738.740 3423.340 ;
        RECT 2738.930 3423.170 2739.100 3423.340 ;
        RECT 2739.290 3423.170 2739.460 3423.340 ;
        RECT 2739.650 3423.170 2739.820 3423.340 ;
        RECT 2741.060 3423.170 2741.230 3423.340 ;
        RECT 2741.420 3423.170 2741.590 3423.340 ;
        RECT 2741.780 3423.170 2741.950 3423.340 ;
        RECT 2742.140 3423.170 2742.310 3423.340 ;
        RECT 2742.500 3423.170 2742.670 3423.340 ;
        RECT 2742.860 3423.170 2743.030 3423.340 ;
        RECT 2743.220 3423.170 2743.390 3423.340 ;
        RECT 2743.580 3423.170 2743.750 3423.340 ;
        RECT 2743.940 3423.170 2744.110 3423.340 ;
        RECT 2744.300 3423.170 2744.470 3423.340 ;
        RECT 2744.660 3423.170 2744.830 3423.340 ;
        RECT 2745.020 3423.170 2745.190 3423.340 ;
        RECT 2745.380 3423.170 2745.550 3423.340 ;
        RECT 2745.740 3423.170 2745.910 3423.340 ;
        RECT 2747.150 3423.170 2747.320 3423.340 ;
        RECT 2747.510 3423.170 2747.680 3423.340 ;
        RECT 2747.870 3423.170 2748.040 3423.340 ;
        RECT 2748.230 3423.170 2748.400 3423.340 ;
        RECT 2748.590 3423.170 2748.760 3423.340 ;
        RECT 2748.950 3423.170 2749.120 3423.340 ;
        RECT 2749.310 3423.170 2749.480 3423.340 ;
        RECT 2749.670 3423.170 2749.840 3423.340 ;
        RECT 2750.030 3423.170 2750.200 3423.340 ;
        RECT 2750.390 3423.170 2750.560 3423.340 ;
        RECT 2750.750 3423.170 2750.920 3423.340 ;
        RECT 2751.110 3423.170 2751.280 3423.340 ;
        RECT 2751.470 3423.170 2751.640 3423.340 ;
        RECT 2751.830 3423.170 2752.000 3423.340 ;
        RECT 2710.610 3422.380 2710.780 3422.550 ;
        RECT 2710.970 3422.380 2711.140 3422.550 ;
        RECT 2711.330 3422.380 2711.500 3422.550 ;
        RECT 2711.690 3422.380 2711.860 3422.550 ;
        RECT 2712.050 3422.380 2712.220 3422.550 ;
        RECT 2712.410 3422.380 2712.580 3422.550 ;
        RECT 2712.770 3422.380 2712.940 3422.550 ;
        RECT 2713.130 3422.380 2713.300 3422.550 ;
        RECT 2713.490 3422.380 2713.660 3422.550 ;
        RECT 2713.850 3422.380 2714.020 3422.550 ;
        RECT 2714.210 3422.380 2714.380 3422.550 ;
        RECT 2714.570 3422.380 2714.740 3422.550 ;
        RECT 2714.930 3422.380 2715.100 3422.550 ;
        RECT 2715.290 3422.380 2715.460 3422.550 ;
        RECT 2716.700 3422.380 2716.870 3422.550 ;
        RECT 2717.060 3422.380 2717.230 3422.550 ;
        RECT 2717.420 3422.380 2717.590 3422.550 ;
        RECT 2717.780 3422.380 2717.950 3422.550 ;
        RECT 2718.140 3422.380 2718.310 3422.550 ;
        RECT 2718.500 3422.380 2718.670 3422.550 ;
        RECT 2718.860 3422.380 2719.030 3422.550 ;
        RECT 2719.220 3422.380 2719.390 3422.550 ;
        RECT 2719.580 3422.380 2719.750 3422.550 ;
        RECT 2719.940 3422.380 2720.110 3422.550 ;
        RECT 2720.300 3422.380 2720.470 3422.550 ;
        RECT 2720.660 3422.380 2720.830 3422.550 ;
        RECT 2721.020 3422.380 2721.190 3422.550 ;
        RECT 2721.380 3422.380 2721.550 3422.550 ;
        RECT 2722.790 3422.380 2722.960 3422.550 ;
        RECT 2723.150 3422.380 2723.320 3422.550 ;
        RECT 2723.510 3422.380 2723.680 3422.550 ;
        RECT 2723.870 3422.380 2724.040 3422.550 ;
        RECT 2724.230 3422.380 2724.400 3422.550 ;
        RECT 2724.590 3422.380 2724.760 3422.550 ;
        RECT 2724.950 3422.380 2725.120 3422.550 ;
        RECT 2725.310 3422.380 2725.480 3422.550 ;
        RECT 2725.670 3422.380 2725.840 3422.550 ;
        RECT 2726.030 3422.380 2726.200 3422.550 ;
        RECT 2726.390 3422.380 2726.560 3422.550 ;
        RECT 2726.750 3422.380 2726.920 3422.550 ;
        RECT 2727.110 3422.380 2727.280 3422.550 ;
        RECT 2727.470 3422.380 2727.640 3422.550 ;
        RECT 2728.880 3422.380 2729.050 3422.550 ;
        RECT 2729.240 3422.380 2729.410 3422.550 ;
        RECT 2729.600 3422.380 2729.770 3422.550 ;
        RECT 2729.960 3422.380 2730.130 3422.550 ;
        RECT 2730.320 3422.380 2730.490 3422.550 ;
        RECT 2730.680 3422.380 2730.850 3422.550 ;
        RECT 2731.040 3422.380 2731.210 3422.550 ;
        RECT 2731.400 3422.380 2731.570 3422.550 ;
        RECT 2731.760 3422.380 2731.930 3422.550 ;
        RECT 2732.120 3422.380 2732.290 3422.550 ;
        RECT 2732.480 3422.380 2732.650 3422.550 ;
        RECT 2732.840 3422.380 2733.010 3422.550 ;
        RECT 2733.200 3422.380 2733.370 3422.550 ;
        RECT 2733.560 3422.380 2733.730 3422.550 ;
        RECT 2734.970 3422.380 2735.140 3422.550 ;
        RECT 2735.330 3422.380 2735.500 3422.550 ;
        RECT 2735.690 3422.380 2735.860 3422.550 ;
        RECT 2736.050 3422.380 2736.220 3422.550 ;
        RECT 2736.410 3422.380 2736.580 3422.550 ;
        RECT 2736.770 3422.380 2736.940 3422.550 ;
        RECT 2737.130 3422.380 2737.300 3422.550 ;
        RECT 2737.490 3422.380 2737.660 3422.550 ;
        RECT 2737.850 3422.380 2738.020 3422.550 ;
        RECT 2738.210 3422.380 2738.380 3422.550 ;
        RECT 2738.570 3422.380 2738.740 3422.550 ;
        RECT 2738.930 3422.380 2739.100 3422.550 ;
        RECT 2739.290 3422.380 2739.460 3422.550 ;
        RECT 2739.650 3422.380 2739.820 3422.550 ;
        RECT 2741.060 3422.380 2741.230 3422.550 ;
        RECT 2741.420 3422.380 2741.590 3422.550 ;
        RECT 2741.780 3422.380 2741.950 3422.550 ;
        RECT 2742.140 3422.380 2742.310 3422.550 ;
        RECT 2742.500 3422.380 2742.670 3422.550 ;
        RECT 2742.860 3422.380 2743.030 3422.550 ;
        RECT 2743.220 3422.380 2743.390 3422.550 ;
        RECT 2743.580 3422.380 2743.750 3422.550 ;
        RECT 2743.940 3422.380 2744.110 3422.550 ;
        RECT 2744.300 3422.380 2744.470 3422.550 ;
        RECT 2744.660 3422.380 2744.830 3422.550 ;
        RECT 2745.020 3422.380 2745.190 3422.550 ;
        RECT 2745.380 3422.380 2745.550 3422.550 ;
        RECT 2745.740 3422.380 2745.910 3422.550 ;
        RECT 2747.150 3422.380 2747.320 3422.550 ;
        RECT 2747.510 3422.380 2747.680 3422.550 ;
        RECT 2747.870 3422.380 2748.040 3422.550 ;
        RECT 2748.230 3422.380 2748.400 3422.550 ;
        RECT 2748.590 3422.380 2748.760 3422.550 ;
        RECT 2748.950 3422.380 2749.120 3422.550 ;
        RECT 2749.310 3422.380 2749.480 3422.550 ;
        RECT 2749.670 3422.380 2749.840 3422.550 ;
        RECT 2750.030 3422.380 2750.200 3422.550 ;
        RECT 2750.390 3422.380 2750.560 3422.550 ;
        RECT 2750.750 3422.380 2750.920 3422.550 ;
        RECT 2751.110 3422.380 2751.280 3422.550 ;
        RECT 2751.470 3422.380 2751.640 3422.550 ;
        RECT 2751.830 3422.380 2752.000 3422.550 ;
        RECT 2710.610 3420.670 2710.780 3420.840 ;
        RECT 2710.970 3420.670 2711.140 3420.840 ;
        RECT 2711.330 3420.670 2711.500 3420.840 ;
        RECT 2711.690 3420.670 2711.860 3420.840 ;
        RECT 2712.050 3420.670 2712.220 3420.840 ;
        RECT 2712.410 3420.670 2712.580 3420.840 ;
        RECT 2712.770 3420.670 2712.940 3420.840 ;
        RECT 2713.130 3420.670 2713.300 3420.840 ;
        RECT 2713.490 3420.670 2713.660 3420.840 ;
        RECT 2713.850 3420.670 2714.020 3420.840 ;
        RECT 2714.210 3420.670 2714.380 3420.840 ;
        RECT 2714.570 3420.670 2714.740 3420.840 ;
        RECT 2714.930 3420.670 2715.100 3420.840 ;
        RECT 2715.290 3420.670 2715.460 3420.840 ;
        RECT 2716.700 3420.670 2716.870 3420.840 ;
        RECT 2717.060 3420.670 2717.230 3420.840 ;
        RECT 2717.420 3420.670 2717.590 3420.840 ;
        RECT 2717.780 3420.670 2717.950 3420.840 ;
        RECT 2718.140 3420.670 2718.310 3420.840 ;
        RECT 2718.500 3420.670 2718.670 3420.840 ;
        RECT 2718.860 3420.670 2719.030 3420.840 ;
        RECT 2719.220 3420.670 2719.390 3420.840 ;
        RECT 2719.580 3420.670 2719.750 3420.840 ;
        RECT 2719.940 3420.670 2720.110 3420.840 ;
        RECT 2720.300 3420.670 2720.470 3420.840 ;
        RECT 2720.660 3420.670 2720.830 3420.840 ;
        RECT 2721.020 3420.670 2721.190 3420.840 ;
        RECT 2721.380 3420.670 2721.550 3420.840 ;
        RECT 2722.790 3420.670 2722.960 3420.840 ;
        RECT 2723.150 3420.670 2723.320 3420.840 ;
        RECT 2723.510 3420.670 2723.680 3420.840 ;
        RECT 2723.870 3420.670 2724.040 3420.840 ;
        RECT 2724.230 3420.670 2724.400 3420.840 ;
        RECT 2724.590 3420.670 2724.760 3420.840 ;
        RECT 2724.950 3420.670 2725.120 3420.840 ;
        RECT 2725.310 3420.670 2725.480 3420.840 ;
        RECT 2725.670 3420.670 2725.840 3420.840 ;
        RECT 2726.030 3420.670 2726.200 3420.840 ;
        RECT 2726.390 3420.670 2726.560 3420.840 ;
        RECT 2726.750 3420.670 2726.920 3420.840 ;
        RECT 2727.110 3420.670 2727.280 3420.840 ;
        RECT 2727.470 3420.670 2727.640 3420.840 ;
        RECT 2728.880 3420.670 2729.050 3420.840 ;
        RECT 2729.240 3420.670 2729.410 3420.840 ;
        RECT 2729.600 3420.670 2729.770 3420.840 ;
        RECT 2729.960 3420.670 2730.130 3420.840 ;
        RECT 2730.320 3420.670 2730.490 3420.840 ;
        RECT 2730.680 3420.670 2730.850 3420.840 ;
        RECT 2731.040 3420.670 2731.210 3420.840 ;
        RECT 2731.400 3420.670 2731.570 3420.840 ;
        RECT 2731.760 3420.670 2731.930 3420.840 ;
        RECT 2732.120 3420.670 2732.290 3420.840 ;
        RECT 2732.480 3420.670 2732.650 3420.840 ;
        RECT 2732.840 3420.670 2733.010 3420.840 ;
        RECT 2733.200 3420.670 2733.370 3420.840 ;
        RECT 2733.560 3420.670 2733.730 3420.840 ;
        RECT 2734.970 3420.670 2735.140 3420.840 ;
        RECT 2735.330 3420.670 2735.500 3420.840 ;
        RECT 2735.690 3420.670 2735.860 3420.840 ;
        RECT 2736.050 3420.670 2736.220 3420.840 ;
        RECT 2736.410 3420.670 2736.580 3420.840 ;
        RECT 2736.770 3420.670 2736.940 3420.840 ;
        RECT 2737.130 3420.670 2737.300 3420.840 ;
        RECT 2737.490 3420.670 2737.660 3420.840 ;
        RECT 2737.850 3420.670 2738.020 3420.840 ;
        RECT 2738.210 3420.670 2738.380 3420.840 ;
        RECT 2738.570 3420.670 2738.740 3420.840 ;
        RECT 2738.930 3420.670 2739.100 3420.840 ;
        RECT 2739.290 3420.670 2739.460 3420.840 ;
        RECT 2739.650 3420.670 2739.820 3420.840 ;
        RECT 2741.060 3420.670 2741.230 3420.840 ;
        RECT 2741.420 3420.670 2741.590 3420.840 ;
        RECT 2741.780 3420.670 2741.950 3420.840 ;
        RECT 2742.140 3420.670 2742.310 3420.840 ;
        RECT 2742.500 3420.670 2742.670 3420.840 ;
        RECT 2742.860 3420.670 2743.030 3420.840 ;
        RECT 2743.220 3420.670 2743.390 3420.840 ;
        RECT 2743.580 3420.670 2743.750 3420.840 ;
        RECT 2743.940 3420.670 2744.110 3420.840 ;
        RECT 2744.300 3420.670 2744.470 3420.840 ;
        RECT 2744.660 3420.670 2744.830 3420.840 ;
        RECT 2745.020 3420.670 2745.190 3420.840 ;
        RECT 2745.380 3420.670 2745.550 3420.840 ;
        RECT 2745.740 3420.670 2745.910 3420.840 ;
        RECT 2747.150 3420.670 2747.320 3420.840 ;
        RECT 2747.510 3420.670 2747.680 3420.840 ;
        RECT 2747.870 3420.670 2748.040 3420.840 ;
        RECT 2748.230 3420.670 2748.400 3420.840 ;
        RECT 2748.590 3420.670 2748.760 3420.840 ;
        RECT 2748.950 3420.670 2749.120 3420.840 ;
        RECT 2749.310 3420.670 2749.480 3420.840 ;
        RECT 2749.670 3420.670 2749.840 3420.840 ;
        RECT 2750.030 3420.670 2750.200 3420.840 ;
        RECT 2750.390 3420.670 2750.560 3420.840 ;
        RECT 2750.750 3420.670 2750.920 3420.840 ;
        RECT 2751.110 3420.670 2751.280 3420.840 ;
        RECT 2751.470 3420.670 2751.640 3420.840 ;
        RECT 2751.830 3420.670 2752.000 3420.840 ;
        RECT 2710.610 3419.880 2710.780 3420.050 ;
        RECT 2710.970 3419.880 2711.140 3420.050 ;
        RECT 2711.330 3419.880 2711.500 3420.050 ;
        RECT 2711.690 3419.880 2711.860 3420.050 ;
        RECT 2712.050 3419.880 2712.220 3420.050 ;
        RECT 2712.410 3419.880 2712.580 3420.050 ;
        RECT 2712.770 3419.880 2712.940 3420.050 ;
        RECT 2713.130 3419.880 2713.300 3420.050 ;
        RECT 2713.490 3419.880 2713.660 3420.050 ;
        RECT 2713.850 3419.880 2714.020 3420.050 ;
        RECT 2714.210 3419.880 2714.380 3420.050 ;
        RECT 2714.570 3419.880 2714.740 3420.050 ;
        RECT 2714.930 3419.880 2715.100 3420.050 ;
        RECT 2715.290 3419.880 2715.460 3420.050 ;
        RECT 2716.700 3419.880 2716.870 3420.050 ;
        RECT 2717.060 3419.880 2717.230 3420.050 ;
        RECT 2717.420 3419.880 2717.590 3420.050 ;
        RECT 2717.780 3419.880 2717.950 3420.050 ;
        RECT 2718.140 3419.880 2718.310 3420.050 ;
        RECT 2718.500 3419.880 2718.670 3420.050 ;
        RECT 2718.860 3419.880 2719.030 3420.050 ;
        RECT 2719.220 3419.880 2719.390 3420.050 ;
        RECT 2719.580 3419.880 2719.750 3420.050 ;
        RECT 2719.940 3419.880 2720.110 3420.050 ;
        RECT 2720.300 3419.880 2720.470 3420.050 ;
        RECT 2720.660 3419.880 2720.830 3420.050 ;
        RECT 2721.020 3419.880 2721.190 3420.050 ;
        RECT 2721.380 3419.880 2721.550 3420.050 ;
        RECT 2722.790 3419.880 2722.960 3420.050 ;
        RECT 2723.150 3419.880 2723.320 3420.050 ;
        RECT 2723.510 3419.880 2723.680 3420.050 ;
        RECT 2723.870 3419.880 2724.040 3420.050 ;
        RECT 2724.230 3419.880 2724.400 3420.050 ;
        RECT 2724.590 3419.880 2724.760 3420.050 ;
        RECT 2724.950 3419.880 2725.120 3420.050 ;
        RECT 2725.310 3419.880 2725.480 3420.050 ;
        RECT 2725.670 3419.880 2725.840 3420.050 ;
        RECT 2726.030 3419.880 2726.200 3420.050 ;
        RECT 2726.390 3419.880 2726.560 3420.050 ;
        RECT 2726.750 3419.880 2726.920 3420.050 ;
        RECT 2727.110 3419.880 2727.280 3420.050 ;
        RECT 2727.470 3419.880 2727.640 3420.050 ;
        RECT 2728.880 3419.880 2729.050 3420.050 ;
        RECT 2729.240 3419.880 2729.410 3420.050 ;
        RECT 2729.600 3419.880 2729.770 3420.050 ;
        RECT 2729.960 3419.880 2730.130 3420.050 ;
        RECT 2730.320 3419.880 2730.490 3420.050 ;
        RECT 2730.680 3419.880 2730.850 3420.050 ;
        RECT 2731.040 3419.880 2731.210 3420.050 ;
        RECT 2731.400 3419.880 2731.570 3420.050 ;
        RECT 2731.760 3419.880 2731.930 3420.050 ;
        RECT 2732.120 3419.880 2732.290 3420.050 ;
        RECT 2732.480 3419.880 2732.650 3420.050 ;
        RECT 2732.840 3419.880 2733.010 3420.050 ;
        RECT 2733.200 3419.880 2733.370 3420.050 ;
        RECT 2733.560 3419.880 2733.730 3420.050 ;
        RECT 2734.970 3419.880 2735.140 3420.050 ;
        RECT 2735.330 3419.880 2735.500 3420.050 ;
        RECT 2735.690 3419.880 2735.860 3420.050 ;
        RECT 2736.050 3419.880 2736.220 3420.050 ;
        RECT 2736.410 3419.880 2736.580 3420.050 ;
        RECT 2736.770 3419.880 2736.940 3420.050 ;
        RECT 2737.130 3419.880 2737.300 3420.050 ;
        RECT 2737.490 3419.880 2737.660 3420.050 ;
        RECT 2737.850 3419.880 2738.020 3420.050 ;
        RECT 2738.210 3419.880 2738.380 3420.050 ;
        RECT 2738.570 3419.880 2738.740 3420.050 ;
        RECT 2738.930 3419.880 2739.100 3420.050 ;
        RECT 2739.290 3419.880 2739.460 3420.050 ;
        RECT 2739.650 3419.880 2739.820 3420.050 ;
        RECT 2741.060 3419.880 2741.230 3420.050 ;
        RECT 2741.420 3419.880 2741.590 3420.050 ;
        RECT 2741.780 3419.880 2741.950 3420.050 ;
        RECT 2742.140 3419.880 2742.310 3420.050 ;
        RECT 2742.500 3419.880 2742.670 3420.050 ;
        RECT 2742.860 3419.880 2743.030 3420.050 ;
        RECT 2743.220 3419.880 2743.390 3420.050 ;
        RECT 2743.580 3419.880 2743.750 3420.050 ;
        RECT 2743.940 3419.880 2744.110 3420.050 ;
        RECT 2744.300 3419.880 2744.470 3420.050 ;
        RECT 2744.660 3419.880 2744.830 3420.050 ;
        RECT 2745.020 3419.880 2745.190 3420.050 ;
        RECT 2745.380 3419.880 2745.550 3420.050 ;
        RECT 2745.740 3419.880 2745.910 3420.050 ;
        RECT 2747.150 3419.880 2747.320 3420.050 ;
        RECT 2747.510 3419.880 2747.680 3420.050 ;
        RECT 2747.870 3419.880 2748.040 3420.050 ;
        RECT 2748.230 3419.880 2748.400 3420.050 ;
        RECT 2748.590 3419.880 2748.760 3420.050 ;
        RECT 2748.950 3419.880 2749.120 3420.050 ;
        RECT 2749.310 3419.880 2749.480 3420.050 ;
        RECT 2749.670 3419.880 2749.840 3420.050 ;
        RECT 2750.030 3419.880 2750.200 3420.050 ;
        RECT 2750.390 3419.880 2750.560 3420.050 ;
        RECT 2750.750 3419.880 2750.920 3420.050 ;
        RECT 2751.110 3419.880 2751.280 3420.050 ;
        RECT 2751.470 3419.880 2751.640 3420.050 ;
        RECT 2751.830 3419.880 2752.000 3420.050 ;
        RECT 2712.975 3417.705 2713.145 3417.875 ;
        RECT 2712.975 3417.345 2713.145 3417.515 ;
        RECT 2718.525 3417.705 2718.695 3417.875 ;
        RECT 2718.525 3417.345 2718.695 3417.515 ;
        RECT 2719.065 3417.705 2719.235 3417.875 ;
        RECT 2719.065 3417.345 2719.235 3417.515 ;
        RECT 2724.615 3417.705 2724.785 3417.875 ;
        RECT 2724.615 3417.345 2724.785 3417.515 ;
        RECT 2725.155 3417.705 2725.325 3417.875 ;
        RECT 2725.155 3417.345 2725.325 3417.515 ;
        RECT 2730.705 3417.705 2730.875 3417.875 ;
        RECT 2730.705 3417.345 2730.875 3417.515 ;
        RECT 2731.245 3417.705 2731.415 3417.875 ;
        RECT 2731.245 3417.345 2731.415 3417.515 ;
        RECT 2736.795 3417.705 2736.965 3417.875 ;
        RECT 2736.795 3417.345 2736.965 3417.515 ;
        RECT 2737.335 3417.705 2737.505 3417.875 ;
        RECT 2737.335 3417.345 2737.505 3417.515 ;
        RECT 2742.885 3417.705 2743.055 3417.875 ;
        RECT 2742.885 3417.345 2743.055 3417.515 ;
        RECT 2743.425 3417.705 2743.595 3417.875 ;
        RECT 2743.425 3417.345 2743.595 3417.515 ;
        RECT 2748.975 3417.705 2749.145 3417.875 ;
        RECT 2748.975 3417.345 2749.145 3417.515 ;
        RECT 2712.975 3414.605 2713.145 3414.775 ;
        RECT 2712.975 3414.245 2713.145 3414.415 ;
        RECT 2718.525 3414.605 2718.695 3414.775 ;
        RECT 2718.525 3414.245 2718.695 3414.415 ;
        RECT 2719.065 3414.605 2719.235 3414.775 ;
        RECT 2719.065 3414.245 2719.235 3414.415 ;
        RECT 2724.615 3414.605 2724.785 3414.775 ;
        RECT 2724.615 3414.245 2724.785 3414.415 ;
        RECT 2725.155 3414.605 2725.325 3414.775 ;
        RECT 2725.155 3414.245 2725.325 3414.415 ;
        RECT 2730.705 3414.605 2730.875 3414.775 ;
        RECT 2730.705 3414.245 2730.875 3414.415 ;
        RECT 2731.245 3414.605 2731.415 3414.775 ;
        RECT 2731.245 3414.245 2731.415 3414.415 ;
        RECT 2736.795 3414.605 2736.965 3414.775 ;
        RECT 2736.795 3414.245 2736.965 3414.415 ;
        RECT 2737.335 3414.605 2737.505 3414.775 ;
        RECT 2737.335 3414.245 2737.505 3414.415 ;
        RECT 2742.885 3414.605 2743.055 3414.775 ;
        RECT 2742.885 3414.245 2743.055 3414.415 ;
        RECT 2743.425 3414.605 2743.595 3414.775 ;
        RECT 2743.425 3414.245 2743.595 3414.415 ;
        RECT 2748.975 3414.605 2749.145 3414.775 ;
        RECT 2748.975 3414.245 2749.145 3414.415 ;
        RECT 2710.175 3411.605 2710.345 3411.775 ;
        RECT 2710.175 3411.245 2710.345 3411.415 ;
        RECT 2715.725 3411.605 2715.895 3411.775 ;
        RECT 2715.725 3411.245 2715.895 3411.415 ;
        RECT 2716.265 3411.605 2716.435 3411.775 ;
        RECT 2716.265 3411.245 2716.435 3411.415 ;
        RECT 2721.815 3411.605 2721.985 3411.775 ;
        RECT 2721.815 3411.245 2721.985 3411.415 ;
        RECT 2722.355 3411.605 2722.525 3411.775 ;
        RECT 2722.355 3411.245 2722.525 3411.415 ;
        RECT 2727.905 3411.605 2728.075 3411.775 ;
        RECT 2727.905 3411.245 2728.075 3411.415 ;
        RECT 2728.445 3411.605 2728.615 3411.775 ;
        RECT 2728.445 3411.245 2728.615 3411.415 ;
        RECT 2733.995 3411.605 2734.165 3411.775 ;
        RECT 2733.995 3411.245 2734.165 3411.415 ;
        RECT 2734.535 3411.605 2734.705 3411.775 ;
        RECT 2734.535 3411.245 2734.705 3411.415 ;
        RECT 2740.085 3411.605 2740.255 3411.775 ;
        RECT 2740.085 3411.245 2740.255 3411.415 ;
        RECT 2740.625 3411.605 2740.795 3411.775 ;
        RECT 2740.625 3411.245 2740.795 3411.415 ;
        RECT 2746.175 3411.605 2746.345 3411.775 ;
        RECT 2746.175 3411.245 2746.345 3411.415 ;
        RECT 2746.715 3411.605 2746.885 3411.775 ;
        RECT 2746.715 3411.245 2746.885 3411.415 ;
        RECT 2752.265 3411.605 2752.435 3411.775 ;
        RECT 2752.265 3411.245 2752.435 3411.415 ;
        RECT 2710.610 3410.780 2710.780 3410.950 ;
        RECT 2710.970 3410.780 2711.140 3410.950 ;
        RECT 2711.330 3410.780 2711.500 3410.950 ;
        RECT 2711.690 3410.780 2711.860 3410.950 ;
        RECT 2712.050 3410.780 2712.220 3410.950 ;
        RECT 2712.410 3410.780 2712.580 3410.950 ;
        RECT 2712.770 3410.780 2712.940 3410.950 ;
        RECT 2713.130 3410.780 2713.300 3410.950 ;
        RECT 2713.490 3410.780 2713.660 3410.950 ;
        RECT 2713.850 3410.780 2714.020 3410.950 ;
        RECT 2714.210 3410.780 2714.380 3410.950 ;
        RECT 2714.570 3410.780 2714.740 3410.950 ;
        RECT 2714.930 3410.780 2715.100 3410.950 ;
        RECT 2715.290 3410.780 2715.460 3410.950 ;
        RECT 2716.700 3410.780 2716.870 3410.950 ;
        RECT 2717.060 3410.780 2717.230 3410.950 ;
        RECT 2717.420 3410.780 2717.590 3410.950 ;
        RECT 2717.780 3410.780 2717.950 3410.950 ;
        RECT 2718.140 3410.780 2718.310 3410.950 ;
        RECT 2718.500 3410.780 2718.670 3410.950 ;
        RECT 2718.860 3410.780 2719.030 3410.950 ;
        RECT 2719.220 3410.780 2719.390 3410.950 ;
        RECT 2719.580 3410.780 2719.750 3410.950 ;
        RECT 2719.940 3410.780 2720.110 3410.950 ;
        RECT 2720.300 3410.780 2720.470 3410.950 ;
        RECT 2720.660 3410.780 2720.830 3410.950 ;
        RECT 2721.020 3410.780 2721.190 3410.950 ;
        RECT 2721.380 3410.780 2721.550 3410.950 ;
        RECT 2722.790 3410.780 2722.960 3410.950 ;
        RECT 2723.150 3410.780 2723.320 3410.950 ;
        RECT 2723.510 3410.780 2723.680 3410.950 ;
        RECT 2723.870 3410.780 2724.040 3410.950 ;
        RECT 2724.230 3410.780 2724.400 3410.950 ;
        RECT 2724.590 3410.780 2724.760 3410.950 ;
        RECT 2724.950 3410.780 2725.120 3410.950 ;
        RECT 2725.310 3410.780 2725.480 3410.950 ;
        RECT 2725.670 3410.780 2725.840 3410.950 ;
        RECT 2726.030 3410.780 2726.200 3410.950 ;
        RECT 2726.390 3410.780 2726.560 3410.950 ;
        RECT 2726.750 3410.780 2726.920 3410.950 ;
        RECT 2727.110 3410.780 2727.280 3410.950 ;
        RECT 2727.470 3410.780 2727.640 3410.950 ;
        RECT 2728.880 3410.780 2729.050 3410.950 ;
        RECT 2729.240 3410.780 2729.410 3410.950 ;
        RECT 2729.600 3410.780 2729.770 3410.950 ;
        RECT 2729.960 3410.780 2730.130 3410.950 ;
        RECT 2730.320 3410.780 2730.490 3410.950 ;
        RECT 2730.680 3410.780 2730.850 3410.950 ;
        RECT 2731.040 3410.780 2731.210 3410.950 ;
        RECT 2731.400 3410.780 2731.570 3410.950 ;
        RECT 2731.760 3410.780 2731.930 3410.950 ;
        RECT 2732.120 3410.780 2732.290 3410.950 ;
        RECT 2732.480 3410.780 2732.650 3410.950 ;
        RECT 2732.840 3410.780 2733.010 3410.950 ;
        RECT 2733.200 3410.780 2733.370 3410.950 ;
        RECT 2733.560 3410.780 2733.730 3410.950 ;
        RECT 2734.970 3410.780 2735.140 3410.950 ;
        RECT 2735.330 3410.780 2735.500 3410.950 ;
        RECT 2735.690 3410.780 2735.860 3410.950 ;
        RECT 2736.050 3410.780 2736.220 3410.950 ;
        RECT 2736.410 3410.780 2736.580 3410.950 ;
        RECT 2736.770 3410.780 2736.940 3410.950 ;
        RECT 2737.130 3410.780 2737.300 3410.950 ;
        RECT 2737.490 3410.780 2737.660 3410.950 ;
        RECT 2737.850 3410.780 2738.020 3410.950 ;
        RECT 2738.210 3410.780 2738.380 3410.950 ;
        RECT 2738.570 3410.780 2738.740 3410.950 ;
        RECT 2738.930 3410.780 2739.100 3410.950 ;
        RECT 2739.290 3410.780 2739.460 3410.950 ;
        RECT 2739.650 3410.780 2739.820 3410.950 ;
        RECT 2741.060 3410.780 2741.230 3410.950 ;
        RECT 2741.420 3410.780 2741.590 3410.950 ;
        RECT 2741.780 3410.780 2741.950 3410.950 ;
        RECT 2742.140 3410.780 2742.310 3410.950 ;
        RECT 2742.500 3410.780 2742.670 3410.950 ;
        RECT 2742.860 3410.780 2743.030 3410.950 ;
        RECT 2743.220 3410.780 2743.390 3410.950 ;
        RECT 2743.580 3410.780 2743.750 3410.950 ;
        RECT 2743.940 3410.780 2744.110 3410.950 ;
        RECT 2744.300 3410.780 2744.470 3410.950 ;
        RECT 2744.660 3410.780 2744.830 3410.950 ;
        RECT 2745.020 3410.780 2745.190 3410.950 ;
        RECT 2745.380 3410.780 2745.550 3410.950 ;
        RECT 2745.740 3410.780 2745.910 3410.950 ;
        RECT 2747.150 3410.780 2747.320 3410.950 ;
        RECT 2747.510 3410.780 2747.680 3410.950 ;
        RECT 2747.870 3410.780 2748.040 3410.950 ;
        RECT 2748.230 3410.780 2748.400 3410.950 ;
        RECT 2748.590 3410.780 2748.760 3410.950 ;
        RECT 2748.950 3410.780 2749.120 3410.950 ;
        RECT 2749.310 3410.780 2749.480 3410.950 ;
        RECT 2749.670 3410.780 2749.840 3410.950 ;
        RECT 2750.030 3410.780 2750.200 3410.950 ;
        RECT 2750.390 3410.780 2750.560 3410.950 ;
        RECT 2750.750 3410.780 2750.920 3410.950 ;
        RECT 2751.110 3410.780 2751.280 3410.950 ;
        RECT 2751.470 3410.780 2751.640 3410.950 ;
        RECT 2751.830 3410.780 2752.000 3410.950 ;
        RECT 2710.175 3408.605 2710.345 3408.775 ;
        RECT 2710.175 3408.245 2710.345 3408.415 ;
        RECT 2715.725 3408.605 2715.895 3408.775 ;
        RECT 2715.725 3408.245 2715.895 3408.415 ;
        RECT 2716.265 3408.605 2716.435 3408.775 ;
        RECT 2716.265 3408.245 2716.435 3408.415 ;
        RECT 2721.815 3408.605 2721.985 3408.775 ;
        RECT 2721.815 3408.245 2721.985 3408.415 ;
        RECT 2722.355 3408.605 2722.525 3408.775 ;
        RECT 2722.355 3408.245 2722.525 3408.415 ;
        RECT 2727.905 3408.605 2728.075 3408.775 ;
        RECT 2727.905 3408.245 2728.075 3408.415 ;
        RECT 2728.445 3408.605 2728.615 3408.775 ;
        RECT 2728.445 3408.245 2728.615 3408.415 ;
        RECT 2733.995 3408.605 2734.165 3408.775 ;
        RECT 2733.995 3408.245 2734.165 3408.415 ;
        RECT 2734.535 3408.605 2734.705 3408.775 ;
        RECT 2734.535 3408.245 2734.705 3408.415 ;
        RECT 2740.085 3408.605 2740.255 3408.775 ;
        RECT 2740.085 3408.245 2740.255 3408.415 ;
        RECT 2740.625 3408.605 2740.795 3408.775 ;
        RECT 2740.625 3408.245 2740.795 3408.415 ;
        RECT 2746.175 3408.605 2746.345 3408.775 ;
        RECT 2746.175 3408.245 2746.345 3408.415 ;
        RECT 2746.715 3408.605 2746.885 3408.775 ;
        RECT 2746.715 3408.245 2746.885 3408.415 ;
        RECT 2752.265 3408.605 2752.435 3408.775 ;
        RECT 2752.265 3408.245 2752.435 3408.415 ;
        RECT 2710.610 3407.780 2710.780 3407.950 ;
        RECT 2710.970 3407.780 2711.140 3407.950 ;
        RECT 2711.330 3407.780 2711.500 3407.950 ;
        RECT 2711.690 3407.780 2711.860 3407.950 ;
        RECT 2712.050 3407.780 2712.220 3407.950 ;
        RECT 2712.410 3407.780 2712.580 3407.950 ;
        RECT 2712.770 3407.780 2712.940 3407.950 ;
        RECT 2713.130 3407.780 2713.300 3407.950 ;
        RECT 2713.490 3407.780 2713.660 3407.950 ;
        RECT 2713.850 3407.780 2714.020 3407.950 ;
        RECT 2714.210 3407.780 2714.380 3407.950 ;
        RECT 2714.570 3407.780 2714.740 3407.950 ;
        RECT 2714.930 3407.780 2715.100 3407.950 ;
        RECT 2715.290 3407.780 2715.460 3407.950 ;
        RECT 2716.700 3407.780 2716.870 3407.950 ;
        RECT 2717.060 3407.780 2717.230 3407.950 ;
        RECT 2717.420 3407.780 2717.590 3407.950 ;
        RECT 2717.780 3407.780 2717.950 3407.950 ;
        RECT 2718.140 3407.780 2718.310 3407.950 ;
        RECT 2718.500 3407.780 2718.670 3407.950 ;
        RECT 2718.860 3407.780 2719.030 3407.950 ;
        RECT 2719.220 3407.780 2719.390 3407.950 ;
        RECT 2719.580 3407.780 2719.750 3407.950 ;
        RECT 2719.940 3407.780 2720.110 3407.950 ;
        RECT 2720.300 3407.780 2720.470 3407.950 ;
        RECT 2720.660 3407.780 2720.830 3407.950 ;
        RECT 2721.020 3407.780 2721.190 3407.950 ;
        RECT 2721.380 3407.780 2721.550 3407.950 ;
        RECT 2722.790 3407.780 2722.960 3407.950 ;
        RECT 2723.150 3407.780 2723.320 3407.950 ;
        RECT 2723.510 3407.780 2723.680 3407.950 ;
        RECT 2723.870 3407.780 2724.040 3407.950 ;
        RECT 2724.230 3407.780 2724.400 3407.950 ;
        RECT 2724.590 3407.780 2724.760 3407.950 ;
        RECT 2724.950 3407.780 2725.120 3407.950 ;
        RECT 2725.310 3407.780 2725.480 3407.950 ;
        RECT 2725.670 3407.780 2725.840 3407.950 ;
        RECT 2726.030 3407.780 2726.200 3407.950 ;
        RECT 2726.390 3407.780 2726.560 3407.950 ;
        RECT 2726.750 3407.780 2726.920 3407.950 ;
        RECT 2727.110 3407.780 2727.280 3407.950 ;
        RECT 2727.470 3407.780 2727.640 3407.950 ;
        RECT 2728.880 3407.780 2729.050 3407.950 ;
        RECT 2729.240 3407.780 2729.410 3407.950 ;
        RECT 2729.600 3407.780 2729.770 3407.950 ;
        RECT 2729.960 3407.780 2730.130 3407.950 ;
        RECT 2730.320 3407.780 2730.490 3407.950 ;
        RECT 2730.680 3407.780 2730.850 3407.950 ;
        RECT 2731.040 3407.780 2731.210 3407.950 ;
        RECT 2731.400 3407.780 2731.570 3407.950 ;
        RECT 2731.760 3407.780 2731.930 3407.950 ;
        RECT 2732.120 3407.780 2732.290 3407.950 ;
        RECT 2732.480 3407.780 2732.650 3407.950 ;
        RECT 2732.840 3407.780 2733.010 3407.950 ;
        RECT 2733.200 3407.780 2733.370 3407.950 ;
        RECT 2733.560 3407.780 2733.730 3407.950 ;
        RECT 2734.970 3407.780 2735.140 3407.950 ;
        RECT 2735.330 3407.780 2735.500 3407.950 ;
        RECT 2735.690 3407.780 2735.860 3407.950 ;
        RECT 2736.050 3407.780 2736.220 3407.950 ;
        RECT 2736.410 3407.780 2736.580 3407.950 ;
        RECT 2736.770 3407.780 2736.940 3407.950 ;
        RECT 2737.130 3407.780 2737.300 3407.950 ;
        RECT 2737.490 3407.780 2737.660 3407.950 ;
        RECT 2737.850 3407.780 2738.020 3407.950 ;
        RECT 2738.210 3407.780 2738.380 3407.950 ;
        RECT 2738.570 3407.780 2738.740 3407.950 ;
        RECT 2738.930 3407.780 2739.100 3407.950 ;
        RECT 2739.290 3407.780 2739.460 3407.950 ;
        RECT 2739.650 3407.780 2739.820 3407.950 ;
        RECT 2741.060 3407.780 2741.230 3407.950 ;
        RECT 2741.420 3407.780 2741.590 3407.950 ;
        RECT 2741.780 3407.780 2741.950 3407.950 ;
        RECT 2742.140 3407.780 2742.310 3407.950 ;
        RECT 2742.500 3407.780 2742.670 3407.950 ;
        RECT 2742.860 3407.780 2743.030 3407.950 ;
        RECT 2743.220 3407.780 2743.390 3407.950 ;
        RECT 2743.580 3407.780 2743.750 3407.950 ;
        RECT 2743.940 3407.780 2744.110 3407.950 ;
        RECT 2744.300 3407.780 2744.470 3407.950 ;
        RECT 2744.660 3407.780 2744.830 3407.950 ;
        RECT 2745.020 3407.780 2745.190 3407.950 ;
        RECT 2745.380 3407.780 2745.550 3407.950 ;
        RECT 2745.740 3407.780 2745.910 3407.950 ;
        RECT 2747.150 3407.780 2747.320 3407.950 ;
        RECT 2747.510 3407.780 2747.680 3407.950 ;
        RECT 2747.870 3407.780 2748.040 3407.950 ;
        RECT 2748.230 3407.780 2748.400 3407.950 ;
        RECT 2748.590 3407.780 2748.760 3407.950 ;
        RECT 2748.950 3407.780 2749.120 3407.950 ;
        RECT 2749.310 3407.780 2749.480 3407.950 ;
        RECT 2749.670 3407.780 2749.840 3407.950 ;
        RECT 2750.030 3407.780 2750.200 3407.950 ;
        RECT 2750.390 3407.780 2750.560 3407.950 ;
        RECT 2750.750 3407.780 2750.920 3407.950 ;
        RECT 2751.110 3407.780 2751.280 3407.950 ;
        RECT 2751.470 3407.780 2751.640 3407.950 ;
        RECT 2751.830 3407.780 2752.000 3407.950 ;
        RECT 2712.900 3403.735 2713.070 3403.905 ;
        RECT 2712.900 3403.375 2713.070 3403.545 ;
        RECT 2718.540 3403.735 2718.710 3403.905 ;
        RECT 2718.540 3403.375 2718.710 3403.545 ;
        RECT 2719.080 3403.735 2719.250 3403.905 ;
        RECT 2719.080 3403.375 2719.250 3403.545 ;
        RECT 2724.720 3403.735 2724.890 3403.905 ;
        RECT 2724.720 3403.375 2724.890 3403.545 ;
        RECT 2725.260 3403.735 2725.430 3403.905 ;
        RECT 2725.260 3403.375 2725.430 3403.545 ;
        RECT 2730.900 3403.735 2731.070 3403.905 ;
        RECT 2730.900 3403.375 2731.070 3403.545 ;
        RECT 2731.440 3403.735 2731.610 3403.905 ;
        RECT 2731.440 3403.375 2731.610 3403.545 ;
        RECT 2737.080 3403.735 2737.250 3403.905 ;
        RECT 2737.080 3403.375 2737.250 3403.545 ;
        RECT 2737.620 3403.735 2737.790 3403.905 ;
        RECT 2737.620 3403.375 2737.790 3403.545 ;
        RECT 2743.260 3403.735 2743.430 3403.905 ;
        RECT 2743.260 3403.375 2743.430 3403.545 ;
        RECT 2743.800 3403.735 2743.970 3403.905 ;
        RECT 2743.800 3403.375 2743.970 3403.545 ;
        RECT 2749.440 3403.735 2749.610 3403.905 ;
        RECT 2749.440 3403.375 2749.610 3403.545 ;
        RECT 2713.380 3402.910 2713.550 3403.080 ;
        RECT 2713.740 3402.910 2713.910 3403.080 ;
        RECT 2714.100 3402.910 2714.270 3403.080 ;
        RECT 2714.460 3402.910 2714.630 3403.080 ;
        RECT 2714.820 3402.910 2714.990 3403.080 ;
        RECT 2715.180 3402.910 2715.350 3403.080 ;
        RECT 2715.540 3402.910 2715.710 3403.080 ;
        RECT 2715.900 3402.910 2716.070 3403.080 ;
        RECT 2716.260 3402.910 2716.430 3403.080 ;
        RECT 2716.620 3402.910 2716.790 3403.080 ;
        RECT 2716.980 3402.910 2717.150 3403.080 ;
        RECT 2717.340 3402.910 2717.510 3403.080 ;
        RECT 2717.700 3402.910 2717.870 3403.080 ;
        RECT 2718.060 3402.910 2718.230 3403.080 ;
        RECT 2719.560 3402.910 2719.730 3403.080 ;
        RECT 2719.920 3402.910 2720.090 3403.080 ;
        RECT 2720.280 3402.910 2720.450 3403.080 ;
        RECT 2720.640 3402.910 2720.810 3403.080 ;
        RECT 2721.000 3402.910 2721.170 3403.080 ;
        RECT 2721.360 3402.910 2721.530 3403.080 ;
        RECT 2721.720 3402.910 2721.890 3403.080 ;
        RECT 2722.080 3402.910 2722.250 3403.080 ;
        RECT 2722.440 3402.910 2722.610 3403.080 ;
        RECT 2722.800 3402.910 2722.970 3403.080 ;
        RECT 2723.160 3402.910 2723.330 3403.080 ;
        RECT 2723.520 3402.910 2723.690 3403.080 ;
        RECT 2723.880 3402.910 2724.050 3403.080 ;
        RECT 2724.240 3402.910 2724.410 3403.080 ;
        RECT 2725.740 3402.910 2725.910 3403.080 ;
        RECT 2726.100 3402.910 2726.270 3403.080 ;
        RECT 2726.460 3402.910 2726.630 3403.080 ;
        RECT 2726.820 3402.910 2726.990 3403.080 ;
        RECT 2727.180 3402.910 2727.350 3403.080 ;
        RECT 2727.540 3402.910 2727.710 3403.080 ;
        RECT 2727.900 3402.910 2728.070 3403.080 ;
        RECT 2728.260 3402.910 2728.430 3403.080 ;
        RECT 2728.620 3402.910 2728.790 3403.080 ;
        RECT 2728.980 3402.910 2729.150 3403.080 ;
        RECT 2729.340 3402.910 2729.510 3403.080 ;
        RECT 2729.700 3402.910 2729.870 3403.080 ;
        RECT 2730.060 3402.910 2730.230 3403.080 ;
        RECT 2730.420 3402.910 2730.590 3403.080 ;
        RECT 2731.920 3402.910 2732.090 3403.080 ;
        RECT 2732.280 3402.910 2732.450 3403.080 ;
        RECT 2732.640 3402.910 2732.810 3403.080 ;
        RECT 2733.000 3402.910 2733.170 3403.080 ;
        RECT 2733.360 3402.910 2733.530 3403.080 ;
        RECT 2733.720 3402.910 2733.890 3403.080 ;
        RECT 2734.080 3402.910 2734.250 3403.080 ;
        RECT 2734.440 3402.910 2734.610 3403.080 ;
        RECT 2734.800 3402.910 2734.970 3403.080 ;
        RECT 2735.160 3402.910 2735.330 3403.080 ;
        RECT 2735.520 3402.910 2735.690 3403.080 ;
        RECT 2735.880 3402.910 2736.050 3403.080 ;
        RECT 2736.240 3402.910 2736.410 3403.080 ;
        RECT 2736.600 3402.910 2736.770 3403.080 ;
        RECT 2738.100 3402.910 2738.270 3403.080 ;
        RECT 2738.460 3402.910 2738.630 3403.080 ;
        RECT 2738.820 3402.910 2738.990 3403.080 ;
        RECT 2739.180 3402.910 2739.350 3403.080 ;
        RECT 2739.540 3402.910 2739.710 3403.080 ;
        RECT 2739.900 3402.910 2740.070 3403.080 ;
        RECT 2740.260 3402.910 2740.430 3403.080 ;
        RECT 2740.620 3402.910 2740.790 3403.080 ;
        RECT 2740.980 3402.910 2741.150 3403.080 ;
        RECT 2741.340 3402.910 2741.510 3403.080 ;
        RECT 2741.700 3402.910 2741.870 3403.080 ;
        RECT 2742.060 3402.910 2742.230 3403.080 ;
        RECT 2742.420 3402.910 2742.590 3403.080 ;
        RECT 2742.780 3402.910 2742.950 3403.080 ;
        RECT 2744.280 3402.910 2744.450 3403.080 ;
        RECT 2744.640 3402.910 2744.810 3403.080 ;
        RECT 2745.000 3402.910 2745.170 3403.080 ;
        RECT 2745.360 3402.910 2745.530 3403.080 ;
        RECT 2745.720 3402.910 2745.890 3403.080 ;
        RECT 2746.080 3402.910 2746.250 3403.080 ;
        RECT 2746.440 3402.910 2746.610 3403.080 ;
        RECT 2746.800 3402.910 2746.970 3403.080 ;
        RECT 2747.160 3402.910 2747.330 3403.080 ;
        RECT 2747.520 3402.910 2747.690 3403.080 ;
        RECT 2747.880 3402.910 2748.050 3403.080 ;
        RECT 2748.240 3402.910 2748.410 3403.080 ;
        RECT 2748.600 3402.910 2748.770 3403.080 ;
        RECT 2748.960 3402.910 2749.130 3403.080 ;
        RECT 2712.900 3400.785 2713.070 3400.955 ;
        RECT 2712.900 3400.425 2713.070 3400.595 ;
        RECT 2718.540 3400.785 2718.710 3400.955 ;
        RECT 2718.540 3400.425 2718.710 3400.595 ;
        RECT 2719.080 3400.785 2719.250 3400.955 ;
        RECT 2719.080 3400.425 2719.250 3400.595 ;
        RECT 2724.720 3400.785 2724.890 3400.955 ;
        RECT 2724.720 3400.425 2724.890 3400.595 ;
        RECT 2725.260 3400.785 2725.430 3400.955 ;
        RECT 2725.260 3400.425 2725.430 3400.595 ;
        RECT 2730.900 3400.785 2731.070 3400.955 ;
        RECT 2730.900 3400.425 2731.070 3400.595 ;
        RECT 2731.440 3400.785 2731.610 3400.955 ;
        RECT 2731.440 3400.425 2731.610 3400.595 ;
        RECT 2737.080 3400.785 2737.250 3400.955 ;
        RECT 2737.080 3400.425 2737.250 3400.595 ;
        RECT 2737.620 3400.785 2737.790 3400.955 ;
        RECT 2737.620 3400.425 2737.790 3400.595 ;
        RECT 2743.260 3400.785 2743.430 3400.955 ;
        RECT 2743.260 3400.425 2743.430 3400.595 ;
        RECT 2743.800 3400.785 2743.970 3400.955 ;
        RECT 2743.800 3400.425 2743.970 3400.595 ;
        RECT 2749.440 3400.785 2749.610 3400.955 ;
        RECT 2749.440 3400.425 2749.610 3400.595 ;
        RECT 2713.380 3399.960 2713.550 3400.130 ;
        RECT 2713.740 3399.960 2713.910 3400.130 ;
        RECT 2714.100 3399.960 2714.270 3400.130 ;
        RECT 2714.460 3399.960 2714.630 3400.130 ;
        RECT 2714.820 3399.960 2714.990 3400.130 ;
        RECT 2715.180 3399.960 2715.350 3400.130 ;
        RECT 2715.540 3399.960 2715.710 3400.130 ;
        RECT 2715.900 3399.960 2716.070 3400.130 ;
        RECT 2716.260 3399.960 2716.430 3400.130 ;
        RECT 2716.620 3399.960 2716.790 3400.130 ;
        RECT 2716.980 3399.960 2717.150 3400.130 ;
        RECT 2717.340 3399.960 2717.510 3400.130 ;
        RECT 2717.700 3399.960 2717.870 3400.130 ;
        RECT 2718.060 3399.960 2718.230 3400.130 ;
        RECT 2719.560 3399.960 2719.730 3400.130 ;
        RECT 2719.920 3399.960 2720.090 3400.130 ;
        RECT 2720.280 3399.960 2720.450 3400.130 ;
        RECT 2720.640 3399.960 2720.810 3400.130 ;
        RECT 2721.000 3399.960 2721.170 3400.130 ;
        RECT 2721.360 3399.960 2721.530 3400.130 ;
        RECT 2721.720 3399.960 2721.890 3400.130 ;
        RECT 2722.080 3399.960 2722.250 3400.130 ;
        RECT 2722.440 3399.960 2722.610 3400.130 ;
        RECT 2722.800 3399.960 2722.970 3400.130 ;
        RECT 2723.160 3399.960 2723.330 3400.130 ;
        RECT 2723.520 3399.960 2723.690 3400.130 ;
        RECT 2723.880 3399.960 2724.050 3400.130 ;
        RECT 2724.240 3399.960 2724.410 3400.130 ;
        RECT 2725.740 3399.960 2725.910 3400.130 ;
        RECT 2726.100 3399.960 2726.270 3400.130 ;
        RECT 2726.460 3399.960 2726.630 3400.130 ;
        RECT 2726.820 3399.960 2726.990 3400.130 ;
        RECT 2727.180 3399.960 2727.350 3400.130 ;
        RECT 2727.540 3399.960 2727.710 3400.130 ;
        RECT 2727.900 3399.960 2728.070 3400.130 ;
        RECT 2728.260 3399.960 2728.430 3400.130 ;
        RECT 2728.620 3399.960 2728.790 3400.130 ;
        RECT 2728.980 3399.960 2729.150 3400.130 ;
        RECT 2729.340 3399.960 2729.510 3400.130 ;
        RECT 2729.700 3399.960 2729.870 3400.130 ;
        RECT 2730.060 3399.960 2730.230 3400.130 ;
        RECT 2730.420 3399.960 2730.590 3400.130 ;
        RECT 2731.920 3399.960 2732.090 3400.130 ;
        RECT 2732.280 3399.960 2732.450 3400.130 ;
        RECT 2732.640 3399.960 2732.810 3400.130 ;
        RECT 2733.000 3399.960 2733.170 3400.130 ;
        RECT 2733.360 3399.960 2733.530 3400.130 ;
        RECT 2733.720 3399.960 2733.890 3400.130 ;
        RECT 2734.080 3399.960 2734.250 3400.130 ;
        RECT 2734.440 3399.960 2734.610 3400.130 ;
        RECT 2734.800 3399.960 2734.970 3400.130 ;
        RECT 2735.160 3399.960 2735.330 3400.130 ;
        RECT 2735.520 3399.960 2735.690 3400.130 ;
        RECT 2735.880 3399.960 2736.050 3400.130 ;
        RECT 2736.240 3399.960 2736.410 3400.130 ;
        RECT 2736.600 3399.960 2736.770 3400.130 ;
        RECT 2738.100 3399.960 2738.270 3400.130 ;
        RECT 2738.460 3399.960 2738.630 3400.130 ;
        RECT 2738.820 3399.960 2738.990 3400.130 ;
        RECT 2739.180 3399.960 2739.350 3400.130 ;
        RECT 2739.540 3399.960 2739.710 3400.130 ;
        RECT 2739.900 3399.960 2740.070 3400.130 ;
        RECT 2740.260 3399.960 2740.430 3400.130 ;
        RECT 2740.620 3399.960 2740.790 3400.130 ;
        RECT 2740.980 3399.960 2741.150 3400.130 ;
        RECT 2741.340 3399.960 2741.510 3400.130 ;
        RECT 2741.700 3399.960 2741.870 3400.130 ;
        RECT 2742.060 3399.960 2742.230 3400.130 ;
        RECT 2742.420 3399.960 2742.590 3400.130 ;
        RECT 2742.780 3399.960 2742.950 3400.130 ;
        RECT 2744.280 3399.960 2744.450 3400.130 ;
        RECT 2744.640 3399.960 2744.810 3400.130 ;
        RECT 2745.000 3399.960 2745.170 3400.130 ;
        RECT 2745.360 3399.960 2745.530 3400.130 ;
        RECT 2745.720 3399.960 2745.890 3400.130 ;
        RECT 2746.080 3399.960 2746.250 3400.130 ;
        RECT 2746.440 3399.960 2746.610 3400.130 ;
        RECT 2746.800 3399.960 2746.970 3400.130 ;
        RECT 2747.160 3399.960 2747.330 3400.130 ;
        RECT 2747.520 3399.960 2747.690 3400.130 ;
        RECT 2747.880 3399.960 2748.050 3400.130 ;
        RECT 2748.240 3399.960 2748.410 3400.130 ;
        RECT 2748.600 3399.960 2748.770 3400.130 ;
        RECT 2748.960 3399.960 2749.130 3400.130 ;
        RECT 2727.290 3397.300 2727.460 3397.470 ;
        RECT 2727.650 3397.300 2727.820 3397.470 ;
        RECT 2728.010 3397.300 2728.180 3397.470 ;
        RECT 2729.630 3397.300 2729.800 3397.470 ;
        RECT 2729.990 3397.300 2730.160 3397.470 ;
        RECT 2730.350 3397.300 2730.520 3397.470 ;
        RECT 2731.970 3397.300 2732.140 3397.470 ;
        RECT 2732.330 3397.300 2732.500 3397.470 ;
        RECT 2732.690 3397.300 2732.860 3397.470 ;
        RECT 2734.310 3397.300 2734.480 3397.470 ;
        RECT 2734.670 3397.300 2734.840 3397.470 ;
        RECT 2735.030 3397.300 2735.200 3397.470 ;
        RECT 2726.750 3396.835 2726.920 3397.005 ;
        RECT 2726.750 3396.475 2726.920 3396.645 ;
        RECT 2728.550 3396.835 2728.720 3397.005 ;
        RECT 2728.550 3396.475 2728.720 3396.645 ;
        RECT 2729.090 3396.835 2729.260 3397.005 ;
        RECT 2729.090 3396.475 2729.260 3396.645 ;
        RECT 2730.890 3396.835 2731.060 3397.005 ;
        RECT 2730.890 3396.475 2731.060 3396.645 ;
        RECT 2731.430 3396.835 2731.600 3397.005 ;
        RECT 2731.430 3396.475 2731.600 3396.645 ;
        RECT 2733.230 3396.835 2733.400 3397.005 ;
        RECT 2733.230 3396.475 2733.400 3396.645 ;
        RECT 2733.770 3396.835 2733.940 3397.005 ;
        RECT 2733.770 3396.475 2733.940 3396.645 ;
        RECT 2735.570 3396.835 2735.740 3397.005 ;
        RECT 2735.570 3396.475 2735.740 3396.645 ;
        RECT 2728.295 3394.175 2728.465 3394.345 ;
        RECT 2728.655 3394.175 2728.825 3394.345 ;
        RECT 2729.015 3394.175 2729.185 3394.345 ;
        RECT 2729.375 3394.175 2729.545 3394.345 ;
        RECT 2729.735 3394.175 2729.905 3394.345 ;
        RECT 2730.095 3394.175 2730.265 3394.345 ;
        RECT 2730.455 3394.175 2730.625 3394.345 ;
        RECT 2731.885 3394.175 2732.055 3394.345 ;
        RECT 2732.245 3394.175 2732.415 3394.345 ;
        RECT 2732.605 3394.175 2732.775 3394.345 ;
        RECT 2732.965 3394.175 2733.135 3394.345 ;
        RECT 2733.325 3394.175 2733.495 3394.345 ;
        RECT 2733.685 3394.175 2733.855 3394.345 ;
        RECT 2734.045 3394.175 2734.215 3394.345 ;
        RECT 2727.850 3393.780 2728.020 3393.950 ;
        RECT 2730.900 3393.780 2731.070 3393.950 ;
        RECT 2731.440 3393.780 2731.610 3393.950 ;
        RECT 2734.490 3393.780 2734.660 3393.950 ;
        RECT 2728.295 3393.385 2728.465 3393.555 ;
        RECT 2728.655 3393.385 2728.825 3393.555 ;
        RECT 2729.015 3393.385 2729.185 3393.555 ;
        RECT 2729.375 3393.385 2729.545 3393.555 ;
        RECT 2729.735 3393.385 2729.905 3393.555 ;
        RECT 2730.095 3393.385 2730.265 3393.555 ;
        RECT 2730.455 3393.385 2730.625 3393.555 ;
        RECT 2731.885 3393.385 2732.055 3393.555 ;
        RECT 2732.245 3393.385 2732.415 3393.555 ;
        RECT 2732.605 3393.385 2732.775 3393.555 ;
        RECT 2732.965 3393.385 2733.135 3393.555 ;
        RECT 2733.325 3393.385 2733.495 3393.555 ;
        RECT 2733.685 3393.385 2733.855 3393.555 ;
        RECT 2734.045 3393.385 2734.215 3393.555 ;
        RECT 2713.610 3391.550 2713.780 3391.720 ;
        RECT 2713.970 3391.550 2714.140 3391.720 ;
        RECT 2714.330 3391.550 2714.500 3391.720 ;
        RECT 2714.690 3391.550 2714.860 3391.720 ;
        RECT 2715.050 3391.550 2715.220 3391.720 ;
        RECT 2715.410 3391.550 2715.580 3391.720 ;
        RECT 2715.770 3391.550 2715.940 3391.720 ;
        RECT 2716.130 3391.550 2716.300 3391.720 ;
        RECT 2716.490 3391.550 2716.660 3391.720 ;
        RECT 2716.850 3391.550 2717.020 3391.720 ;
        RECT 2717.210 3391.550 2717.380 3391.720 ;
        RECT 2717.570 3391.550 2717.740 3391.720 ;
        RECT 2717.930 3391.550 2718.100 3391.720 ;
        RECT 2718.290 3391.550 2718.460 3391.720 ;
        RECT 2719.700 3391.550 2719.870 3391.720 ;
        RECT 2720.060 3391.550 2720.230 3391.720 ;
        RECT 2720.420 3391.550 2720.590 3391.720 ;
        RECT 2720.780 3391.550 2720.950 3391.720 ;
        RECT 2721.140 3391.550 2721.310 3391.720 ;
        RECT 2721.500 3391.550 2721.670 3391.720 ;
        RECT 2721.860 3391.550 2722.030 3391.720 ;
        RECT 2722.220 3391.550 2722.390 3391.720 ;
        RECT 2722.580 3391.550 2722.750 3391.720 ;
        RECT 2722.940 3391.550 2723.110 3391.720 ;
        RECT 2723.300 3391.550 2723.470 3391.720 ;
        RECT 2723.660 3391.550 2723.830 3391.720 ;
        RECT 2724.020 3391.550 2724.190 3391.720 ;
        RECT 2724.380 3391.550 2724.550 3391.720 ;
        RECT 2725.790 3391.550 2725.960 3391.720 ;
        RECT 2726.150 3391.550 2726.320 3391.720 ;
        RECT 2726.510 3391.550 2726.680 3391.720 ;
        RECT 2726.870 3391.550 2727.040 3391.720 ;
        RECT 2727.230 3391.550 2727.400 3391.720 ;
        RECT 2727.590 3391.550 2727.760 3391.720 ;
        RECT 2727.950 3391.550 2728.120 3391.720 ;
        RECT 2728.310 3391.550 2728.480 3391.720 ;
        RECT 2728.670 3391.550 2728.840 3391.720 ;
        RECT 2729.030 3391.550 2729.200 3391.720 ;
        RECT 2729.390 3391.550 2729.560 3391.720 ;
        RECT 2729.750 3391.550 2729.920 3391.720 ;
        RECT 2730.110 3391.550 2730.280 3391.720 ;
        RECT 2730.470 3391.550 2730.640 3391.720 ;
        RECT 2731.880 3391.550 2732.050 3391.720 ;
        RECT 2732.240 3391.550 2732.410 3391.720 ;
        RECT 2732.600 3391.550 2732.770 3391.720 ;
        RECT 2732.960 3391.550 2733.130 3391.720 ;
        RECT 2733.320 3391.550 2733.490 3391.720 ;
        RECT 2733.680 3391.550 2733.850 3391.720 ;
        RECT 2734.040 3391.550 2734.210 3391.720 ;
        RECT 2734.400 3391.550 2734.570 3391.720 ;
        RECT 2734.760 3391.550 2734.930 3391.720 ;
        RECT 2735.120 3391.550 2735.290 3391.720 ;
        RECT 2735.480 3391.550 2735.650 3391.720 ;
        RECT 2735.840 3391.550 2736.010 3391.720 ;
        RECT 2736.200 3391.550 2736.370 3391.720 ;
        RECT 2736.560 3391.550 2736.730 3391.720 ;
        RECT 2737.970 3391.550 2738.140 3391.720 ;
        RECT 2738.330 3391.550 2738.500 3391.720 ;
        RECT 2738.690 3391.550 2738.860 3391.720 ;
        RECT 2739.050 3391.550 2739.220 3391.720 ;
        RECT 2739.410 3391.550 2739.580 3391.720 ;
        RECT 2739.770 3391.550 2739.940 3391.720 ;
        RECT 2740.130 3391.550 2740.300 3391.720 ;
        RECT 2740.490 3391.550 2740.660 3391.720 ;
        RECT 2740.850 3391.550 2741.020 3391.720 ;
        RECT 2741.210 3391.550 2741.380 3391.720 ;
        RECT 2741.570 3391.550 2741.740 3391.720 ;
        RECT 2741.930 3391.550 2742.100 3391.720 ;
        RECT 2742.290 3391.550 2742.460 3391.720 ;
        RECT 2742.650 3391.550 2742.820 3391.720 ;
        RECT 2744.060 3391.550 2744.230 3391.720 ;
        RECT 2744.420 3391.550 2744.590 3391.720 ;
        RECT 2744.780 3391.550 2744.950 3391.720 ;
        RECT 2745.140 3391.550 2745.310 3391.720 ;
        RECT 2745.500 3391.550 2745.670 3391.720 ;
        RECT 2745.860 3391.550 2746.030 3391.720 ;
        RECT 2746.220 3391.550 2746.390 3391.720 ;
        RECT 2746.580 3391.550 2746.750 3391.720 ;
        RECT 2746.940 3391.550 2747.110 3391.720 ;
        RECT 2747.300 3391.550 2747.470 3391.720 ;
        RECT 2747.660 3391.550 2747.830 3391.720 ;
        RECT 2748.020 3391.550 2748.190 3391.720 ;
        RECT 2748.380 3391.550 2748.550 3391.720 ;
        RECT 2748.740 3391.550 2748.910 3391.720 ;
        RECT 2713.175 3391.085 2713.345 3391.255 ;
        RECT 2713.175 3390.725 2713.345 3390.895 ;
        RECT 2718.725 3391.085 2718.895 3391.255 ;
        RECT 2718.725 3390.725 2718.895 3390.895 ;
        RECT 2719.265 3391.085 2719.435 3391.255 ;
        RECT 2719.265 3390.725 2719.435 3390.895 ;
        RECT 2724.815 3391.085 2724.985 3391.255 ;
        RECT 2724.815 3390.725 2724.985 3390.895 ;
        RECT 2725.355 3391.085 2725.525 3391.255 ;
        RECT 2725.355 3390.725 2725.525 3390.895 ;
        RECT 2730.905 3391.085 2731.075 3391.255 ;
        RECT 2730.905 3390.725 2731.075 3390.895 ;
        RECT 2731.445 3391.085 2731.615 3391.255 ;
        RECT 2731.445 3390.725 2731.615 3390.895 ;
        RECT 2736.995 3391.085 2737.165 3391.255 ;
        RECT 2736.995 3390.725 2737.165 3390.895 ;
        RECT 2737.535 3391.085 2737.705 3391.255 ;
        RECT 2737.535 3390.725 2737.705 3390.895 ;
        RECT 2743.085 3391.085 2743.255 3391.255 ;
        RECT 2743.085 3390.725 2743.255 3390.895 ;
        RECT 2743.625 3391.085 2743.795 3391.255 ;
        RECT 2743.625 3390.725 2743.795 3390.895 ;
        RECT 2749.175 3391.085 2749.345 3391.255 ;
        RECT 2749.175 3390.725 2749.345 3390.895 ;
        RECT 2713.610 3390.260 2713.780 3390.430 ;
        RECT 2713.970 3390.260 2714.140 3390.430 ;
        RECT 2714.330 3390.260 2714.500 3390.430 ;
        RECT 2714.690 3390.260 2714.860 3390.430 ;
        RECT 2715.050 3390.260 2715.220 3390.430 ;
        RECT 2715.410 3390.260 2715.580 3390.430 ;
        RECT 2715.770 3390.260 2715.940 3390.430 ;
        RECT 2716.130 3390.260 2716.300 3390.430 ;
        RECT 2716.490 3390.260 2716.660 3390.430 ;
        RECT 2716.850 3390.260 2717.020 3390.430 ;
        RECT 2717.210 3390.260 2717.380 3390.430 ;
        RECT 2717.570 3390.260 2717.740 3390.430 ;
        RECT 2717.930 3390.260 2718.100 3390.430 ;
        RECT 2718.290 3390.260 2718.460 3390.430 ;
        RECT 2719.700 3390.260 2719.870 3390.430 ;
        RECT 2720.060 3390.260 2720.230 3390.430 ;
        RECT 2720.420 3390.260 2720.590 3390.430 ;
        RECT 2720.780 3390.260 2720.950 3390.430 ;
        RECT 2721.140 3390.260 2721.310 3390.430 ;
        RECT 2721.500 3390.260 2721.670 3390.430 ;
        RECT 2721.860 3390.260 2722.030 3390.430 ;
        RECT 2722.220 3390.260 2722.390 3390.430 ;
        RECT 2722.580 3390.260 2722.750 3390.430 ;
        RECT 2722.940 3390.260 2723.110 3390.430 ;
        RECT 2723.300 3390.260 2723.470 3390.430 ;
        RECT 2723.660 3390.260 2723.830 3390.430 ;
        RECT 2724.020 3390.260 2724.190 3390.430 ;
        RECT 2724.380 3390.260 2724.550 3390.430 ;
        RECT 2725.790 3390.260 2725.960 3390.430 ;
        RECT 2726.150 3390.260 2726.320 3390.430 ;
        RECT 2726.510 3390.260 2726.680 3390.430 ;
        RECT 2726.870 3390.260 2727.040 3390.430 ;
        RECT 2727.230 3390.260 2727.400 3390.430 ;
        RECT 2727.590 3390.260 2727.760 3390.430 ;
        RECT 2727.950 3390.260 2728.120 3390.430 ;
        RECT 2728.310 3390.260 2728.480 3390.430 ;
        RECT 2728.670 3390.260 2728.840 3390.430 ;
        RECT 2729.030 3390.260 2729.200 3390.430 ;
        RECT 2729.390 3390.260 2729.560 3390.430 ;
        RECT 2729.750 3390.260 2729.920 3390.430 ;
        RECT 2730.110 3390.260 2730.280 3390.430 ;
        RECT 2730.470 3390.260 2730.640 3390.430 ;
        RECT 2731.880 3390.260 2732.050 3390.430 ;
        RECT 2732.240 3390.260 2732.410 3390.430 ;
        RECT 2732.600 3390.260 2732.770 3390.430 ;
        RECT 2732.960 3390.260 2733.130 3390.430 ;
        RECT 2733.320 3390.260 2733.490 3390.430 ;
        RECT 2733.680 3390.260 2733.850 3390.430 ;
        RECT 2734.040 3390.260 2734.210 3390.430 ;
        RECT 2734.400 3390.260 2734.570 3390.430 ;
        RECT 2734.760 3390.260 2734.930 3390.430 ;
        RECT 2735.120 3390.260 2735.290 3390.430 ;
        RECT 2735.480 3390.260 2735.650 3390.430 ;
        RECT 2735.840 3390.260 2736.010 3390.430 ;
        RECT 2736.200 3390.260 2736.370 3390.430 ;
        RECT 2736.560 3390.260 2736.730 3390.430 ;
        RECT 2737.970 3390.260 2738.140 3390.430 ;
        RECT 2738.330 3390.260 2738.500 3390.430 ;
        RECT 2738.690 3390.260 2738.860 3390.430 ;
        RECT 2739.050 3390.260 2739.220 3390.430 ;
        RECT 2739.410 3390.260 2739.580 3390.430 ;
        RECT 2739.770 3390.260 2739.940 3390.430 ;
        RECT 2740.130 3390.260 2740.300 3390.430 ;
        RECT 2740.490 3390.260 2740.660 3390.430 ;
        RECT 2740.850 3390.260 2741.020 3390.430 ;
        RECT 2741.210 3390.260 2741.380 3390.430 ;
        RECT 2741.570 3390.260 2741.740 3390.430 ;
        RECT 2741.930 3390.260 2742.100 3390.430 ;
        RECT 2742.290 3390.260 2742.460 3390.430 ;
        RECT 2742.650 3390.260 2742.820 3390.430 ;
        RECT 2744.060 3390.260 2744.230 3390.430 ;
        RECT 2744.420 3390.260 2744.590 3390.430 ;
        RECT 2744.780 3390.260 2744.950 3390.430 ;
        RECT 2745.140 3390.260 2745.310 3390.430 ;
        RECT 2745.500 3390.260 2745.670 3390.430 ;
        RECT 2745.860 3390.260 2746.030 3390.430 ;
        RECT 2746.220 3390.260 2746.390 3390.430 ;
        RECT 2746.580 3390.260 2746.750 3390.430 ;
        RECT 2746.940 3390.260 2747.110 3390.430 ;
        RECT 2747.300 3390.260 2747.470 3390.430 ;
        RECT 2747.660 3390.260 2747.830 3390.430 ;
        RECT 2748.020 3390.260 2748.190 3390.430 ;
        RECT 2748.380 3390.260 2748.550 3390.430 ;
        RECT 2748.740 3390.260 2748.910 3390.430 ;
        RECT 2717.125 3385.960 2722.695 3387.930 ;
        RECT 2724.725 3385.960 2730.295 3387.930 ;
        RECT 2732.275 3385.990 2737.845 3387.960 ;
        RECT 2739.825 3385.990 2745.395 3387.960 ;
      LAYER met1 ;
        RECT 2709.645 3451.580 2709.875 3451.690 ;
        RECT 2715.285 3451.630 2715.515 3451.690 ;
        RECT 2715.825 3451.630 2716.055 3451.690 ;
        RECT 2715.285 3451.580 2716.055 3451.630 ;
        RECT 2721.465 3451.630 2721.695 3451.690 ;
        RECT 2722.005 3451.630 2722.235 3451.690 ;
        RECT 2727.645 3451.630 2727.875 3451.690 ;
        RECT 2728.185 3451.630 2728.415 3451.690 ;
        RECT 2721.465 3451.580 2722.235 3451.630 ;
        RECT 2727.635 3451.580 2728.415 3451.630 ;
        RECT 2733.825 3451.630 2734.055 3451.690 ;
        RECT 2734.365 3451.630 2734.595 3451.690 ;
        RECT 2733.825 3451.580 2734.595 3451.630 ;
        RECT 2740.005 3451.630 2740.235 3451.690 ;
        RECT 2740.545 3451.630 2740.775 3451.690 ;
        RECT 2746.185 3451.630 2746.415 3451.690 ;
        RECT 2746.725 3451.630 2746.955 3451.690 ;
        RECT 2740.005 3451.580 2740.785 3451.630 ;
        RECT 2746.185 3451.580 2746.955 3451.630 ;
        RECT 2752.365 3451.580 2752.595 3451.690 ;
        RECT 2709.645 3451.380 2752.595 3451.580 ;
        RECT 2709.585 3450.880 2752.635 3451.380 ;
        RECT 2711.685 3450.680 2712.185 3450.880 ;
        RECT 2712.535 3450.680 2713.035 3450.880 ;
        RECT 2724.285 3450.680 2724.785 3450.880 ;
        RECT 2725.135 3450.680 2725.635 3450.880 ;
        RECT 2736.735 3450.680 2737.235 3450.880 ;
        RECT 2737.585 3450.680 2738.085 3450.880 ;
        RECT 2748.985 3450.680 2749.485 3450.880 ;
        RECT 2749.835 3450.680 2750.335 3450.880 ;
        RECT 2709.645 3448.880 2709.875 3448.990 ;
        RECT 2715.285 3448.930 2715.515 3448.990 ;
        RECT 2715.825 3448.930 2716.055 3448.990 ;
        RECT 2715.285 3448.880 2716.055 3448.930 ;
        RECT 2721.465 3448.930 2721.695 3448.990 ;
        RECT 2722.005 3448.930 2722.235 3448.990 ;
        RECT 2727.645 3448.930 2727.875 3448.990 ;
        RECT 2728.185 3448.930 2728.415 3448.990 ;
        RECT 2721.465 3448.880 2722.235 3448.930 ;
        RECT 2727.635 3448.880 2728.415 3448.930 ;
        RECT 2733.825 3448.930 2734.055 3448.990 ;
        RECT 2734.365 3448.930 2734.595 3448.990 ;
        RECT 2733.825 3448.880 2734.595 3448.930 ;
        RECT 2740.005 3448.930 2740.235 3448.990 ;
        RECT 2740.545 3448.930 2740.775 3448.990 ;
        RECT 2746.185 3448.930 2746.415 3448.990 ;
        RECT 2746.725 3448.930 2746.955 3448.990 ;
        RECT 2740.005 3448.880 2740.785 3448.930 ;
        RECT 2746.185 3448.880 2746.955 3448.930 ;
        RECT 2752.365 3448.880 2752.595 3448.990 ;
        RECT 2709.645 3448.680 2752.595 3448.880 ;
        RECT 2709.635 3448.530 2752.595 3448.680 ;
        RECT 2709.635 3448.180 2752.535 3448.530 ;
        RECT 2711.685 3447.980 2712.185 3448.180 ;
        RECT 2712.535 3447.980 2713.035 3448.180 ;
        RECT 2724.285 3447.980 2724.785 3448.180 ;
        RECT 2725.135 3447.980 2725.635 3448.180 ;
        RECT 2736.735 3447.980 2737.235 3448.180 ;
        RECT 2737.585 3447.980 2738.085 3448.180 ;
        RECT 2748.985 3447.930 2749.485 3448.180 ;
        RECT 2749.835 3447.930 2750.335 3448.180 ;
        RECT 2709.645 3446.180 2709.875 3446.290 ;
        RECT 2715.285 3446.230 2715.515 3446.290 ;
        RECT 2715.825 3446.230 2716.055 3446.290 ;
        RECT 2715.285 3446.180 2716.055 3446.230 ;
        RECT 2721.465 3446.230 2721.695 3446.290 ;
        RECT 2722.005 3446.230 2722.235 3446.290 ;
        RECT 2727.645 3446.230 2727.875 3446.290 ;
        RECT 2728.185 3446.230 2728.415 3446.290 ;
        RECT 2721.465 3446.180 2722.235 3446.230 ;
        RECT 2727.635 3446.180 2728.415 3446.230 ;
        RECT 2733.825 3446.230 2734.055 3446.290 ;
        RECT 2734.365 3446.230 2734.595 3446.290 ;
        RECT 2733.825 3446.180 2734.595 3446.230 ;
        RECT 2740.005 3446.230 2740.235 3446.290 ;
        RECT 2740.545 3446.230 2740.775 3446.290 ;
        RECT 2746.185 3446.230 2746.415 3446.290 ;
        RECT 2746.725 3446.230 2746.955 3446.290 ;
        RECT 2740.005 3446.180 2740.785 3446.230 ;
        RECT 2746.185 3446.180 2746.955 3446.230 ;
        RECT 2752.365 3446.180 2752.595 3446.290 ;
        RECT 2709.645 3445.830 2752.595 3446.180 ;
        RECT 2709.685 3445.480 2752.585 3445.830 ;
        RECT 2711.685 3445.280 2712.185 3445.480 ;
        RECT 2712.535 3445.280 2713.035 3445.480 ;
        RECT 2724.285 3445.280 2724.785 3445.480 ;
        RECT 2725.135 3445.280 2725.635 3445.480 ;
        RECT 2736.735 3445.230 2737.235 3445.480 ;
        RECT 2737.585 3445.230 2738.085 3445.480 ;
        RECT 2748.985 3445.280 2749.485 3445.480 ;
        RECT 2749.835 3445.280 2750.335 3445.480 ;
        RECT 2709.645 3443.480 2709.875 3443.590 ;
        RECT 2715.285 3443.530 2715.515 3443.590 ;
        RECT 2715.825 3443.530 2716.055 3443.590 ;
        RECT 2715.285 3443.480 2716.055 3443.530 ;
        RECT 2721.465 3443.530 2721.695 3443.590 ;
        RECT 2722.005 3443.530 2722.235 3443.590 ;
        RECT 2727.645 3443.530 2727.875 3443.590 ;
        RECT 2728.185 3443.530 2728.415 3443.590 ;
        RECT 2721.465 3443.480 2722.235 3443.530 ;
        RECT 2727.635 3443.480 2728.415 3443.530 ;
        RECT 2733.825 3443.530 2734.055 3443.590 ;
        RECT 2734.365 3443.530 2734.595 3443.590 ;
        RECT 2740.005 3443.530 2740.235 3443.590 ;
        RECT 2740.545 3443.530 2740.775 3443.590 ;
        RECT 2733.825 3443.480 2734.595 3443.530 ;
        RECT 2739.985 3443.480 2740.775 3443.530 ;
        RECT 2746.185 3443.530 2746.415 3443.590 ;
        RECT 2746.725 3443.530 2746.955 3443.590 ;
        RECT 2746.185 3443.480 2746.955 3443.530 ;
        RECT 2752.365 3443.480 2752.595 3443.590 ;
        RECT 2709.645 3443.230 2752.595 3443.480 ;
        RECT 2709.645 3443.130 2709.875 3443.230 ;
        RECT 2715.285 3443.180 2716.055 3443.230 ;
        RECT 2715.285 3443.130 2715.515 3443.180 ;
        RECT 2715.825 3443.130 2716.055 3443.180 ;
        RECT 2721.465 3443.180 2722.235 3443.230 ;
        RECT 2727.635 3443.180 2728.415 3443.230 ;
        RECT 2721.465 3443.130 2721.695 3443.180 ;
        RECT 2722.005 3443.130 2722.235 3443.180 ;
        RECT 2727.645 3443.130 2727.875 3443.180 ;
        RECT 2728.185 3443.130 2728.415 3443.180 ;
        RECT 2733.825 3443.180 2734.595 3443.230 ;
        RECT 2739.985 3443.180 2740.775 3443.230 ;
        RECT 2733.825 3443.130 2734.055 3443.180 ;
        RECT 2734.365 3443.130 2734.595 3443.180 ;
        RECT 2740.005 3443.130 2740.235 3443.180 ;
        RECT 2740.545 3443.130 2740.775 3443.180 ;
        RECT 2746.185 3443.180 2746.955 3443.230 ;
        RECT 2746.185 3443.130 2746.415 3443.180 ;
        RECT 2746.725 3443.130 2746.955 3443.180 ;
        RECT 2752.365 3443.130 2752.595 3443.230 ;
        RECT 2710.080 3442.980 2715.080 3443.080 ;
        RECT 2716.260 3442.980 2721.260 3443.080 ;
        RECT 2722.440 3442.980 2727.440 3443.080 ;
        RECT 2728.620 3442.980 2733.620 3443.080 ;
        RECT 2734.800 3442.980 2739.800 3443.080 ;
        RECT 2740.980 3442.980 2745.980 3443.080 ;
        RECT 2747.160 3442.980 2752.160 3443.080 ;
        RECT 2710.035 3442.780 2752.235 3442.980 ;
        RECT 2711.685 3442.580 2712.185 3442.780 ;
        RECT 2712.535 3442.580 2713.035 3442.780 ;
        RECT 2720.035 3442.480 2721.185 3442.780 ;
        RECT 2724.235 3442.580 2724.735 3442.780 ;
        RECT 2725.085 3442.580 2725.585 3442.780 ;
        RECT 2732.085 3442.580 2733.235 3442.780 ;
        RECT 2736.685 3442.580 2737.185 3442.780 ;
        RECT 2737.535 3442.580 2738.035 3442.780 ;
        RECT 2744.385 3442.480 2745.535 3442.780 ;
        RECT 2749.135 3442.580 2749.635 3442.780 ;
        RECT 2749.985 3442.580 2750.485 3442.780 ;
        RECT 2709.645 3440.580 2709.875 3440.690 ;
        RECT 2715.285 3440.630 2715.515 3440.690 ;
        RECT 2715.825 3440.630 2716.055 3440.690 ;
        RECT 2715.285 3440.580 2716.055 3440.630 ;
        RECT 2721.465 3440.630 2721.695 3440.690 ;
        RECT 2722.005 3440.630 2722.235 3440.690 ;
        RECT 2721.465 3440.580 2722.235 3440.630 ;
        RECT 2727.645 3440.630 2727.875 3440.690 ;
        RECT 2728.185 3440.630 2728.415 3440.690 ;
        RECT 2733.825 3440.630 2734.055 3440.690 ;
        RECT 2734.365 3440.630 2734.595 3440.690 ;
        RECT 2740.005 3440.630 2740.235 3440.690 ;
        RECT 2740.545 3440.630 2740.775 3440.690 ;
        RECT 2727.645 3440.580 2728.435 3440.630 ;
        RECT 2733.825 3440.580 2734.595 3440.630 ;
        RECT 2739.985 3440.580 2740.775 3440.630 ;
        RECT 2746.185 3440.630 2746.415 3440.690 ;
        RECT 2746.725 3440.630 2746.955 3440.690 ;
        RECT 2746.185 3440.580 2746.955 3440.630 ;
        RECT 2752.365 3440.580 2752.595 3440.690 ;
        RECT 2709.645 3440.330 2752.595 3440.580 ;
        RECT 2709.645 3440.230 2709.875 3440.330 ;
        RECT 2715.285 3440.280 2716.055 3440.330 ;
        RECT 2715.285 3440.230 2715.515 3440.280 ;
        RECT 2715.825 3440.230 2716.055 3440.280 ;
        RECT 2721.465 3440.280 2722.235 3440.330 ;
        RECT 2721.465 3440.230 2721.695 3440.280 ;
        RECT 2722.005 3440.230 2722.235 3440.280 ;
        RECT 2727.645 3440.280 2728.435 3440.330 ;
        RECT 2733.825 3440.280 2734.595 3440.330 ;
        RECT 2739.985 3440.280 2740.775 3440.330 ;
        RECT 2727.645 3440.230 2727.875 3440.280 ;
        RECT 2728.185 3440.230 2728.415 3440.280 ;
        RECT 2733.825 3440.230 2734.055 3440.280 ;
        RECT 2734.365 3440.230 2734.595 3440.280 ;
        RECT 2740.005 3440.230 2740.235 3440.280 ;
        RECT 2740.545 3440.230 2740.775 3440.280 ;
        RECT 2746.185 3440.280 2746.955 3440.330 ;
        RECT 2746.185 3440.230 2746.415 3440.280 ;
        RECT 2746.725 3440.230 2746.955 3440.280 ;
        RECT 2752.365 3440.230 2752.595 3440.330 ;
        RECT 2710.080 3440.080 2715.080 3440.180 ;
        RECT 2716.260 3440.080 2721.260 3440.180 ;
        RECT 2722.440 3440.080 2727.440 3440.180 ;
        RECT 2728.620 3440.080 2733.620 3440.180 ;
        RECT 2734.800 3440.080 2739.800 3440.180 ;
        RECT 2740.980 3440.080 2745.980 3440.180 ;
        RECT 2747.160 3440.080 2752.160 3440.180 ;
        RECT 2710.035 3439.880 2752.235 3440.080 ;
        RECT 2711.685 3439.680 2712.185 3439.880 ;
        RECT 2712.535 3439.680 2713.035 3439.880 ;
        RECT 2720.035 3439.530 2721.185 3439.880 ;
        RECT 2724.235 3439.680 2724.735 3439.880 ;
        RECT 2725.085 3439.680 2725.585 3439.880 ;
        RECT 2732.085 3439.580 2733.235 3439.880 ;
        RECT 2736.685 3439.630 2737.185 3439.880 ;
        RECT 2737.535 3439.630 2738.035 3439.880 ;
        RECT 2744.385 3439.580 2745.535 3439.880 ;
        RECT 2749.135 3439.680 2749.635 3439.880 ;
        RECT 2749.985 3439.680 2750.485 3439.880 ;
        RECT 2681.285 3437.855 2683.435 3439.280 ;
        RECT 2778.785 3437.855 2780.935 3440.130 ;
        RECT 2681.285 3432.165 2683.955 3437.855 ;
        RECT 2694.065 3437.330 2696.110 3437.855 ;
        RECT 2709.645 3437.680 2709.875 3437.790 ;
        RECT 2715.285 3437.730 2715.515 3437.790 ;
        RECT 2715.825 3437.730 2716.055 3437.790 ;
        RECT 2715.285 3437.680 2716.055 3437.730 ;
        RECT 2721.465 3437.730 2721.695 3437.790 ;
        RECT 2722.005 3437.730 2722.235 3437.790 ;
        RECT 2727.645 3437.730 2727.875 3437.790 ;
        RECT 2728.185 3437.730 2728.415 3437.790 ;
        RECT 2721.465 3437.680 2722.235 3437.730 ;
        RECT 2727.635 3437.680 2728.415 3437.730 ;
        RECT 2733.825 3437.730 2734.055 3437.790 ;
        RECT 2734.365 3437.730 2734.595 3437.790 ;
        RECT 2740.005 3437.730 2740.235 3437.790 ;
        RECT 2740.545 3437.730 2740.775 3437.790 ;
        RECT 2733.825 3437.680 2734.595 3437.730 ;
        RECT 2739.985 3437.680 2740.775 3437.730 ;
        RECT 2746.185 3437.730 2746.415 3437.790 ;
        RECT 2746.725 3437.730 2746.955 3437.790 ;
        RECT 2746.185 3437.680 2746.955 3437.730 ;
        RECT 2752.365 3437.680 2752.595 3437.790 ;
        RECT 2709.645 3437.430 2752.595 3437.680 ;
        RECT 2709.645 3437.330 2709.875 3437.430 ;
        RECT 2715.285 3437.380 2716.055 3437.430 ;
        RECT 2715.285 3437.330 2715.515 3437.380 ;
        RECT 2715.825 3437.330 2716.055 3437.380 ;
        RECT 2721.465 3437.380 2722.235 3437.430 ;
        RECT 2727.635 3437.380 2728.415 3437.430 ;
        RECT 2721.465 3437.330 2721.695 3437.380 ;
        RECT 2722.005 3437.330 2722.235 3437.380 ;
        RECT 2727.645 3437.330 2727.875 3437.380 ;
        RECT 2728.185 3437.330 2728.415 3437.380 ;
        RECT 2733.825 3437.380 2734.595 3437.430 ;
        RECT 2739.985 3437.380 2740.775 3437.430 ;
        RECT 2733.825 3437.330 2734.055 3437.380 ;
        RECT 2734.365 3437.330 2734.595 3437.380 ;
        RECT 2740.005 3437.330 2740.235 3437.380 ;
        RECT 2740.545 3437.330 2740.775 3437.380 ;
        RECT 2746.185 3437.380 2746.955 3437.430 ;
        RECT 2746.185 3437.330 2746.415 3437.380 ;
        RECT 2746.725 3437.330 2746.955 3437.380 ;
        RECT 2752.365 3437.330 2752.595 3437.430 ;
        RECT 2767.210 3437.330 2769.255 3437.855 ;
        RECT 2693.435 3435.130 2696.110 3437.330 ;
        RECT 2710.080 3437.130 2715.080 3437.280 ;
        RECT 2716.260 3437.130 2721.260 3437.280 ;
        RECT 2722.440 3437.130 2727.440 3437.280 ;
        RECT 2728.620 3437.130 2733.620 3437.280 ;
        RECT 2734.800 3437.130 2739.800 3437.280 ;
        RECT 2740.980 3437.130 2745.980 3437.280 ;
        RECT 2747.160 3437.130 2752.160 3437.280 ;
        RECT 2710.035 3436.930 2752.235 3437.130 ;
        RECT 2711.585 3436.630 2712.085 3436.930 ;
        RECT 2712.635 3436.630 2713.135 3436.930 ;
        RECT 2720.035 3436.680 2721.185 3436.930 ;
        RECT 2724.235 3436.780 2724.735 3436.930 ;
        RECT 2725.085 3436.780 2725.585 3436.930 ;
        RECT 2732.085 3436.680 2733.235 3436.930 ;
        RECT 2736.685 3436.780 2737.185 3436.930 ;
        RECT 2737.535 3436.780 2738.035 3436.930 ;
        RECT 2744.385 3436.680 2745.535 3436.930 ;
        RECT 2749.135 3436.780 2749.635 3436.930 ;
        RECT 2749.985 3436.780 2750.485 3436.930 ;
        RECT 2766.585 3435.130 2769.255 3437.330 ;
        RECT 2693.435 3435.090 2700.635 3435.130 ;
        RECT 2761.735 3435.090 2769.255 3435.130 ;
        RECT 2693.435 3434.980 2700.675 3435.090 ;
        RECT 2706.085 3435.030 2706.315 3435.090 ;
        RECT 2706.625 3435.030 2706.855 3435.090 ;
        RECT 2706.085 3434.980 2706.855 3435.030 ;
        RECT 2712.265 3435.030 2712.495 3435.090 ;
        RECT 2712.805 3435.030 2713.035 3435.090 ;
        RECT 2718.445 3435.030 2718.675 3435.090 ;
        RECT 2718.985 3435.030 2719.215 3435.090 ;
        RECT 2712.265 3434.980 2713.035 3435.030 ;
        RECT 2718.435 3434.980 2719.215 3435.030 ;
        RECT 2724.625 3435.030 2724.855 3435.090 ;
        RECT 2725.165 3435.030 2725.395 3435.090 ;
        RECT 2724.625 3434.980 2725.395 3435.030 ;
        RECT 2730.805 3435.030 2731.035 3435.090 ;
        RECT 2731.345 3435.030 2731.575 3435.090 ;
        RECT 2736.985 3435.030 2737.215 3435.090 ;
        RECT 2737.525 3435.030 2737.755 3435.090 ;
        RECT 2730.805 3434.980 2731.585 3435.030 ;
        RECT 2736.985 3434.980 2737.755 3435.030 ;
        RECT 2743.165 3435.030 2743.395 3435.090 ;
        RECT 2743.705 3435.030 2743.935 3435.090 ;
        RECT 2749.345 3435.030 2749.575 3435.090 ;
        RECT 2749.885 3435.030 2750.115 3435.090 ;
        RECT 2743.165 3434.980 2743.935 3435.030 ;
        RECT 2749.335 3434.980 2750.115 3435.030 ;
        RECT 2755.525 3435.030 2755.755 3435.090 ;
        RECT 2756.065 3435.030 2756.295 3435.090 ;
        RECT 2755.525 3434.980 2756.295 3435.030 ;
        RECT 2761.705 3434.980 2769.255 3435.090 ;
        RECT 2693.435 3434.780 2769.255 3434.980 ;
        RECT 2693.435 3434.630 2700.675 3434.780 ;
        RECT 2706.085 3434.680 2706.855 3434.780 ;
        RECT 2706.085 3434.630 2706.315 3434.680 ;
        RECT 2706.625 3434.630 2706.855 3434.680 ;
        RECT 2712.265 3434.680 2713.035 3434.780 ;
        RECT 2718.435 3434.680 2719.215 3434.780 ;
        RECT 2712.265 3434.630 2712.495 3434.680 ;
        RECT 2712.805 3434.630 2713.035 3434.680 ;
        RECT 2718.445 3434.630 2718.675 3434.680 ;
        RECT 2718.985 3434.630 2719.215 3434.680 ;
        RECT 2724.625 3434.680 2725.395 3434.780 ;
        RECT 2724.625 3434.630 2724.855 3434.680 ;
        RECT 2725.165 3434.630 2725.395 3434.680 ;
        RECT 2730.805 3434.680 2731.585 3434.780 ;
        RECT 2736.985 3434.680 2737.755 3434.780 ;
        RECT 2730.805 3434.630 2731.035 3434.680 ;
        RECT 2731.345 3434.630 2731.575 3434.680 ;
        RECT 2736.985 3434.630 2737.215 3434.680 ;
        RECT 2737.525 3434.630 2737.755 3434.680 ;
        RECT 2743.165 3434.680 2743.935 3434.780 ;
        RECT 2749.335 3434.680 2750.115 3434.780 ;
        RECT 2743.165 3434.630 2743.395 3434.680 ;
        RECT 2743.705 3434.630 2743.935 3434.680 ;
        RECT 2749.345 3434.630 2749.575 3434.680 ;
        RECT 2749.885 3434.630 2750.115 3434.680 ;
        RECT 2755.525 3434.680 2756.295 3434.780 ;
        RECT 2755.525 3434.630 2755.755 3434.680 ;
        RECT 2756.065 3434.630 2756.295 3434.680 ;
        RECT 2761.705 3434.630 2769.255 3434.780 ;
        RECT 2693.435 3432.430 2696.110 3434.630 ;
        RECT 2693.435 3432.390 2700.635 3432.430 ;
        RECT 2693.435 3432.280 2700.675 3432.390 ;
        RECT 2706.085 3432.380 2706.315 3432.390 ;
        RECT 2706.625 3432.380 2706.855 3432.390 ;
        RECT 2706.085 3432.280 2706.855 3432.380 ;
        RECT 2712.265 3432.330 2712.495 3432.390 ;
        RECT 2712.805 3432.330 2713.035 3432.390 ;
        RECT 2718.445 3432.330 2718.675 3432.390 ;
        RECT 2718.985 3432.330 2719.215 3432.390 ;
        RECT 2712.265 3432.280 2713.035 3432.330 ;
        RECT 2718.435 3432.280 2719.215 3432.330 ;
        RECT 2724.625 3432.330 2724.855 3432.390 ;
        RECT 2725.165 3432.330 2725.395 3432.390 ;
        RECT 2724.625 3432.280 2725.395 3432.330 ;
        RECT 2730.805 3432.330 2731.035 3432.390 ;
        RECT 2731.345 3432.330 2731.575 3432.390 ;
        RECT 2736.985 3432.330 2737.215 3432.390 ;
        RECT 2737.525 3432.330 2737.755 3432.390 ;
        RECT 2730.805 3432.280 2731.585 3432.330 ;
        RECT 2736.985 3432.280 2737.755 3432.330 ;
        RECT 2743.165 3432.330 2743.395 3432.390 ;
        RECT 2743.705 3432.330 2743.935 3432.390 ;
        RECT 2749.345 3432.330 2749.575 3432.390 ;
        RECT 2749.885 3432.330 2750.115 3432.390 ;
        RECT 2743.165 3432.280 2743.935 3432.330 ;
        RECT 2749.335 3432.280 2750.115 3432.330 ;
        RECT 2755.525 3432.330 2755.755 3432.390 ;
        RECT 2756.065 3432.330 2756.295 3432.390 ;
        RECT 2755.525 3432.280 2756.295 3432.330 ;
        RECT 2761.705 3432.380 2761.935 3432.390 ;
        RECT 2766.585 3432.380 2769.255 3434.630 ;
        RECT 2761.705 3432.280 2769.255 3432.380 ;
        RECT 2693.435 3432.165 2769.255 3432.280 ;
        RECT 2778.785 3432.165 2781.410 3437.855 ;
        RECT 2681.285 3430.505 2683.435 3432.165 ;
        RECT 2693.435 3432.080 2768.735 3432.165 ;
        RECT 2693.435 3431.930 2700.675 3432.080 ;
        RECT 2706.085 3432.030 2706.855 3432.080 ;
        RECT 2706.085 3431.930 2706.315 3432.030 ;
        RECT 2706.625 3431.930 2706.855 3432.030 ;
        RECT 2712.265 3431.980 2713.035 3432.080 ;
        RECT 2718.435 3431.980 2719.215 3432.080 ;
        RECT 2712.265 3431.930 2712.495 3431.980 ;
        RECT 2712.805 3431.930 2713.035 3431.980 ;
        RECT 2718.445 3431.930 2718.675 3431.980 ;
        RECT 2718.985 3431.930 2719.215 3431.980 ;
        RECT 2724.625 3431.980 2725.395 3432.080 ;
        RECT 2724.625 3431.930 2724.855 3431.980 ;
        RECT 2725.165 3431.930 2725.395 3431.980 ;
        RECT 2730.805 3431.980 2731.585 3432.080 ;
        RECT 2736.985 3431.980 2737.755 3432.080 ;
        RECT 2730.805 3431.930 2731.035 3431.980 ;
        RECT 2731.345 3431.930 2731.575 3431.980 ;
        RECT 2736.985 3431.930 2737.215 3431.980 ;
        RECT 2737.525 3431.930 2737.755 3431.980 ;
        RECT 2743.165 3431.980 2743.935 3432.080 ;
        RECT 2749.335 3431.980 2750.115 3432.080 ;
        RECT 2743.165 3431.930 2743.395 3431.980 ;
        RECT 2743.705 3431.930 2743.935 3431.980 ;
        RECT 2749.345 3431.930 2749.575 3431.980 ;
        RECT 2749.885 3431.930 2750.115 3431.980 ;
        RECT 2755.525 3431.980 2756.295 3432.080 ;
        RECT 2755.525 3431.930 2755.755 3431.980 ;
        RECT 2756.065 3431.930 2756.295 3431.980 ;
        RECT 2761.705 3431.930 2768.735 3432.080 ;
        RECT 2693.435 3431.880 2700.635 3431.930 ;
        RECT 2761.735 3431.880 2768.735 3431.930 ;
        RECT 2693.435 3430.505 2695.585 3431.880 ;
        RECT 2766.585 3430.505 2768.735 3431.880 ;
        RECT 2778.785 3430.505 2780.935 3432.165 ;
        RECT 2681.285 3424.980 2683.955 3430.505 ;
        RECT 2681.910 3424.815 2683.955 3424.980 ;
        RECT 2693.435 3429.730 2696.110 3430.505 ;
        RECT 2766.585 3429.730 2769.255 3430.505 ;
        RECT 2693.435 3429.580 2700.735 3429.730 ;
        RECT 2761.735 3429.690 2769.255 3429.730 ;
        RECT 2706.085 3429.630 2706.315 3429.690 ;
        RECT 2706.625 3429.630 2706.855 3429.690 ;
        RECT 2706.085 3429.580 2706.855 3429.630 ;
        RECT 2712.265 3429.630 2712.495 3429.690 ;
        RECT 2712.805 3429.630 2713.035 3429.690 ;
        RECT 2718.445 3429.630 2718.675 3429.690 ;
        RECT 2718.985 3429.630 2719.215 3429.690 ;
        RECT 2712.265 3429.580 2713.035 3429.630 ;
        RECT 2718.435 3429.580 2719.215 3429.630 ;
        RECT 2724.625 3429.630 2724.855 3429.690 ;
        RECT 2725.165 3429.630 2725.395 3429.690 ;
        RECT 2724.625 3429.580 2725.395 3429.630 ;
        RECT 2730.805 3429.630 2731.035 3429.690 ;
        RECT 2731.345 3429.630 2731.575 3429.690 ;
        RECT 2736.985 3429.630 2737.215 3429.690 ;
        RECT 2737.525 3429.630 2737.755 3429.690 ;
        RECT 2730.805 3429.580 2731.585 3429.630 ;
        RECT 2736.985 3429.580 2737.755 3429.630 ;
        RECT 2743.165 3429.630 2743.395 3429.690 ;
        RECT 2743.705 3429.630 2743.935 3429.690 ;
        RECT 2749.345 3429.630 2749.575 3429.690 ;
        RECT 2749.885 3429.630 2750.115 3429.690 ;
        RECT 2743.165 3429.580 2743.935 3429.630 ;
        RECT 2749.335 3429.580 2750.115 3429.630 ;
        RECT 2755.525 3429.630 2755.755 3429.690 ;
        RECT 2756.065 3429.630 2756.295 3429.690 ;
        RECT 2755.525 3429.580 2756.295 3429.630 ;
        RECT 2761.705 3429.580 2769.255 3429.690 ;
        RECT 2693.435 3429.380 2769.255 3429.580 ;
        RECT 2693.435 3429.180 2700.735 3429.380 ;
        RECT 2706.085 3429.280 2706.855 3429.380 ;
        RECT 2706.085 3429.230 2706.315 3429.280 ;
        RECT 2706.625 3429.230 2706.855 3429.280 ;
        RECT 2712.265 3429.280 2713.035 3429.380 ;
        RECT 2718.435 3429.280 2719.215 3429.380 ;
        RECT 2712.265 3429.230 2712.495 3429.280 ;
        RECT 2712.805 3429.230 2713.035 3429.280 ;
        RECT 2718.445 3429.230 2718.675 3429.280 ;
        RECT 2718.985 3429.230 2719.215 3429.280 ;
        RECT 2724.625 3429.280 2725.395 3429.380 ;
        RECT 2724.625 3429.230 2724.855 3429.280 ;
        RECT 2725.165 3429.230 2725.395 3429.280 ;
        RECT 2730.805 3429.280 2731.585 3429.380 ;
        RECT 2736.985 3429.280 2737.755 3429.380 ;
        RECT 2730.805 3429.230 2731.035 3429.280 ;
        RECT 2731.345 3429.230 2731.575 3429.280 ;
        RECT 2736.985 3429.230 2737.215 3429.280 ;
        RECT 2737.525 3429.230 2737.755 3429.280 ;
        RECT 2743.165 3429.280 2743.935 3429.380 ;
        RECT 2749.335 3429.280 2750.115 3429.380 ;
        RECT 2743.165 3429.230 2743.395 3429.280 ;
        RECT 2743.705 3429.230 2743.935 3429.280 ;
        RECT 2749.345 3429.230 2749.575 3429.280 ;
        RECT 2749.885 3429.230 2750.115 3429.280 ;
        RECT 2755.525 3429.280 2756.295 3429.380 ;
        RECT 2755.525 3429.230 2755.755 3429.280 ;
        RECT 2756.065 3429.230 2756.295 3429.280 ;
        RECT 2761.705 3429.230 2769.255 3429.380 ;
        RECT 2693.435 3427.030 2696.110 3429.180 ;
        RECT 2766.585 3427.030 2769.255 3429.230 ;
        RECT 2693.435 3426.880 2700.685 3427.030 ;
        RECT 2761.735 3426.990 2769.255 3427.030 ;
        RECT 2706.085 3426.930 2706.315 3426.990 ;
        RECT 2706.625 3426.930 2706.855 3426.990 ;
        RECT 2706.085 3426.880 2706.855 3426.930 ;
        RECT 2712.265 3426.930 2712.495 3426.990 ;
        RECT 2712.805 3426.930 2713.035 3426.990 ;
        RECT 2718.445 3426.930 2718.675 3426.990 ;
        RECT 2718.985 3426.930 2719.215 3426.990 ;
        RECT 2712.265 3426.880 2713.035 3426.930 ;
        RECT 2718.435 3426.880 2719.215 3426.930 ;
        RECT 2724.625 3426.930 2724.855 3426.990 ;
        RECT 2725.165 3426.930 2725.395 3426.990 ;
        RECT 2724.625 3426.880 2725.395 3426.930 ;
        RECT 2730.805 3426.930 2731.035 3426.990 ;
        RECT 2731.345 3426.930 2731.575 3426.990 ;
        RECT 2736.985 3426.930 2737.215 3426.990 ;
        RECT 2737.525 3426.930 2737.755 3426.990 ;
        RECT 2730.805 3426.880 2731.585 3426.930 ;
        RECT 2736.985 3426.880 2737.755 3426.930 ;
        RECT 2743.165 3426.930 2743.395 3426.990 ;
        RECT 2743.705 3426.930 2743.935 3426.990 ;
        RECT 2749.345 3426.930 2749.575 3426.990 ;
        RECT 2749.885 3426.930 2750.115 3426.990 ;
        RECT 2743.165 3426.880 2743.935 3426.930 ;
        RECT 2749.335 3426.880 2750.115 3426.930 ;
        RECT 2755.525 3426.930 2755.755 3426.990 ;
        RECT 2756.065 3426.930 2756.295 3426.990 ;
        RECT 2755.525 3426.880 2756.295 3426.930 ;
        RECT 2761.705 3426.880 2769.255 3426.990 ;
        RECT 2693.435 3426.680 2769.255 3426.880 ;
        RECT 2693.435 3426.480 2700.685 3426.680 ;
        RECT 2706.085 3426.580 2706.855 3426.680 ;
        RECT 2706.085 3426.530 2706.315 3426.580 ;
        RECT 2706.625 3426.530 2706.855 3426.580 ;
        RECT 2712.265 3426.580 2713.035 3426.680 ;
        RECT 2718.435 3426.580 2719.215 3426.680 ;
        RECT 2712.265 3426.530 2712.495 3426.580 ;
        RECT 2712.805 3426.530 2713.035 3426.580 ;
        RECT 2718.445 3426.530 2718.675 3426.580 ;
        RECT 2718.985 3426.530 2719.215 3426.580 ;
        RECT 2724.625 3426.580 2725.395 3426.680 ;
        RECT 2724.625 3426.530 2724.855 3426.580 ;
        RECT 2725.165 3426.530 2725.395 3426.580 ;
        RECT 2730.805 3426.580 2731.585 3426.680 ;
        RECT 2736.985 3426.580 2737.755 3426.680 ;
        RECT 2730.805 3426.530 2731.035 3426.580 ;
        RECT 2731.345 3426.530 2731.575 3426.580 ;
        RECT 2736.985 3426.530 2737.215 3426.580 ;
        RECT 2737.525 3426.530 2737.755 3426.580 ;
        RECT 2743.165 3426.580 2743.935 3426.680 ;
        RECT 2749.335 3426.580 2750.115 3426.680 ;
        RECT 2743.165 3426.530 2743.395 3426.580 ;
        RECT 2743.705 3426.530 2743.935 3426.580 ;
        RECT 2749.345 3426.530 2749.575 3426.580 ;
        RECT 2749.885 3426.530 2750.115 3426.580 ;
        RECT 2755.525 3426.580 2756.295 3426.680 ;
        RECT 2755.525 3426.530 2755.755 3426.580 ;
        RECT 2756.065 3426.530 2756.295 3426.580 ;
        RECT 2761.705 3426.530 2769.255 3426.680 ;
        RECT 2693.435 3424.930 2696.110 3426.480 ;
        RECT 2766.585 3424.930 2769.255 3426.530 ;
        RECT 2694.065 3424.815 2696.110 3424.930 ;
        RECT 2767.210 3424.815 2769.255 3424.930 ;
        RECT 2778.785 3424.830 2781.410 3430.505 ;
        RECT 2779.365 3424.815 2781.410 3424.830 ;
        RECT 2712.285 3423.430 2713.035 3423.680 ;
        RECT 2718.885 3423.630 2719.385 3423.680 ;
        RECT 2718.435 3423.430 2719.385 3423.630 ;
        RECT 2720.035 3423.430 2721.185 3423.730 ;
        RECT 2730.985 3423.630 2731.485 3423.780 ;
        RECT 2724.635 3423.430 2725.385 3423.630 ;
        RECT 2730.835 3423.430 2731.585 3423.630 ;
        RECT 2732.085 3423.430 2733.235 3423.780 ;
        RECT 2736.985 3423.430 2737.735 3423.630 ;
        RECT 2743.135 3423.430 2743.935 3423.730 ;
        RECT 2744.385 3423.430 2745.535 3423.780 ;
        RECT 2749.335 3423.430 2750.085 3423.630 ;
        RECT 2710.485 3423.230 2752.135 3423.430 ;
        RECT 2710.535 3423.140 2715.535 3423.230 ;
        RECT 2716.625 3423.140 2721.625 3423.230 ;
        RECT 2722.715 3423.140 2727.715 3423.230 ;
        RECT 2728.805 3423.140 2733.805 3423.230 ;
        RECT 2734.895 3423.140 2739.895 3423.230 ;
        RECT 2740.985 3423.140 2745.985 3423.230 ;
        RECT 2747.075 3423.140 2752.075 3423.230 ;
        RECT 2710.535 3422.480 2715.535 3422.580 ;
        RECT 2716.625 3422.480 2721.625 3422.580 ;
        RECT 2722.715 3422.480 2727.715 3422.580 ;
        RECT 2728.805 3422.480 2733.805 3422.580 ;
        RECT 2734.895 3422.480 2739.895 3422.580 ;
        RECT 2740.985 3422.480 2745.985 3422.580 ;
        RECT 2747.075 3422.480 2752.075 3422.580 ;
        RECT 2710.485 3422.280 2752.135 3422.480 ;
        RECT 2711.985 3421.930 2713.235 3422.280 ;
        RECT 2724.935 3422.030 2725.435 3422.280 ;
        RECT 2737.035 3422.030 2738.285 3422.280 ;
        RECT 2712.035 3421.180 2713.185 3421.930 ;
        RECT 2711.985 3420.930 2713.235 3421.180 ;
        RECT 2718.885 3420.930 2719.385 3421.180 ;
        RECT 2730.985 3420.930 2731.485 3421.280 ;
        RECT 2737.085 3421.130 2738.235 3422.030 ;
        RECT 2749.335 3421.980 2749.835 3422.280 ;
        RECT 2737.035 3420.930 2738.285 3421.130 ;
        RECT 2743.135 3420.930 2743.635 3421.230 ;
        RECT 2710.485 3420.730 2752.135 3420.930 ;
        RECT 2710.535 3420.640 2715.535 3420.730 ;
        RECT 2716.625 3420.640 2721.625 3420.730 ;
        RECT 2722.715 3420.640 2727.715 3420.730 ;
        RECT 2728.805 3420.640 2733.805 3420.730 ;
        RECT 2734.895 3420.640 2739.895 3420.730 ;
        RECT 2740.985 3420.640 2745.985 3420.730 ;
        RECT 2747.075 3420.640 2752.075 3420.730 ;
        RECT 2710.535 3419.980 2715.535 3420.080 ;
        RECT 2716.625 3419.980 2721.625 3420.080 ;
        RECT 2722.715 3419.980 2727.715 3420.080 ;
        RECT 2728.805 3419.980 2733.805 3420.080 ;
        RECT 2734.895 3419.980 2739.895 3420.080 ;
        RECT 2740.985 3419.980 2745.985 3420.080 ;
        RECT 2747.075 3419.980 2752.075 3420.080 ;
        RECT 2710.485 3419.780 2752.135 3419.980 ;
        RECT 2712.685 3419.530 2713.185 3419.780 ;
        RECT 2713.635 3419.480 2714.135 3419.780 ;
        RECT 2714.385 3419.480 2714.885 3419.780 ;
        RECT 2718.435 3419.680 2719.185 3419.780 ;
        RECT 2724.635 3419.630 2725.435 3419.780 ;
        RECT 2724.935 3419.530 2725.435 3419.630 ;
        RECT 2726.085 3419.580 2726.585 3419.780 ;
        RECT 2726.835 3419.580 2727.335 3419.780 ;
        RECT 2730.835 3419.630 2731.585 3419.780 ;
        RECT 2737.135 3419.480 2737.635 3419.780 ;
        RECT 2738.485 3419.580 2738.985 3419.780 ;
        RECT 2739.185 3419.580 2739.685 3419.780 ;
        RECT 2743.185 3419.630 2743.935 3419.780 ;
        RECT 2749.335 3419.630 2750.085 3419.780 ;
        RECT 2749.335 3419.480 2749.835 3419.630 ;
        RECT 2712.945 3417.930 2713.175 3418.090 ;
        RECT 2718.495 3417.930 2718.725 3418.090 ;
        RECT 2719.035 3417.930 2719.265 3418.090 ;
        RECT 2724.585 3417.930 2724.815 3418.090 ;
        RECT 2725.125 3417.930 2725.355 3418.090 ;
        RECT 2730.675 3417.930 2730.905 3418.090 ;
        RECT 2731.215 3417.930 2731.445 3418.090 ;
        RECT 2736.765 3417.930 2736.995 3418.090 ;
        RECT 2737.305 3417.930 2737.535 3418.090 ;
        RECT 2742.855 3417.930 2743.085 3418.090 ;
        RECT 2743.395 3417.930 2743.625 3418.090 ;
        RECT 2748.945 3417.930 2749.175 3418.090 ;
        RECT 2712.885 3417.330 2749.175 3417.930 ;
        RECT 2712.945 3417.130 2713.175 3417.330 ;
        RECT 2718.495 3417.130 2718.725 3417.330 ;
        RECT 2719.035 3417.130 2719.265 3417.330 ;
        RECT 2724.585 3417.130 2724.815 3417.330 ;
        RECT 2725.125 3417.130 2725.355 3417.330 ;
        RECT 2730.675 3417.130 2730.905 3417.330 ;
        RECT 2731.215 3417.130 2731.445 3417.330 ;
        RECT 2736.765 3417.130 2736.995 3417.330 ;
        RECT 2737.305 3417.130 2737.535 3417.330 ;
        RECT 2742.855 3417.130 2743.085 3417.330 ;
        RECT 2743.395 3417.130 2743.625 3417.330 ;
        RECT 2748.945 3417.130 2749.175 3417.330 ;
        RECT 2712.945 3414.830 2713.175 3414.990 ;
        RECT 2718.495 3414.830 2718.725 3414.990 ;
        RECT 2719.035 3414.830 2719.265 3414.990 ;
        RECT 2724.585 3414.830 2724.815 3414.990 ;
        RECT 2725.125 3414.830 2725.355 3414.990 ;
        RECT 2730.675 3414.830 2730.905 3414.990 ;
        RECT 2731.215 3414.830 2731.445 3414.990 ;
        RECT 2736.765 3414.830 2736.995 3414.990 ;
        RECT 2737.305 3414.830 2737.535 3414.990 ;
        RECT 2742.855 3414.830 2743.085 3414.990 ;
        RECT 2743.395 3414.830 2743.625 3414.990 ;
        RECT 2748.945 3414.830 2749.175 3414.990 ;
        RECT 2712.945 3414.780 2749.185 3414.830 ;
        RECT 2712.785 3414.280 2749.185 3414.780 ;
        RECT 2712.945 3414.230 2749.185 3414.280 ;
        RECT 2712.945 3414.030 2713.175 3414.230 ;
        RECT 2718.495 3414.030 2718.725 3414.230 ;
        RECT 2719.035 3414.030 2719.265 3414.230 ;
        RECT 2724.585 3414.030 2724.815 3414.230 ;
        RECT 2725.125 3414.030 2725.355 3414.230 ;
        RECT 2730.675 3414.030 2730.905 3414.230 ;
        RECT 2731.215 3414.030 2731.445 3414.230 ;
        RECT 2736.765 3414.030 2736.995 3414.230 ;
        RECT 2737.305 3414.030 2737.535 3414.230 ;
        RECT 2742.855 3414.030 2743.085 3414.230 ;
        RECT 2743.395 3414.030 2743.625 3414.230 ;
        RECT 2748.945 3414.030 2749.175 3414.230 ;
        RECT 2710.145 3411.830 2710.375 3411.990 ;
        RECT 2715.695 3411.830 2715.925 3411.990 ;
        RECT 2716.235 3411.830 2716.465 3411.990 ;
        RECT 2721.785 3411.830 2722.015 3411.990 ;
        RECT 2722.325 3411.830 2722.555 3411.990 ;
        RECT 2727.875 3411.830 2728.105 3411.990 ;
        RECT 2728.415 3411.830 2728.645 3411.990 ;
        RECT 2733.965 3411.830 2734.195 3411.990 ;
        RECT 2734.505 3411.830 2734.735 3411.990 ;
        RECT 2740.055 3411.830 2740.285 3411.990 ;
        RECT 2740.595 3411.830 2740.825 3411.990 ;
        RECT 2746.145 3411.830 2746.375 3411.990 ;
        RECT 2746.685 3411.830 2746.915 3411.990 ;
        RECT 2752.235 3411.830 2752.465 3411.990 ;
        RECT 2710.085 3411.230 2752.485 3411.830 ;
        RECT 2710.145 3411.030 2710.375 3411.230 ;
        RECT 2715.695 3411.030 2715.925 3411.230 ;
        RECT 2716.235 3411.030 2716.465 3411.230 ;
        RECT 2721.785 3411.030 2722.015 3411.230 ;
        RECT 2722.325 3411.030 2722.555 3411.230 ;
        RECT 2727.875 3411.030 2728.105 3411.230 ;
        RECT 2728.415 3411.030 2728.645 3411.230 ;
        RECT 2733.965 3411.030 2734.195 3411.230 ;
        RECT 2734.505 3411.030 2734.735 3411.230 ;
        RECT 2740.055 3411.030 2740.285 3411.230 ;
        RECT 2740.595 3411.030 2740.825 3411.230 ;
        RECT 2746.145 3411.030 2746.375 3411.230 ;
        RECT 2746.685 3411.030 2746.915 3411.230 ;
        RECT 2752.235 3411.030 2752.465 3411.230 ;
        RECT 2710.535 3410.830 2715.535 3410.980 ;
        RECT 2716.625 3410.830 2721.625 3410.980 ;
        RECT 2722.715 3410.830 2727.715 3410.980 ;
        RECT 2728.805 3410.830 2733.805 3410.980 ;
        RECT 2734.895 3410.830 2739.895 3410.980 ;
        RECT 2740.985 3410.830 2745.985 3410.980 ;
        RECT 2747.075 3410.830 2752.075 3410.980 ;
        RECT 2710.485 3410.630 2752.085 3410.830 ;
        RECT 2711.985 3410.530 2712.535 3410.630 ;
        RECT 2712.685 3410.530 2713.235 3410.630 ;
        RECT 2737.035 3410.530 2737.585 3410.630 ;
        RECT 2737.735 3410.530 2738.285 3410.630 ;
        RECT 2710.145 3408.830 2710.375 3408.990 ;
        RECT 2715.695 3408.830 2715.925 3408.990 ;
        RECT 2716.235 3408.830 2716.465 3408.990 ;
        RECT 2721.785 3408.830 2722.015 3408.990 ;
        RECT 2722.325 3408.830 2722.555 3408.990 ;
        RECT 2727.875 3408.830 2728.105 3408.990 ;
        RECT 2728.415 3408.830 2728.645 3408.990 ;
        RECT 2733.965 3408.830 2734.195 3408.990 ;
        RECT 2734.505 3408.830 2734.735 3408.990 ;
        RECT 2740.055 3408.830 2740.285 3408.990 ;
        RECT 2740.595 3408.830 2740.825 3408.990 ;
        RECT 2746.145 3408.830 2746.375 3408.990 ;
        RECT 2746.685 3408.830 2746.915 3408.990 ;
        RECT 2752.235 3408.830 2752.465 3408.990 ;
        RECT 2710.145 3408.230 2752.485 3408.830 ;
        RECT 2710.145 3408.030 2710.375 3408.230 ;
        RECT 2715.695 3408.030 2715.925 3408.230 ;
        RECT 2716.235 3408.030 2716.465 3408.230 ;
        RECT 2721.785 3408.030 2722.015 3408.230 ;
        RECT 2722.325 3408.030 2722.555 3408.230 ;
        RECT 2727.875 3408.030 2728.105 3408.230 ;
        RECT 2728.415 3408.030 2728.645 3408.230 ;
        RECT 2733.965 3408.030 2734.195 3408.230 ;
        RECT 2734.505 3408.030 2734.735 3408.230 ;
        RECT 2740.055 3408.030 2740.285 3408.230 ;
        RECT 2740.595 3408.030 2740.825 3408.230 ;
        RECT 2746.145 3408.030 2746.375 3408.230 ;
        RECT 2746.685 3408.030 2746.915 3408.230 ;
        RECT 2752.235 3408.030 2752.465 3408.230 ;
        RECT 2710.535 3407.830 2715.535 3407.980 ;
        RECT 2716.625 3407.830 2721.625 3407.980 ;
        RECT 2722.715 3407.830 2727.715 3407.980 ;
        RECT 2728.805 3407.830 2733.805 3407.980 ;
        RECT 2734.895 3407.830 2739.895 3407.980 ;
        RECT 2740.985 3407.830 2745.985 3407.980 ;
        RECT 2747.075 3407.830 2752.075 3407.980 ;
        RECT 2710.485 3407.630 2752.085 3407.830 ;
        RECT 2711.985 3407.430 2712.535 3407.630 ;
        RECT 2712.685 3407.430 2713.235 3407.630 ;
        RECT 2737.035 3407.530 2737.585 3407.630 ;
        RECT 2737.735 3407.530 2738.285 3407.630 ;
        RECT 2712.870 3403.860 2713.100 3404.120 ;
        RECT 2718.510 3403.860 2718.740 3404.120 ;
        RECT 2719.050 3403.860 2719.280 3404.120 ;
        RECT 2724.690 3403.860 2724.920 3404.120 ;
        RECT 2725.230 3403.860 2725.460 3404.120 ;
        RECT 2730.870 3403.860 2731.100 3404.120 ;
        RECT 2731.410 3403.860 2731.640 3404.120 ;
        RECT 2737.050 3403.860 2737.280 3404.120 ;
        RECT 2737.590 3403.860 2737.820 3404.120 ;
        RECT 2743.230 3403.860 2743.460 3404.120 ;
        RECT 2743.770 3403.860 2744.000 3404.120 ;
        RECT 2749.410 3403.860 2749.640 3404.120 ;
        RECT 2712.870 3403.160 2749.640 3403.860 ;
        RECT 2712.870 3402.800 2749.610 3403.160 ;
        RECT 2712.870 3400.910 2713.100 3401.170 ;
        RECT 2718.510 3400.910 2718.740 3401.170 ;
        RECT 2719.050 3400.910 2719.280 3401.170 ;
        RECT 2724.690 3400.910 2724.920 3401.170 ;
        RECT 2725.230 3400.910 2725.460 3401.170 ;
        RECT 2730.870 3400.910 2731.100 3401.170 ;
        RECT 2731.410 3400.910 2731.640 3401.170 ;
        RECT 2737.050 3400.910 2737.280 3401.170 ;
        RECT 2737.590 3400.910 2737.820 3401.170 ;
        RECT 2743.230 3400.910 2743.460 3401.170 ;
        RECT 2743.770 3400.910 2744.000 3401.170 ;
        RECT 2749.410 3400.910 2749.640 3401.170 ;
        RECT 2712.860 3400.460 2749.640 3400.910 ;
        RECT 2712.870 3400.210 2713.100 3400.460 ;
        RECT 2718.510 3400.210 2718.740 3400.460 ;
        RECT 2719.050 3400.210 2719.280 3400.460 ;
        RECT 2724.690 3400.210 2724.920 3400.460 ;
        RECT 2725.230 3400.210 2725.460 3400.460 ;
        RECT 2730.870 3400.210 2731.100 3400.460 ;
        RECT 2731.410 3400.210 2731.640 3400.460 ;
        RECT 2737.050 3400.210 2737.280 3400.460 ;
        RECT 2737.590 3400.210 2737.820 3400.460 ;
        RECT 2743.230 3400.210 2743.460 3400.460 ;
        RECT 2743.770 3400.210 2744.000 3400.460 ;
        RECT 2749.410 3400.210 2749.640 3400.460 ;
        RECT 2713.260 3400.060 2718.305 3400.160 ;
        RECT 2719.485 3400.060 2724.485 3400.160 ;
        RECT 2725.665 3400.060 2730.665 3400.160 ;
        RECT 2731.845 3400.060 2736.845 3400.160 ;
        RECT 2738.025 3400.060 2743.025 3400.160 ;
        RECT 2744.205 3400.060 2749.230 3400.160 ;
        RECT 2713.260 3399.660 2749.230 3400.060 ;
        RECT 2730.240 3397.610 2732.140 3397.650 ;
        RECT 2726.660 3397.220 2735.760 3397.610 ;
        RECT 2726.660 3396.860 2735.770 3397.220 ;
        RECT 2726.720 3396.460 2735.770 3396.860 ;
        RECT 2726.720 3396.260 2726.950 3396.460 ;
        RECT 2728.510 3396.260 2729.310 3396.460 ;
        RECT 2730.860 3396.260 2731.635 3396.460 ;
        RECT 2733.200 3396.260 2733.985 3396.460 ;
        RECT 2735.540 3396.260 2735.770 3396.460 ;
        RECT 2738.460 3394.660 2740.210 3394.760 ;
        RECT 2722.560 3393.760 2740.210 3394.660 ;
        RECT 2722.560 3393.610 2724.210 3393.760 ;
        RECT 2727.820 3393.635 2728.050 3393.760 ;
        RECT 2730.870 3393.635 2731.100 3393.760 ;
        RECT 2731.410 3393.635 2731.640 3393.760 ;
        RECT 2734.460 3393.635 2734.690 3393.760 ;
        RECT 2728.210 3393.485 2730.710 3393.585 ;
        RECT 2731.800 3393.485 2734.300 3393.585 ;
        RECT 2728.185 3393.410 2734.360 3393.485 ;
        RECT 2728.160 3393.060 2734.410 3393.410 ;
        RECT 2713.510 3391.750 2748.960 3391.985 ;
        RECT 2713.510 3391.610 2748.985 3391.750 ;
        RECT 2713.535 3391.520 2718.535 3391.610 ;
        RECT 2719.625 3391.520 2724.625 3391.610 ;
        RECT 2725.715 3391.520 2730.715 3391.610 ;
        RECT 2731.805 3391.520 2736.805 3391.610 ;
        RECT 2737.895 3391.520 2742.895 3391.610 ;
        RECT 2743.985 3391.520 2748.985 3391.610 ;
        RECT 2713.145 3391.235 2713.375 3391.470 ;
        RECT 2718.695 3391.235 2718.925 3391.470 ;
        RECT 2719.235 3391.235 2719.465 3391.470 ;
        RECT 2724.785 3391.235 2725.015 3391.470 ;
        RECT 2725.325 3391.235 2725.555 3391.470 ;
        RECT 2730.875 3391.235 2731.105 3391.470 ;
        RECT 2731.415 3391.235 2731.645 3391.470 ;
        RECT 2736.965 3391.235 2737.195 3391.470 ;
        RECT 2737.505 3391.235 2737.735 3391.470 ;
        RECT 2743.055 3391.235 2743.285 3391.470 ;
        RECT 2743.595 3391.235 2743.825 3391.470 ;
        RECT 2749.145 3391.235 2749.375 3391.470 ;
        RECT 2713.145 3390.810 2749.375 3391.235 ;
        RECT 2713.145 3390.510 2713.375 3390.810 ;
        RECT 2718.695 3390.510 2718.925 3390.810 ;
        RECT 2719.235 3390.510 2719.465 3390.810 ;
        RECT 2724.785 3390.510 2725.015 3390.810 ;
        RECT 2725.325 3390.510 2725.555 3390.810 ;
        RECT 2730.875 3390.510 2731.105 3390.810 ;
        RECT 2731.415 3390.510 2731.645 3390.810 ;
        RECT 2736.965 3390.510 2737.195 3390.810 ;
        RECT 2737.505 3390.510 2737.735 3390.810 ;
        RECT 2743.055 3390.510 2743.285 3390.810 ;
        RECT 2743.595 3390.510 2743.825 3390.810 ;
        RECT 2749.145 3390.510 2749.375 3390.810 ;
        RECT 2713.535 3390.360 2718.535 3390.460 ;
        RECT 2719.625 3390.360 2724.625 3390.460 ;
        RECT 2725.715 3390.360 2730.715 3390.460 ;
        RECT 2731.805 3390.360 2736.805 3390.460 ;
        RECT 2737.895 3390.360 2742.895 3390.460 ;
        RECT 2743.985 3390.360 2748.985 3390.460 ;
        RECT 2713.510 3390.230 2748.985 3390.360 ;
        RECT 2713.510 3389.985 2748.960 3390.230 ;
        RECT 2720.260 3388.510 2722.260 3389.985 ;
        RECT 2727.260 3388.510 2729.260 3389.985 ;
        RECT 2733.760 3388.510 2735.760 3389.985 ;
        RECT 2740.210 3388.510 2742.260 3389.985 ;
        RECT 2716.260 3385.510 2746.260 3388.510 ;
      LAYER via ;
        RECT 2713.755 3451.100 2714.015 3451.360 ;
        RECT 2714.505 3451.100 2714.765 3451.360 ;
        RECT 2715.370 3451.325 2715.630 3451.585 ;
        RECT 2715.690 3451.325 2715.950 3451.585 ;
        RECT 2721.570 3451.325 2721.830 3451.585 ;
        RECT 2721.890 3451.325 2722.150 3451.585 ;
        RECT 2726.205 3451.100 2726.465 3451.360 ;
        RECT 2726.955 3451.100 2727.215 3451.360 ;
        RECT 2727.720 3451.325 2727.980 3451.585 ;
        RECT 2728.040 3451.325 2728.300 3451.585 ;
        RECT 2733.920 3451.325 2734.180 3451.585 ;
        RECT 2734.240 3451.325 2734.500 3451.585 ;
        RECT 2738.605 3451.100 2738.865 3451.360 ;
        RECT 2739.355 3451.100 2739.615 3451.360 ;
        RECT 2740.120 3451.325 2740.380 3451.585 ;
        RECT 2740.440 3451.325 2740.700 3451.585 ;
        RECT 2746.270 3451.325 2746.530 3451.585 ;
        RECT 2746.590 3451.325 2746.850 3451.585 ;
        RECT 2711.805 3450.750 2712.065 3451.010 ;
        RECT 2712.655 3450.750 2712.915 3451.010 ;
        RECT 2724.405 3450.750 2724.665 3451.010 ;
        RECT 2725.255 3450.750 2725.515 3451.010 ;
        RECT 2736.855 3450.750 2737.115 3451.010 ;
        RECT 2737.705 3450.750 2737.965 3451.010 ;
        RECT 2749.105 3450.750 2749.365 3451.010 ;
        RECT 2749.955 3450.750 2750.215 3451.010 ;
        RECT 2713.755 3448.400 2714.015 3448.660 ;
        RECT 2714.505 3448.400 2714.765 3448.660 ;
        RECT 2715.370 3448.625 2715.630 3448.885 ;
        RECT 2715.690 3448.625 2715.950 3448.885 ;
        RECT 2721.570 3448.625 2721.830 3448.885 ;
        RECT 2721.890 3448.625 2722.150 3448.885 ;
        RECT 2726.205 3448.400 2726.465 3448.660 ;
        RECT 2726.955 3448.400 2727.215 3448.660 ;
        RECT 2727.720 3448.625 2727.980 3448.885 ;
        RECT 2728.040 3448.625 2728.300 3448.885 ;
        RECT 2733.920 3448.625 2734.180 3448.885 ;
        RECT 2734.240 3448.625 2734.500 3448.885 ;
        RECT 2738.605 3448.400 2738.865 3448.660 ;
        RECT 2739.355 3448.400 2739.615 3448.660 ;
        RECT 2740.120 3448.625 2740.380 3448.885 ;
        RECT 2740.440 3448.625 2740.700 3448.885 ;
        RECT 2746.270 3448.625 2746.530 3448.885 ;
        RECT 2746.590 3448.625 2746.850 3448.885 ;
        RECT 2711.805 3448.050 2712.065 3448.310 ;
        RECT 2712.655 3448.050 2712.915 3448.310 ;
        RECT 2724.405 3448.050 2724.665 3448.310 ;
        RECT 2725.255 3448.050 2725.515 3448.310 ;
        RECT 2736.855 3448.050 2737.115 3448.310 ;
        RECT 2737.705 3448.050 2737.965 3448.310 ;
        RECT 2749.105 3448.000 2749.365 3448.260 ;
        RECT 2749.955 3448.000 2750.215 3448.260 ;
        RECT 2713.755 3445.700 2714.015 3445.960 ;
        RECT 2714.505 3445.700 2714.765 3445.960 ;
        RECT 2715.370 3445.925 2715.630 3446.185 ;
        RECT 2715.690 3445.925 2715.950 3446.185 ;
        RECT 2721.570 3445.925 2721.830 3446.185 ;
        RECT 2721.890 3445.925 2722.150 3446.185 ;
        RECT 2726.205 3445.700 2726.465 3445.960 ;
        RECT 2726.955 3445.700 2727.215 3445.960 ;
        RECT 2727.720 3445.925 2727.980 3446.185 ;
        RECT 2728.040 3445.925 2728.300 3446.185 ;
        RECT 2733.920 3445.925 2734.180 3446.185 ;
        RECT 2734.240 3445.925 2734.500 3446.185 ;
        RECT 2738.655 3445.700 2738.915 3445.960 ;
        RECT 2739.355 3445.700 2739.615 3445.960 ;
        RECT 2740.120 3445.925 2740.380 3446.185 ;
        RECT 2740.440 3445.925 2740.700 3446.185 ;
        RECT 2746.270 3445.925 2746.530 3446.185 ;
        RECT 2746.590 3445.925 2746.850 3446.185 ;
        RECT 2711.805 3445.350 2712.065 3445.610 ;
        RECT 2712.655 3445.350 2712.915 3445.610 ;
        RECT 2724.405 3445.350 2724.665 3445.610 ;
        RECT 2725.255 3445.350 2725.515 3445.610 ;
        RECT 2736.855 3445.300 2737.115 3445.560 ;
        RECT 2737.705 3445.300 2737.965 3445.560 ;
        RECT 2749.105 3445.350 2749.365 3445.610 ;
        RECT 2749.955 3445.350 2750.215 3445.610 ;
        RECT 2715.370 3443.225 2715.630 3443.485 ;
        RECT 2715.690 3443.225 2715.950 3443.485 ;
        RECT 2721.570 3443.225 2721.830 3443.485 ;
        RECT 2721.890 3443.225 2722.150 3443.485 ;
        RECT 2727.720 3443.225 2727.980 3443.485 ;
        RECT 2728.040 3443.225 2728.300 3443.485 ;
        RECT 2733.920 3443.225 2734.180 3443.485 ;
        RECT 2734.240 3443.225 2734.500 3443.485 ;
        RECT 2740.070 3443.225 2740.330 3443.485 ;
        RECT 2740.390 3443.225 2740.650 3443.485 ;
        RECT 2746.270 3443.225 2746.530 3443.485 ;
        RECT 2746.590 3443.225 2746.850 3443.485 ;
        RECT 2711.805 3442.650 2712.065 3442.910 ;
        RECT 2712.655 3442.650 2712.915 3442.910 ;
        RECT 2720.205 3442.700 2720.465 3442.960 ;
        RECT 2720.755 3442.700 2721.015 3442.960 ;
        RECT 2724.355 3442.650 2724.615 3442.910 ;
        RECT 2725.205 3442.650 2725.465 3442.910 ;
        RECT 2732.255 3442.700 2732.515 3442.960 ;
        RECT 2732.805 3442.700 2733.065 3442.960 ;
        RECT 2736.805 3442.650 2737.065 3442.910 ;
        RECT 2737.655 3442.650 2737.915 3442.910 ;
        RECT 2744.555 3442.650 2744.815 3442.910 ;
        RECT 2745.105 3442.650 2745.365 3442.910 ;
        RECT 2749.255 3442.650 2749.515 3442.910 ;
        RECT 2750.105 3442.650 2750.365 3442.910 ;
        RECT 2715.370 3440.325 2715.630 3440.585 ;
        RECT 2715.690 3440.325 2715.950 3440.585 ;
        RECT 2721.570 3440.325 2721.830 3440.585 ;
        RECT 2721.890 3440.325 2722.150 3440.585 ;
        RECT 2727.770 3440.325 2728.030 3440.585 ;
        RECT 2728.090 3440.325 2728.350 3440.585 ;
        RECT 2733.920 3440.325 2734.180 3440.585 ;
        RECT 2734.240 3440.325 2734.500 3440.585 ;
        RECT 2740.070 3440.325 2740.330 3440.585 ;
        RECT 2740.390 3440.325 2740.650 3440.585 ;
        RECT 2746.270 3440.325 2746.530 3440.585 ;
        RECT 2746.590 3440.325 2746.850 3440.585 ;
        RECT 2711.805 3439.750 2712.065 3440.010 ;
        RECT 2712.655 3439.750 2712.915 3440.010 ;
        RECT 2720.205 3439.650 2720.465 3439.910 ;
        RECT 2720.755 3439.650 2721.015 3439.910 ;
        RECT 2724.355 3439.750 2724.615 3440.010 ;
        RECT 2725.205 3439.750 2725.465 3440.010 ;
        RECT 2732.255 3439.750 2732.515 3440.010 ;
        RECT 2732.805 3439.750 2733.065 3440.010 ;
        RECT 2736.805 3439.700 2737.065 3439.960 ;
        RECT 2737.655 3439.700 2737.915 3439.960 ;
        RECT 2744.555 3439.750 2744.815 3440.010 ;
        RECT 2745.105 3439.750 2745.365 3440.010 ;
        RECT 2749.255 3439.750 2749.515 3440.010 ;
        RECT 2750.105 3439.750 2750.365 3440.010 ;
        RECT 2681.420 3438.040 2682.000 3438.620 ;
        RECT 2682.670 3438.040 2683.250 3438.620 ;
        RECT 2778.920 3438.890 2779.500 3439.470 ;
        RECT 2780.220 3438.890 2780.800 3439.470 ;
        RECT 2715.370 3437.425 2715.630 3437.685 ;
        RECT 2715.690 3437.425 2715.950 3437.685 ;
        RECT 2721.570 3437.425 2721.830 3437.685 ;
        RECT 2721.890 3437.425 2722.150 3437.685 ;
        RECT 2727.720 3437.425 2727.980 3437.685 ;
        RECT 2728.040 3437.425 2728.300 3437.685 ;
        RECT 2733.920 3437.425 2734.180 3437.685 ;
        RECT 2734.240 3437.425 2734.500 3437.685 ;
        RECT 2740.070 3437.425 2740.330 3437.685 ;
        RECT 2740.390 3437.425 2740.650 3437.685 ;
        RECT 2746.270 3437.425 2746.530 3437.685 ;
        RECT 2746.590 3437.425 2746.850 3437.685 ;
        RECT 2711.705 3436.700 2711.965 3436.960 ;
        RECT 2712.755 3436.700 2713.015 3436.960 ;
        RECT 2724.355 3436.850 2724.615 3437.110 ;
        RECT 2725.205 3436.850 2725.465 3437.110 ;
        RECT 2732.255 3436.850 2732.515 3437.110 ;
        RECT 2732.805 3436.850 2733.065 3437.110 ;
        RECT 2736.805 3436.850 2737.065 3437.110 ;
        RECT 2737.655 3436.850 2737.915 3437.110 ;
        RECT 2744.555 3436.850 2744.815 3437.110 ;
        RECT 2745.105 3436.850 2745.365 3437.110 ;
        RECT 2749.255 3436.850 2749.515 3437.110 ;
        RECT 2750.105 3436.850 2750.365 3437.110 ;
        RECT 2706.170 3434.725 2706.430 3434.985 ;
        RECT 2706.490 3434.725 2706.750 3434.985 ;
        RECT 2712.370 3434.725 2712.630 3434.985 ;
        RECT 2712.690 3434.725 2712.950 3434.985 ;
        RECT 2718.520 3434.725 2718.780 3434.985 ;
        RECT 2718.840 3434.725 2719.100 3434.985 ;
        RECT 2724.720 3434.725 2724.980 3434.985 ;
        RECT 2725.040 3434.725 2725.300 3434.985 ;
        RECT 2730.920 3434.725 2731.180 3434.985 ;
        RECT 2731.240 3434.725 2731.500 3434.985 ;
        RECT 2737.070 3434.725 2737.330 3434.985 ;
        RECT 2737.390 3434.725 2737.650 3434.985 ;
        RECT 2743.270 3434.725 2743.530 3434.985 ;
        RECT 2743.590 3434.725 2743.850 3434.985 ;
        RECT 2749.420 3434.725 2749.680 3434.985 ;
        RECT 2749.740 3434.725 2750.000 3434.985 ;
        RECT 2755.620 3434.725 2755.880 3434.985 ;
        RECT 2755.940 3434.725 2756.200 3434.985 ;
        RECT 2706.170 3432.075 2706.430 3432.335 ;
        RECT 2706.490 3432.075 2706.750 3432.335 ;
        RECT 2712.370 3432.025 2712.630 3432.285 ;
        RECT 2712.690 3432.025 2712.950 3432.285 ;
        RECT 2718.520 3432.025 2718.780 3432.285 ;
        RECT 2718.840 3432.025 2719.100 3432.285 ;
        RECT 2724.720 3432.025 2724.980 3432.285 ;
        RECT 2725.040 3432.025 2725.300 3432.285 ;
        RECT 2730.920 3432.025 2731.180 3432.285 ;
        RECT 2731.240 3432.025 2731.500 3432.285 ;
        RECT 2737.070 3432.025 2737.330 3432.285 ;
        RECT 2737.390 3432.025 2737.650 3432.285 ;
        RECT 2743.270 3432.025 2743.530 3432.285 ;
        RECT 2743.590 3432.025 2743.850 3432.285 ;
        RECT 2749.420 3432.025 2749.680 3432.285 ;
        RECT 2749.740 3432.025 2750.000 3432.285 ;
        RECT 2755.620 3432.025 2755.880 3432.285 ;
        RECT 2755.940 3432.025 2756.200 3432.285 ;
        RECT 2706.170 3429.325 2706.430 3429.585 ;
        RECT 2706.490 3429.325 2706.750 3429.585 ;
        RECT 2712.370 3429.325 2712.630 3429.585 ;
        RECT 2712.690 3429.325 2712.950 3429.585 ;
        RECT 2718.520 3429.325 2718.780 3429.585 ;
        RECT 2718.840 3429.325 2719.100 3429.585 ;
        RECT 2724.720 3429.325 2724.980 3429.585 ;
        RECT 2725.040 3429.325 2725.300 3429.585 ;
        RECT 2730.920 3429.325 2731.180 3429.585 ;
        RECT 2731.240 3429.325 2731.500 3429.585 ;
        RECT 2737.070 3429.325 2737.330 3429.585 ;
        RECT 2737.390 3429.325 2737.650 3429.585 ;
        RECT 2743.270 3429.325 2743.530 3429.585 ;
        RECT 2743.590 3429.325 2743.850 3429.585 ;
        RECT 2749.420 3429.325 2749.680 3429.585 ;
        RECT 2749.740 3429.325 2750.000 3429.585 ;
        RECT 2755.620 3429.325 2755.880 3429.585 ;
        RECT 2755.940 3429.325 2756.200 3429.585 ;
        RECT 2706.170 3426.625 2706.430 3426.885 ;
        RECT 2706.490 3426.625 2706.750 3426.885 ;
        RECT 2712.370 3426.625 2712.630 3426.885 ;
        RECT 2712.690 3426.625 2712.950 3426.885 ;
        RECT 2718.520 3426.625 2718.780 3426.885 ;
        RECT 2718.840 3426.625 2719.100 3426.885 ;
        RECT 2724.720 3426.625 2724.980 3426.885 ;
        RECT 2725.040 3426.625 2725.300 3426.885 ;
        RECT 2730.920 3426.625 2731.180 3426.885 ;
        RECT 2731.240 3426.625 2731.500 3426.885 ;
        RECT 2737.070 3426.625 2737.330 3426.885 ;
        RECT 2737.390 3426.625 2737.650 3426.885 ;
        RECT 2743.270 3426.625 2743.530 3426.885 ;
        RECT 2743.590 3426.625 2743.850 3426.885 ;
        RECT 2749.420 3426.625 2749.680 3426.885 ;
        RECT 2749.740 3426.625 2750.000 3426.885 ;
        RECT 2755.620 3426.625 2755.880 3426.885 ;
        RECT 2755.940 3426.625 2756.200 3426.885 ;
        RECT 2712.370 3423.375 2712.630 3423.635 ;
        RECT 2712.690 3423.375 2712.950 3423.635 ;
        RECT 2718.520 3423.325 2718.780 3423.585 ;
        RECT 2718.840 3423.325 2719.100 3423.585 ;
        RECT 2720.205 3423.350 2720.465 3423.610 ;
        RECT 2720.755 3423.350 2721.015 3423.610 ;
        RECT 2724.720 3423.325 2724.980 3423.585 ;
        RECT 2725.040 3423.325 2725.300 3423.585 ;
        RECT 2730.920 3423.325 2731.180 3423.585 ;
        RECT 2731.240 3423.325 2731.500 3423.585 ;
        RECT 2732.255 3423.350 2732.515 3423.610 ;
        RECT 2732.805 3423.350 2733.065 3423.610 ;
        RECT 2737.070 3423.325 2737.330 3423.585 ;
        RECT 2737.390 3423.325 2737.650 3423.585 ;
        RECT 2743.270 3423.425 2743.530 3423.685 ;
        RECT 2743.590 3423.425 2743.850 3423.685 ;
        RECT 2744.555 3423.400 2744.815 3423.660 ;
        RECT 2745.105 3423.400 2745.365 3423.660 ;
        RECT 2749.420 3423.325 2749.680 3423.585 ;
        RECT 2749.740 3423.325 2750.000 3423.585 ;
        RECT 2712.130 3422.000 2712.390 3422.260 ;
        RECT 2712.830 3422.000 2713.090 3422.260 ;
        RECT 2737.180 3422.100 2737.440 3422.360 ;
        RECT 2737.880 3422.100 2738.140 3422.360 ;
        RECT 2712.130 3420.850 2712.390 3421.110 ;
        RECT 2712.830 3420.850 2713.090 3421.110 ;
        RECT 2737.180 3420.800 2737.440 3421.060 ;
        RECT 2737.880 3420.800 2738.140 3421.060 ;
        RECT 2713.755 3419.550 2714.015 3419.810 ;
        RECT 2714.505 3419.550 2714.765 3419.810 ;
        RECT 2726.205 3419.650 2726.465 3419.910 ;
        RECT 2726.955 3419.650 2727.215 3419.910 ;
        RECT 2738.605 3419.650 2738.865 3419.910 ;
        RECT 2739.305 3419.650 2739.565 3419.910 ;
        RECT 2721.905 3417.500 2722.165 3417.760 ;
        RECT 2733.955 3417.500 2734.215 3417.760 ;
        RECT 2718.880 3414.400 2719.140 3414.660 ;
        RECT 2719.480 3414.400 2719.740 3414.660 ;
        RECT 2721.905 3414.400 2722.165 3414.660 ;
        RECT 2731.130 3414.400 2731.390 3414.660 ;
        RECT 2731.730 3414.400 2731.990 3414.660 ;
        RECT 2733.955 3414.400 2734.215 3414.660 ;
        RECT 2743.280 3414.400 2743.540 3414.660 ;
        RECT 2743.880 3414.400 2744.140 3414.660 ;
        RECT 2718.880 3411.400 2719.140 3411.660 ;
        RECT 2719.480 3411.400 2719.740 3411.660 ;
        RECT 2731.130 3411.400 2731.390 3411.660 ;
        RECT 2731.730 3411.400 2731.990 3411.660 ;
        RECT 2743.280 3411.400 2743.540 3411.660 ;
        RECT 2743.880 3411.400 2744.140 3411.660 ;
        RECT 2712.130 3410.600 2712.390 3410.860 ;
        RECT 2712.830 3410.600 2713.090 3410.860 ;
        RECT 2737.180 3410.600 2737.440 3410.860 ;
        RECT 2737.880 3410.600 2738.140 3410.860 ;
        RECT 2718.880 3408.400 2719.140 3408.660 ;
        RECT 2719.480 3408.400 2719.740 3408.660 ;
        RECT 2730.430 3408.395 2730.690 3408.655 ;
        RECT 2731.130 3408.400 2731.390 3408.660 ;
        RECT 2731.730 3408.400 2731.990 3408.660 ;
        RECT 2743.280 3408.400 2743.540 3408.660 ;
        RECT 2743.880 3408.400 2744.140 3408.660 ;
        RECT 2712.130 3407.500 2712.390 3407.760 ;
        RECT 2712.830 3407.500 2713.090 3407.760 ;
        RECT 2737.180 3407.600 2737.440 3407.860 ;
        RECT 2737.880 3407.600 2738.140 3407.860 ;
        RECT 2722.705 3403.505 2722.965 3403.765 ;
        RECT 2723.805 3403.505 2724.065 3403.765 ;
        RECT 2738.605 3403.505 2738.865 3403.765 ;
        RECT 2739.805 3403.505 2740.065 3403.765 ;
        RECT 2722.705 3400.555 2722.965 3400.815 ;
        RECT 2723.805 3400.555 2724.065 3400.815 ;
        RECT 2738.605 3400.555 2738.865 3400.815 ;
        RECT 2739.805 3400.555 2740.065 3400.815 ;
        RECT 2728.505 3399.755 2728.765 3400.015 ;
        RECT 2729.055 3399.755 2729.315 3400.015 ;
        RECT 2733.205 3399.755 2733.465 3400.015 ;
        RECT 2733.755 3399.755 2734.015 3400.015 ;
        RECT 2730.310 3397.370 2730.570 3397.630 ;
        RECT 2730.810 3397.370 2731.070 3397.630 ;
        RECT 2731.310 3397.370 2731.570 3397.630 ;
        RECT 2731.810 3397.370 2732.070 3397.630 ;
        RECT 2728.505 3396.905 2728.765 3397.165 ;
        RECT 2729.055 3396.905 2729.315 3397.165 ;
        RECT 2733.205 3396.955 2733.465 3397.215 ;
        RECT 2733.755 3396.955 2734.015 3397.215 ;
        RECT 2722.705 3394.255 2722.965 3394.515 ;
        RECT 2723.755 3394.255 2724.015 3394.515 ;
        RECT 2738.605 3394.355 2738.865 3394.615 ;
        RECT 2739.805 3394.355 2740.065 3394.615 ;
        RECT 2722.705 3393.805 2722.965 3394.065 ;
        RECT 2723.755 3393.805 2724.015 3394.065 ;
        RECT 2738.605 3393.905 2738.865 3394.165 ;
        RECT 2739.805 3393.905 2740.065 3394.165 ;
        RECT 2728.505 3393.155 2728.765 3393.415 ;
        RECT 2729.055 3393.155 2729.315 3393.415 ;
        RECT 2733.205 3393.155 2733.465 3393.415 ;
        RECT 2733.755 3393.155 2734.015 3393.415 ;
        RECT 2722.705 3391.655 2722.965 3391.915 ;
        RECT 2723.805 3391.655 2724.065 3391.915 ;
        RECT 2738.605 3391.655 2738.865 3391.915 ;
        RECT 2739.805 3391.655 2740.065 3391.915 ;
        RECT 2728.505 3390.905 2728.765 3391.165 ;
        RECT 2729.055 3390.905 2729.315 3391.165 ;
        RECT 2733.205 3390.905 2733.465 3391.165 ;
        RECT 2733.755 3390.905 2734.015 3391.165 ;
      LAYER met2 ;
        RECT 2711.635 3445.180 2713.085 3451.680 ;
        RECT 2713.685 3450.980 2714.085 3451.480 ;
        RECT 2714.435 3450.980 2714.835 3451.480 ;
        RECT 2713.685 3448.280 2714.085 3448.780 ;
        RECT 2714.435 3448.280 2714.835 3448.780 ;
        RECT 2713.685 3445.580 2714.085 3446.080 ;
        RECT 2714.435 3445.580 2714.835 3446.080 ;
        RECT 2681.385 3437.930 2682.035 3438.730 ;
        RECT 2682.635 3437.930 2683.285 3438.730 ;
        RECT 2711.635 3436.630 2713.085 3443.130 ;
        RECT 2715.285 3437.180 2716.035 3451.880 ;
        RECT 2720.135 3442.580 2720.535 3443.080 ;
        RECT 2720.685 3442.580 2721.085 3443.080 ;
        RECT 2720.135 3439.530 2720.535 3440.030 ;
        RECT 2720.685 3439.530 2721.085 3440.030 ;
        RECT 2720.035 3436.780 2721.185 3437.230 ;
        RECT 2721.485 3436.980 2722.235 3451.930 ;
        RECT 2724.235 3445.130 2725.685 3452.080 ;
        RECT 2726.135 3450.980 2726.535 3451.480 ;
        RECT 2726.885 3450.980 2727.285 3451.480 ;
        RECT 2726.135 3448.280 2726.535 3448.780 ;
        RECT 2726.885 3448.280 2727.285 3448.780 ;
        RECT 2726.135 3445.580 2726.535 3446.080 ;
        RECT 2726.885 3445.580 2727.285 3446.080 ;
        RECT 2711.635 3436.580 2712.035 3436.630 ;
        RECT 2712.685 3436.580 2713.085 3436.630 ;
        RECT 2724.145 3436.490 2725.805 3443.230 ;
        RECT 2727.635 3437.230 2728.385 3451.880 ;
        RECT 2732.185 3442.580 2732.585 3443.080 ;
        RECT 2732.735 3442.580 2733.135 3443.080 ;
        RECT 2732.185 3439.630 2732.585 3440.130 ;
        RECT 2732.735 3439.630 2733.135 3440.130 ;
        RECT 2733.835 3437.230 2734.585 3451.880 ;
        RECT 2736.685 3445.130 2738.135 3452.080 ;
        RECT 2738.535 3450.980 2738.935 3451.480 ;
        RECT 2739.285 3450.980 2739.685 3451.480 ;
        RECT 2740.035 3450.180 2740.785 3451.830 ;
        RECT 2738.535 3448.280 2738.935 3448.780 ;
        RECT 2739.285 3448.280 2739.685 3448.780 ;
        RECT 2738.585 3445.580 2738.985 3446.080 ;
        RECT 2739.285 3445.580 2739.685 3446.080 ;
        RECT 2739.985 3445.680 2740.785 3450.180 ;
        RECT 2732.185 3436.730 2732.585 3437.230 ;
        RECT 2732.735 3436.730 2733.135 3437.230 ;
        RECT 2736.635 3436.680 2738.085 3443.180 ;
        RECT 2739.985 3437.180 2740.735 3445.680 ;
        RECT 2744.485 3442.530 2744.885 3443.030 ;
        RECT 2745.035 3442.530 2745.435 3443.030 ;
        RECT 2744.485 3439.630 2744.885 3440.130 ;
        RECT 2745.035 3439.630 2745.435 3440.130 ;
        RECT 2746.185 3437.230 2746.935 3451.780 ;
        RECT 2748.935 3445.230 2750.385 3452.430 ;
        RECT 2744.485 3436.730 2744.885 3437.230 ;
        RECT 2745.035 3436.730 2745.435 3437.230 ;
        RECT 2749.085 3436.680 2750.535 3443.430 ;
        RECT 2778.885 3438.780 2779.535 3439.580 ;
        RECT 2780.185 3438.780 2780.835 3439.580 ;
        RECT 2706.085 3426.380 2706.835 3435.180 ;
        RECT 2712.285 3423.280 2713.035 3435.230 ;
        RECT 2718.435 3423.030 2719.185 3435.180 ;
        RECT 2720.135 3423.230 2720.535 3423.730 ;
        RECT 2720.685 3423.230 2721.085 3423.730 ;
        RECT 2724.635 3422.830 2725.385 3435.180 ;
        RECT 2730.835 3422.930 2731.585 3435.130 ;
        RECT 2732.185 3423.230 2732.585 3423.730 ;
        RECT 2732.735 3423.230 2733.135 3423.730 ;
        RECT 2736.985 3423.230 2737.735 3435.180 ;
        RECT 2743.185 3423.080 2743.935 3435.280 ;
        RECT 2744.485 3423.280 2744.885 3423.780 ;
        RECT 2745.035 3423.280 2745.435 3423.780 ;
        RECT 2749.335 3423.080 2750.085 3435.230 ;
        RECT 2755.535 3426.430 2756.285 3435.230 ;
        RECT 2737.085 3422.430 2737.535 3422.480 ;
        RECT 2737.785 3422.430 2738.235 3422.480 ;
        RECT 2712.035 3422.280 2712.485 3422.380 ;
        RECT 2712.735 3422.280 2713.185 3422.380 ;
        RECT 2712.035 3407.380 2713.185 3422.280 ;
        RECT 2713.585 3419.480 2714.935 3419.930 ;
        RECT 2726.135 3419.530 2726.535 3420.030 ;
        RECT 2726.885 3419.530 2727.285 3420.030 ;
        RECT 2713.685 3419.430 2714.085 3419.480 ;
        RECT 2714.435 3419.430 2714.835 3419.480 ;
        RECT 2718.785 3408.280 2719.835 3414.830 ;
        RECT 2721.835 3414.280 2722.235 3417.980 ;
        RECT 2731.035 3409.000 2732.085 3414.830 ;
        RECT 2733.885 3414.280 2734.285 3417.980 ;
        RECT 2722.560 3391.560 2724.210 3403.810 ;
        RECT 2728.360 3390.510 2729.460 3400.110 ;
        RECT 2730.190 3397.250 2732.190 3409.000 ;
        RECT 2737.085 3407.480 2738.235 3422.430 ;
        RECT 2738.535 3419.530 2738.935 3420.030 ;
        RECT 2739.235 3419.530 2739.635 3420.030 ;
        RECT 2743.185 3408.280 2744.235 3414.830 ;
        RECT 2733.060 3390.560 2734.160 3400.160 ;
        RECT 2738.460 3391.460 2740.210 3403.860 ;
      LAYER via2 ;
        RECT 2713.745 3451.090 2714.025 3451.370 ;
        RECT 2714.495 3451.090 2714.775 3451.370 ;
        RECT 2713.745 3448.390 2714.025 3448.670 ;
        RECT 2714.495 3448.390 2714.775 3448.670 ;
        RECT 2713.745 3445.690 2714.025 3445.970 ;
        RECT 2714.495 3445.690 2714.775 3445.970 ;
        RECT 2681.570 3438.390 2681.850 3438.670 ;
        RECT 2681.570 3437.990 2681.850 3438.270 ;
        RECT 2682.820 3438.390 2683.100 3438.670 ;
        RECT 2682.820 3437.990 2683.100 3438.270 ;
        RECT 2720.195 3442.690 2720.475 3442.970 ;
        RECT 2720.745 3442.690 2721.025 3442.970 ;
        RECT 2720.195 3439.640 2720.475 3439.920 ;
        RECT 2720.745 3439.640 2721.025 3439.920 ;
        RECT 2726.195 3451.090 2726.475 3451.370 ;
        RECT 2726.945 3451.090 2727.225 3451.370 ;
        RECT 2726.195 3448.390 2726.475 3448.670 ;
        RECT 2726.945 3448.390 2727.225 3448.670 ;
        RECT 2726.195 3445.690 2726.475 3445.970 ;
        RECT 2726.945 3445.690 2727.225 3445.970 ;
        RECT 2732.245 3442.690 2732.525 3442.970 ;
        RECT 2732.795 3442.690 2733.075 3442.970 ;
        RECT 2732.245 3439.740 2732.525 3440.020 ;
        RECT 2732.795 3439.740 2733.075 3440.020 ;
        RECT 2738.595 3451.090 2738.875 3451.370 ;
        RECT 2739.345 3451.090 2739.625 3451.370 ;
        RECT 2738.595 3448.390 2738.875 3448.670 ;
        RECT 2739.345 3448.390 2739.625 3448.670 ;
        RECT 2738.645 3445.690 2738.925 3445.970 ;
        RECT 2739.345 3445.690 2739.625 3445.970 ;
        RECT 2732.245 3436.840 2732.525 3437.120 ;
        RECT 2732.795 3436.840 2733.075 3437.120 ;
        RECT 2744.545 3442.640 2744.825 3442.920 ;
        RECT 2745.095 3442.640 2745.375 3442.920 ;
        RECT 2744.545 3439.740 2744.825 3440.020 ;
        RECT 2745.095 3439.740 2745.375 3440.020 ;
        RECT 2744.545 3436.840 2744.825 3437.120 ;
        RECT 2745.095 3436.840 2745.375 3437.120 ;
        RECT 2779.070 3439.240 2779.350 3439.520 ;
        RECT 2779.070 3438.840 2779.350 3439.120 ;
        RECT 2780.370 3439.240 2780.650 3439.520 ;
        RECT 2780.370 3438.840 2780.650 3439.120 ;
        RECT 2720.195 3423.340 2720.475 3423.620 ;
        RECT 2720.745 3423.340 2721.025 3423.620 ;
        RECT 2732.245 3423.340 2732.525 3423.620 ;
        RECT 2732.795 3423.340 2733.075 3423.620 ;
        RECT 2744.545 3423.390 2744.825 3423.670 ;
        RECT 2745.095 3423.390 2745.375 3423.670 ;
        RECT 2713.745 3419.540 2714.025 3419.820 ;
        RECT 2714.495 3419.540 2714.775 3419.820 ;
        RECT 2726.195 3419.640 2726.475 3419.920 ;
        RECT 2726.945 3419.640 2727.225 3419.920 ;
        RECT 2738.595 3419.640 2738.875 3419.920 ;
        RECT 2739.295 3419.640 2739.575 3419.920 ;
      LAYER met3 ;
        RECT 2681.285 3437.880 2683.485 3473.230 ;
        RECT 2694.085 3455.230 2711.085 3472.725 ;
        RECT 2713.085 3455.230 2730.085 3472.725 ;
        RECT 2732.085 3455.230 2749.085 3472.725 ;
        RECT 2751.085 3455.230 2768.085 3472.725 ;
        RECT 2713.585 3450.930 2714.935 3451.530 ;
        RECT 2726.035 3450.930 2727.385 3451.480 ;
        RECT 2738.435 3450.930 2739.785 3451.530 ;
        RECT 2713.585 3448.230 2714.935 3448.830 ;
        RECT 2726.035 3448.230 2727.385 3448.780 ;
        RECT 2738.435 3448.230 2739.785 3448.830 ;
        RECT 2713.585 3445.530 2714.935 3446.180 ;
        RECT 2726.035 3445.530 2727.385 3446.080 ;
        RECT 2738.435 3445.530 2739.785 3446.180 ;
        RECT 2720.035 3442.480 2721.185 3443.130 ;
        RECT 2732.085 3442.580 2733.235 3443.130 ;
        RECT 2744.385 3442.480 2745.535 3443.030 ;
        RECT 2720.035 3439.530 2721.185 3440.030 ;
        RECT 2732.085 3439.580 2733.235 3440.130 ;
        RECT 2744.385 3439.580 2745.535 3440.130 ;
        RECT 2778.785 3438.780 2780.935 3473.280 ;
        RECT 2720.035 3436.680 2721.185 3437.280 ;
        RECT 2732.085 3436.680 2733.235 3437.230 ;
        RECT 2744.385 3436.680 2745.535 3437.230 ;
        RECT 2720.035 3423.230 2721.185 3423.730 ;
        RECT 2732.085 3423.230 2733.235 3423.780 ;
        RECT 2744.385 3423.280 2745.535 3423.780 ;
        RECT 2713.585 3419.330 2714.935 3419.980 ;
        RECT 2726.035 3419.480 2727.385 3420.030 ;
        RECT 2738.435 3419.480 2739.785 3420.030 ;
      LAYER via3 ;
        RECT 2681.525 3472.495 2681.845 3472.815 ;
        RECT 2682.825 3472.495 2683.145 3472.815 ;
        RECT 2694.225 3472.305 2694.545 3472.625 ;
        RECT 2694.625 3472.305 2694.945 3472.625 ;
        RECT 2695.025 3472.305 2695.345 3472.625 ;
        RECT 2695.425 3472.305 2695.745 3472.625 ;
        RECT 2695.825 3472.305 2696.145 3472.625 ;
        RECT 2696.225 3472.305 2696.545 3472.625 ;
        RECT 2696.625 3472.305 2696.945 3472.625 ;
        RECT 2697.025 3472.305 2697.345 3472.625 ;
        RECT 2697.425 3472.305 2697.745 3472.625 ;
        RECT 2697.825 3472.305 2698.145 3472.625 ;
        RECT 2698.225 3472.305 2698.545 3472.625 ;
        RECT 2698.625 3472.305 2698.945 3472.625 ;
        RECT 2699.025 3472.305 2699.345 3472.625 ;
        RECT 2699.425 3472.305 2699.745 3472.625 ;
        RECT 2699.825 3472.305 2700.145 3472.625 ;
        RECT 2700.225 3472.305 2700.545 3472.625 ;
        RECT 2700.625 3472.305 2700.945 3472.625 ;
        RECT 2701.025 3472.305 2701.345 3472.625 ;
        RECT 2701.425 3472.305 2701.745 3472.625 ;
        RECT 2701.825 3472.305 2702.145 3472.625 ;
        RECT 2702.225 3472.305 2702.545 3472.625 ;
        RECT 2702.625 3472.305 2702.945 3472.625 ;
        RECT 2703.025 3472.305 2703.345 3472.625 ;
        RECT 2703.425 3472.305 2703.745 3472.625 ;
        RECT 2703.825 3472.305 2704.145 3472.625 ;
        RECT 2704.225 3472.305 2704.545 3472.625 ;
        RECT 2704.625 3472.305 2704.945 3472.625 ;
        RECT 2705.025 3472.305 2705.345 3472.625 ;
        RECT 2705.425 3472.305 2705.745 3472.625 ;
        RECT 2705.825 3472.305 2706.145 3472.625 ;
        RECT 2706.225 3472.305 2706.545 3472.625 ;
        RECT 2706.625 3472.305 2706.945 3472.625 ;
        RECT 2707.025 3472.305 2707.345 3472.625 ;
        RECT 2707.425 3472.305 2707.745 3472.625 ;
        RECT 2707.825 3472.305 2708.145 3472.625 ;
        RECT 2708.225 3472.305 2708.545 3472.625 ;
        RECT 2708.625 3472.305 2708.945 3472.625 ;
        RECT 2709.025 3472.305 2709.345 3472.625 ;
        RECT 2709.425 3472.305 2709.745 3472.625 ;
        RECT 2709.825 3472.305 2710.145 3472.625 ;
        RECT 2710.225 3472.305 2710.545 3472.625 ;
        RECT 2710.625 3472.305 2710.945 3472.625 ;
        RECT 2713.225 3472.305 2713.545 3472.625 ;
        RECT 2713.625 3472.305 2713.945 3472.625 ;
        RECT 2714.025 3472.305 2714.345 3472.625 ;
        RECT 2714.425 3472.305 2714.745 3472.625 ;
        RECT 2714.825 3472.305 2715.145 3472.625 ;
        RECT 2715.225 3472.305 2715.545 3472.625 ;
        RECT 2715.625 3472.305 2715.945 3472.625 ;
        RECT 2716.025 3472.305 2716.345 3472.625 ;
        RECT 2716.425 3472.305 2716.745 3472.625 ;
        RECT 2716.825 3472.305 2717.145 3472.625 ;
        RECT 2717.225 3472.305 2717.545 3472.625 ;
        RECT 2717.625 3472.305 2717.945 3472.625 ;
        RECT 2718.025 3472.305 2718.345 3472.625 ;
        RECT 2718.425 3472.305 2718.745 3472.625 ;
        RECT 2718.825 3472.305 2719.145 3472.625 ;
        RECT 2719.225 3472.305 2719.545 3472.625 ;
        RECT 2719.625 3472.305 2719.945 3472.625 ;
        RECT 2720.025 3472.305 2720.345 3472.625 ;
        RECT 2720.425 3472.305 2720.745 3472.625 ;
        RECT 2720.825 3472.305 2721.145 3472.625 ;
        RECT 2721.225 3472.305 2721.545 3472.625 ;
        RECT 2721.625 3472.305 2721.945 3472.625 ;
        RECT 2722.025 3472.305 2722.345 3472.625 ;
        RECT 2722.425 3472.305 2722.745 3472.625 ;
        RECT 2722.825 3472.305 2723.145 3472.625 ;
        RECT 2723.225 3472.305 2723.545 3472.625 ;
        RECT 2723.625 3472.305 2723.945 3472.625 ;
        RECT 2724.025 3472.305 2724.345 3472.625 ;
        RECT 2724.425 3472.305 2724.745 3472.625 ;
        RECT 2724.825 3472.305 2725.145 3472.625 ;
        RECT 2725.225 3472.305 2725.545 3472.625 ;
        RECT 2725.625 3472.305 2725.945 3472.625 ;
        RECT 2726.025 3472.305 2726.345 3472.625 ;
        RECT 2726.425 3472.305 2726.745 3472.625 ;
        RECT 2726.825 3472.305 2727.145 3472.625 ;
        RECT 2727.225 3472.305 2727.545 3472.625 ;
        RECT 2727.625 3472.305 2727.945 3472.625 ;
        RECT 2728.025 3472.305 2728.345 3472.625 ;
        RECT 2728.425 3472.305 2728.745 3472.625 ;
        RECT 2728.825 3472.305 2729.145 3472.625 ;
        RECT 2729.225 3472.305 2729.545 3472.625 ;
        RECT 2729.625 3472.305 2729.945 3472.625 ;
        RECT 2732.225 3472.305 2732.545 3472.625 ;
        RECT 2732.625 3472.305 2732.945 3472.625 ;
        RECT 2733.025 3472.305 2733.345 3472.625 ;
        RECT 2733.425 3472.305 2733.745 3472.625 ;
        RECT 2733.825 3472.305 2734.145 3472.625 ;
        RECT 2734.225 3472.305 2734.545 3472.625 ;
        RECT 2734.625 3472.305 2734.945 3472.625 ;
        RECT 2735.025 3472.305 2735.345 3472.625 ;
        RECT 2735.425 3472.305 2735.745 3472.625 ;
        RECT 2735.825 3472.305 2736.145 3472.625 ;
        RECT 2736.225 3472.305 2736.545 3472.625 ;
        RECT 2736.625 3472.305 2736.945 3472.625 ;
        RECT 2737.025 3472.305 2737.345 3472.625 ;
        RECT 2737.425 3472.305 2737.745 3472.625 ;
        RECT 2737.825 3472.305 2738.145 3472.625 ;
        RECT 2738.225 3472.305 2738.545 3472.625 ;
        RECT 2738.625 3472.305 2738.945 3472.625 ;
        RECT 2739.025 3472.305 2739.345 3472.625 ;
        RECT 2739.425 3472.305 2739.745 3472.625 ;
        RECT 2739.825 3472.305 2740.145 3472.625 ;
        RECT 2740.225 3472.305 2740.545 3472.625 ;
        RECT 2740.625 3472.305 2740.945 3472.625 ;
        RECT 2741.025 3472.305 2741.345 3472.625 ;
        RECT 2741.425 3472.305 2741.745 3472.625 ;
        RECT 2741.825 3472.305 2742.145 3472.625 ;
        RECT 2742.225 3472.305 2742.545 3472.625 ;
        RECT 2742.625 3472.305 2742.945 3472.625 ;
        RECT 2743.025 3472.305 2743.345 3472.625 ;
        RECT 2743.425 3472.305 2743.745 3472.625 ;
        RECT 2743.825 3472.305 2744.145 3472.625 ;
        RECT 2744.225 3472.305 2744.545 3472.625 ;
        RECT 2744.625 3472.305 2744.945 3472.625 ;
        RECT 2745.025 3472.305 2745.345 3472.625 ;
        RECT 2745.425 3472.305 2745.745 3472.625 ;
        RECT 2745.825 3472.305 2746.145 3472.625 ;
        RECT 2746.225 3472.305 2746.545 3472.625 ;
        RECT 2746.625 3472.305 2746.945 3472.625 ;
        RECT 2747.025 3472.305 2747.345 3472.625 ;
        RECT 2747.425 3472.305 2747.745 3472.625 ;
        RECT 2747.825 3472.305 2748.145 3472.625 ;
        RECT 2748.225 3472.305 2748.545 3472.625 ;
        RECT 2748.625 3472.305 2748.945 3472.625 ;
        RECT 2751.225 3472.305 2751.545 3472.625 ;
        RECT 2751.625 3472.305 2751.945 3472.625 ;
        RECT 2752.025 3472.305 2752.345 3472.625 ;
        RECT 2752.425 3472.305 2752.745 3472.625 ;
        RECT 2752.825 3472.305 2753.145 3472.625 ;
        RECT 2753.225 3472.305 2753.545 3472.625 ;
        RECT 2753.625 3472.305 2753.945 3472.625 ;
        RECT 2754.025 3472.305 2754.345 3472.625 ;
        RECT 2754.425 3472.305 2754.745 3472.625 ;
        RECT 2754.825 3472.305 2755.145 3472.625 ;
        RECT 2755.225 3472.305 2755.545 3472.625 ;
        RECT 2755.625 3472.305 2755.945 3472.625 ;
        RECT 2756.025 3472.305 2756.345 3472.625 ;
        RECT 2756.425 3472.305 2756.745 3472.625 ;
        RECT 2756.825 3472.305 2757.145 3472.625 ;
        RECT 2757.225 3472.305 2757.545 3472.625 ;
        RECT 2757.625 3472.305 2757.945 3472.625 ;
        RECT 2758.025 3472.305 2758.345 3472.625 ;
        RECT 2758.425 3472.305 2758.745 3472.625 ;
        RECT 2758.825 3472.305 2759.145 3472.625 ;
        RECT 2759.225 3472.305 2759.545 3472.625 ;
        RECT 2759.625 3472.305 2759.945 3472.625 ;
        RECT 2760.025 3472.305 2760.345 3472.625 ;
        RECT 2760.425 3472.305 2760.745 3472.625 ;
        RECT 2760.825 3472.305 2761.145 3472.625 ;
        RECT 2761.225 3472.305 2761.545 3472.625 ;
        RECT 2761.625 3472.305 2761.945 3472.625 ;
        RECT 2762.025 3472.305 2762.345 3472.625 ;
        RECT 2762.425 3472.305 2762.745 3472.625 ;
        RECT 2762.825 3472.305 2763.145 3472.625 ;
        RECT 2763.225 3472.305 2763.545 3472.625 ;
        RECT 2763.625 3472.305 2763.945 3472.625 ;
        RECT 2764.025 3472.305 2764.345 3472.625 ;
        RECT 2764.425 3472.305 2764.745 3472.625 ;
        RECT 2764.825 3472.305 2765.145 3472.625 ;
        RECT 2765.225 3472.305 2765.545 3472.625 ;
        RECT 2765.625 3472.305 2765.945 3472.625 ;
        RECT 2766.025 3472.305 2766.345 3472.625 ;
        RECT 2766.425 3472.305 2766.745 3472.625 ;
        RECT 2766.825 3472.305 2767.145 3472.625 ;
        RECT 2767.225 3472.305 2767.545 3472.625 ;
        RECT 2767.625 3472.305 2767.945 3472.625 ;
        RECT 2779.000 3472.495 2779.320 3472.815 ;
        RECT 2780.300 3472.495 2780.620 3472.815 ;
        RECT 2713.725 3451.070 2714.045 3451.390 ;
        RECT 2714.475 3451.070 2714.795 3451.390 ;
        RECT 2726.175 3451.070 2726.495 3451.390 ;
        RECT 2726.925 3451.070 2727.245 3451.390 ;
        RECT 2738.575 3451.070 2738.895 3451.390 ;
        RECT 2739.325 3451.070 2739.645 3451.390 ;
        RECT 2713.725 3448.370 2714.045 3448.690 ;
        RECT 2714.475 3448.370 2714.795 3448.690 ;
        RECT 2726.175 3448.370 2726.495 3448.690 ;
        RECT 2726.925 3448.370 2727.245 3448.690 ;
        RECT 2738.575 3448.370 2738.895 3448.690 ;
        RECT 2739.325 3448.370 2739.645 3448.690 ;
        RECT 2713.725 3445.670 2714.045 3445.990 ;
        RECT 2714.475 3445.670 2714.795 3445.990 ;
        RECT 2726.175 3445.670 2726.495 3445.990 ;
        RECT 2726.925 3445.670 2727.245 3445.990 ;
        RECT 2738.625 3445.670 2738.945 3445.990 ;
        RECT 2739.325 3445.670 2739.645 3445.990 ;
        RECT 2720.175 3442.670 2720.495 3442.990 ;
        RECT 2720.725 3442.670 2721.045 3442.990 ;
        RECT 2732.225 3442.670 2732.545 3442.990 ;
        RECT 2732.775 3442.670 2733.095 3442.990 ;
        RECT 2744.525 3442.620 2744.845 3442.940 ;
        RECT 2745.075 3442.620 2745.395 3442.940 ;
        RECT 2720.175 3439.620 2720.495 3439.940 ;
        RECT 2720.725 3439.620 2721.045 3439.940 ;
        RECT 2732.225 3439.720 2732.545 3440.040 ;
        RECT 2732.775 3439.720 2733.095 3440.040 ;
        RECT 2744.525 3439.720 2744.845 3440.040 ;
        RECT 2745.075 3439.720 2745.395 3440.040 ;
        RECT 2720.175 3436.820 2720.495 3437.140 ;
        RECT 2720.725 3436.820 2721.045 3437.140 ;
        RECT 2732.225 3436.820 2732.545 3437.140 ;
        RECT 2732.775 3436.820 2733.095 3437.140 ;
        RECT 2744.525 3436.820 2744.845 3437.140 ;
        RECT 2745.075 3436.820 2745.395 3437.140 ;
        RECT 2720.175 3423.320 2720.495 3423.640 ;
        RECT 2720.725 3423.320 2721.045 3423.640 ;
        RECT 2732.225 3423.320 2732.545 3423.640 ;
        RECT 2732.775 3423.320 2733.095 3423.640 ;
        RECT 2744.525 3423.370 2744.845 3423.690 ;
        RECT 2745.075 3423.370 2745.395 3423.690 ;
        RECT 2713.725 3419.520 2714.045 3419.840 ;
        RECT 2714.475 3419.520 2714.795 3419.840 ;
        RECT 2726.175 3419.620 2726.495 3419.940 ;
        RECT 2726.925 3419.620 2727.245 3419.940 ;
        RECT 2738.575 3419.620 2738.895 3419.940 ;
        RECT 2739.275 3419.620 2739.595 3419.940 ;
      LAYER met4 ;
        RECT 2681.235 3472.080 2780.935 3473.280 ;
        RECT 2713.585 3419.330 2714.935 3452.080 ;
        RECT 2720.035 3423.180 2721.185 3443.130 ;
        RECT 2726.035 3419.480 2727.385 3452.330 ;
        RECT 2732.085 3423.180 2733.235 3443.130 ;
        RECT 2738.435 3419.480 2739.785 3452.380 ;
        RECT 2744.385 3423.230 2745.535 3443.180 ;
  END
END MULT_AMPLIFIER
END LIBRARY

