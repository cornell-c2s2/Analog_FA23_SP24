magic
tech sky130A
timestamp 1709331665
<< metal1 >>
rect 280110 343500 285830 343550
rect 280110 343300 283250 343500
rect 283450 343300 283650 343500
rect 283850 343300 284050 343500
rect 284250 343300 284450 343500
rect 284650 343300 284850 343500
rect 285050 343300 285250 343500
rect 285450 343300 285830 343500
rect 280110 343100 285830 343300
rect 280110 342900 283250 343100
rect 283450 342900 283650 343100
rect 283850 342900 284050 343100
rect 284250 342900 284450 343100
rect 284650 342900 284850 343100
rect 285050 342900 285250 343100
rect 285450 342900 285830 343100
rect 280110 342830 285830 342900
rect 280110 342350 280540 342830
rect 275250 342320 280540 342350
rect 275230 342250 280540 342320
rect 275250 342150 280540 342250
rect 275230 342000 281000 342070
rect 275320 341850 280500 342000
rect 280650 341850 280800 342000
rect 280950 341850 281000 342000
rect 275320 341800 281000 341850
rect 280060 341750 281000 341800
rect 280060 341600 280500 341750
rect 280650 341600 280800 341750
rect 280950 341600 281000 341750
rect 280060 341500 281000 341600
rect 280060 341350 280500 341500
rect 280650 341350 280800 341500
rect 280950 341350 281000 341500
rect 280060 341250 281000 341350
rect 280060 341100 280500 341250
rect 280650 341100 280800 341250
rect 280950 341100 281000 341250
rect 280060 341000 281000 341100
rect 280060 340850 280500 341000
rect 280650 340850 280800 341000
rect 280950 340850 281000 341000
rect 280060 340750 281000 340850
rect 280060 340600 280500 340750
rect 280650 340600 280800 340750
rect 280950 340600 281000 340750
rect 280060 340500 281000 340600
rect 280060 340350 280500 340500
rect 280650 340350 280800 340500
rect 280950 340350 281000 340500
rect 280060 340250 281000 340350
rect 280060 340100 280500 340250
rect 280650 340100 280800 340250
rect 280950 340100 281000 340250
rect 280060 340000 281000 340100
rect 280060 339850 280500 340000
rect 280650 339850 280800 340000
rect 280950 339850 281000 340000
rect 280060 339750 281000 339850
rect 280060 339600 280500 339750
rect 280650 339600 280800 339750
rect 280950 339600 281000 339750
rect 280060 339500 281000 339600
rect 280060 339350 280500 339500
rect 280650 339350 280800 339500
rect 280950 339350 281000 339500
rect 280060 339250 281000 339350
rect 280060 339100 280500 339250
rect 280650 339100 280800 339250
rect 280950 339100 281000 339250
rect 280060 338950 281000 339100
<< via1 >>
rect 283250 343300 283450 343500
rect 283650 343300 283850 343500
rect 284050 343300 284250 343500
rect 284450 343300 284650 343500
rect 284850 343300 285050 343500
rect 285250 343300 285450 343500
rect 283250 342900 283450 343100
rect 283650 342900 283850 343100
rect 284050 342900 284250 343100
rect 284450 342900 284650 343100
rect 284850 342900 285050 343100
rect 285250 342900 285450 343100
rect 280500 341850 280650 342000
rect 280800 341850 280950 342000
rect 280500 341600 280650 341750
rect 280800 341600 280950 341750
rect 280500 341350 280650 341500
rect 280800 341350 280950 341500
rect 280500 341100 280650 341250
rect 280800 341100 280950 341250
rect 280500 340850 280650 341000
rect 280800 340850 280950 341000
rect 280500 340600 280650 340750
rect 280800 340600 280950 340750
rect 280500 340350 280650 340500
rect 280800 340350 280950 340500
rect 280500 340100 280650 340250
rect 280800 340100 280950 340250
rect 280500 339850 280650 340000
rect 280800 339850 280950 340000
rect 280500 339600 280650 339750
rect 280800 339600 280950 339750
rect 280500 339350 280650 339500
rect 280800 339350 280950 339500
rect 280500 339100 280650 339250
rect 280800 339100 280950 339250
<< metal2 >>
rect 283250 343500 283450 343505
rect 283250 343295 283450 343300
rect 283650 343500 283850 343505
rect 283650 343295 283850 343300
rect 284050 343500 284250 343505
rect 284050 343295 284250 343300
rect 284450 343500 284650 343505
rect 284450 343295 284650 343300
rect 284850 343500 285050 343505
rect 284850 343295 285050 343300
rect 285250 343500 285450 343505
rect 285250 343295 285450 343300
rect 283250 343100 283450 343105
rect 283250 342895 283450 342900
rect 283650 343100 283850 343105
rect 283650 342895 283850 342900
rect 284050 343100 284250 343105
rect 284050 342895 284250 342900
rect 284450 343100 284650 343105
rect 284450 342895 284650 342900
rect 284850 343100 285050 343105
rect 284850 342895 285050 342900
rect 285250 343100 285450 343105
rect 285250 342895 285450 342900
rect 280500 342000 280650 342005
rect 280500 341845 280650 341850
rect 280800 342000 280950 342005
rect 280800 341845 280950 341850
rect 280500 341750 280650 341755
rect 280500 341595 280650 341600
rect 280800 341750 280950 341755
rect 280800 341595 280950 341600
rect 280500 341500 280650 341505
rect 280500 341345 280650 341350
rect 280800 341500 280950 341505
rect 280800 341345 280950 341350
rect 280500 341250 280650 341255
rect 280500 341095 280650 341100
rect 280800 341250 280950 341255
rect 280800 341095 280950 341100
rect 280500 341000 280650 341005
rect 280500 340845 280650 340850
rect 280800 341000 280950 341005
rect 280800 340845 280950 340850
rect 280500 340750 280650 340755
rect 280500 340595 280650 340600
rect 280800 340750 280950 340755
rect 280800 340595 280950 340600
rect 280500 340500 280650 340505
rect 280500 340345 280650 340350
rect 280800 340500 280950 340505
rect 280800 340345 280950 340350
rect 280500 340250 280650 340255
rect 280500 340095 280650 340100
rect 280800 340250 280950 340255
rect 280800 340095 280950 340100
rect 280500 340000 280650 340005
rect 280500 339845 280650 339850
rect 280800 340000 280950 340005
rect 280800 339845 280950 339850
rect 280500 339750 280650 339755
rect 280500 339595 280650 339600
rect 280800 339750 280950 339755
rect 280800 339595 280950 339600
rect 280500 339500 280650 339505
rect 280500 339345 280650 339350
rect 280800 339500 280950 339505
rect 280800 339345 280950 339350
rect 280500 339250 280650 339255
rect 280500 339095 280650 339100
rect 280800 339250 280950 339255
rect 280800 339095 280950 339100
<< via2 >>
rect 283250 343300 283450 343500
rect 283650 343300 283850 343500
rect 284050 343300 284250 343500
rect 284450 343300 284650 343500
rect 284850 343300 285050 343500
rect 285250 343300 285450 343500
rect 283250 342900 283450 343100
rect 283650 342900 283850 343100
rect 284050 342900 284250 343100
rect 284450 342900 284650 343100
rect 284850 342900 285050 343100
rect 285250 342900 285450 343100
rect 280500 341850 280650 342000
rect 280800 341850 280950 342000
rect 280500 341600 280650 341750
rect 280800 341600 280950 341750
rect 280500 341350 280650 341500
rect 280800 341350 280950 341500
rect 280500 341100 280650 341250
rect 280800 341100 280950 341250
rect 280500 340850 280650 341000
rect 280800 340850 280950 341000
rect 280500 340600 280650 340750
rect 280800 340600 280950 340750
rect 280500 340350 280650 340500
rect 280800 340350 280950 340500
rect 280500 340100 280650 340250
rect 280800 340100 280950 340250
rect 280500 339850 280650 340000
rect 280800 339850 280950 340000
rect 280500 339600 280650 339750
rect 280800 339600 280950 339750
rect 280500 339350 280650 339500
rect 280800 339350 280950 339500
rect 280500 339100 280650 339250
rect 280800 339100 280950 339250
<< metal3 >>
rect 232697 351150 235197 352400
rect 255297 351450 257697 352400
rect 260297 351450 262697 352400
rect 283297 351980 285797 352400
rect 232700 346550 235200 351150
rect 255250 351000 262900 351450
rect 255250 350700 258000 351000
rect 258300 350700 258500 351000
rect 258800 350700 259000 351000
rect 259300 350700 259500 351000
rect 259800 350700 260000 351000
rect 260300 350700 262900 351000
rect 255250 350600 262900 350700
rect 255250 350300 258000 350600
rect 258300 350300 258500 350600
rect 258800 350300 259000 350600
rect 259300 350300 259500 350600
rect 259800 350300 260000 350600
rect 260300 350300 262900 350600
rect 255250 350200 262900 350300
rect 255250 349900 258000 350200
rect 258300 349900 258500 350200
rect 258800 349900 259000 350200
rect 259300 349900 259500 350200
rect 259800 349900 260000 350200
rect 260300 349900 262900 350200
rect 255250 349630 262900 349900
rect 232700 346450 267250 346550
rect 232700 346350 266900 346450
rect 267000 346350 267100 346450
rect 267200 346350 267250 346450
rect 232700 346300 267250 346350
rect 232700 346200 266900 346300
rect 267000 346200 267100 346300
rect 267200 346200 267250 346300
rect 232700 346150 267250 346200
rect 232700 346050 266900 346150
rect 267000 346050 267100 346150
rect 267200 346050 267250 346150
rect 232700 346000 267250 346050
rect 232700 345900 266900 346000
rect 267000 345900 267100 346000
rect 267200 345900 267250 346000
rect 232700 345850 267250 345900
rect 232700 345750 266900 345850
rect 267000 345750 267100 345850
rect 267200 345750 267250 345850
rect 232700 345700 267250 345750
rect 232700 345600 266900 345700
rect 267000 345600 267100 345700
rect 267200 345600 267250 345700
rect 232700 345550 267250 345600
rect 232700 345450 266900 345550
rect 267000 345450 267100 345550
rect 267200 345450 267250 345550
rect 232700 345400 267250 345450
rect 232700 345300 266900 345400
rect 267000 345300 267100 345400
rect 267200 345300 267250 345400
rect 232700 345250 267250 345300
rect 232700 345150 266900 345250
rect 267000 345150 267100 345250
rect 267200 345150 267250 345250
rect 232700 345100 267250 345150
rect 232700 345000 266900 345100
rect 267000 345000 267100 345100
rect 267200 345000 267250 345100
rect 232700 344950 267250 345000
rect 232700 344850 266900 344950
rect 267000 344850 267100 344950
rect 267200 344850 267250 344950
rect 232700 344800 267250 344850
rect 232700 344700 266900 344800
rect 267000 344700 267100 344800
rect 267200 344700 267250 344800
rect 232700 344650 267250 344700
rect 232700 344550 266900 344650
rect 267000 344550 267100 344650
rect 267200 344550 267250 344650
rect 232700 344500 267250 344550
rect 232700 344400 266900 344500
rect 267000 344400 267100 344500
rect 267200 344400 267250 344500
rect 232700 344350 267250 344400
rect 232700 344250 266900 344350
rect 267000 344250 267100 344350
rect 267200 344250 267250 344350
rect 232700 344200 267250 344250
rect 232700 344100 266900 344200
rect 267000 344100 267100 344200
rect 267200 344100 267250 344200
rect 232700 344050 267250 344100
rect 232700 343950 266900 344050
rect 267000 343950 267100 344050
rect 267200 343950 267250 344050
rect 232700 343900 267250 343950
rect 232700 343800 266900 343900
rect 267000 343800 267100 343900
rect 267200 343800 267250 343900
rect 232700 343750 267250 343800
rect 232700 343650 266900 343750
rect 267000 343650 267100 343750
rect 267200 343650 267250 343750
rect 232700 343500 267250 343650
rect 283150 343500 285830 351980
rect 275595 343300 275600 343400
rect 275700 343300 275705 343400
rect 275795 343300 275800 343400
rect 275900 343300 275905 343400
rect 275995 343300 276000 343400
rect 276100 343300 276105 343400
rect 276195 343300 276200 343400
rect 276300 343300 276305 343400
rect 276395 343300 276400 343400
rect 276500 343300 276505 343400
rect 283150 343300 283250 343500
rect 283450 343300 283650 343500
rect 283850 343300 284050 343500
rect 284250 343300 284450 343500
rect 284650 343300 284850 343500
rect 285050 343300 285250 343500
rect 285450 343300 285830 343500
rect 283150 343100 285830 343300
rect 283150 342900 283250 343100
rect 283450 342900 283650 343100
rect 283850 342900 284050 343100
rect 284250 342900 284450 343100
rect 284650 342900 284850 343100
rect 285050 342900 285250 343100
rect 285450 342900 285830 343100
rect 275595 342750 275600 342850
rect 275700 342750 275705 342850
rect 275795 342750 275800 342850
rect 275900 342750 275905 342850
rect 275995 342750 276000 342850
rect 276100 342750 276105 342850
rect 276195 342750 276200 342850
rect 276300 342750 276305 342850
rect 283150 342830 285830 342900
rect 257850 342200 270850 342250
rect 257850 341900 258000 342200
rect 258300 341900 258500 342200
rect 258800 341900 259000 342200
rect 259300 341900 259500 342200
rect 259800 341900 260000 342200
rect 260300 341900 270850 342200
rect 257850 341700 270850 341900
rect 257850 341400 258000 341700
rect 258300 341400 258500 341700
rect 258800 341400 259000 341700
rect 259300 341400 259500 341700
rect 259800 341400 260000 341700
rect 260300 341400 270850 341700
rect 257850 341200 270850 341400
rect 257850 340900 258000 341200
rect 258300 340900 258500 341200
rect 258800 340900 259000 341200
rect 259300 340900 259500 341200
rect 259800 340900 260000 341200
rect 260300 340900 270850 341200
rect 257850 340750 270850 340900
rect 280450 342000 281000 342070
rect 280450 341850 280500 342000
rect 280650 341850 280800 342000
rect 280950 341850 281000 342000
rect 280450 341750 281000 341850
rect 280450 341600 280500 341750
rect 280650 341600 280800 341750
rect 280950 341600 281000 341750
rect 280450 341550 281000 341600
rect 280450 341500 292000 341550
rect 280450 341350 280500 341500
rect 280650 341350 280800 341500
rect 280950 341492 292000 341500
rect 280950 341350 292400 341492
rect 280450 341250 292400 341350
rect 280450 341100 280500 341250
rect 280650 341100 280800 341250
rect 280950 341100 292400 341250
rect 280450 341000 292400 341100
rect 280450 340850 280500 341000
rect 280650 340850 280800 341000
rect 280950 340850 292400 341000
rect 280450 340750 292400 340850
rect 280450 340600 280500 340750
rect 280650 340600 280800 340750
rect 280950 340600 292400 340750
rect 280450 340500 292400 340600
rect 273495 340400 273500 340500
rect 273600 340400 273605 340500
rect 273695 340400 273700 340500
rect 273800 340400 273805 340500
rect 273895 340400 273900 340500
rect 274000 340400 274005 340500
rect 274095 340400 274100 340500
rect 274200 340400 274205 340500
rect 274295 340400 274300 340500
rect 274400 340400 274405 340500
rect 274495 340400 274500 340500
rect 274600 340400 274605 340500
rect 280450 340350 280500 340500
rect 280650 340350 280800 340500
rect 280950 340350 292400 340500
rect 273495 340250 273500 340350
rect 273600 340250 273605 340350
rect 273695 340250 273700 340350
rect 273800 340250 273805 340350
rect 273895 340250 273900 340350
rect 274000 340250 274005 340350
rect 274095 340250 274100 340350
rect 274200 340250 274205 340350
rect 274295 340250 274300 340350
rect 274400 340250 274405 340350
rect 280450 340250 292400 340350
rect 280450 340100 280500 340250
rect 280650 340100 280800 340250
rect 280950 340100 292400 340250
rect 280450 340000 292400 340100
rect 280450 339850 280500 340000
rect 280650 339850 280800 340000
rect 280950 339850 292400 340000
rect 280450 339750 292400 339850
rect 257850 339400 271800 339650
rect 275490 339600 275880 339620
rect 257850 339100 258000 339400
rect 258300 339100 258500 339400
rect 258800 339100 259000 339400
rect 259300 339100 259500 339400
rect 259800 339100 260000 339400
rect 260300 339100 271800 339400
rect 274750 339260 275880 339600
rect 280450 339600 280500 339750
rect 280650 339600 280800 339750
rect 280950 339600 292400 339750
rect 280450 339500 292400 339600
rect 280450 339350 280500 339500
rect 280650 339350 280800 339500
rect 280950 339350 292400 339500
rect 274750 339250 275550 339260
rect 280450 339250 292400 339350
rect 257850 338900 271800 339100
rect 280450 339100 280500 339250
rect 280650 339100 280800 339250
rect 280950 339100 292400 339250
rect 280450 338992 292400 339100
rect 280450 338950 292000 338992
rect 257850 338600 258000 338900
rect 258300 338600 258500 338900
rect 258800 338600 259000 338900
rect 259300 338600 259500 338900
rect 259800 338600 260000 338900
rect 260300 338600 271800 338900
rect 257850 338400 271800 338600
rect 257850 338100 258000 338400
rect 258300 338100 258500 338400
rect 258800 338100 259000 338400
rect 259300 338100 259500 338400
rect 259800 338100 260000 338400
rect 260300 338100 271800 338400
rect 257850 338000 271800 338100
rect 289500 322300 291200 322350
rect 275500 322292 291200 322300
rect 275500 321800 292400 322292
rect 275500 321400 275600 321800
rect 276000 321400 276500 321800
rect 276900 321400 292400 321800
rect 275500 321000 292400 321400
rect 275500 320600 275600 321000
rect 276000 320600 276500 321000
rect 276900 320600 292400 321000
rect 275500 320200 292400 320600
rect 275500 319800 275600 320200
rect 276000 319800 276500 320200
rect 276900 319892 292400 320200
rect 276900 319800 291200 319892
rect 275500 319400 291200 319800
rect 275500 319000 275600 319400
rect 276000 319000 276500 319400
rect 276900 319000 291200 319400
rect 275500 318600 291200 319000
rect 275500 318200 275600 318600
rect 276000 318200 276500 318600
rect 276900 318200 291200 318600
rect 275500 317800 291200 318200
rect 275500 317400 275600 317800
rect 276000 317400 276500 317800
rect 276900 317400 291200 317800
rect 275500 317292 291200 317400
rect 275500 317000 292400 317292
rect 275500 316600 275600 317000
rect 276000 316600 276500 317000
rect 276900 316600 292400 317000
rect 275500 316200 292400 316600
rect 275500 315800 275600 316200
rect 276000 315800 276500 316200
rect 276900 315800 292400 316200
rect 275500 315400 292400 315800
rect 275500 315000 275600 315400
rect 276000 315000 276500 315400
rect 276900 315000 292400 315400
rect 275500 314900 292400 315000
rect 275500 314850 289900 314900
rect 291170 314892 292400 314900
<< via3 >>
rect 258000 350700 258300 351000
rect 258500 350700 258800 351000
rect 259000 350700 259300 351000
rect 259500 350700 259800 351000
rect 260000 350700 260300 351000
rect 258000 350300 258300 350600
rect 258500 350300 258800 350600
rect 259000 350300 259300 350600
rect 259500 350300 259800 350600
rect 260000 350300 260300 350600
rect 258000 349900 258300 350200
rect 258500 349900 258800 350200
rect 259000 349900 259300 350200
rect 259500 349900 259800 350200
rect 260000 349900 260300 350200
rect 266900 346350 267000 346450
rect 267100 346350 267200 346450
rect 266900 346200 267000 346300
rect 267100 346200 267200 346300
rect 266900 346050 267000 346150
rect 267100 346050 267200 346150
rect 266900 345900 267000 346000
rect 267100 345900 267200 346000
rect 266900 345750 267000 345850
rect 267100 345750 267200 345850
rect 266900 345600 267000 345700
rect 267100 345600 267200 345700
rect 266900 345450 267000 345550
rect 267100 345450 267200 345550
rect 266900 345300 267000 345400
rect 267100 345300 267200 345400
rect 266900 345150 267000 345250
rect 267100 345150 267200 345250
rect 266900 345000 267000 345100
rect 267100 345000 267200 345100
rect 266900 344850 267000 344950
rect 267100 344850 267200 344950
rect 266900 344700 267000 344800
rect 267100 344700 267200 344800
rect 266900 344550 267000 344650
rect 267100 344550 267200 344650
rect 266900 344400 267000 344500
rect 267100 344400 267200 344500
rect 266900 344250 267000 344350
rect 267100 344250 267200 344350
rect 266900 344100 267000 344200
rect 267100 344100 267200 344200
rect 266900 343950 267000 344050
rect 267100 343950 267200 344050
rect 266900 343800 267000 343900
rect 267100 343800 267200 343900
rect 266900 343650 267000 343750
rect 267100 343650 267200 343750
rect 275600 343300 275700 343400
rect 275800 343300 275900 343400
rect 276000 343300 276100 343400
rect 276200 343300 276300 343400
rect 276400 343300 276500 343400
rect 275600 342750 275700 342850
rect 275800 342750 275900 342850
rect 276000 342750 276100 342850
rect 276200 342750 276300 342850
rect 258000 341900 258300 342200
rect 258500 341900 258800 342200
rect 259000 341900 259300 342200
rect 259500 341900 259800 342200
rect 260000 341900 260300 342200
rect 258000 341400 258300 341700
rect 258500 341400 258800 341700
rect 259000 341400 259300 341700
rect 259500 341400 259800 341700
rect 260000 341400 260300 341700
rect 258000 340900 258300 341200
rect 258500 340900 258800 341200
rect 259000 340900 259300 341200
rect 259500 340900 259800 341200
rect 260000 340900 260300 341200
rect 273500 340400 273600 340500
rect 273700 340400 273800 340500
rect 273900 340400 274000 340500
rect 274100 340400 274200 340500
rect 274300 340400 274400 340500
rect 274500 340400 274600 340500
rect 273500 340250 273600 340350
rect 273700 340250 273800 340350
rect 273900 340250 274000 340350
rect 274100 340250 274200 340350
rect 274300 340250 274400 340350
rect 258000 339100 258300 339400
rect 258500 339100 258800 339400
rect 259000 339100 259300 339400
rect 259500 339100 259800 339400
rect 260000 339100 260300 339400
rect 258000 338600 258300 338900
rect 258500 338600 258800 338900
rect 259000 338600 259300 338900
rect 259500 338600 259800 338900
rect 260000 338600 260300 338900
rect 258000 338100 258300 338400
rect 258500 338100 258800 338400
rect 259000 338100 259300 338400
rect 259500 338100 259800 338400
rect 260000 338100 260300 338400
rect 275600 321400 276000 321800
rect 276500 321400 276900 321800
rect 275600 320600 276000 321000
rect 276500 320600 276900 321000
rect 275600 319800 276000 320200
rect 276500 319800 276900 320200
rect 275600 319000 276000 319400
rect 276500 319000 276900 319400
rect 275600 318200 276000 318600
rect 276500 318200 276900 318600
rect 275600 317400 276000 317800
rect 276500 317400 276900 317800
rect 275600 316600 276000 317000
rect 276500 316600 276900 317000
rect 275600 315800 276000 316200
rect 276500 315800 276900 316200
rect 275600 315000 276000 315400
rect 276500 315000 276900 315400
<< metal4 >>
rect 257850 351000 260410 351100
rect 257850 350700 258000 351000
rect 258300 350700 258500 351000
rect 258800 350700 259000 351000
rect 259300 350700 259500 351000
rect 259800 350700 260000 351000
rect 260300 350700 260410 351000
rect 257850 350600 260400 350700
rect 257850 350300 258000 350600
rect 258300 350300 258500 350600
rect 258800 350300 259000 350600
rect 259300 350300 259500 350600
rect 259800 350300 260000 350600
rect 260300 350300 260400 350600
rect 257850 350200 260400 350300
rect 257850 349900 258000 350200
rect 258300 349900 258500 350200
rect 258800 349900 259000 350200
rect 259300 349900 259500 350200
rect 259800 349900 260000 350200
rect 260300 349900 260400 350200
rect 257850 342200 260400 349900
rect 266850 346450 267250 346550
rect 266850 346350 266900 346450
rect 267000 346350 267100 346450
rect 267200 346350 267250 346450
rect 266850 346300 267250 346350
rect 266850 346200 266900 346300
rect 267000 346200 267100 346300
rect 267200 346200 267250 346300
rect 266850 346150 267250 346200
rect 266850 346050 266900 346150
rect 267000 346050 267100 346150
rect 267200 346050 267250 346150
rect 266850 346000 267250 346050
rect 266850 345900 266900 346000
rect 267000 345900 267100 346000
rect 267200 345900 267250 346000
rect 266850 345850 267250 345900
rect 266850 345750 266900 345850
rect 267000 345750 267100 345850
rect 267200 345750 267250 345850
rect 266850 345700 267250 345750
rect 266850 345600 266900 345700
rect 267000 345600 267100 345700
rect 267200 345600 267250 345700
rect 266850 345550 267250 345600
rect 266850 345450 266900 345550
rect 267000 345450 267100 345550
rect 267200 345450 267250 345550
rect 266850 345400 267250 345450
rect 266850 345300 266900 345400
rect 267000 345300 267100 345400
rect 267200 345300 267250 345400
rect 266850 345250 267250 345300
rect 266850 345150 266900 345250
rect 267000 345150 267100 345250
rect 267200 345170 267250 345250
rect 267200 345150 270380 345170
rect 266850 345100 270380 345150
rect 266850 345000 266900 345100
rect 267000 345000 267100 345100
rect 267200 345000 270380 345100
rect 266850 344950 270380 345000
rect 266850 344850 266900 344950
rect 267000 344850 267100 344950
rect 267200 344850 270380 344950
rect 266850 344800 270380 344850
rect 266850 344700 266900 344800
rect 267000 344700 267100 344800
rect 267200 344700 270380 344800
rect 266850 344650 270380 344700
rect 266850 344550 266900 344650
rect 267000 344550 267100 344650
rect 267200 344550 270380 344650
rect 266850 344500 270380 344550
rect 266850 344400 266900 344500
rect 267000 344400 267100 344500
rect 267200 344480 270380 344500
rect 267200 344400 267250 344480
rect 266850 344350 267250 344400
rect 266850 344250 266900 344350
rect 267000 344250 267100 344350
rect 267200 344250 267250 344350
rect 266850 344200 267250 344250
rect 266850 344100 266900 344200
rect 267000 344100 267100 344200
rect 267200 344100 267250 344200
rect 266850 344050 267250 344100
rect 266850 343950 266900 344050
rect 267000 343950 267100 344050
rect 267200 343950 267250 344050
rect 266850 343900 267250 343950
rect 266850 343800 266900 343900
rect 267000 343800 267100 343900
rect 267200 343800 267250 343900
rect 266850 343750 267250 343800
rect 266850 343650 266900 343750
rect 267000 343650 267100 343750
rect 267200 343650 267250 343750
rect 266850 343500 267250 343650
rect 257850 341900 258000 342200
rect 258300 341900 258500 342200
rect 258800 341900 259000 342200
rect 259300 341900 259500 342200
rect 259800 341900 260000 342200
rect 260300 341900 260400 342200
rect 257850 341700 260400 341900
rect 257850 341400 258000 341700
rect 258300 341400 258500 341700
rect 258800 341400 259000 341700
rect 259300 341400 259500 341700
rect 259800 341400 260000 341700
rect 260300 341400 260400 341700
rect 257850 341200 260400 341400
rect 257850 340900 258000 341200
rect 258300 340900 258500 341200
rect 258800 340900 259000 341200
rect 259300 340900 259500 341200
rect 259800 340900 260000 341200
rect 260300 340900 260400 341200
rect 257850 339400 260400 340900
rect 275500 343400 277000 343450
rect 275500 343300 275600 343400
rect 275700 343300 275800 343400
rect 275900 343300 276000 343400
rect 276100 343300 276200 343400
rect 276300 343300 276400 343400
rect 276500 343300 277000 343400
rect 275500 342850 277000 343300
rect 275500 342750 275600 342850
rect 275700 342750 275800 342850
rect 275900 342750 276000 342850
rect 276100 342750 276200 342850
rect 276300 342750 277000 342850
rect 275500 340550 277000 342750
rect 273350 340500 277000 340550
rect 273350 340400 273500 340500
rect 273600 340400 273700 340500
rect 273800 340400 273900 340500
rect 274000 340400 274100 340500
rect 274200 340400 274300 340500
rect 274400 340400 274500 340500
rect 274600 340400 277000 340500
rect 273350 340350 277000 340400
rect 273350 340250 273500 340350
rect 273600 340250 273700 340350
rect 273800 340250 273900 340350
rect 274000 340250 274100 340350
rect 274200 340250 274300 340350
rect 274400 340250 277000 340350
rect 273350 340200 277000 340250
rect 257850 339100 258000 339400
rect 258300 339100 258500 339400
rect 258800 339100 259000 339400
rect 259300 339100 259500 339400
rect 259800 339100 260000 339400
rect 260300 339100 260400 339400
rect 257850 338900 260400 339100
rect 257850 338600 258000 338900
rect 258300 338600 258500 338900
rect 258800 338600 259000 338900
rect 259300 338600 259500 338900
rect 259800 338600 260000 338900
rect 260300 338600 260400 338900
rect 257850 338400 260400 338600
rect 257850 338100 258000 338400
rect 258300 338100 258500 338400
rect 258800 338100 259000 338400
rect 259300 338100 259500 338400
rect 259800 338100 260000 338400
rect 260300 338100 260400 338400
rect 257850 338000 260400 338100
rect 275500 321800 277000 340200
rect 275500 321400 275600 321800
rect 276000 321400 276500 321800
rect 276900 321400 277000 321800
rect 275500 321000 277000 321400
rect 275500 320600 275600 321000
rect 276000 320600 276500 321000
rect 276900 320600 277000 321000
rect 275500 320200 277000 320600
rect 275500 319800 275600 320200
rect 276000 319800 276500 320200
rect 276900 319800 277000 320200
rect 275500 319400 277000 319800
rect 275500 319000 275600 319400
rect 276000 319000 276500 319400
rect 276900 319000 277000 319400
rect 275500 318600 277000 319000
rect 275500 318200 275600 318600
rect 276000 318200 276500 318600
rect 276900 318200 277000 318600
rect 275500 317800 277000 318200
rect 275500 317400 275600 317800
rect 276000 317400 276500 317800
rect 276900 317400 277000 317800
rect 275500 317000 277000 317400
rect 275500 316600 275600 317000
rect 276000 316600 276500 317000
rect 276900 316600 277000 317000
rect 275500 316200 277000 316600
rect 275500 315800 275600 316200
rect 276000 315800 276500 316200
rect 276900 315800 277000 316200
rect 275500 315400 277000 315800
rect 275500 315000 275600 315400
rect 276000 315000 276500 315400
rect 276900 315000 277000 315400
rect 275500 314850 277000 315000
use MULT_Amp  MULT_Amp_0
timestamp 1709331665
transform 1 0 268107 0 1 331446
box 0 -5 10118 15882
<< labels >>
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 560 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 960 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 960 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 560 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 560 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 960 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 960 180 0 0 vssa1
port 563 nsew signal bidirectional
<< end >>
