magic
tech sky130A
magscale 1 2
timestamp 1712803619
<< error_s >>
rect 866 765 907 797
rect 1456 717 1497 749
rect 1954 669 1995 701
rect 5034 381 5075 413
rect 5624 333 5665 365
rect 6306 285 6347 317
rect 6988 237 7029 269
rect 7670 189 7711 221
rect 8352 141 8393 173
rect 8850 93 8891 125
rect 9938 -3 9979 29
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
use sky130_fd_sc_hd__or4_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 314 0 1 552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  x2
timestamp 1701704242
transform 1 0 904 0 1 504
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 9976 0 1 -264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1494 0 1 456
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1701704242
transform 1 0 10290 0 1 -312
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1701704242
transform 1 0 10604 0 1 -360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1701704242
transform 1 0 10918 0 1 -408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1992 0 1 408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1701704242
transform 1 0 0 0 1 600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x10
timestamp 1701704242
transform 1 0 2490 0 1 360
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x11
timestamp 1701704242
transform 1 0 2988 0 1 312
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x12
timestamp 1701704242
transform 1 0 3486 0 1 264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x13
timestamp 1701704242
transform 1 0 3984 0 1 216
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x14
timestamp 1701704242
transform 1 0 4482 0 1 168
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5662 0 1 72
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x16
timestamp 1701704242
transform 1 0 6344 0 1 24
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  x17
timestamp 1701704242
transform 1 0 5072 0 1 120
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x18
timestamp 1701704242
transform 1 0 7026 0 1 -24
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x19
timestamp 1701704242
transform 1 0 7708 0 1 -72
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8390 0 1 -120
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x21
timestamp 1701704242
transform 1 0 8888 0 1 -168
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x22
timestamp 1701704242
transform 1 0 9386 0 1 -216
box -38 -48 590 592
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 I1
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 I5
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 I3
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 I0
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 I2
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 I6
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 I7
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 I4
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 EO
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 GS
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 A2
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 A1
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 A0
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 EI
port 13 nsew
<< end >>
