magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< pwell >>
rect -5086 -13686 5086 13686
<< psubdiff >>
rect -5050 13616 -4954 13650
rect 4954 13616 5050 13650
rect -5050 13554 -5016 13616
rect 5016 13554 5050 13616
rect -5050 -13616 -5016 -13554
rect 5016 -13616 5050 -13554
rect -5050 -13650 -4954 -13616
rect 4954 -13650 5050 -13616
<< psubdiffcont >>
rect -4954 13616 4954 13650
rect -5050 -13554 -5016 13554
rect 5016 -13554 5050 13554
rect -4954 -13650 4954 -13616
<< xpolycontact >>
rect -4920 13088 -3774 13520
rect -4920 12116 -3774 12548
rect -3678 13088 -2532 13520
rect -3678 12116 -2532 12548
rect -2436 13088 -1290 13520
rect -2436 12116 -1290 12548
rect -1194 13088 -48 13520
rect -1194 12116 -48 12548
rect 48 13088 1194 13520
rect 48 12116 1194 12548
rect 1290 13088 2436 13520
rect 1290 12116 2436 12548
rect 2532 13088 3678 13520
rect 2532 12116 3678 12548
rect 3774 13088 4920 13520
rect 3774 12116 4920 12548
rect -4920 11580 -3774 12012
rect -4920 10608 -3774 11040
rect -3678 11580 -2532 12012
rect -3678 10608 -2532 11040
rect -2436 11580 -1290 12012
rect -2436 10608 -1290 11040
rect -1194 11580 -48 12012
rect -1194 10608 -48 11040
rect 48 11580 1194 12012
rect 48 10608 1194 11040
rect 1290 11580 2436 12012
rect 1290 10608 2436 11040
rect 2532 11580 3678 12012
rect 2532 10608 3678 11040
rect 3774 11580 4920 12012
rect 3774 10608 4920 11040
rect -4920 10072 -3774 10504
rect -4920 9100 -3774 9532
rect -3678 10072 -2532 10504
rect -3678 9100 -2532 9532
rect -2436 10072 -1290 10504
rect -2436 9100 -1290 9532
rect -1194 10072 -48 10504
rect -1194 9100 -48 9532
rect 48 10072 1194 10504
rect 48 9100 1194 9532
rect 1290 10072 2436 10504
rect 1290 9100 2436 9532
rect 2532 10072 3678 10504
rect 2532 9100 3678 9532
rect 3774 10072 4920 10504
rect 3774 9100 4920 9532
rect -4920 8564 -3774 8996
rect -4920 7592 -3774 8024
rect -3678 8564 -2532 8996
rect -3678 7592 -2532 8024
rect -2436 8564 -1290 8996
rect -2436 7592 -1290 8024
rect -1194 8564 -48 8996
rect -1194 7592 -48 8024
rect 48 8564 1194 8996
rect 48 7592 1194 8024
rect 1290 8564 2436 8996
rect 1290 7592 2436 8024
rect 2532 8564 3678 8996
rect 2532 7592 3678 8024
rect 3774 8564 4920 8996
rect 3774 7592 4920 8024
rect -4920 7056 -3774 7488
rect -4920 6084 -3774 6516
rect -3678 7056 -2532 7488
rect -3678 6084 -2532 6516
rect -2436 7056 -1290 7488
rect -2436 6084 -1290 6516
rect -1194 7056 -48 7488
rect -1194 6084 -48 6516
rect 48 7056 1194 7488
rect 48 6084 1194 6516
rect 1290 7056 2436 7488
rect 1290 6084 2436 6516
rect 2532 7056 3678 7488
rect 2532 6084 3678 6516
rect 3774 7056 4920 7488
rect 3774 6084 4920 6516
rect -4920 5548 -3774 5980
rect -4920 4576 -3774 5008
rect -3678 5548 -2532 5980
rect -3678 4576 -2532 5008
rect -2436 5548 -1290 5980
rect -2436 4576 -1290 5008
rect -1194 5548 -48 5980
rect -1194 4576 -48 5008
rect 48 5548 1194 5980
rect 48 4576 1194 5008
rect 1290 5548 2436 5980
rect 1290 4576 2436 5008
rect 2532 5548 3678 5980
rect 2532 4576 3678 5008
rect 3774 5548 4920 5980
rect 3774 4576 4920 5008
rect -4920 4040 -3774 4472
rect -4920 3068 -3774 3500
rect -3678 4040 -2532 4472
rect -3678 3068 -2532 3500
rect -2436 4040 -1290 4472
rect -2436 3068 -1290 3500
rect -1194 4040 -48 4472
rect -1194 3068 -48 3500
rect 48 4040 1194 4472
rect 48 3068 1194 3500
rect 1290 4040 2436 4472
rect 1290 3068 2436 3500
rect 2532 4040 3678 4472
rect 2532 3068 3678 3500
rect 3774 4040 4920 4472
rect 3774 3068 4920 3500
rect -4920 2532 -3774 2964
rect -4920 1560 -3774 1992
rect -3678 2532 -2532 2964
rect -3678 1560 -2532 1992
rect -2436 2532 -1290 2964
rect -2436 1560 -1290 1992
rect -1194 2532 -48 2964
rect -1194 1560 -48 1992
rect 48 2532 1194 2964
rect 48 1560 1194 1992
rect 1290 2532 2436 2964
rect 1290 1560 2436 1992
rect 2532 2532 3678 2964
rect 2532 1560 3678 1992
rect 3774 2532 4920 2964
rect 3774 1560 4920 1992
rect -4920 1024 -3774 1456
rect -4920 52 -3774 484
rect -3678 1024 -2532 1456
rect -3678 52 -2532 484
rect -2436 1024 -1290 1456
rect -2436 52 -1290 484
rect -1194 1024 -48 1456
rect -1194 52 -48 484
rect 48 1024 1194 1456
rect 48 52 1194 484
rect 1290 1024 2436 1456
rect 1290 52 2436 484
rect 2532 1024 3678 1456
rect 2532 52 3678 484
rect 3774 1024 4920 1456
rect 3774 52 4920 484
rect -4920 -484 -3774 -52
rect -4920 -1456 -3774 -1024
rect -3678 -484 -2532 -52
rect -3678 -1456 -2532 -1024
rect -2436 -484 -1290 -52
rect -2436 -1456 -1290 -1024
rect -1194 -484 -48 -52
rect -1194 -1456 -48 -1024
rect 48 -484 1194 -52
rect 48 -1456 1194 -1024
rect 1290 -484 2436 -52
rect 1290 -1456 2436 -1024
rect 2532 -484 3678 -52
rect 2532 -1456 3678 -1024
rect 3774 -484 4920 -52
rect 3774 -1456 4920 -1024
rect -4920 -1992 -3774 -1560
rect -4920 -2964 -3774 -2532
rect -3678 -1992 -2532 -1560
rect -3678 -2964 -2532 -2532
rect -2436 -1992 -1290 -1560
rect -2436 -2964 -1290 -2532
rect -1194 -1992 -48 -1560
rect -1194 -2964 -48 -2532
rect 48 -1992 1194 -1560
rect 48 -2964 1194 -2532
rect 1290 -1992 2436 -1560
rect 1290 -2964 2436 -2532
rect 2532 -1992 3678 -1560
rect 2532 -2964 3678 -2532
rect 3774 -1992 4920 -1560
rect 3774 -2964 4920 -2532
rect -4920 -3500 -3774 -3068
rect -4920 -4472 -3774 -4040
rect -3678 -3500 -2532 -3068
rect -3678 -4472 -2532 -4040
rect -2436 -3500 -1290 -3068
rect -2436 -4472 -1290 -4040
rect -1194 -3500 -48 -3068
rect -1194 -4472 -48 -4040
rect 48 -3500 1194 -3068
rect 48 -4472 1194 -4040
rect 1290 -3500 2436 -3068
rect 1290 -4472 2436 -4040
rect 2532 -3500 3678 -3068
rect 2532 -4472 3678 -4040
rect 3774 -3500 4920 -3068
rect 3774 -4472 4920 -4040
rect -4920 -5008 -3774 -4576
rect -4920 -5980 -3774 -5548
rect -3678 -5008 -2532 -4576
rect -3678 -5980 -2532 -5548
rect -2436 -5008 -1290 -4576
rect -2436 -5980 -1290 -5548
rect -1194 -5008 -48 -4576
rect -1194 -5980 -48 -5548
rect 48 -5008 1194 -4576
rect 48 -5980 1194 -5548
rect 1290 -5008 2436 -4576
rect 1290 -5980 2436 -5548
rect 2532 -5008 3678 -4576
rect 2532 -5980 3678 -5548
rect 3774 -5008 4920 -4576
rect 3774 -5980 4920 -5548
rect -4920 -6516 -3774 -6084
rect -4920 -7488 -3774 -7056
rect -3678 -6516 -2532 -6084
rect -3678 -7488 -2532 -7056
rect -2436 -6516 -1290 -6084
rect -2436 -7488 -1290 -7056
rect -1194 -6516 -48 -6084
rect -1194 -7488 -48 -7056
rect 48 -6516 1194 -6084
rect 48 -7488 1194 -7056
rect 1290 -6516 2436 -6084
rect 1290 -7488 2436 -7056
rect 2532 -6516 3678 -6084
rect 2532 -7488 3678 -7056
rect 3774 -6516 4920 -6084
rect 3774 -7488 4920 -7056
rect -4920 -8024 -3774 -7592
rect -4920 -8996 -3774 -8564
rect -3678 -8024 -2532 -7592
rect -3678 -8996 -2532 -8564
rect -2436 -8024 -1290 -7592
rect -2436 -8996 -1290 -8564
rect -1194 -8024 -48 -7592
rect -1194 -8996 -48 -8564
rect 48 -8024 1194 -7592
rect 48 -8996 1194 -8564
rect 1290 -8024 2436 -7592
rect 1290 -8996 2436 -8564
rect 2532 -8024 3678 -7592
rect 2532 -8996 3678 -8564
rect 3774 -8024 4920 -7592
rect 3774 -8996 4920 -8564
rect -4920 -9532 -3774 -9100
rect -4920 -10504 -3774 -10072
rect -3678 -9532 -2532 -9100
rect -3678 -10504 -2532 -10072
rect -2436 -9532 -1290 -9100
rect -2436 -10504 -1290 -10072
rect -1194 -9532 -48 -9100
rect -1194 -10504 -48 -10072
rect 48 -9532 1194 -9100
rect 48 -10504 1194 -10072
rect 1290 -9532 2436 -9100
rect 1290 -10504 2436 -10072
rect 2532 -9532 3678 -9100
rect 2532 -10504 3678 -10072
rect 3774 -9532 4920 -9100
rect 3774 -10504 4920 -10072
rect -4920 -11040 -3774 -10608
rect -4920 -12012 -3774 -11580
rect -3678 -11040 -2532 -10608
rect -3678 -12012 -2532 -11580
rect -2436 -11040 -1290 -10608
rect -2436 -12012 -1290 -11580
rect -1194 -11040 -48 -10608
rect -1194 -12012 -48 -11580
rect 48 -11040 1194 -10608
rect 48 -12012 1194 -11580
rect 1290 -11040 2436 -10608
rect 1290 -12012 2436 -11580
rect 2532 -11040 3678 -10608
rect 2532 -12012 3678 -11580
rect 3774 -11040 4920 -10608
rect 3774 -12012 4920 -11580
rect -4920 -12548 -3774 -12116
rect -4920 -13520 -3774 -13088
rect -3678 -12548 -2532 -12116
rect -3678 -13520 -2532 -13088
rect -2436 -12548 -1290 -12116
rect -2436 -13520 -1290 -13088
rect -1194 -12548 -48 -12116
rect -1194 -13520 -48 -13088
rect 48 -12548 1194 -12116
rect 48 -13520 1194 -13088
rect 1290 -12548 2436 -12116
rect 1290 -13520 2436 -13088
rect 2532 -12548 3678 -12116
rect 2532 -13520 3678 -13088
rect 3774 -12548 4920 -12116
rect 3774 -13520 4920 -13088
<< xpolyres >>
rect -4920 12548 -3774 13088
rect -3678 12548 -2532 13088
rect -2436 12548 -1290 13088
rect -1194 12548 -48 13088
rect 48 12548 1194 13088
rect 1290 12548 2436 13088
rect 2532 12548 3678 13088
rect 3774 12548 4920 13088
rect -4920 11040 -3774 11580
rect -3678 11040 -2532 11580
rect -2436 11040 -1290 11580
rect -1194 11040 -48 11580
rect 48 11040 1194 11580
rect 1290 11040 2436 11580
rect 2532 11040 3678 11580
rect 3774 11040 4920 11580
rect -4920 9532 -3774 10072
rect -3678 9532 -2532 10072
rect -2436 9532 -1290 10072
rect -1194 9532 -48 10072
rect 48 9532 1194 10072
rect 1290 9532 2436 10072
rect 2532 9532 3678 10072
rect 3774 9532 4920 10072
rect -4920 8024 -3774 8564
rect -3678 8024 -2532 8564
rect -2436 8024 -1290 8564
rect -1194 8024 -48 8564
rect 48 8024 1194 8564
rect 1290 8024 2436 8564
rect 2532 8024 3678 8564
rect 3774 8024 4920 8564
rect -4920 6516 -3774 7056
rect -3678 6516 -2532 7056
rect -2436 6516 -1290 7056
rect -1194 6516 -48 7056
rect 48 6516 1194 7056
rect 1290 6516 2436 7056
rect 2532 6516 3678 7056
rect 3774 6516 4920 7056
rect -4920 5008 -3774 5548
rect -3678 5008 -2532 5548
rect -2436 5008 -1290 5548
rect -1194 5008 -48 5548
rect 48 5008 1194 5548
rect 1290 5008 2436 5548
rect 2532 5008 3678 5548
rect 3774 5008 4920 5548
rect -4920 3500 -3774 4040
rect -3678 3500 -2532 4040
rect -2436 3500 -1290 4040
rect -1194 3500 -48 4040
rect 48 3500 1194 4040
rect 1290 3500 2436 4040
rect 2532 3500 3678 4040
rect 3774 3500 4920 4040
rect -4920 1992 -3774 2532
rect -3678 1992 -2532 2532
rect -2436 1992 -1290 2532
rect -1194 1992 -48 2532
rect 48 1992 1194 2532
rect 1290 1992 2436 2532
rect 2532 1992 3678 2532
rect 3774 1992 4920 2532
rect -4920 484 -3774 1024
rect -3678 484 -2532 1024
rect -2436 484 -1290 1024
rect -1194 484 -48 1024
rect 48 484 1194 1024
rect 1290 484 2436 1024
rect 2532 484 3678 1024
rect 3774 484 4920 1024
rect -4920 -1024 -3774 -484
rect -3678 -1024 -2532 -484
rect -2436 -1024 -1290 -484
rect -1194 -1024 -48 -484
rect 48 -1024 1194 -484
rect 1290 -1024 2436 -484
rect 2532 -1024 3678 -484
rect 3774 -1024 4920 -484
rect -4920 -2532 -3774 -1992
rect -3678 -2532 -2532 -1992
rect -2436 -2532 -1290 -1992
rect -1194 -2532 -48 -1992
rect 48 -2532 1194 -1992
rect 1290 -2532 2436 -1992
rect 2532 -2532 3678 -1992
rect 3774 -2532 4920 -1992
rect -4920 -4040 -3774 -3500
rect -3678 -4040 -2532 -3500
rect -2436 -4040 -1290 -3500
rect -1194 -4040 -48 -3500
rect 48 -4040 1194 -3500
rect 1290 -4040 2436 -3500
rect 2532 -4040 3678 -3500
rect 3774 -4040 4920 -3500
rect -4920 -5548 -3774 -5008
rect -3678 -5548 -2532 -5008
rect -2436 -5548 -1290 -5008
rect -1194 -5548 -48 -5008
rect 48 -5548 1194 -5008
rect 1290 -5548 2436 -5008
rect 2532 -5548 3678 -5008
rect 3774 -5548 4920 -5008
rect -4920 -7056 -3774 -6516
rect -3678 -7056 -2532 -6516
rect -2436 -7056 -1290 -6516
rect -1194 -7056 -48 -6516
rect 48 -7056 1194 -6516
rect 1290 -7056 2436 -6516
rect 2532 -7056 3678 -6516
rect 3774 -7056 4920 -6516
rect -4920 -8564 -3774 -8024
rect -3678 -8564 -2532 -8024
rect -2436 -8564 -1290 -8024
rect -1194 -8564 -48 -8024
rect 48 -8564 1194 -8024
rect 1290 -8564 2436 -8024
rect 2532 -8564 3678 -8024
rect 3774 -8564 4920 -8024
rect -4920 -10072 -3774 -9532
rect -3678 -10072 -2532 -9532
rect -2436 -10072 -1290 -9532
rect -1194 -10072 -48 -9532
rect 48 -10072 1194 -9532
rect 1290 -10072 2436 -9532
rect 2532 -10072 3678 -9532
rect 3774 -10072 4920 -9532
rect -4920 -11580 -3774 -11040
rect -3678 -11580 -2532 -11040
rect -2436 -11580 -1290 -11040
rect -1194 -11580 -48 -11040
rect 48 -11580 1194 -11040
rect 1290 -11580 2436 -11040
rect 2532 -11580 3678 -11040
rect 3774 -11580 4920 -11040
rect -4920 -13088 -3774 -12548
rect -3678 -13088 -2532 -12548
rect -2436 -13088 -1290 -12548
rect -1194 -13088 -48 -12548
rect 48 -13088 1194 -12548
rect 1290 -13088 2436 -12548
rect 2532 -13088 3678 -12548
rect 3774 -13088 4920 -12548
<< locali >>
rect -5050 13616 -4954 13650
rect 4954 13616 5050 13650
rect -5050 13554 -5016 13616
rect 5016 13554 5050 13616
rect -5050 -13616 -5016 -13554
rect 5016 -13616 5050 -13554
rect -5050 -13650 -4954 -13616
rect 4954 -13650 5050 -13616
<< viali >>
rect -4904 13105 -3790 13502
rect -3662 13105 -2548 13502
rect -2420 13105 -1306 13502
rect -1178 13105 -64 13502
rect 64 13105 1178 13502
rect 1306 13105 2420 13502
rect 2548 13105 3662 13502
rect 3790 13105 4904 13502
rect -4904 12134 -3790 12531
rect -3662 12134 -2548 12531
rect -2420 12134 -1306 12531
rect -1178 12134 -64 12531
rect 64 12134 1178 12531
rect 1306 12134 2420 12531
rect 2548 12134 3662 12531
rect 3790 12134 4904 12531
rect -4904 11597 -3790 11994
rect -3662 11597 -2548 11994
rect -2420 11597 -1306 11994
rect -1178 11597 -64 11994
rect 64 11597 1178 11994
rect 1306 11597 2420 11994
rect 2548 11597 3662 11994
rect 3790 11597 4904 11994
rect -4904 10626 -3790 11023
rect -3662 10626 -2548 11023
rect -2420 10626 -1306 11023
rect -1178 10626 -64 11023
rect 64 10626 1178 11023
rect 1306 10626 2420 11023
rect 2548 10626 3662 11023
rect 3790 10626 4904 11023
rect -4904 10089 -3790 10486
rect -3662 10089 -2548 10486
rect -2420 10089 -1306 10486
rect -1178 10089 -64 10486
rect 64 10089 1178 10486
rect 1306 10089 2420 10486
rect 2548 10089 3662 10486
rect 3790 10089 4904 10486
rect -4904 9118 -3790 9515
rect -3662 9118 -2548 9515
rect -2420 9118 -1306 9515
rect -1178 9118 -64 9515
rect 64 9118 1178 9515
rect 1306 9118 2420 9515
rect 2548 9118 3662 9515
rect 3790 9118 4904 9515
rect -4904 8581 -3790 8978
rect -3662 8581 -2548 8978
rect -2420 8581 -1306 8978
rect -1178 8581 -64 8978
rect 64 8581 1178 8978
rect 1306 8581 2420 8978
rect 2548 8581 3662 8978
rect 3790 8581 4904 8978
rect -4904 7610 -3790 8007
rect -3662 7610 -2548 8007
rect -2420 7610 -1306 8007
rect -1178 7610 -64 8007
rect 64 7610 1178 8007
rect 1306 7610 2420 8007
rect 2548 7610 3662 8007
rect 3790 7610 4904 8007
rect -4904 7073 -3790 7470
rect -3662 7073 -2548 7470
rect -2420 7073 -1306 7470
rect -1178 7073 -64 7470
rect 64 7073 1178 7470
rect 1306 7073 2420 7470
rect 2548 7073 3662 7470
rect 3790 7073 4904 7470
rect -4904 6102 -3790 6499
rect -3662 6102 -2548 6499
rect -2420 6102 -1306 6499
rect -1178 6102 -64 6499
rect 64 6102 1178 6499
rect 1306 6102 2420 6499
rect 2548 6102 3662 6499
rect 3790 6102 4904 6499
rect -4904 5565 -3790 5962
rect -3662 5565 -2548 5962
rect -2420 5565 -1306 5962
rect -1178 5565 -64 5962
rect 64 5565 1178 5962
rect 1306 5565 2420 5962
rect 2548 5565 3662 5962
rect 3790 5565 4904 5962
rect -4904 4594 -3790 4991
rect -3662 4594 -2548 4991
rect -2420 4594 -1306 4991
rect -1178 4594 -64 4991
rect 64 4594 1178 4991
rect 1306 4594 2420 4991
rect 2548 4594 3662 4991
rect 3790 4594 4904 4991
rect -4904 4057 -3790 4454
rect -3662 4057 -2548 4454
rect -2420 4057 -1306 4454
rect -1178 4057 -64 4454
rect 64 4057 1178 4454
rect 1306 4057 2420 4454
rect 2548 4057 3662 4454
rect 3790 4057 4904 4454
rect -4904 3086 -3790 3483
rect -3662 3086 -2548 3483
rect -2420 3086 -1306 3483
rect -1178 3086 -64 3483
rect 64 3086 1178 3483
rect 1306 3086 2420 3483
rect 2548 3086 3662 3483
rect 3790 3086 4904 3483
rect -4904 2549 -3790 2946
rect -3662 2549 -2548 2946
rect -2420 2549 -1306 2946
rect -1178 2549 -64 2946
rect 64 2549 1178 2946
rect 1306 2549 2420 2946
rect 2548 2549 3662 2946
rect 3790 2549 4904 2946
rect -4904 1578 -3790 1975
rect -3662 1578 -2548 1975
rect -2420 1578 -1306 1975
rect -1178 1578 -64 1975
rect 64 1578 1178 1975
rect 1306 1578 2420 1975
rect 2548 1578 3662 1975
rect 3790 1578 4904 1975
rect -4904 1041 -3790 1438
rect -3662 1041 -2548 1438
rect -2420 1041 -1306 1438
rect -1178 1041 -64 1438
rect 64 1041 1178 1438
rect 1306 1041 2420 1438
rect 2548 1041 3662 1438
rect 3790 1041 4904 1438
rect -4904 70 -3790 467
rect -3662 70 -2548 467
rect -2420 70 -1306 467
rect -1178 70 -64 467
rect 64 70 1178 467
rect 1306 70 2420 467
rect 2548 70 3662 467
rect 3790 70 4904 467
rect -4904 -467 -3790 -70
rect -3662 -467 -2548 -70
rect -2420 -467 -1306 -70
rect -1178 -467 -64 -70
rect 64 -467 1178 -70
rect 1306 -467 2420 -70
rect 2548 -467 3662 -70
rect 3790 -467 4904 -70
rect -4904 -1438 -3790 -1041
rect -3662 -1438 -2548 -1041
rect -2420 -1438 -1306 -1041
rect -1178 -1438 -64 -1041
rect 64 -1438 1178 -1041
rect 1306 -1438 2420 -1041
rect 2548 -1438 3662 -1041
rect 3790 -1438 4904 -1041
rect -4904 -1975 -3790 -1578
rect -3662 -1975 -2548 -1578
rect -2420 -1975 -1306 -1578
rect -1178 -1975 -64 -1578
rect 64 -1975 1178 -1578
rect 1306 -1975 2420 -1578
rect 2548 -1975 3662 -1578
rect 3790 -1975 4904 -1578
rect -4904 -2946 -3790 -2549
rect -3662 -2946 -2548 -2549
rect -2420 -2946 -1306 -2549
rect -1178 -2946 -64 -2549
rect 64 -2946 1178 -2549
rect 1306 -2946 2420 -2549
rect 2548 -2946 3662 -2549
rect 3790 -2946 4904 -2549
rect -4904 -3483 -3790 -3086
rect -3662 -3483 -2548 -3086
rect -2420 -3483 -1306 -3086
rect -1178 -3483 -64 -3086
rect 64 -3483 1178 -3086
rect 1306 -3483 2420 -3086
rect 2548 -3483 3662 -3086
rect 3790 -3483 4904 -3086
rect -4904 -4454 -3790 -4057
rect -3662 -4454 -2548 -4057
rect -2420 -4454 -1306 -4057
rect -1178 -4454 -64 -4057
rect 64 -4454 1178 -4057
rect 1306 -4454 2420 -4057
rect 2548 -4454 3662 -4057
rect 3790 -4454 4904 -4057
rect -4904 -4991 -3790 -4594
rect -3662 -4991 -2548 -4594
rect -2420 -4991 -1306 -4594
rect -1178 -4991 -64 -4594
rect 64 -4991 1178 -4594
rect 1306 -4991 2420 -4594
rect 2548 -4991 3662 -4594
rect 3790 -4991 4904 -4594
rect -4904 -5962 -3790 -5565
rect -3662 -5962 -2548 -5565
rect -2420 -5962 -1306 -5565
rect -1178 -5962 -64 -5565
rect 64 -5962 1178 -5565
rect 1306 -5962 2420 -5565
rect 2548 -5962 3662 -5565
rect 3790 -5962 4904 -5565
rect -4904 -6499 -3790 -6102
rect -3662 -6499 -2548 -6102
rect -2420 -6499 -1306 -6102
rect -1178 -6499 -64 -6102
rect 64 -6499 1178 -6102
rect 1306 -6499 2420 -6102
rect 2548 -6499 3662 -6102
rect 3790 -6499 4904 -6102
rect -4904 -7470 -3790 -7073
rect -3662 -7470 -2548 -7073
rect -2420 -7470 -1306 -7073
rect -1178 -7470 -64 -7073
rect 64 -7470 1178 -7073
rect 1306 -7470 2420 -7073
rect 2548 -7470 3662 -7073
rect 3790 -7470 4904 -7073
rect -4904 -8007 -3790 -7610
rect -3662 -8007 -2548 -7610
rect -2420 -8007 -1306 -7610
rect -1178 -8007 -64 -7610
rect 64 -8007 1178 -7610
rect 1306 -8007 2420 -7610
rect 2548 -8007 3662 -7610
rect 3790 -8007 4904 -7610
rect -4904 -8978 -3790 -8581
rect -3662 -8978 -2548 -8581
rect -2420 -8978 -1306 -8581
rect -1178 -8978 -64 -8581
rect 64 -8978 1178 -8581
rect 1306 -8978 2420 -8581
rect 2548 -8978 3662 -8581
rect 3790 -8978 4904 -8581
rect -4904 -9515 -3790 -9118
rect -3662 -9515 -2548 -9118
rect -2420 -9515 -1306 -9118
rect -1178 -9515 -64 -9118
rect 64 -9515 1178 -9118
rect 1306 -9515 2420 -9118
rect 2548 -9515 3662 -9118
rect 3790 -9515 4904 -9118
rect -4904 -10486 -3790 -10089
rect -3662 -10486 -2548 -10089
rect -2420 -10486 -1306 -10089
rect -1178 -10486 -64 -10089
rect 64 -10486 1178 -10089
rect 1306 -10486 2420 -10089
rect 2548 -10486 3662 -10089
rect 3790 -10486 4904 -10089
rect -4904 -11023 -3790 -10626
rect -3662 -11023 -2548 -10626
rect -2420 -11023 -1306 -10626
rect -1178 -11023 -64 -10626
rect 64 -11023 1178 -10626
rect 1306 -11023 2420 -10626
rect 2548 -11023 3662 -10626
rect 3790 -11023 4904 -10626
rect -4904 -11994 -3790 -11597
rect -3662 -11994 -2548 -11597
rect -2420 -11994 -1306 -11597
rect -1178 -11994 -64 -11597
rect 64 -11994 1178 -11597
rect 1306 -11994 2420 -11597
rect 2548 -11994 3662 -11597
rect 3790 -11994 4904 -11597
rect -4904 -12531 -3790 -12134
rect -3662 -12531 -2548 -12134
rect -2420 -12531 -1306 -12134
rect -1178 -12531 -64 -12134
rect 64 -12531 1178 -12134
rect 1306 -12531 2420 -12134
rect 2548 -12531 3662 -12134
rect 3790 -12531 4904 -12134
rect -4904 -13502 -3790 -13105
rect -3662 -13502 -2548 -13105
rect -2420 -13502 -1306 -13105
rect -1178 -13502 -64 -13105
rect 64 -13502 1178 -13105
rect 1306 -13502 2420 -13105
rect 2548 -13502 3662 -13105
rect 3790 -13502 4904 -13105
<< metal1 >>
rect -4916 13502 -3778 13508
rect -4916 13105 -4904 13502
rect -3790 13105 -3778 13502
rect -4916 13099 -3778 13105
rect -3674 13502 -2536 13508
rect -3674 13105 -3662 13502
rect -2548 13105 -2536 13502
rect -3674 13099 -2536 13105
rect -2432 13502 -1294 13508
rect -2432 13105 -2420 13502
rect -1306 13105 -1294 13502
rect -2432 13099 -1294 13105
rect -1190 13502 -52 13508
rect -1190 13105 -1178 13502
rect -64 13105 -52 13502
rect -1190 13099 -52 13105
rect 52 13502 1190 13508
rect 52 13105 64 13502
rect 1178 13105 1190 13502
rect 52 13099 1190 13105
rect 1294 13502 2432 13508
rect 1294 13105 1306 13502
rect 2420 13105 2432 13502
rect 1294 13099 2432 13105
rect 2536 13502 3674 13508
rect 2536 13105 2548 13502
rect 3662 13105 3674 13502
rect 2536 13099 3674 13105
rect 3778 13502 4916 13508
rect 3778 13105 3790 13502
rect 4904 13105 4916 13502
rect 3778 13099 4916 13105
rect -4916 12531 -3778 12537
rect -4916 12134 -4904 12531
rect -3790 12134 -3778 12531
rect -4916 12128 -3778 12134
rect -3674 12531 -2536 12537
rect -3674 12134 -3662 12531
rect -2548 12134 -2536 12531
rect -3674 12128 -2536 12134
rect -2432 12531 -1294 12537
rect -2432 12134 -2420 12531
rect -1306 12134 -1294 12531
rect -2432 12128 -1294 12134
rect -1190 12531 -52 12537
rect -1190 12134 -1178 12531
rect -64 12134 -52 12531
rect -1190 12128 -52 12134
rect 52 12531 1190 12537
rect 52 12134 64 12531
rect 1178 12134 1190 12531
rect 52 12128 1190 12134
rect 1294 12531 2432 12537
rect 1294 12134 1306 12531
rect 2420 12134 2432 12531
rect 1294 12128 2432 12134
rect 2536 12531 3674 12537
rect 2536 12134 2548 12531
rect 3662 12134 3674 12531
rect 2536 12128 3674 12134
rect 3778 12531 4916 12537
rect 3778 12134 3790 12531
rect 4904 12134 4916 12531
rect 3778 12128 4916 12134
rect -4916 11994 -3778 12000
rect -4916 11597 -4904 11994
rect -3790 11597 -3778 11994
rect -4916 11591 -3778 11597
rect -3674 11994 -2536 12000
rect -3674 11597 -3662 11994
rect -2548 11597 -2536 11994
rect -3674 11591 -2536 11597
rect -2432 11994 -1294 12000
rect -2432 11597 -2420 11994
rect -1306 11597 -1294 11994
rect -2432 11591 -1294 11597
rect -1190 11994 -52 12000
rect -1190 11597 -1178 11994
rect -64 11597 -52 11994
rect -1190 11591 -52 11597
rect 52 11994 1190 12000
rect 52 11597 64 11994
rect 1178 11597 1190 11994
rect 52 11591 1190 11597
rect 1294 11994 2432 12000
rect 1294 11597 1306 11994
rect 2420 11597 2432 11994
rect 1294 11591 2432 11597
rect 2536 11994 3674 12000
rect 2536 11597 2548 11994
rect 3662 11597 3674 11994
rect 2536 11591 3674 11597
rect 3778 11994 4916 12000
rect 3778 11597 3790 11994
rect 4904 11597 4916 11994
rect 3778 11591 4916 11597
rect -4916 11023 -3778 11029
rect -4916 10626 -4904 11023
rect -3790 10626 -3778 11023
rect -4916 10620 -3778 10626
rect -3674 11023 -2536 11029
rect -3674 10626 -3662 11023
rect -2548 10626 -2536 11023
rect -3674 10620 -2536 10626
rect -2432 11023 -1294 11029
rect -2432 10626 -2420 11023
rect -1306 10626 -1294 11023
rect -2432 10620 -1294 10626
rect -1190 11023 -52 11029
rect -1190 10626 -1178 11023
rect -64 10626 -52 11023
rect -1190 10620 -52 10626
rect 52 11023 1190 11029
rect 52 10626 64 11023
rect 1178 10626 1190 11023
rect 52 10620 1190 10626
rect 1294 11023 2432 11029
rect 1294 10626 1306 11023
rect 2420 10626 2432 11023
rect 1294 10620 2432 10626
rect 2536 11023 3674 11029
rect 2536 10626 2548 11023
rect 3662 10626 3674 11023
rect 2536 10620 3674 10626
rect 3778 11023 4916 11029
rect 3778 10626 3790 11023
rect 4904 10626 4916 11023
rect 3778 10620 4916 10626
rect -4916 10486 -3778 10492
rect -4916 10089 -4904 10486
rect -3790 10089 -3778 10486
rect -4916 10083 -3778 10089
rect -3674 10486 -2536 10492
rect -3674 10089 -3662 10486
rect -2548 10089 -2536 10486
rect -3674 10083 -2536 10089
rect -2432 10486 -1294 10492
rect -2432 10089 -2420 10486
rect -1306 10089 -1294 10486
rect -2432 10083 -1294 10089
rect -1190 10486 -52 10492
rect -1190 10089 -1178 10486
rect -64 10089 -52 10486
rect -1190 10083 -52 10089
rect 52 10486 1190 10492
rect 52 10089 64 10486
rect 1178 10089 1190 10486
rect 52 10083 1190 10089
rect 1294 10486 2432 10492
rect 1294 10089 1306 10486
rect 2420 10089 2432 10486
rect 1294 10083 2432 10089
rect 2536 10486 3674 10492
rect 2536 10089 2548 10486
rect 3662 10089 3674 10486
rect 2536 10083 3674 10089
rect 3778 10486 4916 10492
rect 3778 10089 3790 10486
rect 4904 10089 4916 10486
rect 3778 10083 4916 10089
rect -4916 9515 -3778 9521
rect -4916 9118 -4904 9515
rect -3790 9118 -3778 9515
rect -4916 9112 -3778 9118
rect -3674 9515 -2536 9521
rect -3674 9118 -3662 9515
rect -2548 9118 -2536 9515
rect -3674 9112 -2536 9118
rect -2432 9515 -1294 9521
rect -2432 9118 -2420 9515
rect -1306 9118 -1294 9515
rect -2432 9112 -1294 9118
rect -1190 9515 -52 9521
rect -1190 9118 -1178 9515
rect -64 9118 -52 9515
rect -1190 9112 -52 9118
rect 52 9515 1190 9521
rect 52 9118 64 9515
rect 1178 9118 1190 9515
rect 52 9112 1190 9118
rect 1294 9515 2432 9521
rect 1294 9118 1306 9515
rect 2420 9118 2432 9515
rect 1294 9112 2432 9118
rect 2536 9515 3674 9521
rect 2536 9118 2548 9515
rect 3662 9118 3674 9515
rect 2536 9112 3674 9118
rect 3778 9515 4916 9521
rect 3778 9118 3790 9515
rect 4904 9118 4916 9515
rect 3778 9112 4916 9118
rect -4916 8978 -3778 8984
rect -4916 8581 -4904 8978
rect -3790 8581 -3778 8978
rect -4916 8575 -3778 8581
rect -3674 8978 -2536 8984
rect -3674 8581 -3662 8978
rect -2548 8581 -2536 8978
rect -3674 8575 -2536 8581
rect -2432 8978 -1294 8984
rect -2432 8581 -2420 8978
rect -1306 8581 -1294 8978
rect -2432 8575 -1294 8581
rect -1190 8978 -52 8984
rect -1190 8581 -1178 8978
rect -64 8581 -52 8978
rect -1190 8575 -52 8581
rect 52 8978 1190 8984
rect 52 8581 64 8978
rect 1178 8581 1190 8978
rect 52 8575 1190 8581
rect 1294 8978 2432 8984
rect 1294 8581 1306 8978
rect 2420 8581 2432 8978
rect 1294 8575 2432 8581
rect 2536 8978 3674 8984
rect 2536 8581 2548 8978
rect 3662 8581 3674 8978
rect 2536 8575 3674 8581
rect 3778 8978 4916 8984
rect 3778 8581 3790 8978
rect 4904 8581 4916 8978
rect 3778 8575 4916 8581
rect -4916 8007 -3778 8013
rect -4916 7610 -4904 8007
rect -3790 7610 -3778 8007
rect -4916 7604 -3778 7610
rect -3674 8007 -2536 8013
rect -3674 7610 -3662 8007
rect -2548 7610 -2536 8007
rect -3674 7604 -2536 7610
rect -2432 8007 -1294 8013
rect -2432 7610 -2420 8007
rect -1306 7610 -1294 8007
rect -2432 7604 -1294 7610
rect -1190 8007 -52 8013
rect -1190 7610 -1178 8007
rect -64 7610 -52 8007
rect -1190 7604 -52 7610
rect 52 8007 1190 8013
rect 52 7610 64 8007
rect 1178 7610 1190 8007
rect 52 7604 1190 7610
rect 1294 8007 2432 8013
rect 1294 7610 1306 8007
rect 2420 7610 2432 8007
rect 1294 7604 2432 7610
rect 2536 8007 3674 8013
rect 2536 7610 2548 8007
rect 3662 7610 3674 8007
rect 2536 7604 3674 7610
rect 3778 8007 4916 8013
rect 3778 7610 3790 8007
rect 4904 7610 4916 8007
rect 3778 7604 4916 7610
rect -4916 7470 -3778 7476
rect -4916 7073 -4904 7470
rect -3790 7073 -3778 7470
rect -4916 7067 -3778 7073
rect -3674 7470 -2536 7476
rect -3674 7073 -3662 7470
rect -2548 7073 -2536 7470
rect -3674 7067 -2536 7073
rect -2432 7470 -1294 7476
rect -2432 7073 -2420 7470
rect -1306 7073 -1294 7470
rect -2432 7067 -1294 7073
rect -1190 7470 -52 7476
rect -1190 7073 -1178 7470
rect -64 7073 -52 7470
rect -1190 7067 -52 7073
rect 52 7470 1190 7476
rect 52 7073 64 7470
rect 1178 7073 1190 7470
rect 52 7067 1190 7073
rect 1294 7470 2432 7476
rect 1294 7073 1306 7470
rect 2420 7073 2432 7470
rect 1294 7067 2432 7073
rect 2536 7470 3674 7476
rect 2536 7073 2548 7470
rect 3662 7073 3674 7470
rect 2536 7067 3674 7073
rect 3778 7470 4916 7476
rect 3778 7073 3790 7470
rect 4904 7073 4916 7470
rect 3778 7067 4916 7073
rect -4916 6499 -3778 6505
rect -4916 6102 -4904 6499
rect -3790 6102 -3778 6499
rect -4916 6096 -3778 6102
rect -3674 6499 -2536 6505
rect -3674 6102 -3662 6499
rect -2548 6102 -2536 6499
rect -3674 6096 -2536 6102
rect -2432 6499 -1294 6505
rect -2432 6102 -2420 6499
rect -1306 6102 -1294 6499
rect -2432 6096 -1294 6102
rect -1190 6499 -52 6505
rect -1190 6102 -1178 6499
rect -64 6102 -52 6499
rect -1190 6096 -52 6102
rect 52 6499 1190 6505
rect 52 6102 64 6499
rect 1178 6102 1190 6499
rect 52 6096 1190 6102
rect 1294 6499 2432 6505
rect 1294 6102 1306 6499
rect 2420 6102 2432 6499
rect 1294 6096 2432 6102
rect 2536 6499 3674 6505
rect 2536 6102 2548 6499
rect 3662 6102 3674 6499
rect 2536 6096 3674 6102
rect 3778 6499 4916 6505
rect 3778 6102 3790 6499
rect 4904 6102 4916 6499
rect 3778 6096 4916 6102
rect -4916 5962 -3778 5968
rect -4916 5565 -4904 5962
rect -3790 5565 -3778 5962
rect -4916 5559 -3778 5565
rect -3674 5962 -2536 5968
rect -3674 5565 -3662 5962
rect -2548 5565 -2536 5962
rect -3674 5559 -2536 5565
rect -2432 5962 -1294 5968
rect -2432 5565 -2420 5962
rect -1306 5565 -1294 5962
rect -2432 5559 -1294 5565
rect -1190 5962 -52 5968
rect -1190 5565 -1178 5962
rect -64 5565 -52 5962
rect -1190 5559 -52 5565
rect 52 5962 1190 5968
rect 52 5565 64 5962
rect 1178 5565 1190 5962
rect 52 5559 1190 5565
rect 1294 5962 2432 5968
rect 1294 5565 1306 5962
rect 2420 5565 2432 5962
rect 1294 5559 2432 5565
rect 2536 5962 3674 5968
rect 2536 5565 2548 5962
rect 3662 5565 3674 5962
rect 2536 5559 3674 5565
rect 3778 5962 4916 5968
rect 3778 5565 3790 5962
rect 4904 5565 4916 5962
rect 3778 5559 4916 5565
rect -4916 4991 -3778 4997
rect -4916 4594 -4904 4991
rect -3790 4594 -3778 4991
rect -4916 4588 -3778 4594
rect -3674 4991 -2536 4997
rect -3674 4594 -3662 4991
rect -2548 4594 -2536 4991
rect -3674 4588 -2536 4594
rect -2432 4991 -1294 4997
rect -2432 4594 -2420 4991
rect -1306 4594 -1294 4991
rect -2432 4588 -1294 4594
rect -1190 4991 -52 4997
rect -1190 4594 -1178 4991
rect -64 4594 -52 4991
rect -1190 4588 -52 4594
rect 52 4991 1190 4997
rect 52 4594 64 4991
rect 1178 4594 1190 4991
rect 52 4588 1190 4594
rect 1294 4991 2432 4997
rect 1294 4594 1306 4991
rect 2420 4594 2432 4991
rect 1294 4588 2432 4594
rect 2536 4991 3674 4997
rect 2536 4594 2548 4991
rect 3662 4594 3674 4991
rect 2536 4588 3674 4594
rect 3778 4991 4916 4997
rect 3778 4594 3790 4991
rect 4904 4594 4916 4991
rect 3778 4588 4916 4594
rect -4916 4454 -3778 4460
rect -4916 4057 -4904 4454
rect -3790 4057 -3778 4454
rect -4916 4051 -3778 4057
rect -3674 4454 -2536 4460
rect -3674 4057 -3662 4454
rect -2548 4057 -2536 4454
rect -3674 4051 -2536 4057
rect -2432 4454 -1294 4460
rect -2432 4057 -2420 4454
rect -1306 4057 -1294 4454
rect -2432 4051 -1294 4057
rect -1190 4454 -52 4460
rect -1190 4057 -1178 4454
rect -64 4057 -52 4454
rect -1190 4051 -52 4057
rect 52 4454 1190 4460
rect 52 4057 64 4454
rect 1178 4057 1190 4454
rect 52 4051 1190 4057
rect 1294 4454 2432 4460
rect 1294 4057 1306 4454
rect 2420 4057 2432 4454
rect 1294 4051 2432 4057
rect 2536 4454 3674 4460
rect 2536 4057 2548 4454
rect 3662 4057 3674 4454
rect 2536 4051 3674 4057
rect 3778 4454 4916 4460
rect 3778 4057 3790 4454
rect 4904 4057 4916 4454
rect 3778 4051 4916 4057
rect -4916 3483 -3778 3489
rect -4916 3086 -4904 3483
rect -3790 3086 -3778 3483
rect -4916 3080 -3778 3086
rect -3674 3483 -2536 3489
rect -3674 3086 -3662 3483
rect -2548 3086 -2536 3483
rect -3674 3080 -2536 3086
rect -2432 3483 -1294 3489
rect -2432 3086 -2420 3483
rect -1306 3086 -1294 3483
rect -2432 3080 -1294 3086
rect -1190 3483 -52 3489
rect -1190 3086 -1178 3483
rect -64 3086 -52 3483
rect -1190 3080 -52 3086
rect 52 3483 1190 3489
rect 52 3086 64 3483
rect 1178 3086 1190 3483
rect 52 3080 1190 3086
rect 1294 3483 2432 3489
rect 1294 3086 1306 3483
rect 2420 3086 2432 3483
rect 1294 3080 2432 3086
rect 2536 3483 3674 3489
rect 2536 3086 2548 3483
rect 3662 3086 3674 3483
rect 2536 3080 3674 3086
rect 3778 3483 4916 3489
rect 3778 3086 3790 3483
rect 4904 3086 4916 3483
rect 3778 3080 4916 3086
rect -4916 2946 -3778 2952
rect -4916 2549 -4904 2946
rect -3790 2549 -3778 2946
rect -4916 2543 -3778 2549
rect -3674 2946 -2536 2952
rect -3674 2549 -3662 2946
rect -2548 2549 -2536 2946
rect -3674 2543 -2536 2549
rect -2432 2946 -1294 2952
rect -2432 2549 -2420 2946
rect -1306 2549 -1294 2946
rect -2432 2543 -1294 2549
rect -1190 2946 -52 2952
rect -1190 2549 -1178 2946
rect -64 2549 -52 2946
rect -1190 2543 -52 2549
rect 52 2946 1190 2952
rect 52 2549 64 2946
rect 1178 2549 1190 2946
rect 52 2543 1190 2549
rect 1294 2946 2432 2952
rect 1294 2549 1306 2946
rect 2420 2549 2432 2946
rect 1294 2543 2432 2549
rect 2536 2946 3674 2952
rect 2536 2549 2548 2946
rect 3662 2549 3674 2946
rect 2536 2543 3674 2549
rect 3778 2946 4916 2952
rect 3778 2549 3790 2946
rect 4904 2549 4916 2946
rect 3778 2543 4916 2549
rect -4916 1975 -3778 1981
rect -4916 1578 -4904 1975
rect -3790 1578 -3778 1975
rect -4916 1572 -3778 1578
rect -3674 1975 -2536 1981
rect -3674 1578 -3662 1975
rect -2548 1578 -2536 1975
rect -3674 1572 -2536 1578
rect -2432 1975 -1294 1981
rect -2432 1578 -2420 1975
rect -1306 1578 -1294 1975
rect -2432 1572 -1294 1578
rect -1190 1975 -52 1981
rect -1190 1578 -1178 1975
rect -64 1578 -52 1975
rect -1190 1572 -52 1578
rect 52 1975 1190 1981
rect 52 1578 64 1975
rect 1178 1578 1190 1975
rect 52 1572 1190 1578
rect 1294 1975 2432 1981
rect 1294 1578 1306 1975
rect 2420 1578 2432 1975
rect 1294 1572 2432 1578
rect 2536 1975 3674 1981
rect 2536 1578 2548 1975
rect 3662 1578 3674 1975
rect 2536 1572 3674 1578
rect 3778 1975 4916 1981
rect 3778 1578 3790 1975
rect 4904 1578 4916 1975
rect 3778 1572 4916 1578
rect -4916 1438 -3778 1444
rect -4916 1041 -4904 1438
rect -3790 1041 -3778 1438
rect -4916 1035 -3778 1041
rect -3674 1438 -2536 1444
rect -3674 1041 -3662 1438
rect -2548 1041 -2536 1438
rect -3674 1035 -2536 1041
rect -2432 1438 -1294 1444
rect -2432 1041 -2420 1438
rect -1306 1041 -1294 1438
rect -2432 1035 -1294 1041
rect -1190 1438 -52 1444
rect -1190 1041 -1178 1438
rect -64 1041 -52 1438
rect -1190 1035 -52 1041
rect 52 1438 1190 1444
rect 52 1041 64 1438
rect 1178 1041 1190 1438
rect 52 1035 1190 1041
rect 1294 1438 2432 1444
rect 1294 1041 1306 1438
rect 2420 1041 2432 1438
rect 1294 1035 2432 1041
rect 2536 1438 3674 1444
rect 2536 1041 2548 1438
rect 3662 1041 3674 1438
rect 2536 1035 3674 1041
rect 3778 1438 4916 1444
rect 3778 1041 3790 1438
rect 4904 1041 4916 1438
rect 3778 1035 4916 1041
rect -4916 467 -3778 473
rect -4916 70 -4904 467
rect -3790 70 -3778 467
rect -4916 64 -3778 70
rect -3674 467 -2536 473
rect -3674 70 -3662 467
rect -2548 70 -2536 467
rect -3674 64 -2536 70
rect -2432 467 -1294 473
rect -2432 70 -2420 467
rect -1306 70 -1294 467
rect -2432 64 -1294 70
rect -1190 467 -52 473
rect -1190 70 -1178 467
rect -64 70 -52 467
rect -1190 64 -52 70
rect 52 467 1190 473
rect 52 70 64 467
rect 1178 70 1190 467
rect 52 64 1190 70
rect 1294 467 2432 473
rect 1294 70 1306 467
rect 2420 70 2432 467
rect 1294 64 2432 70
rect 2536 467 3674 473
rect 2536 70 2548 467
rect 3662 70 3674 467
rect 2536 64 3674 70
rect 3778 467 4916 473
rect 3778 70 3790 467
rect 4904 70 4916 467
rect 3778 64 4916 70
rect -4916 -70 -3778 -64
rect -4916 -467 -4904 -70
rect -3790 -467 -3778 -70
rect -4916 -473 -3778 -467
rect -3674 -70 -2536 -64
rect -3674 -467 -3662 -70
rect -2548 -467 -2536 -70
rect -3674 -473 -2536 -467
rect -2432 -70 -1294 -64
rect -2432 -467 -2420 -70
rect -1306 -467 -1294 -70
rect -2432 -473 -1294 -467
rect -1190 -70 -52 -64
rect -1190 -467 -1178 -70
rect -64 -467 -52 -70
rect -1190 -473 -52 -467
rect 52 -70 1190 -64
rect 52 -467 64 -70
rect 1178 -467 1190 -70
rect 52 -473 1190 -467
rect 1294 -70 2432 -64
rect 1294 -467 1306 -70
rect 2420 -467 2432 -70
rect 1294 -473 2432 -467
rect 2536 -70 3674 -64
rect 2536 -467 2548 -70
rect 3662 -467 3674 -70
rect 2536 -473 3674 -467
rect 3778 -70 4916 -64
rect 3778 -467 3790 -70
rect 4904 -467 4916 -70
rect 3778 -473 4916 -467
rect -4916 -1041 -3778 -1035
rect -4916 -1438 -4904 -1041
rect -3790 -1438 -3778 -1041
rect -4916 -1444 -3778 -1438
rect -3674 -1041 -2536 -1035
rect -3674 -1438 -3662 -1041
rect -2548 -1438 -2536 -1041
rect -3674 -1444 -2536 -1438
rect -2432 -1041 -1294 -1035
rect -2432 -1438 -2420 -1041
rect -1306 -1438 -1294 -1041
rect -2432 -1444 -1294 -1438
rect -1190 -1041 -52 -1035
rect -1190 -1438 -1178 -1041
rect -64 -1438 -52 -1041
rect -1190 -1444 -52 -1438
rect 52 -1041 1190 -1035
rect 52 -1438 64 -1041
rect 1178 -1438 1190 -1041
rect 52 -1444 1190 -1438
rect 1294 -1041 2432 -1035
rect 1294 -1438 1306 -1041
rect 2420 -1438 2432 -1041
rect 1294 -1444 2432 -1438
rect 2536 -1041 3674 -1035
rect 2536 -1438 2548 -1041
rect 3662 -1438 3674 -1041
rect 2536 -1444 3674 -1438
rect 3778 -1041 4916 -1035
rect 3778 -1438 3790 -1041
rect 4904 -1438 4916 -1041
rect 3778 -1444 4916 -1438
rect -4916 -1578 -3778 -1572
rect -4916 -1975 -4904 -1578
rect -3790 -1975 -3778 -1578
rect -4916 -1981 -3778 -1975
rect -3674 -1578 -2536 -1572
rect -3674 -1975 -3662 -1578
rect -2548 -1975 -2536 -1578
rect -3674 -1981 -2536 -1975
rect -2432 -1578 -1294 -1572
rect -2432 -1975 -2420 -1578
rect -1306 -1975 -1294 -1578
rect -2432 -1981 -1294 -1975
rect -1190 -1578 -52 -1572
rect -1190 -1975 -1178 -1578
rect -64 -1975 -52 -1578
rect -1190 -1981 -52 -1975
rect 52 -1578 1190 -1572
rect 52 -1975 64 -1578
rect 1178 -1975 1190 -1578
rect 52 -1981 1190 -1975
rect 1294 -1578 2432 -1572
rect 1294 -1975 1306 -1578
rect 2420 -1975 2432 -1578
rect 1294 -1981 2432 -1975
rect 2536 -1578 3674 -1572
rect 2536 -1975 2548 -1578
rect 3662 -1975 3674 -1578
rect 2536 -1981 3674 -1975
rect 3778 -1578 4916 -1572
rect 3778 -1975 3790 -1578
rect 4904 -1975 4916 -1578
rect 3778 -1981 4916 -1975
rect -4916 -2549 -3778 -2543
rect -4916 -2946 -4904 -2549
rect -3790 -2946 -3778 -2549
rect -4916 -2952 -3778 -2946
rect -3674 -2549 -2536 -2543
rect -3674 -2946 -3662 -2549
rect -2548 -2946 -2536 -2549
rect -3674 -2952 -2536 -2946
rect -2432 -2549 -1294 -2543
rect -2432 -2946 -2420 -2549
rect -1306 -2946 -1294 -2549
rect -2432 -2952 -1294 -2946
rect -1190 -2549 -52 -2543
rect -1190 -2946 -1178 -2549
rect -64 -2946 -52 -2549
rect -1190 -2952 -52 -2946
rect 52 -2549 1190 -2543
rect 52 -2946 64 -2549
rect 1178 -2946 1190 -2549
rect 52 -2952 1190 -2946
rect 1294 -2549 2432 -2543
rect 1294 -2946 1306 -2549
rect 2420 -2946 2432 -2549
rect 1294 -2952 2432 -2946
rect 2536 -2549 3674 -2543
rect 2536 -2946 2548 -2549
rect 3662 -2946 3674 -2549
rect 2536 -2952 3674 -2946
rect 3778 -2549 4916 -2543
rect 3778 -2946 3790 -2549
rect 4904 -2946 4916 -2549
rect 3778 -2952 4916 -2946
rect -4916 -3086 -3778 -3080
rect -4916 -3483 -4904 -3086
rect -3790 -3483 -3778 -3086
rect -4916 -3489 -3778 -3483
rect -3674 -3086 -2536 -3080
rect -3674 -3483 -3662 -3086
rect -2548 -3483 -2536 -3086
rect -3674 -3489 -2536 -3483
rect -2432 -3086 -1294 -3080
rect -2432 -3483 -2420 -3086
rect -1306 -3483 -1294 -3086
rect -2432 -3489 -1294 -3483
rect -1190 -3086 -52 -3080
rect -1190 -3483 -1178 -3086
rect -64 -3483 -52 -3086
rect -1190 -3489 -52 -3483
rect 52 -3086 1190 -3080
rect 52 -3483 64 -3086
rect 1178 -3483 1190 -3086
rect 52 -3489 1190 -3483
rect 1294 -3086 2432 -3080
rect 1294 -3483 1306 -3086
rect 2420 -3483 2432 -3086
rect 1294 -3489 2432 -3483
rect 2536 -3086 3674 -3080
rect 2536 -3483 2548 -3086
rect 3662 -3483 3674 -3086
rect 2536 -3489 3674 -3483
rect 3778 -3086 4916 -3080
rect 3778 -3483 3790 -3086
rect 4904 -3483 4916 -3086
rect 3778 -3489 4916 -3483
rect -4916 -4057 -3778 -4051
rect -4916 -4454 -4904 -4057
rect -3790 -4454 -3778 -4057
rect -4916 -4460 -3778 -4454
rect -3674 -4057 -2536 -4051
rect -3674 -4454 -3662 -4057
rect -2548 -4454 -2536 -4057
rect -3674 -4460 -2536 -4454
rect -2432 -4057 -1294 -4051
rect -2432 -4454 -2420 -4057
rect -1306 -4454 -1294 -4057
rect -2432 -4460 -1294 -4454
rect -1190 -4057 -52 -4051
rect -1190 -4454 -1178 -4057
rect -64 -4454 -52 -4057
rect -1190 -4460 -52 -4454
rect 52 -4057 1190 -4051
rect 52 -4454 64 -4057
rect 1178 -4454 1190 -4057
rect 52 -4460 1190 -4454
rect 1294 -4057 2432 -4051
rect 1294 -4454 1306 -4057
rect 2420 -4454 2432 -4057
rect 1294 -4460 2432 -4454
rect 2536 -4057 3674 -4051
rect 2536 -4454 2548 -4057
rect 3662 -4454 3674 -4057
rect 2536 -4460 3674 -4454
rect 3778 -4057 4916 -4051
rect 3778 -4454 3790 -4057
rect 4904 -4454 4916 -4057
rect 3778 -4460 4916 -4454
rect -4916 -4594 -3778 -4588
rect -4916 -4991 -4904 -4594
rect -3790 -4991 -3778 -4594
rect -4916 -4997 -3778 -4991
rect -3674 -4594 -2536 -4588
rect -3674 -4991 -3662 -4594
rect -2548 -4991 -2536 -4594
rect -3674 -4997 -2536 -4991
rect -2432 -4594 -1294 -4588
rect -2432 -4991 -2420 -4594
rect -1306 -4991 -1294 -4594
rect -2432 -4997 -1294 -4991
rect -1190 -4594 -52 -4588
rect -1190 -4991 -1178 -4594
rect -64 -4991 -52 -4594
rect -1190 -4997 -52 -4991
rect 52 -4594 1190 -4588
rect 52 -4991 64 -4594
rect 1178 -4991 1190 -4594
rect 52 -4997 1190 -4991
rect 1294 -4594 2432 -4588
rect 1294 -4991 1306 -4594
rect 2420 -4991 2432 -4594
rect 1294 -4997 2432 -4991
rect 2536 -4594 3674 -4588
rect 2536 -4991 2548 -4594
rect 3662 -4991 3674 -4594
rect 2536 -4997 3674 -4991
rect 3778 -4594 4916 -4588
rect 3778 -4991 3790 -4594
rect 4904 -4991 4916 -4594
rect 3778 -4997 4916 -4991
rect -4916 -5565 -3778 -5559
rect -4916 -5962 -4904 -5565
rect -3790 -5962 -3778 -5565
rect -4916 -5968 -3778 -5962
rect -3674 -5565 -2536 -5559
rect -3674 -5962 -3662 -5565
rect -2548 -5962 -2536 -5565
rect -3674 -5968 -2536 -5962
rect -2432 -5565 -1294 -5559
rect -2432 -5962 -2420 -5565
rect -1306 -5962 -1294 -5565
rect -2432 -5968 -1294 -5962
rect -1190 -5565 -52 -5559
rect -1190 -5962 -1178 -5565
rect -64 -5962 -52 -5565
rect -1190 -5968 -52 -5962
rect 52 -5565 1190 -5559
rect 52 -5962 64 -5565
rect 1178 -5962 1190 -5565
rect 52 -5968 1190 -5962
rect 1294 -5565 2432 -5559
rect 1294 -5962 1306 -5565
rect 2420 -5962 2432 -5565
rect 1294 -5968 2432 -5962
rect 2536 -5565 3674 -5559
rect 2536 -5962 2548 -5565
rect 3662 -5962 3674 -5565
rect 2536 -5968 3674 -5962
rect 3778 -5565 4916 -5559
rect 3778 -5962 3790 -5565
rect 4904 -5962 4916 -5565
rect 3778 -5968 4916 -5962
rect -4916 -6102 -3778 -6096
rect -4916 -6499 -4904 -6102
rect -3790 -6499 -3778 -6102
rect -4916 -6505 -3778 -6499
rect -3674 -6102 -2536 -6096
rect -3674 -6499 -3662 -6102
rect -2548 -6499 -2536 -6102
rect -3674 -6505 -2536 -6499
rect -2432 -6102 -1294 -6096
rect -2432 -6499 -2420 -6102
rect -1306 -6499 -1294 -6102
rect -2432 -6505 -1294 -6499
rect -1190 -6102 -52 -6096
rect -1190 -6499 -1178 -6102
rect -64 -6499 -52 -6102
rect -1190 -6505 -52 -6499
rect 52 -6102 1190 -6096
rect 52 -6499 64 -6102
rect 1178 -6499 1190 -6102
rect 52 -6505 1190 -6499
rect 1294 -6102 2432 -6096
rect 1294 -6499 1306 -6102
rect 2420 -6499 2432 -6102
rect 1294 -6505 2432 -6499
rect 2536 -6102 3674 -6096
rect 2536 -6499 2548 -6102
rect 3662 -6499 3674 -6102
rect 2536 -6505 3674 -6499
rect 3778 -6102 4916 -6096
rect 3778 -6499 3790 -6102
rect 4904 -6499 4916 -6102
rect 3778 -6505 4916 -6499
rect -4916 -7073 -3778 -7067
rect -4916 -7470 -4904 -7073
rect -3790 -7470 -3778 -7073
rect -4916 -7476 -3778 -7470
rect -3674 -7073 -2536 -7067
rect -3674 -7470 -3662 -7073
rect -2548 -7470 -2536 -7073
rect -3674 -7476 -2536 -7470
rect -2432 -7073 -1294 -7067
rect -2432 -7470 -2420 -7073
rect -1306 -7470 -1294 -7073
rect -2432 -7476 -1294 -7470
rect -1190 -7073 -52 -7067
rect -1190 -7470 -1178 -7073
rect -64 -7470 -52 -7073
rect -1190 -7476 -52 -7470
rect 52 -7073 1190 -7067
rect 52 -7470 64 -7073
rect 1178 -7470 1190 -7073
rect 52 -7476 1190 -7470
rect 1294 -7073 2432 -7067
rect 1294 -7470 1306 -7073
rect 2420 -7470 2432 -7073
rect 1294 -7476 2432 -7470
rect 2536 -7073 3674 -7067
rect 2536 -7470 2548 -7073
rect 3662 -7470 3674 -7073
rect 2536 -7476 3674 -7470
rect 3778 -7073 4916 -7067
rect 3778 -7470 3790 -7073
rect 4904 -7470 4916 -7073
rect 3778 -7476 4916 -7470
rect -4916 -7610 -3778 -7604
rect -4916 -8007 -4904 -7610
rect -3790 -8007 -3778 -7610
rect -4916 -8013 -3778 -8007
rect -3674 -7610 -2536 -7604
rect -3674 -8007 -3662 -7610
rect -2548 -8007 -2536 -7610
rect -3674 -8013 -2536 -8007
rect -2432 -7610 -1294 -7604
rect -2432 -8007 -2420 -7610
rect -1306 -8007 -1294 -7610
rect -2432 -8013 -1294 -8007
rect -1190 -7610 -52 -7604
rect -1190 -8007 -1178 -7610
rect -64 -8007 -52 -7610
rect -1190 -8013 -52 -8007
rect 52 -7610 1190 -7604
rect 52 -8007 64 -7610
rect 1178 -8007 1190 -7610
rect 52 -8013 1190 -8007
rect 1294 -7610 2432 -7604
rect 1294 -8007 1306 -7610
rect 2420 -8007 2432 -7610
rect 1294 -8013 2432 -8007
rect 2536 -7610 3674 -7604
rect 2536 -8007 2548 -7610
rect 3662 -8007 3674 -7610
rect 2536 -8013 3674 -8007
rect 3778 -7610 4916 -7604
rect 3778 -8007 3790 -7610
rect 4904 -8007 4916 -7610
rect 3778 -8013 4916 -8007
rect -4916 -8581 -3778 -8575
rect -4916 -8978 -4904 -8581
rect -3790 -8978 -3778 -8581
rect -4916 -8984 -3778 -8978
rect -3674 -8581 -2536 -8575
rect -3674 -8978 -3662 -8581
rect -2548 -8978 -2536 -8581
rect -3674 -8984 -2536 -8978
rect -2432 -8581 -1294 -8575
rect -2432 -8978 -2420 -8581
rect -1306 -8978 -1294 -8581
rect -2432 -8984 -1294 -8978
rect -1190 -8581 -52 -8575
rect -1190 -8978 -1178 -8581
rect -64 -8978 -52 -8581
rect -1190 -8984 -52 -8978
rect 52 -8581 1190 -8575
rect 52 -8978 64 -8581
rect 1178 -8978 1190 -8581
rect 52 -8984 1190 -8978
rect 1294 -8581 2432 -8575
rect 1294 -8978 1306 -8581
rect 2420 -8978 2432 -8581
rect 1294 -8984 2432 -8978
rect 2536 -8581 3674 -8575
rect 2536 -8978 2548 -8581
rect 3662 -8978 3674 -8581
rect 2536 -8984 3674 -8978
rect 3778 -8581 4916 -8575
rect 3778 -8978 3790 -8581
rect 4904 -8978 4916 -8581
rect 3778 -8984 4916 -8978
rect -4916 -9118 -3778 -9112
rect -4916 -9515 -4904 -9118
rect -3790 -9515 -3778 -9118
rect -4916 -9521 -3778 -9515
rect -3674 -9118 -2536 -9112
rect -3674 -9515 -3662 -9118
rect -2548 -9515 -2536 -9118
rect -3674 -9521 -2536 -9515
rect -2432 -9118 -1294 -9112
rect -2432 -9515 -2420 -9118
rect -1306 -9515 -1294 -9118
rect -2432 -9521 -1294 -9515
rect -1190 -9118 -52 -9112
rect -1190 -9515 -1178 -9118
rect -64 -9515 -52 -9118
rect -1190 -9521 -52 -9515
rect 52 -9118 1190 -9112
rect 52 -9515 64 -9118
rect 1178 -9515 1190 -9118
rect 52 -9521 1190 -9515
rect 1294 -9118 2432 -9112
rect 1294 -9515 1306 -9118
rect 2420 -9515 2432 -9118
rect 1294 -9521 2432 -9515
rect 2536 -9118 3674 -9112
rect 2536 -9515 2548 -9118
rect 3662 -9515 3674 -9118
rect 2536 -9521 3674 -9515
rect 3778 -9118 4916 -9112
rect 3778 -9515 3790 -9118
rect 4904 -9515 4916 -9118
rect 3778 -9521 4916 -9515
rect -4916 -10089 -3778 -10083
rect -4916 -10486 -4904 -10089
rect -3790 -10486 -3778 -10089
rect -4916 -10492 -3778 -10486
rect -3674 -10089 -2536 -10083
rect -3674 -10486 -3662 -10089
rect -2548 -10486 -2536 -10089
rect -3674 -10492 -2536 -10486
rect -2432 -10089 -1294 -10083
rect -2432 -10486 -2420 -10089
rect -1306 -10486 -1294 -10089
rect -2432 -10492 -1294 -10486
rect -1190 -10089 -52 -10083
rect -1190 -10486 -1178 -10089
rect -64 -10486 -52 -10089
rect -1190 -10492 -52 -10486
rect 52 -10089 1190 -10083
rect 52 -10486 64 -10089
rect 1178 -10486 1190 -10089
rect 52 -10492 1190 -10486
rect 1294 -10089 2432 -10083
rect 1294 -10486 1306 -10089
rect 2420 -10486 2432 -10089
rect 1294 -10492 2432 -10486
rect 2536 -10089 3674 -10083
rect 2536 -10486 2548 -10089
rect 3662 -10486 3674 -10089
rect 2536 -10492 3674 -10486
rect 3778 -10089 4916 -10083
rect 3778 -10486 3790 -10089
rect 4904 -10486 4916 -10089
rect 3778 -10492 4916 -10486
rect -4916 -10626 -3778 -10620
rect -4916 -11023 -4904 -10626
rect -3790 -11023 -3778 -10626
rect -4916 -11029 -3778 -11023
rect -3674 -10626 -2536 -10620
rect -3674 -11023 -3662 -10626
rect -2548 -11023 -2536 -10626
rect -3674 -11029 -2536 -11023
rect -2432 -10626 -1294 -10620
rect -2432 -11023 -2420 -10626
rect -1306 -11023 -1294 -10626
rect -2432 -11029 -1294 -11023
rect -1190 -10626 -52 -10620
rect -1190 -11023 -1178 -10626
rect -64 -11023 -52 -10626
rect -1190 -11029 -52 -11023
rect 52 -10626 1190 -10620
rect 52 -11023 64 -10626
rect 1178 -11023 1190 -10626
rect 52 -11029 1190 -11023
rect 1294 -10626 2432 -10620
rect 1294 -11023 1306 -10626
rect 2420 -11023 2432 -10626
rect 1294 -11029 2432 -11023
rect 2536 -10626 3674 -10620
rect 2536 -11023 2548 -10626
rect 3662 -11023 3674 -10626
rect 2536 -11029 3674 -11023
rect 3778 -10626 4916 -10620
rect 3778 -11023 3790 -10626
rect 4904 -11023 4916 -10626
rect 3778 -11029 4916 -11023
rect -4916 -11597 -3778 -11591
rect -4916 -11994 -4904 -11597
rect -3790 -11994 -3778 -11597
rect -4916 -12000 -3778 -11994
rect -3674 -11597 -2536 -11591
rect -3674 -11994 -3662 -11597
rect -2548 -11994 -2536 -11597
rect -3674 -12000 -2536 -11994
rect -2432 -11597 -1294 -11591
rect -2432 -11994 -2420 -11597
rect -1306 -11994 -1294 -11597
rect -2432 -12000 -1294 -11994
rect -1190 -11597 -52 -11591
rect -1190 -11994 -1178 -11597
rect -64 -11994 -52 -11597
rect -1190 -12000 -52 -11994
rect 52 -11597 1190 -11591
rect 52 -11994 64 -11597
rect 1178 -11994 1190 -11597
rect 52 -12000 1190 -11994
rect 1294 -11597 2432 -11591
rect 1294 -11994 1306 -11597
rect 2420 -11994 2432 -11597
rect 1294 -12000 2432 -11994
rect 2536 -11597 3674 -11591
rect 2536 -11994 2548 -11597
rect 3662 -11994 3674 -11597
rect 2536 -12000 3674 -11994
rect 3778 -11597 4916 -11591
rect 3778 -11994 3790 -11597
rect 4904 -11994 4916 -11597
rect 3778 -12000 4916 -11994
rect -4916 -12134 -3778 -12128
rect -4916 -12531 -4904 -12134
rect -3790 -12531 -3778 -12134
rect -4916 -12537 -3778 -12531
rect -3674 -12134 -2536 -12128
rect -3674 -12531 -3662 -12134
rect -2548 -12531 -2536 -12134
rect -3674 -12537 -2536 -12531
rect -2432 -12134 -1294 -12128
rect -2432 -12531 -2420 -12134
rect -1306 -12531 -1294 -12134
rect -2432 -12537 -1294 -12531
rect -1190 -12134 -52 -12128
rect -1190 -12531 -1178 -12134
rect -64 -12531 -52 -12134
rect -1190 -12537 -52 -12531
rect 52 -12134 1190 -12128
rect 52 -12531 64 -12134
rect 1178 -12531 1190 -12134
rect 52 -12537 1190 -12531
rect 1294 -12134 2432 -12128
rect 1294 -12531 1306 -12134
rect 2420 -12531 2432 -12134
rect 1294 -12537 2432 -12531
rect 2536 -12134 3674 -12128
rect 2536 -12531 2548 -12134
rect 3662 -12531 3674 -12134
rect 2536 -12537 3674 -12531
rect 3778 -12134 4916 -12128
rect 3778 -12531 3790 -12134
rect 4904 -12531 4916 -12134
rect 3778 -12537 4916 -12531
rect -4916 -13105 -3778 -13099
rect -4916 -13502 -4904 -13105
rect -3790 -13502 -3778 -13105
rect -4916 -13508 -3778 -13502
rect -3674 -13105 -2536 -13099
rect -3674 -13502 -3662 -13105
rect -2548 -13502 -2536 -13105
rect -3674 -13508 -2536 -13502
rect -2432 -13105 -1294 -13099
rect -2432 -13502 -2420 -13105
rect -1306 -13502 -1294 -13105
rect -2432 -13508 -1294 -13502
rect -1190 -13105 -52 -13099
rect -1190 -13502 -1178 -13105
rect -64 -13502 -52 -13105
rect -1190 -13508 -52 -13502
rect 52 -13105 1190 -13099
rect 52 -13502 64 -13105
rect 1178 -13502 1190 -13105
rect 52 -13508 1190 -13502
rect 1294 -13105 2432 -13099
rect 1294 -13502 1306 -13105
rect 2420 -13502 2432 -13105
rect 1294 -13508 2432 -13502
rect 2536 -13105 3674 -13099
rect 2536 -13502 2548 -13105
rect 3662 -13502 3674 -13105
rect 2536 -13508 3674 -13502
rect 3778 -13105 4916 -13099
rect 3778 -13502 3790 -13105
rect 4904 -13502 4916 -13105
rect 3778 -13508 4916 -13502
<< properties >>
string FIXED_BBOX -5033 -13633 5033 13633
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 2.857 m 18 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 1.062k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
