magic
tech sky130A
magscale 1 2
timestamp 1709390584
<< metal3 >>
rect -1000 7550 1000 7607
rect -1000 -7607 1000 -7550
<< rmetal3 >>
rect -1000 -7550 1000 7550
<< properties >>
string gencell sky130_fd_pr__res_generic_m3
string library sky130
string parameters w 10.0 l 75.5 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 354.849m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
