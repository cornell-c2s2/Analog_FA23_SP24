magic
tech sky130A
magscale 1 2
timestamp 1716869746
<< pwell >>
rect -5086 -850 5086 850
<< psubdiff >>
rect -5050 780 -4954 814
rect 4954 780 5050 814
rect -5050 718 -5016 780
rect 5016 718 5050 780
rect -5050 -780 -5016 -718
rect 5016 -780 5050 -718
rect -5050 -814 -4954 -780
rect 4954 -814 5050 -780
<< psubdiffcont >>
rect -4954 780 4954 814
rect -5050 -718 -5016 718
rect 5016 -718 5050 718
rect -4954 -814 4954 -780
<< xpolycontact >>
rect -4920 252 -3774 684
rect -4920 -684 -3774 -252
rect -3678 252 -2532 684
rect -3678 -684 -2532 -252
rect -2436 252 -1290 684
rect -2436 -684 -1290 -252
rect -1194 252 -48 684
rect -1194 -684 -48 -252
rect 48 252 1194 684
rect 48 -684 1194 -252
rect 1290 252 2436 684
rect 1290 -684 2436 -252
rect 2532 252 3678 684
rect 2532 -684 3678 -252
rect 3774 252 4920 684
rect 3774 -684 4920 -252
<< xpolyres >>
rect -4920 -252 -3774 252
rect -3678 -252 -2532 252
rect -2436 -252 -1290 252
rect -1194 -252 -48 252
rect 48 -252 1194 252
rect 1290 -252 2436 252
rect 2532 -252 3678 252
rect 3774 -252 4920 252
<< locali >>
rect -5050 780 -4954 814
rect 4954 780 5050 814
rect -5050 718 -5016 780
rect 5016 718 5050 780
rect -5050 -780 -5016 -718
rect 5016 -780 5050 -718
rect -5050 -814 -4954 -780
rect 4954 -814 5050 -780
<< viali >>
rect -4904 269 -3790 666
rect -3662 269 -2548 666
rect -2420 269 -1306 666
rect -1178 269 -64 666
rect 64 269 1178 666
rect 1306 269 2420 666
rect 2548 269 3662 666
rect 3790 269 4904 666
rect -4904 -666 -3790 -269
rect -3662 -666 -2548 -269
rect -2420 -666 -1306 -269
rect -1178 -666 -64 -269
rect 64 -666 1178 -269
rect 1306 -666 2420 -269
rect 2548 -666 3662 -269
rect 3790 -666 4904 -269
<< metal1 >>
rect -4916 666 -3778 672
rect -4916 269 -4904 666
rect -3790 269 -3778 666
rect -4916 263 -3778 269
rect -3674 666 -2536 672
rect -3674 269 -3662 666
rect -2548 269 -2536 666
rect -3674 263 -2536 269
rect -2432 666 -1294 672
rect -2432 269 -2420 666
rect -1306 269 -1294 666
rect -2432 263 -1294 269
rect -1190 666 -52 672
rect -1190 269 -1178 666
rect -64 269 -52 666
rect -1190 263 -52 269
rect 52 666 1190 672
rect 52 269 64 666
rect 1178 269 1190 666
rect 52 263 1190 269
rect 1294 666 2432 672
rect 1294 269 1306 666
rect 2420 269 2432 666
rect 1294 263 2432 269
rect 2536 666 3674 672
rect 2536 269 2548 666
rect 3662 269 3674 666
rect 2536 263 3674 269
rect 3778 666 4916 672
rect 3778 269 3790 666
rect 4904 269 4916 666
rect 3778 263 4916 269
rect -4916 -269 -3778 -263
rect -4916 -666 -4904 -269
rect -3790 -666 -3778 -269
rect -4916 -672 -3778 -666
rect -3674 -269 -2536 -263
rect -3674 -666 -3662 -269
rect -2548 -666 -2536 -269
rect -3674 -672 -2536 -666
rect -2432 -269 -1294 -263
rect -2432 -666 -2420 -269
rect -1306 -666 -1294 -269
rect -2432 -672 -1294 -666
rect -1190 -269 -52 -263
rect -1190 -666 -1178 -269
rect -64 -666 -52 -269
rect -1190 -672 -52 -666
rect 52 -269 1190 -263
rect 52 -666 64 -269
rect 1178 -666 1190 -269
rect 52 -672 1190 -666
rect 1294 -269 2432 -263
rect 1294 -666 1306 -269
rect 2420 -666 2432 -269
rect 1294 -672 2432 -666
rect 2536 -269 3674 -263
rect 2536 -666 2548 -269
rect 3662 -666 3674 -269
rect 2536 -672 3674 -666
rect 3778 -269 4916 -263
rect 3778 -666 3790 -269
rect 4904 -666 4916 -269
rect 3778 -672 4916 -666
<< properties >>
string FIXED_BBOX -5033 -797 5033 797
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 2.677 m 1 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 1.0k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
