magic
tech sky130A
timestamp 1717029187
<< metal1 >>
rect 19800 2400 20000 2600
rect 26600 2400 26800 2600
rect 32200 2400 32400 2600
rect 39000 2400 39200 2600
rect 47200 2400 47400 2600
rect 54000 2400 54200 2600
rect 60800 2400 61000 2600
rect 66400 2400 66600 2600
rect 73200 2400 73400 2600
rect 81400 2400 81600 2600
rect 18200 2600 18400 2800
rect 33800 2600 34000 2800
rect 40600 2600 40800 2800
rect 52400 2600 52600 2800
rect 68000 2600 68200 2800
rect 24800 2800 25000 3000
rect 27200 2800 27400 3000
rect 59000 2800 59200 3000
rect 61400 2800 61600 3000
rect 34200 3000 34400 3200
rect 52000 3000 52200 3200
rect 68400 3000 68600 3200
rect 38200 3200 38400 3400
rect 48000 3200 48200 3400
rect 72400 3200 72600 3400
rect 82200 3200 82400 3400
rect 17600 3400 17800 3600
rect 34400 3400 34600 3600
rect 51800 3400 52000 3600
rect 68600 3400 68800 3600
rect 27600 3600 27800 3800
rect 31200 3600 31400 3800
rect 65400 3600 65600 3800
rect 20800 3800 21000 4000
rect 31200 3800 31400 4000
rect 55000 3800 55200 4000
rect 65400 3800 65600 4000
rect 20800 4000 21000 4200
rect 38000 4000 38200 4200
rect 72200 4000 72400 4200
rect 82400 4000 82600 4200
rect 20800 4200 21000 4400
rect 38000 4200 38200 4400
rect 72200 4200 72400 4400
rect 82400 4200 82600 4400
rect 20800 4400 21000 4600
rect 38000 4400 38200 4600
rect 72200 4400 72400 4600
rect 82400 4400 82600 4600
rect 20800 4600 21000 4800
rect 38000 4600 38200 4800
rect 72200 4600 72400 4800
rect 82400 4600 82600 4800
rect 20800 4800 21000 5000
rect 38000 4800 38200 5000
rect 72200 4800 72400 5000
rect 82400 4800 82600 5000
rect 20800 5000 21000 5200
rect 38000 5000 38200 5200
rect 72200 5000 72400 5200
rect 82400 5000 82600 5200
rect 20800 5200 21000 5400
rect 38000 5200 38200 5400
rect 72200 5200 72400 5400
rect 82400 5200 82600 5400
rect 20800 5400 21000 5600
rect 38000 5400 38200 5600
rect 72200 5400 72400 5600
rect 82400 5400 82600 5600
rect 20800 5600 21000 5800
rect 38000 5600 38200 5800
rect 72200 5600 72400 5800
rect 82400 5600 82600 5800
rect 20800 5800 21000 6000
rect 38000 5800 38200 6000
rect 72200 5800 72400 6000
rect 82400 5800 82600 6000
rect 20800 6000 21000 6200
rect 38000 6000 38200 6200
rect 72200 6000 72400 6200
rect 82400 6000 82600 6200
rect 20800 6200 21000 6400
rect 38000 6200 38200 6400
rect 72200 6200 72400 6400
rect 82400 6200 82600 6400
rect 20800 6400 21000 6600
rect 38000 6400 38200 6600
rect 72200 6400 72400 6600
rect 82400 6400 82600 6600
rect 20800 6600 21000 6800
rect 38000 6600 38200 6800
rect 72200 6600 72400 6800
rect 82400 6600 82600 6800
rect 20800 6800 21000 7000
rect 38000 6800 38200 7000
rect 72200 6800 72400 7000
rect 82400 6800 82600 7000
rect 20800 7000 21000 7200
rect 38000 7000 38200 7200
rect 72200 7000 72400 7200
rect 82400 7000 82600 7200
rect 20800 7200 21000 7400
rect 38000 7200 38200 7400
rect 72200 7200 72400 7400
rect 82400 7200 82600 7400
rect 20800 7400 21000 7600
rect 38000 7400 38200 7600
rect 72200 7400 72400 7600
rect 82400 7400 82600 7600
rect 20800 7600 21000 7800
rect 38000 7600 38200 7800
rect 72200 7600 72400 7800
rect 82400 7600 82600 7800
rect 20800 7800 21000 8000
rect 38000 7800 38200 8000
rect 72200 7800 72400 8000
rect 82400 7800 82600 8000
rect 20800 8000 21000 8200
rect 38000 8000 38200 8200
rect 72200 8000 72400 8200
rect 82400 8000 82600 8200
rect 20800 8200 21000 8400
rect 38000 8200 38200 8400
rect 72200 8200 72400 8400
rect 82400 8200 82600 8400
rect 20800 8400 21000 8600
rect 38000 8400 38200 8600
rect 72200 8400 72400 8600
rect 82400 8400 82600 8600
rect 20800 8600 21000 8800
rect 38000 8600 38200 8800
rect 72200 8600 72400 8800
rect 82400 8600 82600 8800
rect 20800 8800 21000 9000
rect 38000 8800 38200 9000
rect 72200 8800 72400 9000
rect 82400 8800 82600 9000
rect 20800 9000 21000 9200
rect 38000 9000 38200 9200
rect 72200 9000 72400 9200
rect 82400 9000 82600 9200
rect 20800 9200 21000 9400
rect 38000 9200 38200 9400
rect 72200 9200 72400 9400
rect 82400 9200 82600 9400
rect 20800 9400 21000 9600
rect 38000 9400 38200 9600
rect 72200 9400 72400 9600
rect 82400 9400 82600 9600
rect 20800 9600 21000 9800
rect 38000 9600 38200 9800
rect 72200 9600 72400 9800
rect 82400 9600 82600 9800
rect 20800 9800 21000 10000
rect 38000 9800 38200 10000
rect 72200 9800 72400 10000
rect 82400 9800 82600 10000
rect 20800 10000 21000 10200
rect 38000 10000 38200 10200
rect 72200 10000 72400 10200
rect 82400 10000 82600 10200
rect 20800 10200 21000 10400
rect 38000 10200 38200 10400
rect 72200 10200 72400 10400
rect 82400 10200 82600 10400
rect 20800 10400 21000 10600
rect 38000 10400 38200 10600
rect 72200 10400 72400 10600
rect 82400 10400 82600 10600
rect 20800 10600 21000 10800
rect 38000 10600 38200 10800
rect 72200 10600 72400 10800
rect 82400 10600 82600 10800
rect 20800 10800 21000 11000
rect 38000 10800 38200 11000
rect 72200 10800 72400 11000
rect 82400 10800 82600 11000
rect 20800 11000 21000 11200
rect 38000 11000 38200 11200
rect 72200 11000 72400 11200
rect 82400 11000 82600 11200
rect 20800 11200 21000 11400
rect 38000 11200 38200 11400
rect 72200 11200 72400 11400
rect 82400 11200 82600 11400
rect 20800 11400 21000 11600
rect 38000 11400 38200 11600
rect 72200 11400 72400 11600
rect 82400 11400 82600 11600
rect 20800 11600 21000 11800
rect 38000 11600 38200 11800
rect 72200 11600 72400 11800
rect 82400 11600 82600 11800
rect 20800 11800 21000 12000
rect 38000 11800 38200 12000
rect 72200 11800 72400 12000
rect 82400 11800 82600 12000
rect 20800 12000 21000 12200
rect 38000 12000 38200 12200
rect 72200 12000 72400 12200
rect 82400 12000 82600 12200
rect 20800 12200 21000 12400
rect 38000 12200 38200 12400
rect 72200 12200 72400 12400
rect 82400 12200 82600 12400
rect 20800 12400 21000 12600
rect 38000 12400 38200 12600
rect 72200 12400 72400 12600
rect 82400 12400 82600 12600
rect 20800 12600 21000 12800
rect 38000 12600 38200 12800
rect 72200 12600 72400 12800
rect 82400 12600 82600 12800
rect 20800 12800 21000 13000
rect 38000 12800 38200 13000
rect 72200 12800 72400 13000
rect 82400 12800 82600 13000
rect 20800 13000 21000 13200
rect 38000 13000 38200 13200
rect 72200 13000 72400 13200
rect 82400 13000 82600 13200
rect 20800 13200 21000 13400
rect 38000 13200 38200 13400
rect 72200 13200 72400 13400
rect 82400 13200 82600 13400
rect 20800 13400 21000 13600
rect 38000 13400 38200 13600
rect 72200 13400 72400 13600
rect 82400 13400 82600 13600
rect 20800 13600 21000 13800
rect 38000 13600 38200 13800
rect 72200 13600 72400 13800
rect 82400 13600 82600 13800
rect 20800 13800 21000 14000
rect 38000 13800 38200 14000
rect 72200 13800 72400 14000
rect 82400 13800 82600 14000
rect 20800 14000 21000 14200
rect 38000 14000 38200 14200
rect 72200 14000 72400 14200
rect 82400 14000 82600 14200
rect 17400 14200 17600 14400
rect 41400 14200 41600 14400
rect 44800 14200 45000 14400
rect 48200 14200 48400 14400
rect 75600 14200 75800 14400
rect 79000 14200 79200 14400
rect 84800 14400 85000 14600
rect 85800 15800 86000 16000
rect 85800 16000 86000 16200
rect 85800 16200 86000 16400
rect 85800 16400 86000 16600
rect 85800 16600 86000 16800
rect 85800 16800 86000 17000
rect 85800 17000 86000 17200
rect 85800 17200 86000 17400
rect 85800 17400 86000 17600
rect 2800 18000 3000 18200
rect 2400 18400 2600 18600
rect 97600 18600 97800 18800
rect 2200 18800 2400 19000
rect 18600 19200 18800 19400
rect 43800 19200 44000 19400
rect 18600 19400 18800 19600
rect 18600 19600 18800 19800
rect 18600 19800 18800 20000
rect 18600 20000 18800 20200
rect 18600 20200 18800 20400
rect 18600 20400 18800 20600
rect 46200 20400 46400 20600
rect 97400 20400 97600 20600
rect 18600 20600 18800 20800
rect 97200 20600 97400 20800
rect 3000 20800 3200 21000
rect 18600 20800 18800 21000
rect 3600 21000 14000 21200
rect 18600 21000 18800 21200
rect 86000 21000 96400 21200
rect 18600 21200 18800 21400
rect 85800 21200 86000 21400
rect 18600 21400 18800 21600
rect 47200 21400 47400 21600
rect 85800 21400 86000 21600
rect 18600 21600 18800 21800
rect 85800 21600 86000 21800
rect 18600 21800 18800 22000
rect 85800 21800 86000 22000
rect 18600 22000 18800 22200
rect 47600 22000 47800 22200
rect 85800 22000 86000 22200
rect 18600 22200 18800 22400
rect 85800 22200 86000 22400
rect 18600 22400 18800 22600
rect 85800 22400 86000 22600
rect 18600 22600 18800 22800
rect 85800 22600 86000 22800
rect 18600 22800 18800 23000
rect 85800 22800 86000 23000
rect 18600 23000 18800 23200
rect 85800 23000 86000 23200
rect 18600 23200 18800 23400
rect 48200 23200 48400 23400
rect 85800 23200 86000 23400
rect 18600 23400 18800 23600
rect 85800 23400 86000 23600
rect 18600 23600 18800 23800
rect 85800 23600 86000 23800
rect 18600 23800 18800 24000
rect 85800 23800 86000 24000
rect 18600 24000 18800 24200
rect 48400 24000 48600 24200
rect 85800 24000 86000 24200
rect 18600 24200 18800 24400
rect 85800 24200 86000 24400
rect 18600 24400 18800 24600
rect 85800 24400 86000 24600
rect 3200 24600 3400 24800
rect 18600 24600 18800 24800
rect 96600 24600 96800 24800
rect 18600 24800 18800 25000
rect 97000 24800 97200 25000
rect 2600 25000 2800 25200
rect 18600 25000 18800 25200
rect 57400 25200 57600 25400
rect 57400 25400 57600 25600
rect 2200 25600 2400 25800
rect 57400 25600 57600 25800
rect 57400 25800 57600 26000
rect 57400 26000 57600 26200
rect 57400 26200 57600 26400
rect 57400 26400 57600 26600
rect 57400 26600 57600 26800
rect 2200 26800 2400 27000
rect 57400 26800 57600 27000
rect 57400 27000 57600 27200
rect 57400 27200 57600 27400
rect 2600 27400 2800 27600
rect 57400 27400 57600 27600
rect 57400 27600 57600 27800
rect 97000 27600 97200 27800
rect 3400 27800 3600 28000
rect 57400 27800 57600 28000
rect 96400 27800 96600 28000
rect 57400 28000 57600 28200
rect 85800 28000 86000 28200
rect 57400 28200 57600 28400
rect 85800 28200 86000 28400
rect 57400 28400 57600 28600
rect 85800 28400 86000 28600
rect 57400 28600 57600 28800
rect 85800 28600 86000 28800
rect 57400 28800 57600 29000
rect 85800 28800 86000 29000
rect 57400 29000 57600 29200
rect 85800 29000 86000 29200
rect 57400 29200 57600 29400
rect 85800 29200 86000 29400
rect 57400 29400 57600 29600
rect 85800 29400 86000 29600
rect 57400 29600 57600 29800
rect 85800 29600 86000 29800
rect 57400 29800 57600 30000
rect 85800 29800 86000 30000
rect 57400 30000 57600 30200
rect 85800 30000 86000 30200
rect 57400 30200 57600 30400
rect 85800 30200 86000 30400
rect 57400 30400 57600 30600
rect 85800 30400 86000 30600
rect 57400 30600 57600 30800
rect 85800 30600 86000 30800
rect 57400 30800 57600 31000
rect 85800 30800 86000 31000
rect 24000 31000 24600 31200
rect 75400 31000 76000 31200
rect 85800 31000 86000 31200
rect 23000 31200 23200 31400
rect 76800 31200 77000 31400
rect 85800 31200 86000 31400
rect 3400 31400 14000 31600
rect 22400 31400 22600 31600
rect 77400 31400 77600 31600
rect 86000 31400 96600 31600
rect 22000 31600 22200 31800
rect 21600 31800 21800 32000
rect 51400 31800 51600 32000
rect 78200 31800 78400 32000
rect 97200 31800 97400 32000
rect 48400 32000 48600 32200
rect 97400 32000 97600 32200
rect 21000 32200 21200 32400
rect 78800 32200 79000 32400
rect 20800 32400 21000 32600
rect 48200 32800 48400 33000
rect 20000 33200 20200 33400
rect 19800 33400 20000 33600
rect 48000 33400 48200 33600
rect 80000 33400 80200 33600
rect 2200 33600 2400 33800
rect 2400 34000 2600 34200
rect 80400 34000 80600 34200
rect 2800 34400 3000 34600
rect 19200 34400 19400 34600
rect 52400 34400 52600 34600
rect 3200 34600 3400 34800
rect 96600 34600 96800 34800
rect 19000 34800 19200 35000
rect 85800 35000 86000 35200
rect 85800 35200 86000 35400
rect 18800 35400 19000 35600
rect 85800 35400 86000 35600
rect 85800 35600 86000 35800
rect 85800 35800 86000 36000
rect 45800 36000 46000 36200
rect 54000 36000 54200 36200
rect 85800 36000 86000 36200
rect 54400 36200 54600 36400
rect 85800 36200 86000 36400
rect 81200 36400 81400 36600
rect 85800 36400 86000 36600
rect 18600 36600 18800 36800
rect 85800 36600 86000 36800
rect 18600 36800 18800 37000
rect 55800 36800 56000 37000
rect 85800 36800 86000 37000
rect 18600 37000 18800 37200
rect 42800 37000 43200 37200
rect 56800 37000 57200 37200
rect 85800 37000 86000 37200
rect 18600 37200 18800 37400
rect 75200 37200 75400 37400
rect 85800 37200 86000 37400
rect 18600 37400 18800 37600
rect 75200 37400 75400 37600
rect 85800 37400 86000 37600
rect 18600 37600 18800 37800
rect 75200 37600 75400 37800
rect 85800 37600 86000 37800
rect 18600 37800 18800 38000
rect 75200 37800 75400 38000
rect 85800 37800 86000 38000
rect 18600 38000 18800 38200
rect 75200 38000 75400 38200
rect 85800 38000 86000 38200
rect 14000 38200 14200 38400
rect 18600 38200 18800 38400
rect 75200 38200 75400 38400
rect 3000 38400 3200 38600
rect 18600 38400 18800 38600
rect 75200 38400 75400 38600
rect 18600 38600 18800 38800
rect 75200 38600 75400 38800
rect 18600 38800 18800 39000
rect 75200 38800 75400 39000
rect 18600 39000 18800 39200
rect 75200 39000 75400 39200
rect 18600 39200 18800 39400
rect 75200 39200 75400 39400
rect 97600 39200 97800 39400
rect 18600 39400 18800 39600
rect 75200 39400 75400 39600
rect 18600 39600 18800 39800
rect 75200 39600 75400 39800
rect 18600 39800 18800 40000
rect 75200 39800 75400 40000
rect 18600 40000 18800 40200
rect 75200 40000 75400 40200
rect 18600 40200 18800 40400
rect 75200 40200 75400 40400
rect 18600 40400 18800 40600
rect 75200 40400 75400 40600
rect 18600 40600 18800 40800
rect 75200 40600 75400 40800
rect 97600 40600 97800 40800
rect 18600 40800 18800 41000
rect 75200 40800 75400 41000
rect 18600 41000 18800 41200
rect 75200 41000 75400 41200
rect 18600 41200 18800 41400
rect 75200 41200 75400 41400
rect 18600 41400 18800 41600
rect 75200 41400 75400 41600
rect 96800 41400 97000 41600
rect 14000 41600 14200 41800
rect 18600 41600 18800 41800
rect 75200 41600 75400 41800
rect 18600 41800 18800 42000
rect 75200 41800 75400 42000
rect 85800 41800 86000 42000
rect 18600 42000 18800 42200
rect 75200 42000 75400 42200
rect 85800 42000 86000 42200
rect 18600 42200 18800 42400
rect 75200 42200 75400 42400
rect 85800 42200 86000 42400
rect 18600 42400 18800 42600
rect 75200 42400 75400 42600
rect 85800 42400 86000 42600
rect 18600 42600 18800 42800
rect 75200 42600 75400 42800
rect 85800 42600 86000 42800
rect 18600 42800 18800 43000
rect 75200 42800 75400 43000
rect 85800 42800 86000 43000
rect 18600 43000 18800 43200
rect 85800 43000 86000 43200
rect 18600 43200 18800 43400
rect 85800 43200 86000 43400
rect 18600 43400 18800 43600
rect 81200 43400 81400 43600
rect 85800 43400 86000 43600
rect 81200 43600 81400 43800
rect 85800 43600 86000 43800
rect 85800 43800 86000 44000
rect 85800 44000 86000 44200
rect 85800 44200 86000 44400
rect 85800 44400 86000 44600
rect 81000 44600 81200 44800
rect 85800 44600 86000 44800
rect 85800 44800 86000 45000
rect 14000 45000 14200 45200
rect 80800 45200 81000 45400
rect 2800 45400 3000 45600
rect 80600 45600 80800 45800
rect 2400 45800 2600 46000
rect 97600 46000 97800 46200
rect 2200 46200 2400 46400
rect 79800 46800 80000 47000
rect 20200 47000 20400 47200
rect 79600 47000 79800 47200
rect 20400 47200 20600 47400
rect 20600 47400 20800 47600
rect 79200 47400 79400 47600
rect 97400 47800 97600 48000
rect 21400 48000 21600 48200
rect 78400 48000 78600 48200
rect 97200 48000 97400 48200
rect 3000 48200 3200 48400
rect 21800 48200 22000 48400
rect 3600 48400 14000 48600
rect 86000 48400 96400 48600
rect 22600 48600 22800 48800
rect 77200 48600 77400 48800
rect 85800 48600 86000 48800
rect 76600 48800 76800 49000
rect 85800 48800 86000 49000
rect 85800 49000 86000 49200
rect 85800 49200 86000 49400
rect 85800 49400 86000 49600
rect 85800 49600 86000 49800
rect 85800 49800 86000 50000
rect 85800 50000 86000 50200
rect 85800 50200 86000 50400
rect 85800 50400 86000 50600
rect 85800 50600 86000 50800
rect 85800 50800 86000 51000
rect 22600 51000 22800 51200
rect 85800 51000 86000 51200
rect 85800 51200 86000 51400
rect 21800 51400 22000 51600
rect 85800 51400 86000 51600
rect 21400 51600 21600 51800
rect 85800 51600 86000 51800
rect 3200 52000 3400 52200
rect 96600 52000 96800 52200
rect 97000 52200 97200 52400
rect 2600 52400 2800 52600
rect 20400 52400 20600 52600
rect 20200 52600 20400 52800
rect 2200 53000 2400 53200
rect 2200 54200 2400 54400
rect 2600 54800 2800 55000
rect 97000 55000 97200 55200
rect 3400 55200 3600 55400
rect 18800 55200 19000 55400
rect 96400 55200 96600 55400
rect 85800 55400 86000 55600
rect 85800 55600 86000 55800
rect 85800 55800 86000 56000
rect 85800 56000 86000 56200
rect 18600 56200 18800 56400
rect 85800 56200 86000 56400
rect 18600 56400 18800 56600
rect 85800 56400 86000 56600
rect 18600 56600 18800 56800
rect 85800 56600 86000 56800
rect 18600 56800 18800 57000
rect 57400 56800 57600 57000
rect 85800 56800 86000 57000
rect 18600 57000 18800 57200
rect 57400 57000 57600 57200
rect 85800 57000 86000 57200
rect 18600 57200 18800 57400
rect 57400 57200 57600 57400
rect 85800 57200 86000 57400
rect 18600 57400 18800 57600
rect 57400 57400 57600 57600
rect 85800 57400 86000 57600
rect 18600 57600 18800 57800
rect 57400 57600 57600 57800
rect 85800 57600 86000 57800
rect 18600 57800 18800 58000
rect 57400 57800 57600 58000
rect 85800 57800 86000 58000
rect 18600 58000 18800 58200
rect 57400 58000 57600 58200
rect 85800 58000 86000 58200
rect 18600 58200 18800 58400
rect 57400 58200 57600 58400
rect 85800 58200 86000 58400
rect 18600 58400 18800 58600
rect 57400 58400 57600 58600
rect 85800 58400 86000 58600
rect 18600 58600 18800 58800
rect 57400 58600 57600 58800
rect 85800 58600 86000 58800
rect 3400 58800 3600 59000
rect 18600 58800 18800 59000
rect 57400 58800 57600 59000
rect 96400 58800 96600 59000
rect 18600 59000 18800 59200
rect 57400 59000 57600 59200
rect 18600 59200 18800 59400
rect 57400 59200 57600 59400
rect 97200 59200 97400 59400
rect 18600 59400 18800 59600
rect 57400 59400 57600 59600
rect 97400 59400 97600 59600
rect 18600 59600 18800 59800
rect 57400 59600 57600 59800
rect 18600 59800 18800 60000
rect 57400 59800 57600 60000
rect 18600 60000 18800 60200
rect 57400 60000 57600 60200
rect 18600 60200 18800 60400
rect 57400 60200 57600 60400
rect 18600 60400 18800 60600
rect 57400 60400 57600 60600
rect 18600 60600 18800 60800
rect 57400 60600 57600 60800
rect 18600 60800 18800 61000
rect 57400 60800 57600 61000
rect 2200 61000 2400 61200
rect 18600 61000 18800 61200
rect 57400 61000 57600 61200
rect 18600 61200 18800 61400
rect 57400 61200 57600 61400
rect 2400 61400 2600 61600
rect 18600 61400 18800 61600
rect 57400 61400 57600 61600
rect 18600 61600 18800 61800
rect 57400 61600 57600 61800
rect 2800 61800 3000 62000
rect 18600 61800 18800 62000
rect 57400 61800 57600 62000
rect 3200 62000 3400 62200
rect 18600 62000 18800 62200
rect 57400 62000 57600 62200
rect 96600 62000 96800 62200
rect 18600 62200 18800 62400
rect 57400 62200 57600 62400
rect 18600 62400 18800 62600
rect 57400 62400 57600 62600
rect 85800 62400 86000 62600
rect 18600 62600 18800 62800
rect 75400 62600 76000 62800
rect 85800 62600 86000 62800
rect 18600 62800 18800 63000
rect 76800 62800 77000 63000
rect 85800 62800 86000 63000
rect 18600 63000 18800 63200
rect 77400 63000 77600 63200
rect 85800 63000 86000 63200
rect 18600 63200 18800 63400
rect 85800 63200 86000 63400
rect 18600 63400 18800 63600
rect 51400 63400 51600 63600
rect 78200 63400 78400 63600
rect 85800 63400 86000 63600
rect 18600 63600 18800 63800
rect 85800 63600 86000 63800
rect 18600 63800 18800 64000
rect 78800 63800 79000 64000
rect 85800 63800 86000 64000
rect 18600 64000 18800 64200
rect 85800 64000 86000 64200
rect 18600 64200 18800 64400
rect 85800 64200 86000 64400
rect 18600 64400 18800 64600
rect 85800 64400 86000 64600
rect 18600 64600 18800 64800
rect 85800 64600 86000 64800
rect 18600 64800 18800 65000
rect 85800 64800 86000 65000
rect 18600 65000 18800 65200
rect 80000 65000 80200 65200
rect 85800 65000 86000 65200
rect 18600 65200 18800 65400
rect 85800 65200 86000 65400
rect 18600 65400 18800 65600
rect 85800 65400 86000 65600
rect 3400 65600 14000 65800
rect 18600 65600 18800 65800
rect 80400 65600 80600 65800
rect 86000 65600 96600 65800
rect 18600 65800 18800 66000
rect 18600 66000 18800 66200
rect 52400 66000 52600 66200
rect 97200 66000 97400 66200
rect 18600 66200 18800 66400
rect 97400 66200 97600 66400
rect 18600 66400 18800 66600
rect 18600 66600 18800 66800
rect 18600 66800 18800 67000
rect 18600 67000 18800 67200
rect 18600 67200 18800 67400
rect 18600 67400 18800 67600
rect 18600 67600 18800 67800
rect 54000 67600 54200 67800
rect 18600 67800 18800 68000
rect 54400 67800 54600 68000
rect 18600 68000 18800 68200
rect 81200 68000 81400 68200
rect 97600 68000 97800 68200
rect 18600 68200 18800 68400
rect 18600 68400 18800 68600
rect 55800 68400 56000 68600
rect 18600 68600 18800 68800
rect 56800 68600 57200 68800
rect 18600 68800 18800 69000
rect 75200 68800 75400 69000
rect 96800 68800 97000 69000
rect 14000 69000 14200 69200
rect 18600 69000 18800 69200
rect 75200 69000 75400 69200
rect 18600 69200 18800 69400
rect 75200 69200 75400 69400
rect 85800 69200 86000 69400
rect 18600 69400 18800 69600
rect 75200 69400 75400 69600
rect 85800 69400 86000 69600
rect 18600 69600 18800 69800
rect 75200 69600 75400 69800
rect 85800 69600 86000 69800
rect 18600 69800 18800 70000
rect 75200 69800 75400 70000
rect 85800 69800 86000 70000
rect 18600 70000 18800 70200
rect 75200 70000 75400 70200
rect 85800 70000 86000 70200
rect 18600 70200 18800 70400
rect 75200 70200 75400 70400
rect 85800 70200 86000 70400
rect 18600 70400 18800 70600
rect 75200 70400 75400 70600
rect 85800 70400 86000 70600
rect 18600 70600 18800 70800
rect 75200 70600 75400 70800
rect 85800 70600 86000 70800
rect 18600 70800 18800 71000
rect 75200 70800 75400 71000
rect 85800 70800 86000 71000
rect 18600 71000 18800 71200
rect 75200 71000 75400 71200
rect 85800 71000 86000 71200
rect 18600 71200 18800 71400
rect 75200 71200 75400 71400
rect 85800 71200 86000 71400
rect 18600 71400 18800 71600
rect 75200 71400 75400 71600
rect 85800 71400 86000 71600
rect 18600 71600 18800 71800
rect 75200 71600 75400 71800
rect 85800 71600 86000 71800
rect 18600 71800 18800 72000
rect 75200 71800 75400 72000
rect 85800 71800 86000 72000
rect 18600 72000 18800 72200
rect 75200 72000 75400 72200
rect 85800 72000 86000 72200
rect 18600 72200 18800 72400
rect 75200 72200 75400 72400
rect 85800 72200 86000 72400
rect 14000 72400 14200 72600
rect 18600 72400 18800 72600
rect 75200 72400 75400 72600
rect 3000 72600 3200 72800
rect 18600 72600 18800 72800
rect 75200 72600 75400 72800
rect 18600 72800 18800 73000
rect 75200 72800 75400 73000
rect 18600 73000 18800 73200
rect 75200 73000 75400 73200
rect 18600 73200 18800 73400
rect 75200 73200 75400 73400
rect 18600 73400 18800 73600
rect 75200 73400 75400 73600
rect 97600 73400 97800 73600
rect 18600 73600 18800 73800
rect 75200 73600 75400 73800
rect 18600 73800 18800 74000
rect 75200 73800 75400 74000
rect 18600 74000 18800 74200
rect 75200 74000 75400 74200
rect 18600 74200 18800 74400
rect 75200 74200 75400 74400
rect 18600 74400 18800 74600
rect 75200 74400 75400 74600
rect 18600 74600 18800 74800
rect 18600 74800 18800 75000
rect 18600 75000 18800 75200
rect 81200 75000 81400 75200
rect 81200 75200 81400 75400
rect 97400 75200 97600 75400
rect 97200 75400 97400 75600
rect 3000 75600 3200 75800
rect 3600 75800 14000 76000
rect 86000 75800 96400 76000
rect 85800 76000 86000 76200
rect 81000 76200 81200 76400
rect 85800 76200 86000 76400
rect 85800 76400 86000 76600
rect 85800 76600 86000 76800
rect 80800 76800 81000 77000
rect 85800 76800 86000 77000
rect 85800 77000 86000 77200
rect 80600 77200 80800 77400
rect 85800 77200 86000 77400
rect 85800 77400 86000 77600
rect 85800 77600 86000 77800
rect 85800 77800 86000 78000
rect 85800 78000 86000 78200
rect 85800 78200 86000 78400
rect 79800 78400 80000 78600
rect 85800 78400 86000 78600
rect 20200 78600 20400 78800
rect 79600 78600 79800 78800
rect 85800 78600 86000 78800
rect 20400 78800 20600 79000
rect 85800 78800 86000 79000
rect 20600 79000 20800 79200
rect 79200 79000 79400 79200
rect 85800 79000 86000 79200
rect 2800 79600 3000 79800
rect 21400 79600 21600 79800
rect 78400 79600 78600 79800
rect 21800 79800 22000 80000
rect 2400 80000 2600 80200
rect 22600 80200 22800 80400
rect 77200 80200 77400 80400
rect 97600 80200 97800 80400
rect 2200 80400 2400 80600
rect 76600 80400 76800 80600
rect 2200 81600 2400 81800
rect 2600 82200 2800 82400
rect 97000 82400 97200 82600
rect 3400 82600 3600 82800
rect 96400 82600 96600 82800
rect 85800 82800 86000 83000
rect 85800 83000 86000 83200
rect 85800 83200 86000 83400
rect 85800 83400 86000 83600
rect 85800 83600 86000 83800
rect 85800 83800 86000 84000
rect 85800 84000 86000 84200
rect 85800 84200 86000 84400
rect 85800 84400 86000 84600
rect 14400 85400 14600 85600
rect 14600 85600 14800 85800
rect 85000 85800 85200 86000
rect 15400 86000 15600 86200
rect 84400 86000 84600 86200
rect 20800 86200 21000 86400
rect 38000 86200 38200 86400
rect 72200 86200 72400 86400
rect 82400 86200 82600 86400
rect 20800 86400 21000 86600
rect 38000 86400 38200 86600
rect 72200 86400 72400 86600
rect 82400 86400 82600 86600
rect 20800 86600 21000 86800
rect 38000 86600 38200 86800
rect 72200 86600 72400 86800
rect 82400 86600 82600 86800
rect 20800 86800 21000 87000
rect 38000 86800 38200 87000
rect 72200 86800 72400 87000
rect 82400 86800 82600 87000
rect 20800 87000 21000 87200
rect 38000 87000 38200 87200
rect 72200 87000 72400 87200
rect 82400 87000 82600 87200
rect 20800 87200 21000 87400
rect 38000 87200 38200 87400
rect 72200 87200 72400 87400
rect 82400 87200 82600 87400
rect 20800 87400 21000 87600
rect 38000 87400 38200 87600
rect 72200 87400 72400 87600
rect 82400 87400 82600 87600
rect 20800 87600 21000 87800
rect 38000 87600 38200 87800
rect 72200 87600 72400 87800
rect 82400 87600 82600 87800
rect 20800 87800 21000 88000
rect 38000 87800 38200 88000
rect 72200 87800 72400 88000
rect 82400 87800 82600 88000
rect 20800 88000 21000 88200
rect 38000 88000 38200 88200
rect 72200 88000 72400 88200
rect 82400 88000 82600 88200
rect 20800 88200 21000 88400
rect 38000 88200 38200 88400
rect 72200 88200 72400 88400
rect 82400 88200 82600 88400
rect 20800 88400 21000 88600
rect 38000 88400 38200 88600
rect 72200 88400 72400 88600
rect 82400 88400 82600 88600
rect 20800 88600 21000 88800
rect 38000 88600 38200 88800
rect 72200 88600 72400 88800
rect 82400 88600 82600 88800
rect 20800 88800 21000 89000
rect 38000 88800 38200 89000
rect 72200 88800 72400 89000
rect 82400 88800 82600 89000
rect 20800 89000 21000 89200
rect 38000 89000 38200 89200
rect 72200 89000 72400 89200
rect 82400 89000 82600 89200
rect 20800 89200 21000 89400
rect 38000 89200 38200 89400
rect 72200 89200 72400 89400
rect 82400 89200 82600 89400
rect 20800 89400 21000 89600
rect 38000 89400 38200 89600
rect 72200 89400 72400 89600
rect 82400 89400 82600 89600
rect 20800 89600 21000 89800
rect 38000 89600 38200 89800
rect 72200 89600 72400 89800
rect 82400 89600 82600 89800
rect 20800 89800 21000 90000
rect 38000 89800 38200 90000
rect 72200 89800 72400 90000
rect 82400 89800 82600 90000
rect 20800 90000 21000 90200
rect 38000 90000 38200 90200
rect 72200 90000 72400 90200
rect 82400 90000 82600 90200
rect 20800 90200 21000 90400
rect 38000 90200 38200 90400
rect 72200 90200 72400 90400
rect 82400 90200 82600 90400
rect 20800 90400 21000 90600
rect 38000 90400 38200 90600
rect 72200 90400 72400 90600
rect 82400 90400 82600 90600
rect 20800 90600 21000 90800
rect 38000 90600 38200 90800
rect 72200 90600 72400 90800
rect 82400 90600 82600 90800
rect 20800 90800 21000 91000
rect 38000 90800 38200 91000
rect 72200 90800 72400 91000
rect 82400 90800 82600 91000
rect 20800 91000 21000 91200
rect 38000 91000 38200 91200
rect 72200 91000 72400 91200
rect 82400 91000 82600 91200
rect 20800 91200 21000 91400
rect 38000 91200 38200 91400
rect 72200 91200 72400 91400
rect 82400 91200 82600 91400
rect 20800 91400 21000 91600
rect 38000 91400 38200 91600
rect 72200 91400 72400 91600
rect 82400 91400 82600 91600
rect 20800 91600 21000 91800
rect 38000 91600 38200 91800
rect 72200 91600 72400 91800
rect 82400 91600 82600 91800
rect 20800 91800 21000 92000
rect 38000 91800 38200 92000
rect 72200 91800 72400 92000
rect 82400 91800 82600 92000
rect 20800 92000 21000 92200
rect 38000 92000 38200 92200
rect 72200 92000 72400 92200
rect 82400 92000 82600 92200
rect 20800 92200 21000 92400
rect 38000 92200 38200 92400
rect 72200 92200 72400 92400
rect 82400 92200 82600 92400
rect 20800 92400 21000 92600
rect 38000 92400 38200 92600
rect 72200 92400 72400 92600
rect 82400 92400 82600 92600
rect 20800 92600 21000 92800
rect 38000 92600 38200 92800
rect 72200 92600 72400 92800
rect 82400 92600 82600 92800
rect 20800 92800 21000 93000
rect 38000 92800 38200 93000
rect 72200 92800 72400 93000
rect 82400 92800 82600 93000
rect 20800 93000 21000 93200
rect 38000 93000 38200 93200
rect 72200 93000 72400 93200
rect 82400 93000 82600 93200
rect 20800 93200 21000 93400
rect 38000 93200 38200 93400
rect 72200 93200 72400 93400
rect 82400 93200 82600 93400
rect 20800 93400 21000 93600
rect 38000 93400 38200 93600
rect 72200 93400 72400 93600
rect 82400 93400 82600 93600
rect 20800 93600 21000 93800
rect 38000 93600 38200 93800
rect 72200 93600 72400 93800
rect 82400 93600 82600 93800
rect 20800 93800 21000 94000
rect 38000 93800 38200 94000
rect 72200 93800 72400 94000
rect 82400 93800 82600 94000
rect 20800 94000 21000 94200
rect 38000 94000 38200 94200
rect 72200 94000 72400 94200
rect 82400 94000 82600 94200
rect 20800 94200 21000 94400
rect 38000 94200 38200 94400
rect 72200 94200 72400 94400
rect 82400 94200 82600 94400
rect 20800 94400 21000 94600
rect 38000 94400 38200 94600
rect 72200 94400 72400 94600
rect 82400 94400 82600 94600
rect 20800 94600 21000 94800
rect 38000 94600 38200 94800
rect 72200 94600 72400 94800
rect 82400 94600 82600 94800
rect 20800 94800 21000 95000
rect 38000 94800 38200 95000
rect 72200 94800 72400 95000
rect 82400 94800 82600 95000
rect 20800 95000 21000 95200
rect 38000 95000 38200 95200
rect 72200 95000 72400 95200
rect 82400 95000 82600 95200
rect 20800 95200 21000 95400
rect 38000 95200 38200 95400
rect 72200 95200 72400 95400
rect 82400 95200 82600 95400
rect 20800 95400 21000 95600
rect 38000 95400 38200 95600
rect 72200 95400 72400 95600
rect 82400 95400 82600 95600
rect 20800 95600 21000 95800
rect 38000 95600 38200 95800
rect 72200 95600 72400 95800
rect 82400 95600 82600 95800
rect 20800 95800 21000 96000
rect 38000 95800 38200 96000
rect 72200 95800 72400 96000
rect 82400 95800 82600 96000
rect 20800 96000 21000 96200
rect 38000 96000 38200 96200
rect 72200 96000 72400 96200
rect 82400 96000 82600 96200
rect 20800 96200 21000 96400
rect 38000 96200 38200 96400
rect 72200 96200 72400 96400
rect 82400 96200 82600 96400
rect 20800 96400 21000 96600
rect 38000 96400 38200 96600
rect 55000 96400 55200 96600
rect 20800 96600 21000 96800
rect 31200 96600 31400 96800
rect 55000 96600 55200 96800
rect 65400 96600 65600 96800
rect 27600 96800 27800 97000
rect 31200 96800 31400 97000
rect 61800 96800 62000 97000
rect 17600 97000 17800 97200
rect 41200 97000 41400 97200
rect 51800 97000 52000 97200
rect 75400 97000 75600 97200
rect 20600 97200 20800 97400
rect 38200 97200 38400 97400
rect 54800 97200 55000 97400
rect 17800 97400 18000 97600
rect 41000 97400 41200 97600
rect 45200 97400 45400 97600
rect 75200 97400 75400 97600
rect 79400 97400 79600 97600
rect 18000 97600 18200 97800
rect 40800 97600 41000 97800
rect 52200 97600 52400 97800
rect 68200 97600 68400 97800
rect 75000 97600 75200 97800
rect 79600 97600 79800 97800
rect 20000 97800 20200 98000
rect 38800 97800 39000 98000
rect 47400 97800 47600 98000
rect 54200 97800 54400 98000
rect 66200 97800 66400 98000
rect 73000 97800 73200 98000
rect 81600 97800 81800 98000
rect 18800 98000 19000 98200
rect 19400 98000 19600 98200
rect 25600 98000 25800 98200
rect 26400 98000 26600 98200
rect 32400 98000 32600 98200
rect 33200 98000 33400 98200
rect 39400 98000 39600 98200
rect 40000 98000 40200 98200
rect 46200 98000 46400 98200
rect 46800 98000 47000 98200
rect 53000 98000 53200 98200
rect 53600 98000 53800 98200
rect 59800 98000 60000 98200
rect 60600 98000 60800 98200
rect 67400 98000 67600 98200
rect 73600 98000 73800 98200
rect 74200 98000 74400 98200
rect 80400 98000 80600 98200
rect 81000 98000 81200 98200
<< metal2 >>
rect 18400 2400 18600 2600
rect 40400 2400 40600 2600
rect 45800 2400 46000 2600
rect 52600 2400 52800 2600
rect 74600 2400 74800 2600
rect 80000 2400 80200 2600
rect 25000 2600 25200 2800
rect 27000 2600 27200 2800
rect 31800 2600 32000 2800
rect 59200 2600 59400 2800
rect 61200 2600 61400 2800
rect 20400 2800 20600 3000
rect 31600 2800 31800 3000
rect 54600 2800 54800 3000
rect 65800 2800 66000 3000
rect 24600 3000 24800 3200
rect 27400 3000 27600 3200
rect 58800 3000 59000 3200
rect 61600 3000 61800 3200
rect 41200 3200 41400 3400
rect 45000 3200 45200 3400
rect 75400 3200 75600 3400
rect 79200 3200 79400 3400
rect 24400 3400 24600 3600
rect 27600 3400 27800 3600
rect 58600 3400 58800 3600
rect 61800 3400 62000 3600
rect 20800 3600 21000 3800
rect 38000 3600 38200 3800
rect 55000 3600 55200 3800
rect 38000 3800 38200 4000
rect 48200 3800 48400 4000
rect 72200 3800 72400 4000
rect 82400 3800 82600 4000
rect 44800 4000 45000 4200
rect 48200 4000 48400 4200
rect 44800 4200 45000 4400
rect 48200 4200 48400 4400
rect 75600 4200 75800 4400
rect 44800 4400 45000 4600
rect 48200 4400 48400 4600
rect 75600 4400 75800 4600
rect 44800 4600 45000 4800
rect 48200 4600 48400 4800
rect 75600 4600 75800 4800
rect 44800 4800 45000 5000
rect 48200 4800 48400 5000
rect 75600 4800 75800 5000
rect 44800 5000 45000 5200
rect 48200 5000 48400 5200
rect 75600 5000 75800 5200
rect 44800 5200 45000 5400
rect 48200 5200 48400 5400
rect 75600 5200 75800 5400
rect 44800 5400 45000 5600
rect 48200 5400 48400 5600
rect 75600 5400 75800 5600
rect 44800 5600 45000 5800
rect 48200 5600 48400 5800
rect 75600 5600 75800 5800
rect 44800 5800 45000 6000
rect 48200 5800 48400 6000
rect 75600 5800 75800 6000
rect 44800 6000 45000 6200
rect 48200 6000 48400 6200
rect 75600 6000 75800 6200
rect 44800 6200 45000 6400
rect 48200 6200 48400 6400
rect 75600 6200 75800 6400
rect 44800 6400 45000 6600
rect 48200 6400 48400 6600
rect 75600 6400 75800 6600
rect 44800 6600 45000 6800
rect 48200 6600 48400 6800
rect 75600 6600 75800 6800
rect 44800 6800 45000 7000
rect 48200 6800 48400 7000
rect 75600 6800 75800 7000
rect 44800 7000 45000 7200
rect 48200 7000 48400 7200
rect 75600 7000 75800 7200
rect 44800 7200 45000 7400
rect 48200 7200 48400 7400
rect 75600 7200 75800 7400
rect 44800 7400 45000 7600
rect 48200 7400 48400 7600
rect 75600 7400 75800 7600
rect 44800 7600 45000 7800
rect 48200 7600 48400 7800
rect 75600 7600 75800 7800
rect 44800 7800 45000 8000
rect 48200 7800 48400 8000
rect 75600 7800 75800 8000
rect 44800 8000 45000 8200
rect 48200 8000 48400 8200
rect 75600 8000 75800 8200
rect 44800 8200 45000 8400
rect 48200 8200 48400 8400
rect 75600 8200 75800 8400
rect 44800 8400 45000 8600
rect 48200 8400 48400 8600
rect 75600 8400 75800 8600
rect 44800 8600 45000 8800
rect 48200 8600 48400 8800
rect 75600 8600 75800 8800
rect 44800 8800 45000 9000
rect 48200 8800 48400 9000
rect 75600 8800 75800 9000
rect 44800 9000 45000 9200
rect 48200 9000 48400 9200
rect 75600 9000 75800 9200
rect 44800 9200 45000 9400
rect 48200 9200 48400 9400
rect 75600 9200 75800 9400
rect 44800 9400 45000 9600
rect 48200 9400 48400 9600
rect 75600 9400 75800 9600
rect 44800 9600 45000 9800
rect 48200 9600 48400 9800
rect 75600 9600 75800 9800
rect 44800 9800 45000 10000
rect 48200 9800 48400 10000
rect 75600 9800 75800 10000
rect 44800 10000 45000 10200
rect 48200 10000 48400 10200
rect 75600 10000 75800 10200
rect 44800 10200 45000 10400
rect 48200 10200 48400 10400
rect 75600 10200 75800 10400
rect 44800 10400 45000 10600
rect 48200 10400 48400 10600
rect 75600 10400 75800 10600
rect 44800 10600 45000 10800
rect 48200 10600 48400 10800
rect 75600 10600 75800 10800
rect 44800 10800 45000 11000
rect 48200 10800 48400 11000
rect 75600 10800 75800 11000
rect 44800 11000 45000 11200
rect 48200 11000 48400 11200
rect 75600 11000 75800 11200
rect 44800 11200 45000 11400
rect 48200 11200 48400 11400
rect 75600 11200 75800 11400
rect 44800 11400 45000 11600
rect 48200 11400 48400 11600
rect 75600 11400 75800 11600
rect 44800 11600 45000 11800
rect 48200 11600 48400 11800
rect 75600 11600 75800 11800
rect 44800 11800 45000 12000
rect 48200 11800 48400 12000
rect 75600 11800 75800 12000
rect 44800 12000 45000 12200
rect 48200 12000 48400 12200
rect 75600 12000 75800 12200
rect 44800 12200 45000 12400
rect 48200 12200 48400 12400
rect 75600 12200 75800 12400
rect 44800 12400 45000 12600
rect 48200 12400 48400 12600
rect 75600 12400 75800 12600
rect 44800 12600 45000 12800
rect 48200 12600 48400 12800
rect 75600 12600 75800 12800
rect 44800 12800 45000 13000
rect 48200 12800 48400 13000
rect 75600 12800 75800 13000
rect 44800 13000 45000 13200
rect 48200 13000 48400 13200
rect 75600 13000 75800 13200
rect 44800 13200 45000 13400
rect 48200 13200 48400 13400
rect 75600 13200 75800 13400
rect 44800 13400 45000 13600
rect 48200 13400 48400 13600
rect 75600 13400 75800 13600
rect 44800 13600 45000 13800
rect 48200 13600 48400 13800
rect 75600 13600 75800 13800
rect 44800 13800 45000 14000
rect 48200 13800 48400 14000
rect 75600 13800 75800 14000
rect 44800 14000 45000 14200
rect 48200 14000 48400 14200
rect 75600 14000 75800 14200
rect 15800 14200 17400 14400
rect 21000 14200 24400 14400
rect 27800 14200 31200 14400
rect 34600 14200 38000 14400
rect 41600 14200 44800 14400
rect 48400 14200 51800 14400
rect 55200 14200 58600 14400
rect 62000 14200 65400 14400
rect 68800 14200 72200 14400
rect 75800 14200 79000 14400
rect 82600 14200 84400 14400
rect 15000 14400 15200 14600
rect 14200 15200 14400 15400
rect 85800 15600 86000 15800
rect 14000 17600 14200 17800
rect 3000 17800 3200 18000
rect 96800 17800 97000 18000
rect 43600 19200 43800 19400
rect 81200 19200 81400 19400
rect 44400 19400 44600 19600
rect 81200 19400 81400 19600
rect 81200 19600 81400 19800
rect 81200 19800 81400 20000
rect 2200 20000 2400 20200
rect 45600 20000 45800 20200
rect 81200 20000 81400 20200
rect 81200 20200 81400 20400
rect 81200 20400 81400 20600
rect 2600 20600 2800 20800
rect 46400 20600 46600 20800
rect 81200 20600 81400 20800
rect 81200 20800 81400 21000
rect 3400 21000 3600 21200
rect 81200 21000 81400 21200
rect 96400 21000 96600 21200
rect 47000 21200 47200 21400
rect 81200 21200 81400 21400
rect 81200 21400 81400 21600
rect 81200 21600 81400 21800
rect 81200 21800 81400 22000
rect 81200 22000 81400 22200
rect 81200 22200 81400 22400
rect 47800 22400 48000 22600
rect 81200 22400 81400 22600
rect 81200 22600 81400 22800
rect 48000 22800 48200 23000
rect 81200 22800 81400 23000
rect 81200 23000 81400 23200
rect 81200 23200 81400 23400
rect 48200 23400 48400 23600
rect 81200 23400 81400 23600
rect 81200 23600 81400 23800
rect 81200 23800 81400 24000
rect 81200 24000 81400 24200
rect 48400 24200 48600 24400
rect 81200 24200 81400 24400
rect 48400 24400 48600 24600
rect 81200 24400 81400 24600
rect 81200 24600 81400 24800
rect 2800 24800 3000 25000
rect 81200 24800 81400 25000
rect 81200 25000 81400 25200
rect 2400 25200 2600 25400
rect 97600 25400 97800 25600
rect 97600 27000 97800 27200
rect 2400 27200 2600 27400
rect 2800 27600 3000 27800
rect 96600 27800 96800 28000
rect 24600 31000 42600 31200
rect 57400 31000 75400 31200
rect 23200 31200 23400 31400
rect 51400 31200 51600 31400
rect 51400 31400 51600 31600
rect 96600 31400 96800 31600
rect 51400 31600 51600 31800
rect 77800 31600 78000 31800
rect 97000 31600 97200 31800
rect 2600 31800 2800 32000
rect 48400 31800 48600 32000
rect 2200 32400 2400 32600
rect 79000 32400 79200 32600
rect 20600 32600 20800 32800
rect 51600 32600 51800 32800
rect 20200 33000 20400 33200
rect 51800 33200 52000 33400
rect 79800 33200 80000 33400
rect 52000 33600 52200 33800
rect 97600 33800 97800 34000
rect 52200 34000 52400 34200
rect 47400 34400 47600 34600
rect 80600 34400 80800 34600
rect 52600 34600 52800 34800
rect 14000 34800 14200 35000
rect 80800 34800 81000 35000
rect 81000 35400 81200 35600
rect 18800 35600 19000 35800
rect 46000 35800 46200 36000
rect 53800 35800 54000 36000
rect 45400 36200 45600 36400
rect 45000 36400 45200 36600
rect 54800 36400 55000 36600
rect 44600 36600 44800 36800
rect 55200 36600 55400 36800
rect 81200 36600 81400 36800
rect 44000 36800 44200 37000
rect 81200 36800 81400 37000
rect 24800 37000 42800 37200
rect 57200 37000 75200 37200
rect 81200 37000 81400 37200
rect 24600 37200 24800 37400
rect 81200 37200 81400 37400
rect 24600 37400 24800 37600
rect 81200 37400 81400 37600
rect 24600 37600 24800 37800
rect 81200 37600 81400 37800
rect 24600 37800 24800 38000
rect 81200 37800 81400 38000
rect 24600 38000 24800 38200
rect 81200 38000 81400 38200
rect 3400 38200 14000 38400
rect 24600 38200 24800 38400
rect 81200 38200 81400 38400
rect 86000 38200 96600 38400
rect 24600 38400 24800 38600
rect 81200 38400 81400 38600
rect 24600 38600 24800 38800
rect 81200 38600 81400 38800
rect 97200 38600 97400 38800
rect 24600 38800 24800 39000
rect 81200 38800 81400 39000
rect 97400 38800 97600 39000
rect 24600 39000 24800 39200
rect 81200 39000 81400 39200
rect 2200 39200 2400 39400
rect 24600 39200 24800 39400
rect 81200 39200 81400 39400
rect 24600 39400 24800 39600
rect 81200 39400 81400 39600
rect 24600 39600 24800 39800
rect 81200 39600 81400 39800
rect 24600 39800 24800 40000
rect 81200 39800 81400 40000
rect 24600 40000 24800 40200
rect 81200 40000 81400 40200
rect 24600 40200 24800 40400
rect 81200 40200 81400 40400
rect 24600 40400 24800 40600
rect 81200 40400 81400 40600
rect 2200 40600 2400 40800
rect 24600 40600 24800 40800
rect 81200 40600 81400 40800
rect 24600 40800 24800 41000
rect 81200 40800 81400 41000
rect 24600 41000 24800 41200
rect 81200 41000 81400 41200
rect 97400 41000 97600 41200
rect 24600 41200 24800 41400
rect 81200 41200 81400 41400
rect 97200 41200 97400 41400
rect 3000 41400 3200 41600
rect 24600 41400 24800 41600
rect 81200 41400 81400 41600
rect 3800 41600 14000 41800
rect 24600 41600 24800 41800
rect 81200 41600 81400 41800
rect 86000 41600 96200 41800
rect 24600 41800 24800 42000
rect 81200 41800 81400 42000
rect 24600 42000 24800 42200
rect 81200 42000 81400 42200
rect 24600 42200 24800 42400
rect 81200 42200 81400 42400
rect 24600 42400 24800 42600
rect 81200 42400 81400 42600
rect 24600 42600 24800 42800
rect 81200 42600 81400 42800
rect 24600 42800 24800 43000
rect 81200 42800 81400 43000
rect 51400 43000 51600 43200
rect 81200 43000 81400 43200
rect 81200 43200 81400 43400
rect 18800 44400 19000 44600
rect 81000 44400 81200 44600
rect 3800 45000 14000 45200
rect 19000 45000 19200 45200
rect 86000 45000 96200 45200
rect 3000 45200 3200 45400
rect 96800 45200 97000 45400
rect 19400 45800 19600 46000
rect 19600 46200 19800 46400
rect 79400 47200 79600 47400
rect 2200 47400 2400 47600
rect 2600 48000 2800 48200
rect 78000 48200 78200 48400
rect 3400 48400 3600 48600
rect 22200 48400 22400 48600
rect 77600 48400 77800 48600
rect 96400 48400 96600 48600
rect 23400 48800 23600 49000
rect 76400 48800 76600 49000
rect 23400 50800 23600 51000
rect 81200 50800 81400 51000
rect 81200 51000 81400 51200
rect 22200 51200 22400 51400
rect 81200 51200 81400 51400
rect 81200 51400 81400 51600
rect 81200 51600 81400 51800
rect 14000 51800 14200 52000
rect 81200 51800 81400 52000
rect 81200 52000 81400 52200
rect 2800 52200 3000 52400
rect 81200 52200 81400 52400
rect 81200 52400 81400 52600
rect 2400 52600 2600 52800
rect 81200 52600 81400 52800
rect 81200 52800 81400 53000
rect 97600 52800 97800 53000
rect 81200 53000 81400 53200
rect 81200 53200 81400 53400
rect 19600 53400 19800 53600
rect 81200 53400 81400 53600
rect 81200 53600 81400 53800
rect 19400 53800 19600 54000
rect 81200 53800 81400 54000
rect 81200 54000 81400 54200
rect 81200 54200 81400 54400
rect 81200 54400 81400 54600
rect 97600 54400 97800 54600
rect 2400 54600 2600 54800
rect 19000 54600 19200 54800
rect 81200 54600 81400 54800
rect 81200 54800 81400 55000
rect 2800 55000 3000 55200
rect 81200 55000 81400 55200
rect 81200 55200 81400 55400
rect 96600 55200 96800 55400
rect 81200 55400 81400 55600
rect 81200 55600 81400 55800
rect 81200 55800 81400 56000
rect 81200 56000 81400 56200
rect 81200 56200 81400 56400
rect 81200 56400 81400 56600
rect 81200 56600 81400 56800
rect 24600 56800 24800 57000
rect 24600 57000 24800 57200
rect 24600 57200 24800 57400
rect 24600 57400 24800 57600
rect 24600 57600 24800 57800
rect 24600 57800 24800 58000
rect 24600 58000 24800 58200
rect 24600 58200 24800 58400
rect 24600 58400 24800 58600
rect 24600 58600 24800 58800
rect 24600 58800 24800 59000
rect 96600 58800 96800 59000
rect 24600 59000 24800 59200
rect 97000 59000 97200 59200
rect 2600 59200 2800 59400
rect 24600 59200 24800 59400
rect 24600 59400 24800 59600
rect 24600 59600 24800 59800
rect 2200 59800 2400 60000
rect 24600 59800 24800 60000
rect 24600 60000 24800 60200
rect 24600 60200 24800 60400
rect 24600 60400 24800 60600
rect 24600 60600 24800 60800
rect 24600 60800 24800 61000
rect 24600 61000 24800 61200
rect 24600 61200 24800 61400
rect 97600 61200 97800 61400
rect 24600 61400 24800 61600
rect 24600 61600 24800 61800
rect 24600 61800 24800 62000
rect 24600 62000 24800 62200
rect 14000 62200 14200 62400
rect 24600 62200 24800 62400
rect 24600 62400 24800 62600
rect 24600 62600 24800 62800
rect 57400 62600 75400 62800
rect 24600 62800 24800 63000
rect 51400 62800 51600 63000
rect 24600 63000 24800 63200
rect 51400 63000 51600 63200
rect 24600 63200 24800 63400
rect 51400 63200 51600 63400
rect 77800 63200 78000 63400
rect 24600 63400 24800 63600
rect 24600 63600 24800 63800
rect 24600 63800 24800 64000
rect 24600 64000 24800 64200
rect 79000 64000 79200 64200
rect 24600 64200 24800 64400
rect 51600 64200 51800 64400
rect 24600 64400 24800 64600
rect 24600 64600 24800 64800
rect 24600 64800 24800 65000
rect 51800 64800 52000 65000
rect 79800 64800 80000 65000
rect 24600 65000 24800 65200
rect 24600 65200 24800 65400
rect 52000 65200 52200 65400
rect 24600 65400 24800 65600
rect 24600 65600 24800 65800
rect 52200 65600 52400 65800
rect 96600 65600 96800 65800
rect 24600 65800 24800 66000
rect 97000 65800 97200 66000
rect 2600 66000 2800 66200
rect 24600 66000 24800 66200
rect 80600 66000 80800 66200
rect 24600 66200 24800 66400
rect 52600 66200 52800 66400
rect 24600 66400 24800 66600
rect 80800 66400 81000 66600
rect 2200 66600 2400 66800
rect 24600 66600 24800 66800
rect 24600 66800 24800 67000
rect 24600 67000 24800 67200
rect 81000 67000 81200 67200
rect 24600 67200 24800 67400
rect 24600 67400 24800 67600
rect 53800 67400 54000 67600
rect 24600 67600 24800 67800
rect 24600 67800 24800 68000
rect 2200 68000 2400 68200
rect 24600 68000 24800 68200
rect 54800 68000 55000 68200
rect 24600 68200 24800 68400
rect 55200 68200 55400 68400
rect 81200 68200 81400 68400
rect 24600 68400 24800 68600
rect 81200 68400 81400 68600
rect 97400 68400 97600 68600
rect 24600 68600 24800 68800
rect 57200 68600 75200 68800
rect 81200 68600 81400 68800
rect 97200 68600 97400 68800
rect 3000 68800 3200 69000
rect 24600 68800 24800 69000
rect 81200 68800 81400 69000
rect 3800 69000 14000 69200
rect 24600 69000 24800 69200
rect 81200 69000 81400 69200
rect 86000 69000 96200 69200
rect 24600 69200 24800 69400
rect 81200 69200 81400 69400
rect 24600 69400 24800 69600
rect 81200 69400 81400 69600
rect 24600 69600 24800 69800
rect 81200 69600 81400 69800
rect 24600 69800 24800 70000
rect 81200 69800 81400 70000
rect 24600 70000 24800 70200
rect 81200 70000 81400 70200
rect 24600 70200 24800 70400
rect 81200 70200 81400 70400
rect 24600 70400 24800 70600
rect 81200 70400 81400 70600
rect 24600 70600 24800 70800
rect 81200 70600 81400 70800
rect 24600 70800 24800 71000
rect 81200 70800 81400 71000
rect 24600 71000 24800 71200
rect 81200 71000 81400 71200
rect 24600 71200 24800 71400
rect 81200 71200 81400 71400
rect 24600 71400 24800 71600
rect 81200 71400 81400 71600
rect 24600 71600 24800 71800
rect 81200 71600 81400 71800
rect 24600 71800 24800 72000
rect 81200 71800 81400 72000
rect 24600 72000 24800 72200
rect 81200 72000 81400 72200
rect 24600 72200 24800 72400
rect 81200 72200 81400 72400
rect 3400 72400 14000 72600
rect 24600 72400 24800 72600
rect 81200 72400 81400 72600
rect 86000 72400 96600 72600
rect 24600 72600 24800 72800
rect 81200 72600 81400 72800
rect 24600 72800 24800 73000
rect 81200 72800 81400 73000
rect 97200 72800 97400 73000
rect 24600 73000 24800 73200
rect 81200 73000 81400 73200
rect 97400 73000 97600 73200
rect 24600 73200 24800 73400
rect 81200 73200 81400 73400
rect 2200 73400 2400 73600
rect 24600 73400 24800 73600
rect 81200 73400 81400 73600
rect 24600 73600 24800 73800
rect 81200 73600 81400 73800
rect 24600 73800 24800 74000
rect 81200 73800 81400 74000
rect 24600 74000 24800 74200
rect 81200 74000 81400 74200
rect 24600 74200 24800 74400
rect 81200 74200 81400 74400
rect 24600 74400 24800 74600
rect 81200 74400 81400 74600
rect 51400 74600 51600 74800
rect 81200 74600 81400 74800
rect 2200 74800 2400 75000
rect 81200 74800 81400 75000
rect 2600 75400 2800 75600
rect 3400 75800 3600 76000
rect 96400 75800 96600 76000
rect 18800 76000 19000 76200
rect 81000 76000 81200 76200
rect 19000 76600 19200 76800
rect 19400 77400 19600 77600
rect 19600 77800 19800 78000
rect 79400 78800 79600 79000
rect 14000 79200 14200 79400
rect 3000 79400 3200 79600
rect 96800 79400 97000 79600
rect 78000 79800 78200 80000
rect 22200 80000 22400 80200
rect 77600 80000 77800 80200
rect 23400 80400 23600 80600
rect 76400 80400 76600 80600
rect 97600 81800 97800 82000
rect 2400 82000 2600 82200
rect 2800 82400 3000 82600
rect 96600 82600 96800 82800
rect 85800 84600 86000 84800
rect 85600 85200 85800 85400
rect 14800 85800 15000 86000
rect 15200 86000 15400 86200
rect 84600 86000 84800 86200
rect 44800 86200 45000 86400
rect 48200 86200 48400 86400
rect 75600 86200 75800 86400
rect 44800 86400 45000 86600
rect 48200 86400 48400 86600
rect 75600 86400 75800 86600
rect 44800 86600 45000 86800
rect 48200 86600 48400 86800
rect 75600 86600 75800 86800
rect 44800 86800 45000 87000
rect 48200 86800 48400 87000
rect 75600 86800 75800 87000
rect 44800 87000 45000 87200
rect 48200 87000 48400 87200
rect 75600 87000 75800 87200
rect 44800 87200 45000 87400
rect 48200 87200 48400 87400
rect 75600 87200 75800 87400
rect 44800 87400 45000 87600
rect 48200 87400 48400 87600
rect 75600 87400 75800 87600
rect 44800 87600 45000 87800
rect 48200 87600 48400 87800
rect 75600 87600 75800 87800
rect 44800 87800 45000 88000
rect 48200 87800 48400 88000
rect 75600 87800 75800 88000
rect 44800 88000 45000 88200
rect 48200 88000 48400 88200
rect 75600 88000 75800 88200
rect 44800 88200 45000 88400
rect 48200 88200 48400 88400
rect 75600 88200 75800 88400
rect 44800 88400 45000 88600
rect 48200 88400 48400 88600
rect 75600 88400 75800 88600
rect 44800 88600 45000 88800
rect 48200 88600 48400 88800
rect 75600 88600 75800 88800
rect 44800 88800 45000 89000
rect 48200 88800 48400 89000
rect 75600 88800 75800 89000
rect 44800 89000 45000 89200
rect 48200 89000 48400 89200
rect 75600 89000 75800 89200
rect 44800 89200 45000 89400
rect 48200 89200 48400 89400
rect 75600 89200 75800 89400
rect 44800 89400 45000 89600
rect 48200 89400 48400 89600
rect 75600 89400 75800 89600
rect 44800 89600 45000 89800
rect 48200 89600 48400 89800
rect 75600 89600 75800 89800
rect 44800 89800 45000 90000
rect 48200 89800 48400 90000
rect 75600 89800 75800 90000
rect 44800 90000 45000 90200
rect 48200 90000 48400 90200
rect 75600 90000 75800 90200
rect 44800 90200 45000 90400
rect 48200 90200 48400 90400
rect 75600 90200 75800 90400
rect 44800 90400 45000 90600
rect 48200 90400 48400 90600
rect 75600 90400 75800 90600
rect 44800 90600 45000 90800
rect 48200 90600 48400 90800
rect 75600 90600 75800 90800
rect 44800 90800 45000 91000
rect 48200 90800 48400 91000
rect 75600 90800 75800 91000
rect 44800 91000 45000 91200
rect 48200 91000 48400 91200
rect 75600 91000 75800 91200
rect 44800 91200 45000 91400
rect 48200 91200 48400 91400
rect 75600 91200 75800 91400
rect 44800 91400 45000 91600
rect 48200 91400 48400 91600
rect 75600 91400 75800 91600
rect 44800 91600 45000 91800
rect 48200 91600 48400 91800
rect 75600 91600 75800 91800
rect 44800 91800 45000 92000
rect 48200 91800 48400 92000
rect 75600 91800 75800 92000
rect 44800 92000 45000 92200
rect 48200 92000 48400 92200
rect 75600 92000 75800 92200
rect 44800 92200 45000 92400
rect 48200 92200 48400 92400
rect 75600 92200 75800 92400
rect 44800 92400 45000 92600
rect 48200 92400 48400 92600
rect 75600 92400 75800 92600
rect 44800 92600 45000 92800
rect 48200 92600 48400 92800
rect 75600 92600 75800 92800
rect 44800 92800 45000 93000
rect 48200 92800 48400 93000
rect 75600 92800 75800 93000
rect 44800 93000 45000 93200
rect 48200 93000 48400 93200
rect 75600 93000 75800 93200
rect 44800 93200 45000 93400
rect 48200 93200 48400 93400
rect 75600 93200 75800 93400
rect 44800 93400 45000 93600
rect 48200 93400 48400 93600
rect 75600 93400 75800 93600
rect 44800 93600 45000 93800
rect 48200 93600 48400 93800
rect 75600 93600 75800 93800
rect 44800 93800 45000 94000
rect 48200 93800 48400 94000
rect 75600 93800 75800 94000
rect 44800 94000 45000 94200
rect 48200 94000 48400 94200
rect 75600 94000 75800 94200
rect 44800 94200 45000 94400
rect 48200 94200 48400 94400
rect 75600 94200 75800 94400
rect 44800 94400 45000 94600
rect 48200 94400 48400 94600
rect 75600 94400 75800 94600
rect 44800 94600 45000 94800
rect 48200 94600 48400 94800
rect 75600 94600 75800 94800
rect 44800 94800 45000 95000
rect 48200 94800 48400 95000
rect 75600 94800 75800 95000
rect 44800 95000 45000 95200
rect 48200 95000 48400 95200
rect 75600 95000 75800 95200
rect 44800 95200 45000 95400
rect 48200 95200 48400 95400
rect 75600 95200 75800 95400
rect 44800 95400 45000 95600
rect 48200 95400 48400 95600
rect 75600 95400 75800 95600
rect 44800 95600 45000 95800
rect 48200 95600 48400 95800
rect 75600 95600 75800 95800
rect 44800 95800 45000 96000
rect 48200 95800 48400 96000
rect 75600 95800 75800 96000
rect 44800 96000 45000 96200
rect 48200 96000 48400 96200
rect 75600 96000 75800 96200
rect 44800 96200 45000 96400
rect 48200 96200 48400 96400
rect 75600 96200 75800 96400
rect 44800 96400 45000 96600
rect 48200 96400 48400 96600
rect 72200 96400 72400 96600
rect 82400 96400 82600 96600
rect 38000 96600 38200 96800
rect 48200 96600 48400 96800
rect 72200 96600 72400 96800
rect 82400 96600 82600 96800
rect 20800 96800 21000 97000
rect 55000 96800 55200 97000
rect 65400 96800 65600 97000
rect 24400 97000 24600 97200
rect 34400 97000 34600 97200
rect 58600 97000 58800 97200
rect 68600 97000 68800 97200
rect 48000 97200 48200 97400
rect 72400 97200 72600 97400
rect 82200 97200 82400 97400
rect 34200 97400 34400 97600
rect 52000 97400 52200 97600
rect 68400 97400 68600 97600
rect 24800 97600 25000 97800
rect 34000 97600 34200 97800
rect 59000 97600 59200 97800
rect 18200 97800 18400 98000
rect 40600 97800 40800 98000
rect 45600 97800 45800 98000
rect 52400 97800 52600 98000
rect 74800 97800 75000 98000
rect 79800 97800 80000 98000
rect 19600 98000 19800 98200
rect 39200 98000 39400 98200
rect 40200 98000 40400 98200
rect 46000 98000 46200 98200
rect 47000 98000 47200 98200
rect 53800 98000 54000 98200
rect 66600 98000 66800 98200
rect 73400 98000 73600 98200
rect 74400 98000 74600 98200
rect 80200 98000 80400 98200
rect 81200 98000 81400 98200
<< metal3 >>
rect 25200 2400 25400 2600
rect 33600 2400 33800 2600
rect 59400 2400 59600 2600
rect 67800 2400 68000 2600
rect 20200 2600 20400 2800
rect 38600 2600 38800 2800
rect 54400 2600 54600 2800
rect 66000 2600 66200 2800
rect 38400 2800 38600 3000
rect 47800 2800 48000 3000
rect 72600 2800 72800 3000
rect 82000 2800 82200 3000
rect 20600 3000 20800 3200
rect 31400 3000 31600 3200
rect 54800 3000 55000 3200
rect 65600 3000 65800 3200
rect 17600 3200 17800 3400
rect 51800 3200 52000 3400
rect 68600 3200 68800 3400
rect 20800 3400 21000 3600
rect 31200 3400 31400 3600
rect 55000 3400 55200 3600
rect 65400 3400 65600 3600
rect 44800 3600 45000 3800
rect 48200 3600 48400 3800
rect 72200 3600 72400 3800
rect 82400 3600 82600 3800
rect 41400 3800 41600 4000
rect 44800 3800 45000 4000
rect 75600 3800 75800 4000
rect 79000 3800 79200 4000
rect 17400 4000 17600 4200
rect 41400 4000 41600 4200
rect 75600 4000 75800 4200
rect 79000 4000 79200 4200
rect 17400 4200 17600 4400
rect 41400 4200 41600 4400
rect 79000 4200 79200 4400
rect 17400 4400 17600 4600
rect 41400 4400 41600 4600
rect 79000 4400 79200 4600
rect 17400 4600 17600 4800
rect 41400 4600 41600 4800
rect 79000 4600 79200 4800
rect 17400 4800 17600 5000
rect 41400 4800 41600 5000
rect 79000 4800 79200 5000
rect 17400 5000 17600 5200
rect 41400 5000 41600 5200
rect 79000 5000 79200 5200
rect 17400 5200 17600 5400
rect 41400 5200 41600 5400
rect 79000 5200 79200 5400
rect 17400 5400 17600 5600
rect 41400 5400 41600 5600
rect 79000 5400 79200 5600
rect 17400 5600 17600 5800
rect 41400 5600 41600 5800
rect 79000 5600 79200 5800
rect 17400 5800 17600 6000
rect 41400 5800 41600 6000
rect 79000 5800 79200 6000
rect 17400 6000 17600 6200
rect 41400 6000 41600 6200
rect 79000 6000 79200 6200
rect 17400 6200 17600 6400
rect 41400 6200 41600 6400
rect 79000 6200 79200 6400
rect 17400 6400 17600 6600
rect 41400 6400 41600 6600
rect 79000 6400 79200 6600
rect 17400 6600 17600 6800
rect 41400 6600 41600 6800
rect 79000 6600 79200 6800
rect 17400 6800 17600 7000
rect 41400 6800 41600 7000
rect 79000 6800 79200 7000
rect 17400 7000 17600 7200
rect 41400 7000 41600 7200
rect 79000 7000 79200 7200
rect 17400 7200 17600 7400
rect 41400 7200 41600 7400
rect 79000 7200 79200 7400
rect 17400 7400 17600 7600
rect 41400 7400 41600 7600
rect 79000 7400 79200 7600
rect 17400 7600 17600 7800
rect 41400 7600 41600 7800
rect 79000 7600 79200 7800
rect 17400 7800 17600 8000
rect 41400 7800 41600 8000
rect 79000 7800 79200 8000
rect 17400 8000 17600 8200
rect 41400 8000 41600 8200
rect 79000 8000 79200 8200
rect 17400 8200 17600 8400
rect 41400 8200 41600 8400
rect 79000 8200 79200 8400
rect 17400 8400 17600 8600
rect 41400 8400 41600 8600
rect 79000 8400 79200 8600
rect 17400 8600 17600 8800
rect 41400 8600 41600 8800
rect 79000 8600 79200 8800
rect 17400 8800 17600 9000
rect 41400 8800 41600 9000
rect 79000 8800 79200 9000
rect 17400 9000 17600 9200
rect 41400 9000 41600 9200
rect 79000 9000 79200 9200
rect 17400 9200 17600 9400
rect 41400 9200 41600 9400
rect 79000 9200 79200 9400
rect 17400 9400 17600 9600
rect 41400 9400 41600 9600
rect 79000 9400 79200 9600
rect 17400 9600 17600 9800
rect 41400 9600 41600 9800
rect 79000 9600 79200 9800
rect 17400 9800 17600 10000
rect 41400 9800 41600 10000
rect 79000 9800 79200 10000
rect 17400 10000 17600 10200
rect 41400 10000 41600 10200
rect 79000 10000 79200 10200
rect 17400 10200 17600 10400
rect 41400 10200 41600 10400
rect 79000 10200 79200 10400
rect 17400 10400 17600 10600
rect 41400 10400 41600 10600
rect 79000 10400 79200 10600
rect 17400 10600 17600 10800
rect 41400 10600 41600 10800
rect 79000 10600 79200 10800
rect 17400 10800 17600 11000
rect 41400 10800 41600 11000
rect 79000 10800 79200 11000
rect 17400 11000 17600 11200
rect 41400 11000 41600 11200
rect 79000 11000 79200 11200
rect 17400 11200 17600 11400
rect 41400 11200 41600 11400
rect 79000 11200 79200 11400
rect 17400 11400 17600 11600
rect 41400 11400 41600 11600
rect 79000 11400 79200 11600
rect 17400 11600 17600 11800
rect 41400 11600 41600 11800
rect 79000 11600 79200 11800
rect 17400 11800 17600 12000
rect 41400 11800 41600 12000
rect 79000 11800 79200 12000
rect 17400 12000 17600 12200
rect 41400 12000 41600 12200
rect 79000 12000 79200 12200
rect 17400 12200 17600 12400
rect 41400 12200 41600 12400
rect 79000 12200 79200 12400
rect 17400 12400 17600 12600
rect 41400 12400 41600 12600
rect 79000 12400 79200 12600
rect 17400 12600 17600 12800
rect 41400 12600 41600 12800
rect 79000 12600 79200 12800
rect 17400 12800 17600 13000
rect 41400 12800 41600 13000
rect 79000 12800 79200 13000
rect 17400 13000 17600 13200
rect 41400 13000 41600 13200
rect 79000 13000 79200 13200
rect 17400 13200 17600 13400
rect 41400 13200 41600 13400
rect 79000 13200 79200 13400
rect 17400 13400 17600 13600
rect 41400 13400 41600 13600
rect 79000 13400 79200 13600
rect 17400 13600 17600 13800
rect 41400 13600 41600 13800
rect 79000 13600 79200 13800
rect 17400 13800 17600 14000
rect 41400 13800 41600 14000
rect 79000 13800 79200 14000
rect 17400 14000 17600 14200
rect 41400 14000 41600 14200
rect 79000 14000 79200 14200
rect 15600 14200 15800 14400
rect 84400 14200 84600 14400
rect 85200 14600 85400 14800
rect 85400 14800 85600 15000
rect 14000 15800 14200 16000
rect 14000 16000 14200 16200
rect 14000 16200 14200 16400
rect 14000 16400 14200 16600
rect 14000 16600 14200 16800
rect 14000 16800 14200 17000
rect 14000 17000 14200 17200
rect 14000 17200 14200 17400
rect 14000 17400 14200 17600
rect 97400 18200 97600 18400
rect 2200 18600 2400 18800
rect 43400 19200 43600 19400
rect 51400 19200 51600 19400
rect 97800 19200 98000 19400
rect 44200 19400 44400 19600
rect 51400 19400 51600 19600
rect 97800 19400 98000 19600
rect 44800 19600 45000 19800
rect 51400 19600 51600 19800
rect 97800 19600 98000 19800
rect 45200 19800 45400 20000
rect 51400 19800 51600 20000
rect 51400 20000 51600 20200
rect 51400 20200 51600 20400
rect 97600 20200 97800 20400
rect 2400 20400 2600 20600
rect 51400 20400 51600 20600
rect 51400 20600 51600 20800
rect 46600 20800 46800 21000
rect 51400 20800 51600 21000
rect 97000 20800 97200 21000
rect 46800 21000 47000 21200
rect 51400 21000 51600 21200
rect 96600 21000 96800 21200
rect 14000 21200 14200 21400
rect 51400 21200 51600 21400
rect 14000 21400 14200 21600
rect 51400 21400 51600 21600
rect 14000 21600 14200 21800
rect 51400 21600 51600 21800
rect 14000 21800 14200 22000
rect 51400 21800 51600 22000
rect 14000 22000 14200 22200
rect 51400 22000 51600 22200
rect 14000 22200 14200 22400
rect 51400 22200 51600 22400
rect 14000 22400 14200 22600
rect 51400 22400 51600 22600
rect 14000 22600 14200 22800
rect 51400 22600 51600 22800
rect 14000 22800 14200 23000
rect 51400 22800 51600 23000
rect 14000 23000 14200 23200
rect 51400 23000 51600 23200
rect 14000 23200 14200 23400
rect 51400 23200 51600 23400
rect 14000 23400 14200 23600
rect 51400 23400 51600 23600
rect 14000 23600 14200 23800
rect 51400 23600 51600 23800
rect 14000 23800 14200 24000
rect 51400 23800 51600 24000
rect 14000 24000 14200 24200
rect 51400 24000 51600 24200
rect 14000 24200 14200 24400
rect 51400 24200 51600 24400
rect 14000 24400 14200 24600
rect 51400 24400 51600 24600
rect 48400 24600 48600 24800
rect 51400 24600 51600 24800
rect 96800 24600 97000 24800
rect 48400 24800 48600 25000
rect 51400 24800 51600 25000
rect 48400 25000 48600 25200
rect 51400 25000 51600 25200
rect 48400 25200 48600 25400
rect 51400 25200 51600 25400
rect 48400 25400 48600 25600
rect 51400 25400 51600 25600
rect 48400 25600 48600 25800
rect 51400 25600 51600 25800
rect 48400 25800 48600 26000
rect 51400 25800 51600 26000
rect 48400 26000 48600 26200
rect 51400 26000 51600 26200
rect 97800 26000 98000 26200
rect 48400 26200 48600 26400
rect 51400 26200 51600 26400
rect 97800 26200 98000 26400
rect 48400 26400 48600 26600
rect 51400 26400 51600 26600
rect 97800 26400 98000 26600
rect 48400 26600 48600 26800
rect 51400 26600 51600 26800
rect 48400 26800 48600 27000
rect 51400 26800 51600 27000
rect 48400 27000 48600 27200
rect 51400 27000 51600 27200
rect 48400 27200 48600 27400
rect 51400 27200 51600 27400
rect 48400 27400 48600 27600
rect 51400 27400 51600 27600
rect 48400 27600 48600 27800
rect 51400 27600 51600 27800
rect 3200 27800 3400 28000
rect 48400 27800 48600 28000
rect 51400 27800 51600 28000
rect 14000 28000 14200 28200
rect 48400 28000 48600 28200
rect 51400 28000 51600 28200
rect 14000 28200 14200 28400
rect 48400 28200 48600 28400
rect 51400 28200 51600 28400
rect 14000 28400 14200 28600
rect 48400 28400 48600 28600
rect 51400 28400 51600 28600
rect 14000 28600 14200 28800
rect 48400 28600 48600 28800
rect 51400 28600 51600 28800
rect 14000 28800 14200 29000
rect 48400 28800 48600 29000
rect 51400 28800 51600 29000
rect 14000 29000 14200 29200
rect 48400 29000 48600 29200
rect 51400 29000 51600 29200
rect 14000 29200 14200 29400
rect 48400 29200 48600 29400
rect 51400 29200 51600 29400
rect 14000 29400 14200 29600
rect 48400 29400 48600 29600
rect 51400 29400 51600 29600
rect 14000 29600 14200 29800
rect 48400 29600 48600 29800
rect 51400 29600 51600 29800
rect 14000 29800 14200 30000
rect 48400 29800 48600 30000
rect 51400 29800 51600 30000
rect 14000 30000 14200 30200
rect 48400 30000 48600 30200
rect 51400 30000 51600 30200
rect 14000 30200 14200 30400
rect 48400 30200 48600 30400
rect 51400 30200 51600 30400
rect 14000 30400 14200 30600
rect 48400 30400 48600 30600
rect 51400 30400 51600 30600
rect 14000 30600 14200 30800
rect 48400 30600 48600 30800
rect 51400 30600 51600 30800
rect 14000 30800 14200 31000
rect 48400 30800 48600 31000
rect 51400 30800 51600 31000
rect 14000 31000 14200 31200
rect 48400 31000 48600 31200
rect 51400 31000 51600 31200
rect 14000 31200 14200 31400
rect 48400 31200 48600 31400
rect 76600 31200 76800 31400
rect 3200 31400 3400 31600
rect 22600 31400 22800 31600
rect 48400 31400 48600 31600
rect 77200 31400 77400 31600
rect 48400 31600 48600 31800
rect 21800 31800 22000 32000
rect 2400 32000 2600 32200
rect 21400 32000 21600 32200
rect 78400 32000 78600 32200
rect 97600 32200 97800 32400
rect 51600 32400 51800 32600
rect 48200 32600 48400 32800
rect 79200 32600 79400 32800
rect 20400 32800 20600 33000
rect 97800 32800 98000 33000
rect 79600 33000 79800 33200
rect 97800 33000 98000 33200
rect 48000 33200 48200 33400
rect 97800 33200 98000 33400
rect 47800 33600 48000 33800
rect 2200 33800 2400 34000
rect 19600 33800 19800 34000
rect 47600 34000 47800 34200
rect 19400 34200 19600 34400
rect 97400 34200 97600 34400
rect 3000 34600 3200 34800
rect 47200 34600 47400 34800
rect 96800 34600 97000 34800
rect 47000 34800 47200 35000
rect 52800 34800 53000 35000
rect 14000 35000 14200 35200
rect 19000 35000 19200 35200
rect 80800 35000 81000 35200
rect 14000 35200 14200 35400
rect 14000 35400 14200 35600
rect 53400 35400 53600 35600
rect 14000 35600 14200 35800
rect 46200 35600 46400 35800
rect 53600 35600 53800 35800
rect 81000 35600 81200 35800
rect 14000 35800 14200 36000
rect 18800 35800 19000 36000
rect 14000 36000 14200 36200
rect 14000 36200 14200 36400
rect 14000 36400 14200 36600
rect 14000 36600 14200 36800
rect 14000 36800 14200 37000
rect 43800 36800 44000 37000
rect 56000 36800 56200 37000
rect 14000 37000 14200 37200
rect 24600 37000 24800 37200
rect 75200 37000 75400 37200
rect 14000 37200 14200 37400
rect 14000 37400 14200 37600
rect 14000 37600 14200 37800
rect 14000 37800 14200 38000
rect 14000 38000 14200 38200
rect 97800 39600 98000 39800
rect 97800 39800 98000 40000
rect 97800 40000 98000 40200
rect 3600 41600 3800 41800
rect 96200 41600 96600 41800
rect 14000 41800 14200 42000
rect 14000 42000 14200 42200
rect 14000 42200 14200 42400
rect 14000 42400 14200 42600
rect 14000 42600 14200 42800
rect 14000 42800 14200 43000
rect 14000 43000 14200 43200
rect 48400 43000 48600 43200
rect 14000 43200 14200 43400
rect 48400 43200 48600 43400
rect 51400 43200 51600 43400
rect 14000 43400 14200 43600
rect 48400 43400 48600 43600
rect 51400 43400 51600 43600
rect 14000 43600 14200 43800
rect 48400 43600 48600 43800
rect 51400 43600 51600 43800
rect 14000 43800 14200 44000
rect 48400 43800 48600 44000
rect 51400 43800 51600 44000
rect 14000 44000 14200 44200
rect 48400 44000 48600 44200
rect 51400 44000 51600 44200
rect 14000 44200 14200 44400
rect 18800 44200 19000 44400
rect 48400 44200 48600 44400
rect 51400 44200 51600 44400
rect 14000 44400 14200 44600
rect 48400 44400 48600 44600
rect 51400 44400 51600 44600
rect 14000 44600 14200 44800
rect 48400 44600 48600 44800
rect 51400 44600 51600 44800
rect 14000 44800 14200 45000
rect 48400 44800 48600 45000
rect 51400 44800 51600 45000
rect 3600 45000 3800 45200
rect 48400 45000 48600 45200
rect 51400 45000 51600 45200
rect 80800 45000 81000 45200
rect 96200 45000 96600 45200
rect 48400 45200 48600 45400
rect 51400 45200 51600 45400
rect 19200 45400 19400 45600
rect 48400 45400 48600 45600
rect 51400 45400 51600 45600
rect 80600 45400 80800 45600
rect 48400 45600 48600 45800
rect 51400 45600 51600 45800
rect 97400 45600 97600 45800
rect 48400 45800 48600 46000
rect 51400 45800 51600 46000
rect 80400 45800 80600 46000
rect 2200 46000 2400 46200
rect 48400 46000 48600 46200
rect 51400 46000 51600 46200
rect 48400 46200 48600 46400
rect 51400 46200 51600 46400
rect 80200 46200 80400 46400
rect 19800 46400 20000 46600
rect 48400 46400 48600 46600
rect 51400 46400 51600 46600
rect 48400 46600 48600 46800
rect 51400 46600 51600 46800
rect 97800 46600 98000 46800
rect 48400 46800 48600 47000
rect 51400 46800 51600 47000
rect 97800 46800 98000 47000
rect 48400 47000 48600 47200
rect 51400 47000 51600 47200
rect 97800 47000 98000 47200
rect 48400 47200 48600 47400
rect 51400 47200 51600 47400
rect 48400 47400 48600 47600
rect 51400 47400 51600 47600
rect 48400 47600 48600 47800
rect 51400 47600 51600 47800
rect 97600 47600 97800 47800
rect 2400 47800 2600 48000
rect 21200 47800 21400 48000
rect 48400 47800 48600 48000
rect 51400 47800 51600 48000
rect 48400 48000 48600 48200
rect 51400 48000 51600 48200
rect 48400 48200 48600 48400
rect 51400 48200 51600 48400
rect 97000 48200 97200 48400
rect 48400 48400 48600 48600
rect 51400 48400 51600 48600
rect 96600 48400 96800 48600
rect 14000 48600 14200 48800
rect 22800 48600 23000 48800
rect 48400 48600 48600 48800
rect 51400 48600 51600 48800
rect 77000 48600 77200 48800
rect 14000 48800 14200 49000
rect 23600 48800 24000 49000
rect 48400 48800 48600 49000
rect 51400 48800 51600 49000
rect 76200 48800 76400 49000
rect 14000 49000 14200 49200
rect 14000 49200 14200 49400
rect 14000 49400 14200 49600
rect 14000 49600 14200 49800
rect 14000 49800 14200 50000
rect 14000 50000 14200 50200
rect 14000 50200 14200 50400
rect 14000 50400 14200 50600
rect 14000 50600 14200 50800
rect 14000 50800 14200 51000
rect 23600 50800 24000 51000
rect 48400 50800 48600 51000
rect 51400 50800 51600 51000
rect 14000 51000 14200 51200
rect 22800 51000 23000 51200
rect 48400 51000 48600 51200
rect 51400 51000 51600 51200
rect 14000 51200 14200 51400
rect 48400 51200 48600 51400
rect 51400 51200 51600 51400
rect 14000 51400 14200 51600
rect 48400 51400 48600 51600
rect 51400 51400 51600 51600
rect 14000 51600 14200 51800
rect 48400 51600 48600 51800
rect 51400 51600 51600 51800
rect 21200 51800 21400 52000
rect 48400 51800 48600 52000
rect 51400 51800 51600 52000
rect 48400 52000 48600 52200
rect 51400 52000 51600 52200
rect 96800 52000 97000 52200
rect 48400 52200 48600 52400
rect 51400 52200 51600 52400
rect 48400 52400 48600 52600
rect 51400 52400 51600 52600
rect 48400 52600 48600 52800
rect 51400 52600 51600 52800
rect 48400 52800 48600 53000
rect 51400 52800 51600 53000
rect 48400 53000 48600 53200
rect 51400 53000 51600 53200
rect 19800 53200 20000 53400
rect 48400 53200 48600 53400
rect 51400 53200 51600 53400
rect 48400 53400 48600 53600
rect 51400 53400 51600 53600
rect 97800 53400 98000 53600
rect 48400 53600 48600 53800
rect 51400 53600 51600 53800
rect 97800 53600 98000 53800
rect 48400 53800 48600 54000
rect 51400 53800 51600 54000
rect 97800 53800 98000 54000
rect 48400 54000 48600 54200
rect 51400 54000 51600 54200
rect 19200 54200 19400 54400
rect 48400 54200 48600 54400
rect 51400 54200 51600 54400
rect 48400 54400 48600 54600
rect 51400 54400 51600 54600
rect 48400 54600 48600 54800
rect 51400 54600 51600 54800
rect 48400 54800 48600 55000
rect 51400 54800 51600 55000
rect 48400 55000 48600 55200
rect 51400 55000 51600 55200
rect 3200 55200 3400 55400
rect 48400 55200 48600 55400
rect 51400 55200 51600 55400
rect 14000 55400 14200 55600
rect 18800 55400 19000 55600
rect 48400 55400 48600 55600
rect 51400 55400 51600 55600
rect 14000 55600 14200 55800
rect 48400 55600 48600 55800
rect 51400 55600 51600 55800
rect 14000 55800 14200 56000
rect 48400 55800 48600 56000
rect 51400 55800 51600 56000
rect 14000 56000 14200 56200
rect 48400 56000 48600 56200
rect 51400 56000 51600 56200
rect 14000 56200 14200 56400
rect 48400 56200 48600 56400
rect 51400 56200 51600 56400
rect 14000 56400 14200 56600
rect 48400 56400 48600 56600
rect 51400 56400 51600 56600
rect 14000 56600 14200 56800
rect 48400 56600 48600 56800
rect 51400 56600 51600 56800
rect 14000 56800 14200 57000
rect 51400 56800 51600 57000
rect 14000 57000 14200 57200
rect 51400 57000 51600 57200
rect 14000 57200 14200 57400
rect 51400 57200 51600 57400
rect 14000 57400 14200 57600
rect 51400 57400 51600 57600
rect 14000 57600 14200 57800
rect 51400 57600 51600 57800
rect 14000 57800 14200 58000
rect 51400 57800 51600 58000
rect 14000 58000 14200 58200
rect 51400 58000 51600 58200
rect 14000 58200 14200 58400
rect 51400 58200 51600 58400
rect 14000 58400 14200 58600
rect 51400 58400 51600 58600
rect 14000 58600 14200 58800
rect 51400 58600 51600 58800
rect 3200 58800 3400 59000
rect 51400 58800 51600 59000
rect 51400 59000 51600 59200
rect 51400 59200 51600 59400
rect 2400 59400 2600 59600
rect 51400 59400 51600 59600
rect 51400 59600 51600 59800
rect 97600 59600 97800 59800
rect 51400 59800 51600 60000
rect 51400 60000 51600 60200
rect 51400 60200 51600 60400
rect 97800 60200 98000 60400
rect 51400 60400 51600 60600
rect 97800 60400 98000 60600
rect 51400 60600 51600 60800
rect 97800 60600 98000 60800
rect 51400 60800 51600 61000
rect 51400 61000 51600 61200
rect 2200 61200 2400 61400
rect 51400 61200 51600 61400
rect 51400 61400 51600 61600
rect 51400 61600 51600 61800
rect 97400 61600 97600 61800
rect 51400 61800 51600 62000
rect 3000 62000 3200 62200
rect 51400 62000 51600 62200
rect 96800 62000 97000 62200
rect 51400 62200 51600 62400
rect 14000 62400 14200 62600
rect 51400 62400 51600 62600
rect 14000 62600 14200 62800
rect 51400 62600 51600 62800
rect 14000 62800 14200 63000
rect 76600 62800 76800 63000
rect 14000 63000 14200 63200
rect 77200 63000 77400 63200
rect 14000 63200 14200 63400
rect 14000 63400 14200 63600
rect 14000 63600 14200 63800
rect 78400 63600 78600 63800
rect 14000 63800 14200 64000
rect 14000 64000 14200 64200
rect 51600 64000 51800 64200
rect 14000 64200 14200 64400
rect 79200 64200 79400 64400
rect 14000 64400 14200 64600
rect 14000 64600 14200 64800
rect 79600 64600 79800 64800
rect 14000 64800 14200 65000
rect 14000 65000 14200 65200
rect 14000 65200 14200 65400
rect 14000 65400 14200 65600
rect 3200 65600 3400 65800
rect 2400 66200 2600 66400
rect 52800 66400 53000 66600
rect 97600 66400 97800 66600
rect 80800 66600 81000 66800
rect 53400 67000 53600 67200
rect 97800 67000 98000 67200
rect 53600 67200 53800 67400
rect 81000 67200 81200 67400
rect 97800 67200 98000 67400
rect 97800 67400 98000 67600
rect 56000 68400 56200 68600
rect 75200 68600 75400 68800
rect 3600 69000 3800 69200
rect 96200 69000 96600 69200
rect 14000 69200 14200 69400
rect 14000 69400 14200 69600
rect 14000 69600 14200 69800
rect 14000 69800 14200 70000
rect 14000 70000 14200 70200
rect 14000 70200 14200 70400
rect 14000 70400 14200 70600
rect 14000 70600 14200 70800
rect 14000 70800 14200 71000
rect 14000 71000 14200 71200
rect 14000 71200 14200 71400
rect 14000 71400 14200 71600
rect 14000 71600 14200 71800
rect 14000 71800 14200 72000
rect 14000 72000 14200 72200
rect 14000 72200 14200 72400
rect 97800 73800 98000 74000
rect 97800 74000 98000 74200
rect 97800 74200 98000 74400
rect 97800 74400 98000 74600
rect 48400 74600 48600 74800
rect 48400 74800 48600 75000
rect 51400 74800 51600 75000
rect 48400 75000 48600 75200
rect 51400 75000 51600 75200
rect 97600 75000 97800 75200
rect 2400 75200 2600 75400
rect 48400 75200 48600 75400
rect 51400 75200 51600 75400
rect 48400 75400 48600 75600
rect 51400 75400 51600 75600
rect 48400 75600 48600 75800
rect 51400 75600 51600 75800
rect 97000 75600 97200 75800
rect 18800 75800 19000 76000
rect 48400 75800 48600 76000
rect 51400 75800 51600 76000
rect 96600 75800 96800 76000
rect 14000 76000 14200 76200
rect 48400 76000 48600 76200
rect 51400 76000 51600 76200
rect 14000 76200 14200 76400
rect 48400 76200 48600 76400
rect 51400 76200 51600 76400
rect 14000 76400 14200 76600
rect 48400 76400 48600 76600
rect 51400 76400 51600 76600
rect 14000 76600 14200 76800
rect 48400 76600 48600 76800
rect 51400 76600 51600 76800
rect 80800 76600 81000 76800
rect 14000 76800 14200 77000
rect 48400 76800 48600 77000
rect 51400 76800 51600 77000
rect 14000 77000 14200 77200
rect 19200 77000 19400 77200
rect 48400 77000 48600 77200
rect 51400 77000 51600 77200
rect 80600 77000 80800 77200
rect 14000 77200 14200 77400
rect 48400 77200 48600 77400
rect 51400 77200 51600 77400
rect 14000 77400 14200 77600
rect 48400 77400 48600 77600
rect 51400 77400 51600 77600
rect 80400 77400 80600 77600
rect 14000 77600 14200 77800
rect 48400 77600 48600 77800
rect 51400 77600 51600 77800
rect 14000 77800 14200 78000
rect 48400 77800 48600 78000
rect 51400 77800 51600 78000
rect 80200 77800 80400 78000
rect 14000 78000 14200 78200
rect 19800 78000 20000 78200
rect 48400 78000 48600 78200
rect 51400 78000 51600 78200
rect 14000 78200 14200 78400
rect 48400 78200 48600 78400
rect 51400 78200 51600 78400
rect 14000 78400 14200 78600
rect 48400 78400 48600 78600
rect 51400 78400 51600 78600
rect 14000 78600 14200 78800
rect 48400 78600 48600 78800
rect 51400 78600 51600 78800
rect 14000 78800 14200 79000
rect 48400 78800 48600 79000
rect 51400 78800 51600 79000
rect 14000 79000 14200 79200
rect 48400 79000 48600 79200
rect 51400 79000 51600 79200
rect 48400 79200 48600 79400
rect 51400 79200 51600 79400
rect 21200 79400 21400 79600
rect 48400 79400 48600 79600
rect 51400 79400 51600 79600
rect 48400 79600 48600 79800
rect 51400 79600 51600 79800
rect 48400 79800 48600 80000
rect 51400 79800 51600 80000
rect 97400 79800 97600 80000
rect 48400 80000 48600 80200
rect 51400 80000 51600 80200
rect 2200 80200 2400 80400
rect 22800 80200 23000 80400
rect 48400 80200 48600 80400
rect 51400 80200 51600 80400
rect 77000 80200 77200 80400
rect 23600 80400 24000 80600
rect 48400 80400 48600 80600
rect 51400 80400 51600 80600
rect 76200 80400 76400 80600
rect 97800 80800 98000 81000
rect 97800 81000 98000 81200
rect 97800 81200 98000 81400
rect 3200 82600 3400 82800
rect 14000 82800 14200 83000
rect 14000 83000 14200 83200
rect 14000 83200 14200 83400
rect 14000 83400 14200 83600
rect 14000 83600 14200 83800
rect 14000 83800 14200 84000
rect 14000 84000 14200 84200
rect 14000 84200 14200 84400
rect 14000 84400 14200 84600
rect 14000 84600 14200 84800
rect 85800 84800 86000 85000
rect 14200 85200 14400 85400
rect 17400 86200 17600 86400
rect 41400 86200 41600 86400
rect 79000 86200 79200 86400
rect 17400 86400 17600 86600
rect 41400 86400 41600 86600
rect 79000 86400 79200 86600
rect 17400 86600 17600 86800
rect 41400 86600 41600 86800
rect 79000 86600 79200 86800
rect 17400 86800 17600 87000
rect 41400 86800 41600 87000
rect 79000 86800 79200 87000
rect 17400 87000 17600 87200
rect 41400 87000 41600 87200
rect 79000 87000 79200 87200
rect 17400 87200 17600 87400
rect 41400 87200 41600 87400
rect 79000 87200 79200 87400
rect 17400 87400 17600 87600
rect 41400 87400 41600 87600
rect 79000 87400 79200 87600
rect 17400 87600 17600 87800
rect 41400 87600 41600 87800
rect 79000 87600 79200 87800
rect 17400 87800 17600 88000
rect 41400 87800 41600 88000
rect 79000 87800 79200 88000
rect 17400 88000 17600 88200
rect 41400 88000 41600 88200
rect 79000 88000 79200 88200
rect 17400 88200 17600 88400
rect 41400 88200 41600 88400
rect 79000 88200 79200 88400
rect 17400 88400 17600 88600
rect 41400 88400 41600 88600
rect 79000 88400 79200 88600
rect 17400 88600 17600 88800
rect 41400 88600 41600 88800
rect 79000 88600 79200 88800
rect 17400 88800 17600 89000
rect 41400 88800 41600 89000
rect 79000 88800 79200 89000
rect 17400 89000 17600 89200
rect 41400 89000 41600 89200
rect 79000 89000 79200 89200
rect 17400 89200 17600 89400
rect 41400 89200 41600 89400
rect 79000 89200 79200 89400
rect 17400 89400 17600 89600
rect 41400 89400 41600 89600
rect 79000 89400 79200 89600
rect 17400 89600 17600 89800
rect 41400 89600 41600 89800
rect 79000 89600 79200 89800
rect 17400 89800 17600 90000
rect 41400 89800 41600 90000
rect 79000 89800 79200 90000
rect 17400 90000 17600 90200
rect 41400 90000 41600 90200
rect 79000 90000 79200 90200
rect 17400 90200 17600 90400
rect 41400 90200 41600 90400
rect 79000 90200 79200 90400
rect 17400 90400 17600 90600
rect 41400 90400 41600 90600
rect 79000 90400 79200 90600
rect 17400 90600 17600 90800
rect 41400 90600 41600 90800
rect 79000 90600 79200 90800
rect 17400 90800 17600 91000
rect 41400 90800 41600 91000
rect 79000 90800 79200 91000
rect 17400 91000 17600 91200
rect 41400 91000 41600 91200
rect 79000 91000 79200 91200
rect 17400 91200 17600 91400
rect 41400 91200 41600 91400
rect 79000 91200 79200 91400
rect 17400 91400 17600 91600
rect 41400 91400 41600 91600
rect 79000 91400 79200 91600
rect 17400 91600 17600 91800
rect 41400 91600 41600 91800
rect 79000 91600 79200 91800
rect 17400 91800 17600 92000
rect 41400 91800 41600 92000
rect 79000 91800 79200 92000
rect 17400 92000 17600 92200
rect 41400 92000 41600 92200
rect 79000 92000 79200 92200
rect 17400 92200 17600 92400
rect 41400 92200 41600 92400
rect 79000 92200 79200 92400
rect 17400 92400 17600 92600
rect 41400 92400 41600 92600
rect 79000 92400 79200 92600
rect 17400 92600 17600 92800
rect 41400 92600 41600 92800
rect 79000 92600 79200 92800
rect 17400 92800 17600 93000
rect 41400 92800 41600 93000
rect 79000 92800 79200 93000
rect 17400 93000 17600 93200
rect 41400 93000 41600 93200
rect 79000 93000 79200 93200
rect 17400 93200 17600 93400
rect 41400 93200 41600 93400
rect 79000 93200 79200 93400
rect 17400 93400 17600 93600
rect 41400 93400 41600 93600
rect 79000 93400 79200 93600
rect 17400 93600 17600 93800
rect 41400 93600 41600 93800
rect 79000 93600 79200 93800
rect 17400 93800 17600 94000
rect 41400 93800 41600 94000
rect 79000 93800 79200 94000
rect 17400 94000 17600 94200
rect 41400 94000 41600 94200
rect 79000 94000 79200 94200
rect 17400 94200 17600 94400
rect 41400 94200 41600 94400
rect 79000 94200 79200 94400
rect 17400 94400 17600 94600
rect 41400 94400 41600 94600
rect 79000 94400 79200 94600
rect 17400 94600 17600 94800
rect 41400 94600 41600 94800
rect 79000 94600 79200 94800
rect 17400 94800 17600 95000
rect 41400 94800 41600 95000
rect 79000 94800 79200 95000
rect 17400 95000 17600 95200
rect 41400 95000 41600 95200
rect 79000 95000 79200 95200
rect 17400 95200 17600 95400
rect 41400 95200 41600 95400
rect 79000 95200 79200 95400
rect 17400 95400 17600 95600
rect 41400 95400 41600 95600
rect 79000 95400 79200 95600
rect 17400 95600 17600 95800
rect 41400 95600 41600 95800
rect 79000 95600 79200 95800
rect 17400 95800 17600 96000
rect 41400 95800 41600 96000
rect 79000 95800 79200 96000
rect 17400 96000 17600 96200
rect 41400 96000 41600 96200
rect 79000 96000 79200 96200
rect 17400 96200 17600 96400
rect 41400 96200 41600 96400
rect 79000 96200 79200 96400
rect 17400 96400 17600 96600
rect 41400 96400 41600 96600
rect 75600 96400 75800 96600
rect 79000 96400 79200 96600
rect 44800 96600 45000 96800
rect 75600 96600 75800 96800
rect 79000 96600 79200 96800
rect 38000 96800 38200 97000
rect 48200 96800 48400 97000
rect 72200 96800 72400 97000
rect 82400 96800 82600 97000
rect 27600 97000 27800 97200
rect 31200 97000 31400 97200
rect 61800 97000 62000 97200
rect 65400 97000 65600 97200
rect 17600 97200 17800 97400
rect 41200 97200 41400 97400
rect 45000 97200 45200 97400
rect 75400 97200 75600 97400
rect 79200 97200 79400 97400
rect 24600 97400 24800 97600
rect 27400 97400 27600 97600
rect 58800 97400 59000 97600
rect 61600 97400 61800 97600
rect 27200 97600 27400 97800
rect 31600 97600 31800 97800
rect 54600 97600 54800 97800
rect 61400 97600 61600 97800
rect 65800 97600 66000 97800
rect 25000 97800 25200 98000
rect 33800 97800 34000 98000
rect 59200 97800 59400 98000
rect 61200 97800 61400 98000
rect 68000 97800 68200 98000
rect 18600 98000 18800 98200
rect 25400 98000 25600 98200
rect 26600 98000 26800 98200
rect 32200 98000 32400 98200
rect 33400 98000 33600 98200
rect 52800 98000 53000 98200
rect 59600 98000 59800 98200
rect 60800 98000 61000 98200
rect 66400 98000 66600 98200
rect 67600 98000 67800 98200
<< metal4 >>
rect 18800 2200 19600 2400
rect 25600 2200 26600 2400
rect 32400 2200 33400 2400
rect 39400 2200 40200 2400
rect 46200 2200 47000 2400
rect 53000 2200 53800 2400
rect 59800 2200 60800 2400
rect 66600 2200 67600 2400
rect 73600 2200 74400 2400
rect 80400 2200 81200 2400
rect 20000 2400 20200 2600
rect 26800 2400 27000 2600
rect 32000 2400 32200 2600
rect 38800 2400 39000 2600
rect 54200 2400 54400 2600
rect 61000 2400 61200 2600
rect 66200 2400 66400 2600
rect 73000 2400 73200 2600
rect 18000 2600 18200 2800
rect 40800 2600 41000 2800
rect 45400 2600 45600 2800
rect 47600 2600 47800 2800
rect 72800 2600 73000 2800
rect 75000 2600 75200 2800
rect 79600 2600 79800 2800
rect 81800 2600 82000 2800
rect 17800 2800 18000 3000
rect 41000 2800 41200 3000
rect 45200 2800 45400 3000
rect 52000 2800 52200 3000
rect 75200 2800 75400 3000
rect 79400 2800 79600 3000
rect 38200 3000 38400 3200
rect 48000 3000 48200 3200
rect 72400 3000 72600 3200
rect 82200 3000 82400 3200
rect 24400 3200 24600 3400
rect 27600 3200 27800 3400
rect 34400 3200 34600 3400
rect 58600 3200 58800 3400
rect 61800 3200 62000 3400
rect 38000 3400 38200 3600
rect 48200 3400 48400 3600
rect 72200 3400 72400 3600
rect 82400 3400 82600 3600
rect 17400 3600 17600 3800
rect 41400 3600 41600 3800
rect 75600 3600 75800 3800
rect 79000 3600 79200 3800
rect 17400 3800 17600 4000
rect 34600 3800 34800 4000
rect 51600 3800 51800 4000
rect 68800 3800 69000 4000
rect 24200 4000 24400 4200
rect 34600 4000 34800 4200
rect 51600 4000 51800 4200
rect 68800 4000 69000 4200
rect 24200 4200 24400 4400
rect 34600 4200 34800 4400
rect 51600 4200 51800 4400
rect 68800 4200 69000 4400
rect 24200 4400 24400 4600
rect 34600 4400 34800 4600
rect 51600 4400 51800 4600
rect 68800 4400 69000 4600
rect 24200 4600 24400 4800
rect 34600 4600 34800 4800
rect 51600 4600 51800 4800
rect 68800 4600 69000 4800
rect 24200 4800 24400 5000
rect 34600 4800 34800 5000
rect 51600 4800 51800 5000
rect 68800 4800 69000 5000
rect 24200 5000 24400 5200
rect 34600 5000 34800 5200
rect 51600 5000 51800 5200
rect 68800 5000 69000 5200
rect 24200 5200 24400 5400
rect 34600 5200 34800 5400
rect 51600 5200 51800 5400
rect 68800 5200 69000 5400
rect 24200 5400 24400 5600
rect 34600 5400 34800 5600
rect 51600 5400 51800 5600
rect 68800 5400 69000 5600
rect 24200 5600 24400 5800
rect 34600 5600 34800 5800
rect 51600 5600 51800 5800
rect 68800 5600 69000 5800
rect 24200 5800 24400 6000
rect 34600 5800 34800 6000
rect 51600 5800 51800 6000
rect 68800 5800 69000 6000
rect 24200 6000 24400 6200
rect 34600 6000 34800 6200
rect 51600 6000 51800 6200
rect 68800 6000 69000 6200
rect 24200 6200 24400 6400
rect 34600 6200 34800 6400
rect 51600 6200 51800 6400
rect 68800 6200 69000 6400
rect 24200 6400 24400 6600
rect 34600 6400 34800 6600
rect 51600 6400 51800 6600
rect 68800 6400 69000 6600
rect 24200 6600 24400 6800
rect 34600 6600 34800 6800
rect 51600 6600 51800 6800
rect 68800 6600 69000 6800
rect 24200 6800 24400 7000
rect 34600 6800 34800 7000
rect 51600 6800 51800 7000
rect 68800 6800 69000 7000
rect 24200 7000 24400 7200
rect 34600 7000 34800 7200
rect 51600 7000 51800 7200
rect 68800 7000 69000 7200
rect 24200 7200 24400 7400
rect 34600 7200 34800 7400
rect 51600 7200 51800 7400
rect 68800 7200 69000 7400
rect 24200 7400 24400 7600
rect 34600 7400 34800 7600
rect 51600 7400 51800 7600
rect 68800 7400 69000 7600
rect 24200 7600 24400 7800
rect 34600 7600 34800 7800
rect 51600 7600 51800 7800
rect 68800 7600 69000 7800
rect 24200 7800 24400 8000
rect 34600 7800 34800 8000
rect 51600 7800 51800 8000
rect 68800 7800 69000 8000
rect 24200 8000 24400 8200
rect 34600 8000 34800 8200
rect 51600 8000 51800 8200
rect 68800 8000 69000 8200
rect 24200 8200 24400 8400
rect 34600 8200 34800 8400
rect 51600 8200 51800 8400
rect 68800 8200 69000 8400
rect 24200 8400 24400 8600
rect 34600 8400 34800 8600
rect 51600 8400 51800 8600
rect 68800 8400 69000 8600
rect 24200 8600 24400 8800
rect 34600 8600 34800 8800
rect 51600 8600 51800 8800
rect 68800 8600 69000 8800
rect 24200 8800 24400 9000
rect 34600 8800 34800 9000
rect 51600 8800 51800 9000
rect 68800 8800 69000 9000
rect 24200 9000 24400 9200
rect 34600 9000 34800 9200
rect 51600 9000 51800 9200
rect 68800 9000 69000 9200
rect 24200 9200 24400 9400
rect 34600 9200 34800 9400
rect 51600 9200 51800 9400
rect 68800 9200 69000 9400
rect 24200 9400 24400 9600
rect 34600 9400 34800 9600
rect 51600 9400 51800 9600
rect 68800 9400 69000 9600
rect 24200 9600 24400 9800
rect 34600 9600 34800 9800
rect 51600 9600 51800 9800
rect 68800 9600 69000 9800
rect 24200 9800 24400 10000
rect 34600 9800 34800 10000
rect 51600 9800 51800 10000
rect 68800 9800 69000 10000
rect 24200 10000 24400 10200
rect 34600 10000 34800 10200
rect 51600 10000 51800 10200
rect 68800 10000 69000 10200
rect 24200 10200 24400 10400
rect 34600 10200 34800 10400
rect 51600 10200 51800 10400
rect 68800 10200 69000 10400
rect 24200 10400 24400 10600
rect 34600 10400 34800 10600
rect 51600 10400 51800 10600
rect 68800 10400 69000 10600
rect 24200 10600 24400 10800
rect 34600 10600 34800 10800
rect 51600 10600 51800 10800
rect 68800 10600 69000 10800
rect 24200 10800 24400 11000
rect 34600 10800 34800 11000
rect 51600 10800 51800 11000
rect 68800 10800 69000 11000
rect 24200 11000 24400 11200
rect 34600 11000 34800 11200
rect 51600 11000 51800 11200
rect 68800 11000 69000 11200
rect 24200 11200 24400 11400
rect 34600 11200 34800 11400
rect 51600 11200 51800 11400
rect 68800 11200 69000 11400
rect 24200 11400 24400 11600
rect 34600 11400 34800 11600
rect 51600 11400 51800 11600
rect 68800 11400 69000 11600
rect 24200 11600 24400 11800
rect 34600 11600 34800 11800
rect 51600 11600 51800 11800
rect 68800 11600 69000 11800
rect 24200 11800 24400 12000
rect 34600 11800 34800 12000
rect 51600 11800 51800 12000
rect 68800 11800 69000 12000
rect 24200 12000 24400 12200
rect 34600 12000 34800 12200
rect 51600 12000 51800 12200
rect 68800 12000 69000 12200
rect 24200 12200 24400 12400
rect 34600 12200 34800 12400
rect 51600 12200 51800 12400
rect 68800 12200 69000 12400
rect 24200 12400 24400 12600
rect 34600 12400 34800 12600
rect 51600 12400 51800 12600
rect 68800 12400 69000 12600
rect 24200 12600 24400 12800
rect 34600 12600 34800 12800
rect 51600 12600 51800 12800
rect 68800 12600 69000 12800
rect 24200 12800 24400 13000
rect 34600 12800 34800 13000
rect 51600 12800 51800 13000
rect 68800 12800 69000 13000
rect 24200 13000 24400 13200
rect 34600 13000 34800 13200
rect 51600 13000 51800 13200
rect 68800 13000 69000 13200
rect 24200 13200 24400 13400
rect 34600 13200 34800 13400
rect 51600 13200 51800 13400
rect 68800 13200 69000 13400
rect 24200 13400 24400 13600
rect 34600 13400 34800 13600
rect 51600 13400 51800 13600
rect 68800 13400 69000 13600
rect 24200 13600 24400 13800
rect 34600 13600 34800 13800
rect 51600 13600 51800 13800
rect 68800 13600 69000 13800
rect 24200 13800 24400 14000
rect 34600 13800 34800 14000
rect 51600 13800 51800 14000
rect 68800 13800 69000 14000
rect 24200 14000 24400 14200
rect 34600 14000 34800 14200
rect 51600 14000 51800 14200
rect 68800 14000 69000 14200
rect 15400 14200 15600 14400
rect 85000 14400 85200 14600
rect 14600 14600 14800 14800
rect 14400 14800 14600 15000
rect 85600 15000 85800 15200
rect 85800 15400 86000 15600
rect 14000 15600 14200 15800
rect 3400 17600 14000 17800
rect 86000 17600 96600 17800
rect 2600 18000 2800 18200
rect 97200 18000 97400 18200
rect 2400 18200 2600 18400
rect 97600 18400 97800 18600
rect 97800 19000 98000 19200
rect 2000 19200 2200 19400
rect 43000 19200 43400 19400
rect 2000 19400 2200 19600
rect 2000 19600 2200 19800
rect 97800 19800 98000 20000
rect 2200 20200 2400 20400
rect 45800 20200 46000 20400
rect 2800 20800 3000 21000
rect 3200 21000 3400 21200
rect 47400 21800 47600 22000
rect 47600 22200 47800 22400
rect 48000 23000 48200 23200
rect 48200 23600 48400 23800
rect 3000 24600 3200 24800
rect 18800 25000 42600 25200
rect 57400 25000 81200 25200
rect 97400 25000 97600 25200
rect 2200 25400 2400 25600
rect 97800 25800 98000 26000
rect 2000 26000 2200 26200
rect 2000 26200 2200 26400
rect 2000 26400 2200 26600
rect 97800 26600 98000 26800
rect 2200 27000 2400 27200
rect 97400 27400 97600 27600
rect 96800 27800 97000 28000
rect 23400 31200 23600 31400
rect 76400 31200 76600 31400
rect 96800 31400 97000 31600
rect 2800 31600 3000 31800
rect 22200 31600 22400 31800
rect 77600 31600 77800 31800
rect 78000 31800 78200 32000
rect 2200 32200 2400 32400
rect 21200 32200 21400 32400
rect 48200 32400 48400 32600
rect 97800 32600 98000 32800
rect 2000 32800 2200 33000
rect 79400 32800 79600 33000
rect 2000 33000 2200 33200
rect 51800 33000 52000 33200
rect 2000 33200 2200 33400
rect 2000 33400 2200 33600
rect 97800 33400 98000 33600
rect 19800 33600 20000 33800
rect 52200 33800 52400 34000
rect 80200 33800 80400 34000
rect 97600 34000 97800 34200
rect 2400 34200 2600 34400
rect 52400 34200 52600 34400
rect 80400 34200 80600 34400
rect 97200 34400 97400 34600
rect 19200 34600 19400 34800
rect 80600 34600 80800 34800
rect 3600 34800 14000 35000
rect 86000 34800 96400 35000
rect 46800 35000 47000 35200
rect 53000 35000 53200 35200
rect 19000 35200 19200 35400
rect 53200 35200 53400 35400
rect 46400 35400 46600 35600
rect 81000 35800 81200 36000
rect 18800 36000 19000 36200
rect 45600 36000 45800 36200
rect 54200 36000 54400 36200
rect 54600 36200 54800 36400
rect 44400 36600 44600 36800
rect 55400 36600 55600 36800
rect 43600 36800 43800 37000
rect 56200 36800 56400 37000
rect 3200 38200 3400 38400
rect 96600 38200 96800 38400
rect 2800 38400 3000 38600
rect 97000 38400 97200 38600
rect 2600 38600 2800 38800
rect 2400 38800 2600 39000
rect 97600 39000 97800 39200
rect 97800 39400 98000 39600
rect 2000 39600 2200 39800
rect 2000 39800 2200 40000
rect 2000 40000 2200 40200
rect 2000 40200 2200 40400
rect 97800 40200 98000 40400
rect 97600 40800 97800 41000
rect 2400 41000 2600 41200
rect 2600 41200 2800 41400
rect 97000 41400 97200 41600
rect 3400 41600 3600 41800
rect 24600 43000 48400 43200
rect 51600 43000 75400 43200
rect 18800 44000 19000 44200
rect 81000 44200 81200 44400
rect 19000 44800 19200 45000
rect 3400 45000 3600 45200
rect 2600 45400 2800 45600
rect 97200 45400 97400 45600
rect 2400 45600 2600 45800
rect 97600 45800 97800 46000
rect 19600 46000 19800 46200
rect 80000 46400 80200 46600
rect 97800 46400 98000 46600
rect 2000 46600 2200 46800
rect 20000 46600 20200 46800
rect 79800 46600 80000 46800
rect 2000 46800 2200 47000
rect 20200 46800 20400 47000
rect 2000 47000 2200 47200
rect 97800 47200 98000 47400
rect 20800 47400 21000 47600
rect 2200 47600 2400 47800
rect 21000 47600 21200 47800
rect 78800 47600 79000 47800
rect 78600 47800 78800 48000
rect 21600 48000 21800 48200
rect 78200 48000 78400 48200
rect 2800 48200 3000 48400
rect 22000 48200 22200 48400
rect 3200 48400 3400 48600
rect 22400 48400 22600 48600
rect 23000 48600 23200 48800
rect 24000 48800 24200 49000
rect 75800 48800 76200 49000
rect 24000 50800 24400 51000
rect 23000 51000 23200 51200
rect 22400 51200 22600 51400
rect 22000 51400 22200 51600
rect 21600 51600 21800 51800
rect 3600 51800 14000 52000
rect 86000 51800 96400 52000
rect 3000 52000 3200 52200
rect 21000 52000 21200 52200
rect 20800 52200 21000 52400
rect 97400 52400 97600 52600
rect 2200 52800 2400 53000
rect 20200 52800 20400 53000
rect 20000 53000 20200 53200
rect 97800 53200 98000 53400
rect 2000 53400 2200 53600
rect 2000 53600 2200 53800
rect 19600 53600 19800 53800
rect 2000 53800 2200 54000
rect 97800 54000 98000 54200
rect 2200 54400 2400 54600
rect 19000 54800 19200 55000
rect 97400 54800 97600 55000
rect 96800 55200 97000 55400
rect 18800 55600 19000 55800
rect 24600 56600 48400 56800
rect 57400 56600 81200 56800
rect 96800 58800 97000 59000
rect 2800 59000 3000 59200
rect 2200 59600 2400 59800
rect 97800 60000 98000 60200
rect 2000 60200 2200 60400
rect 2000 60400 2200 60600
rect 2000 60600 2200 60800
rect 2000 60800 2200 61000
rect 97800 60800 98000 61000
rect 97600 61400 97800 61600
rect 2400 61600 2600 61800
rect 97200 61800 97400 62000
rect 3600 62200 14000 62400
rect 86000 62200 96400 62400
rect 76400 62800 76600 63000
rect 77600 63200 77800 63400
rect 78000 63400 78200 63600
rect 79400 64400 79600 64600
rect 51800 64600 52000 64800
rect 52200 65400 52400 65600
rect 80200 65400 80400 65600
rect 96800 65600 97000 65800
rect 2800 65800 3000 66000
rect 52400 65800 52600 66000
rect 80400 65800 80600 66000
rect 80600 66200 80800 66400
rect 2200 66400 2400 66600
rect 53000 66600 53200 66800
rect 53200 66800 53400 67000
rect 97800 66800 98000 67000
rect 2000 67000 2200 67200
rect 2000 67200 2200 67400
rect 2000 67400 2200 67600
rect 81000 67400 81200 67600
rect 2000 67600 2200 67800
rect 54200 67600 54400 67800
rect 97800 67600 98000 67800
rect 54600 67800 54800 68000
rect 55400 68200 55600 68400
rect 97600 68200 97800 68400
rect 2400 68400 2600 68600
rect 56200 68400 56400 68600
rect 2600 68600 2800 68800
rect 97000 68800 97200 69000
rect 3400 69000 3600 69200
rect 3200 72400 3400 72600
rect 96600 72400 96800 72600
rect 2800 72600 3000 72800
rect 97000 72600 97200 72800
rect 2600 72800 2800 73000
rect 2400 73000 2600 73200
rect 97600 73200 97800 73400
rect 97800 73600 98000 73800
rect 2000 73800 2200 74000
rect 2000 74000 2200 74200
rect 2000 74200 2200 74400
rect 2000 74400 2200 74600
rect 24600 74600 48400 74800
rect 51600 74600 75400 74800
rect 97800 74600 98000 74800
rect 2200 75000 2400 75200
rect 2800 75600 3000 75800
rect 18800 75600 19000 75800
rect 3200 75800 3400 76000
rect 81000 75800 81200 76000
rect 19000 76400 19200 76600
rect 19600 77600 19800 77800
rect 80000 78000 80200 78200
rect 20000 78200 20200 78400
rect 79800 78200 80000 78400
rect 20200 78400 20400 78600
rect 20800 79000 21000 79200
rect 3400 79200 14000 79400
rect 21000 79200 21200 79400
rect 78800 79200 79000 79400
rect 86000 79200 96600 79400
rect 78600 79400 78800 79600
rect 2600 79600 2800 79800
rect 21600 79600 21800 79800
rect 78200 79600 78400 79800
rect 97200 79600 97400 79800
rect 2400 79800 2600 80000
rect 22000 79800 22200 80000
rect 22400 80000 22600 80200
rect 97600 80000 97800 80200
rect 23000 80200 23200 80400
rect 24000 80400 24200 80600
rect 75800 80400 76200 80600
rect 97800 80600 98000 80800
rect 2000 80800 2200 81000
rect 2000 81000 2200 81200
rect 2000 81200 2200 81400
rect 97800 81400 98000 81600
rect 2200 81800 2400 82000
rect 97400 82200 97600 82400
rect 96800 82600 97000 82800
rect 14000 84800 14200 85000
rect 85800 85000 86000 85200
rect 85600 85400 85800 85600
rect 85400 85600 85600 85800
rect 85200 85800 85400 86000
rect 15000 86000 15200 86200
rect 84800 86000 85000 86200
rect 24200 86200 24400 86400
rect 34600 86200 34800 86400
rect 51600 86200 51800 86400
rect 68800 86200 69000 86400
rect 24200 86400 24400 86600
rect 34600 86400 34800 86600
rect 51600 86400 51800 86600
rect 68800 86400 69000 86600
rect 24200 86600 24400 86800
rect 34600 86600 34800 86800
rect 51600 86600 51800 86800
rect 68800 86600 69000 86800
rect 24200 86800 24400 87000
rect 34600 86800 34800 87000
rect 51600 86800 51800 87000
rect 68800 86800 69000 87000
rect 24200 87000 24400 87200
rect 34600 87000 34800 87200
rect 51600 87000 51800 87200
rect 68800 87000 69000 87200
rect 24200 87200 24400 87400
rect 34600 87200 34800 87400
rect 51600 87200 51800 87400
rect 68800 87200 69000 87400
rect 24200 87400 24400 87600
rect 34600 87400 34800 87600
rect 51600 87400 51800 87600
rect 68800 87400 69000 87600
rect 24200 87600 24400 87800
rect 34600 87600 34800 87800
rect 51600 87600 51800 87800
rect 68800 87600 69000 87800
rect 24200 87800 24400 88000
rect 34600 87800 34800 88000
rect 51600 87800 51800 88000
rect 68800 87800 69000 88000
rect 24200 88000 24400 88200
rect 34600 88000 34800 88200
rect 51600 88000 51800 88200
rect 68800 88000 69000 88200
rect 24200 88200 24400 88400
rect 34600 88200 34800 88400
rect 51600 88200 51800 88400
rect 68800 88200 69000 88400
rect 24200 88400 24400 88600
rect 34600 88400 34800 88600
rect 51600 88400 51800 88600
rect 68800 88400 69000 88600
rect 24200 88600 24400 88800
rect 34600 88600 34800 88800
rect 51600 88600 51800 88800
rect 68800 88600 69000 88800
rect 24200 88800 24400 89000
rect 34600 88800 34800 89000
rect 51600 88800 51800 89000
rect 68800 88800 69000 89000
rect 24200 89000 24400 89200
rect 34600 89000 34800 89200
rect 51600 89000 51800 89200
rect 68800 89000 69000 89200
rect 24200 89200 24400 89400
rect 34600 89200 34800 89400
rect 51600 89200 51800 89400
rect 68800 89200 69000 89400
rect 24200 89400 24400 89600
rect 34600 89400 34800 89600
rect 51600 89400 51800 89600
rect 68800 89400 69000 89600
rect 24200 89600 24400 89800
rect 34600 89600 34800 89800
rect 51600 89600 51800 89800
rect 68800 89600 69000 89800
rect 24200 89800 24400 90000
rect 34600 89800 34800 90000
rect 51600 89800 51800 90000
rect 68800 89800 69000 90000
rect 24200 90000 24400 90200
rect 34600 90000 34800 90200
rect 51600 90000 51800 90200
rect 68800 90000 69000 90200
rect 24200 90200 24400 90400
rect 34600 90200 34800 90400
rect 51600 90200 51800 90400
rect 68800 90200 69000 90400
rect 24200 90400 24400 90600
rect 34600 90400 34800 90600
rect 51600 90400 51800 90600
rect 68800 90400 69000 90600
rect 24200 90600 24400 90800
rect 34600 90600 34800 90800
rect 51600 90600 51800 90800
rect 68800 90600 69000 90800
rect 24200 90800 24400 91000
rect 34600 90800 34800 91000
rect 51600 90800 51800 91000
rect 68800 90800 69000 91000
rect 24200 91000 24400 91200
rect 34600 91000 34800 91200
rect 51600 91000 51800 91200
rect 68800 91000 69000 91200
rect 24200 91200 24400 91400
rect 34600 91200 34800 91400
rect 51600 91200 51800 91400
rect 68800 91200 69000 91400
rect 24200 91400 24400 91600
rect 34600 91400 34800 91600
rect 51600 91400 51800 91600
rect 68800 91400 69000 91600
rect 24200 91600 24400 91800
rect 34600 91600 34800 91800
rect 51600 91600 51800 91800
rect 68800 91600 69000 91800
rect 24200 91800 24400 92000
rect 34600 91800 34800 92000
rect 51600 91800 51800 92000
rect 68800 91800 69000 92000
rect 24200 92000 24400 92200
rect 34600 92000 34800 92200
rect 51600 92000 51800 92200
rect 68800 92000 69000 92200
rect 24200 92200 24400 92400
rect 34600 92200 34800 92400
rect 51600 92200 51800 92400
rect 68800 92200 69000 92400
rect 24200 92400 24400 92600
rect 34600 92400 34800 92600
rect 51600 92400 51800 92600
rect 68800 92400 69000 92600
rect 24200 92600 24400 92800
rect 34600 92600 34800 92800
rect 51600 92600 51800 92800
rect 68800 92600 69000 92800
rect 24200 92800 24400 93000
rect 34600 92800 34800 93000
rect 51600 92800 51800 93000
rect 68800 92800 69000 93000
rect 24200 93000 24400 93200
rect 34600 93000 34800 93200
rect 51600 93000 51800 93200
rect 68800 93000 69000 93200
rect 24200 93200 24400 93400
rect 34600 93200 34800 93400
rect 51600 93200 51800 93400
rect 68800 93200 69000 93400
rect 24200 93400 24400 93600
rect 34600 93400 34800 93600
rect 51600 93400 51800 93600
rect 68800 93400 69000 93600
rect 24200 93600 24400 93800
rect 34600 93600 34800 93800
rect 51600 93600 51800 93800
rect 68800 93600 69000 93800
rect 24200 93800 24400 94000
rect 34600 93800 34800 94000
rect 51600 93800 51800 94000
rect 68800 93800 69000 94000
rect 24200 94000 24400 94200
rect 34600 94000 34800 94200
rect 51600 94000 51800 94200
rect 68800 94000 69000 94200
rect 24200 94200 24400 94400
rect 34600 94200 34800 94400
rect 51600 94200 51800 94400
rect 68800 94200 69000 94400
rect 24200 94400 24400 94600
rect 34600 94400 34800 94600
rect 51600 94400 51800 94600
rect 68800 94400 69000 94600
rect 24200 94600 24400 94800
rect 34600 94600 34800 94800
rect 51600 94600 51800 94800
rect 68800 94600 69000 94800
rect 24200 94800 24400 95000
rect 34600 94800 34800 95000
rect 51600 94800 51800 95000
rect 68800 94800 69000 95000
rect 24200 95000 24400 95200
rect 34600 95000 34800 95200
rect 51600 95000 51800 95200
rect 68800 95000 69000 95200
rect 24200 95200 24400 95400
rect 34600 95200 34800 95400
rect 51600 95200 51800 95400
rect 68800 95200 69000 95400
rect 24200 95400 24400 95600
rect 34600 95400 34800 95600
rect 51600 95400 51800 95600
rect 68800 95400 69000 95600
rect 24200 95600 24400 95800
rect 34600 95600 34800 95800
rect 51600 95600 51800 95800
rect 68800 95600 69000 95800
rect 24200 95800 24400 96000
rect 34600 95800 34800 96000
rect 51600 95800 51800 96000
rect 68800 95800 69000 96000
rect 24200 96000 24400 96200
rect 34600 96000 34800 96200
rect 51600 96000 51800 96200
rect 68800 96000 69000 96200
rect 24200 96200 24400 96400
rect 34600 96200 34800 96400
rect 51600 96200 51800 96400
rect 68800 96200 69000 96400
rect 34600 96400 34800 96600
rect 51600 96400 51800 96600
rect 68800 96400 69000 96600
rect 17400 96600 17600 96800
rect 41400 96600 41600 96800
rect 51600 96600 51800 96800
rect 68800 96600 69000 96800
rect 17400 96800 17600 97000
rect 41400 96800 41600 97000
rect 44800 96800 45000 97000
rect 75600 96800 75800 97000
rect 79000 96800 79200 97000
rect 20800 97000 21000 97200
rect 38000 97000 38200 97200
rect 55000 97000 55200 97200
rect 72200 97000 72400 97200
rect 24400 97200 24600 97400
rect 34400 97200 34600 97400
rect 51800 97200 52000 97400
rect 68600 97200 68800 97400
rect 20600 97400 20800 97600
rect 31400 97400 31600 97600
rect 38200 97400 38400 97600
rect 54800 97400 55000 97600
rect 65600 97400 65800 97600
rect 72400 97400 72600 97600
rect 20400 97600 20600 97800
rect 38400 97600 38600 97800
rect 45200 97600 45400 97800
rect 47800 97600 48000 97800
rect 72600 97600 72800 97800
rect 82000 97600 82200 97800
rect 20200 97800 20400 98000
rect 27000 97800 27200 98000
rect 31800 97800 32000 98000
rect 38600 97800 38800 98000
rect 54400 97800 54600 98000
rect 66000 97800 66200 98000
rect 72800 97800 73000 98000
rect 19800 98000 20000 98200
rect 39000 98000 39200 98200
rect 40400 98000 40600 98200
rect 45800 98000 46000 98200
rect 47200 98000 47400 98200
rect 54000 98000 54200 98200
rect 73200 98000 73400 98200
rect 74600 98000 74800 98200
rect 80000 98000 80200 98200
rect 81400 98000 81600 98200
rect -600 0 -500 100000
rect 100500 0 100600 100000
<< metal5 >>
rect 0 0 100000 200
rect 0 200 100000 400
rect 0 400 100000 600
rect 0 600 100000 800
rect 0 800 100000 1000
rect 0 1000 100000 1200
rect 0 1200 100000 1400
rect 0 1400 100000 1600
rect 0 1600 100000 1800
rect 0 1800 100000 2000
rect 0 2000 100000 2200
rect 0 2200 18800 2400
rect 19600 2200 25600 2400
rect 26600 2200 32400 2400
rect 33400 2200 39400 2400
rect 40200 2200 46200 2400
rect 47000 2200 53000 2400
rect 53800 2200 59800 2400
rect 60800 2200 66600 2400
rect 67600 2200 73600 2400
rect 74400 2200 80400 2400
rect 81200 2200 100000 2400
rect 0 2400 18400 2600
rect 20200 2400 25200 2600
rect 27000 2400 32000 2600
rect 33800 2400 38800 2600
rect 40600 2400 45800 2600
rect 47400 2400 52600 2600
rect 54400 2400 59400 2600
rect 61200 2400 66200 2600
rect 68000 2400 73000 2600
rect 74800 2400 80000 2600
rect 81600 2400 100000 2600
rect 0 2600 18000 2800
rect 20400 2600 25000 2800
rect 27200 2600 31800 2800
rect 34000 2600 38600 2800
rect 41000 2600 45400 2800
rect 47800 2600 52400 2800
rect 54600 2600 59200 2800
rect 61400 2600 66000 2800
rect 68200 2600 72800 2800
rect 75200 2600 79600 2800
rect 82000 2600 100000 2800
rect 0 2800 17800 3000
rect 20600 2800 24800 3000
rect 27400 2800 31600 3000
rect 34200 2800 38400 3000
rect 41200 2800 45200 3000
rect 48000 2800 52000 3000
rect 54800 2800 59000 3000
rect 61600 2800 65800 3000
rect 68400 2800 72600 3000
rect 75400 2800 79400 3000
rect 82200 2800 100000 3000
rect 0 3000 17800 3200
rect 20800 3000 24600 3200
rect 27600 3000 31400 3200
rect 34400 3000 38200 3200
rect 41200 3000 45200 3200
rect 48200 3000 52000 3200
rect 55000 3000 58800 3200
rect 61800 3000 65600 3200
rect 68600 3000 72400 3200
rect 75400 3000 79400 3200
rect 82400 3000 100000 3200
rect 0 3200 17600 3400
rect 20800 3200 24400 3400
rect 27800 3200 31400 3400
rect 34600 3200 38200 3400
rect 41400 3200 45000 3400
rect 48200 3200 51800 3400
rect 55000 3200 58600 3400
rect 62000 3200 65600 3400
rect 68800 3200 72400 3400
rect 75600 3200 79200 3400
rect 82400 3200 100000 3400
rect 0 3400 17600 3600
rect 21000 3400 24400 3600
rect 27800 3400 31200 3600
rect 34600 3400 38000 3600
rect 41400 3400 45000 3600
rect 48400 3400 51800 3600
rect 55200 3400 58600 3600
rect 62000 3400 65400 3600
rect 68800 3400 72200 3600
rect 75600 3400 79200 3600
rect 82600 3400 100000 3600
rect 0 3600 17400 3800
rect 21000 3600 24400 3800
rect 27800 3600 31200 3800
rect 34600 3600 38000 3800
rect 41600 3600 44800 3800
rect 48400 3600 51800 3800
rect 55200 3600 58600 3800
rect 62000 3600 65400 3800
rect 68800 3600 72200 3800
rect 75800 3600 79000 3800
rect 82600 3600 100000 3800
rect 0 3800 17400 4000
rect 21000 3800 24400 4000
rect 27800 3800 31200 4000
rect 34800 3800 38000 4000
rect 41600 3800 44800 4000
rect 48400 3800 51600 4000
rect 55200 3800 58600 4000
rect 62000 3800 65400 4000
rect 69000 3800 72200 4000
rect 75800 3800 79000 4000
rect 82600 3800 100000 4000
rect 0 4000 17400 4200
rect 21000 4000 24200 4200
rect 27800 4000 31200 4200
rect 34800 4000 38000 4200
rect 41600 4000 44800 4200
rect 48400 4000 51600 4200
rect 55200 4000 58600 4200
rect 62000 4000 65400 4200
rect 69000 4000 72200 4200
rect 75800 4000 79000 4200
rect 82600 4000 100000 4200
rect 0 4200 17400 4400
rect 21000 4200 24200 4400
rect 27800 4200 31200 4400
rect 34800 4200 38000 4400
rect 41600 4200 44800 4400
rect 48400 4200 51600 4400
rect 55200 4200 58600 4400
rect 62000 4200 65400 4400
rect 69000 4200 72200 4400
rect 75800 4200 79000 4400
rect 82600 4200 100000 4400
rect 0 4400 17400 4600
rect 21000 4400 24200 4600
rect 27800 4400 31200 4600
rect 34800 4400 38000 4600
rect 41600 4400 44800 4600
rect 48400 4400 51600 4600
rect 55200 4400 58600 4600
rect 62000 4400 65400 4600
rect 69000 4400 72200 4600
rect 75800 4400 79000 4600
rect 82600 4400 100000 4600
rect 0 4600 17400 4800
rect 21000 4600 24200 4800
rect 27800 4600 31200 4800
rect 34800 4600 38000 4800
rect 41600 4600 44800 4800
rect 48400 4600 51600 4800
rect 55200 4600 58600 4800
rect 62000 4600 65400 4800
rect 69000 4600 72200 4800
rect 75800 4600 79000 4800
rect 82600 4600 100000 4800
rect 0 4800 17400 5000
rect 21000 4800 24200 5000
rect 27800 4800 31200 5000
rect 34800 4800 38000 5000
rect 41600 4800 44800 5000
rect 48400 4800 51600 5000
rect 55200 4800 58600 5000
rect 62000 4800 65400 5000
rect 69000 4800 72200 5000
rect 75800 4800 79000 5000
rect 82600 4800 100000 5000
rect 0 5000 17400 5200
rect 21000 5000 24200 5200
rect 27800 5000 31200 5200
rect 34800 5000 38000 5200
rect 41600 5000 44800 5200
rect 48400 5000 51600 5200
rect 55200 5000 58600 5200
rect 62000 5000 65400 5200
rect 69000 5000 72200 5200
rect 75800 5000 79000 5200
rect 82600 5000 100000 5200
rect 0 5200 17400 5400
rect 21000 5200 24200 5400
rect 27800 5200 31200 5400
rect 34800 5200 38000 5400
rect 41600 5200 44800 5400
rect 48400 5200 51600 5400
rect 55200 5200 58600 5400
rect 62000 5200 65400 5400
rect 69000 5200 72200 5400
rect 75800 5200 79000 5400
rect 82600 5200 100000 5400
rect 0 5400 17400 5600
rect 21000 5400 24200 5600
rect 27800 5400 31200 5600
rect 34800 5400 38000 5600
rect 41600 5400 44800 5600
rect 48400 5400 51600 5600
rect 55200 5400 58600 5600
rect 62000 5400 65400 5600
rect 69000 5400 72200 5600
rect 75800 5400 79000 5600
rect 82600 5400 100000 5600
rect 0 5600 17400 5800
rect 21000 5600 24200 5800
rect 27800 5600 31200 5800
rect 34800 5600 38000 5800
rect 41600 5600 44800 5800
rect 48400 5600 51600 5800
rect 55200 5600 58600 5800
rect 62000 5600 65400 5800
rect 69000 5600 72200 5800
rect 75800 5600 79000 5800
rect 82600 5600 100000 5800
rect 0 5800 17400 6000
rect 21000 5800 24200 6000
rect 27800 5800 31200 6000
rect 34800 5800 38000 6000
rect 41600 5800 44800 6000
rect 48400 5800 51600 6000
rect 55200 5800 58600 6000
rect 62000 5800 65400 6000
rect 69000 5800 72200 6000
rect 75800 5800 79000 6000
rect 82600 5800 100000 6000
rect 0 6000 17400 6200
rect 21000 6000 24200 6200
rect 27800 6000 31200 6200
rect 34800 6000 38000 6200
rect 41600 6000 44800 6200
rect 48400 6000 51600 6200
rect 55200 6000 58600 6200
rect 62000 6000 65400 6200
rect 69000 6000 72200 6200
rect 75800 6000 79000 6200
rect 82600 6000 100000 6200
rect 0 6200 17400 6400
rect 21000 6200 24200 6400
rect 27800 6200 31200 6400
rect 34800 6200 38000 6400
rect 41600 6200 44800 6400
rect 48400 6200 51600 6400
rect 55200 6200 58600 6400
rect 62000 6200 65400 6400
rect 69000 6200 72200 6400
rect 75800 6200 79000 6400
rect 82600 6200 100000 6400
rect 0 6400 17400 6600
rect 21000 6400 24200 6600
rect 27800 6400 31200 6600
rect 34800 6400 38000 6600
rect 41600 6400 44800 6600
rect 48400 6400 51600 6600
rect 55200 6400 58600 6600
rect 62000 6400 65400 6600
rect 69000 6400 72200 6600
rect 75800 6400 79000 6600
rect 82600 6400 100000 6600
rect 0 6600 17400 6800
rect 21000 6600 24200 6800
rect 27800 6600 31200 6800
rect 34800 6600 38000 6800
rect 41600 6600 44800 6800
rect 48400 6600 51600 6800
rect 55200 6600 58600 6800
rect 62000 6600 65400 6800
rect 69000 6600 72200 6800
rect 75800 6600 79000 6800
rect 82600 6600 100000 6800
rect 0 6800 17400 7000
rect 21000 6800 24200 7000
rect 27800 6800 31200 7000
rect 34800 6800 38000 7000
rect 41600 6800 44800 7000
rect 48400 6800 51600 7000
rect 55200 6800 58600 7000
rect 62000 6800 65400 7000
rect 69000 6800 72200 7000
rect 75800 6800 79000 7000
rect 82600 6800 100000 7000
rect 0 7000 17400 7200
rect 21000 7000 24200 7200
rect 27800 7000 31200 7200
rect 34800 7000 38000 7200
rect 41600 7000 44800 7200
rect 48400 7000 51600 7200
rect 55200 7000 58600 7200
rect 62000 7000 65400 7200
rect 69000 7000 72200 7200
rect 75800 7000 79000 7200
rect 82600 7000 100000 7200
rect 0 7200 17400 7400
rect 21000 7200 24200 7400
rect 27800 7200 31200 7400
rect 34800 7200 38000 7400
rect 41600 7200 44800 7400
rect 48400 7200 51600 7400
rect 55200 7200 58600 7400
rect 62000 7200 65400 7400
rect 69000 7200 72200 7400
rect 75800 7200 79000 7400
rect 82600 7200 100000 7400
rect 0 7400 17400 7600
rect 21000 7400 24200 7600
rect 27800 7400 31200 7600
rect 34800 7400 38000 7600
rect 41600 7400 44800 7600
rect 48400 7400 51600 7600
rect 55200 7400 58600 7600
rect 62000 7400 65400 7600
rect 69000 7400 72200 7600
rect 75800 7400 79000 7600
rect 82600 7400 100000 7600
rect 0 7600 17400 7800
rect 21000 7600 24200 7800
rect 27800 7600 31200 7800
rect 34800 7600 38000 7800
rect 41600 7600 44800 7800
rect 48400 7600 51600 7800
rect 55200 7600 58600 7800
rect 62000 7600 65400 7800
rect 69000 7600 72200 7800
rect 75800 7600 79000 7800
rect 82600 7600 100000 7800
rect 0 7800 17400 8000
rect 21000 7800 24200 8000
rect 27800 7800 31200 8000
rect 34800 7800 38000 8000
rect 41600 7800 44800 8000
rect 48400 7800 51600 8000
rect 55200 7800 58600 8000
rect 62000 7800 65400 8000
rect 69000 7800 72200 8000
rect 75800 7800 79000 8000
rect 82600 7800 100000 8000
rect 0 8000 17400 8200
rect 21000 8000 24200 8200
rect 27800 8000 31200 8200
rect 34800 8000 38000 8200
rect 41600 8000 44800 8200
rect 48400 8000 51600 8200
rect 55200 8000 58600 8200
rect 62000 8000 65400 8200
rect 69000 8000 72200 8200
rect 75800 8000 79000 8200
rect 82600 8000 100000 8200
rect 0 8200 17400 8400
rect 21000 8200 24200 8400
rect 27800 8200 31200 8400
rect 34800 8200 38000 8400
rect 41600 8200 44800 8400
rect 48400 8200 51600 8400
rect 55200 8200 58600 8400
rect 62000 8200 65400 8400
rect 69000 8200 72200 8400
rect 75800 8200 79000 8400
rect 82600 8200 100000 8400
rect 0 8400 17400 8600
rect 21000 8400 24200 8600
rect 27800 8400 31200 8600
rect 34800 8400 38000 8600
rect 41600 8400 44800 8600
rect 48400 8400 51600 8600
rect 55200 8400 58600 8600
rect 62000 8400 65400 8600
rect 69000 8400 72200 8600
rect 75800 8400 79000 8600
rect 82600 8400 100000 8600
rect 0 8600 17400 8800
rect 21000 8600 24200 8800
rect 27800 8600 31200 8800
rect 34800 8600 38000 8800
rect 41600 8600 44800 8800
rect 48400 8600 51600 8800
rect 55200 8600 58600 8800
rect 62000 8600 65400 8800
rect 69000 8600 72200 8800
rect 75800 8600 79000 8800
rect 82600 8600 100000 8800
rect 0 8800 17400 9000
rect 21000 8800 24200 9000
rect 27800 8800 31200 9000
rect 34800 8800 38000 9000
rect 41600 8800 44800 9000
rect 48400 8800 51600 9000
rect 55200 8800 58600 9000
rect 62000 8800 65400 9000
rect 69000 8800 72200 9000
rect 75800 8800 79000 9000
rect 82600 8800 100000 9000
rect 0 9000 17400 9200
rect 21000 9000 24200 9200
rect 27800 9000 31200 9200
rect 34800 9000 38000 9200
rect 41600 9000 44800 9200
rect 48400 9000 51600 9200
rect 55200 9000 58600 9200
rect 62000 9000 65400 9200
rect 69000 9000 72200 9200
rect 75800 9000 79000 9200
rect 82600 9000 100000 9200
rect 0 9200 17400 9400
rect 21000 9200 24200 9400
rect 27800 9200 31200 9400
rect 34800 9200 38000 9400
rect 41600 9200 44800 9400
rect 48400 9200 51600 9400
rect 55200 9200 58600 9400
rect 62000 9200 65400 9400
rect 69000 9200 72200 9400
rect 75800 9200 79000 9400
rect 82600 9200 100000 9400
rect 0 9400 17400 9600
rect 21000 9400 24200 9600
rect 27800 9400 31200 9600
rect 34800 9400 38000 9600
rect 41600 9400 44800 9600
rect 48400 9400 51600 9600
rect 55200 9400 58600 9600
rect 62000 9400 65400 9600
rect 69000 9400 72200 9600
rect 75800 9400 79000 9600
rect 82600 9400 100000 9600
rect 0 9600 17400 9800
rect 21000 9600 24200 9800
rect 27800 9600 31200 9800
rect 34800 9600 38000 9800
rect 41600 9600 44800 9800
rect 48400 9600 51600 9800
rect 55200 9600 58600 9800
rect 62000 9600 65400 9800
rect 69000 9600 72200 9800
rect 75800 9600 79000 9800
rect 82600 9600 100000 9800
rect 0 9800 17400 10000
rect 21000 9800 24200 10000
rect 27800 9800 31200 10000
rect 34800 9800 38000 10000
rect 41600 9800 44800 10000
rect 48400 9800 51600 10000
rect 55200 9800 58600 10000
rect 62000 9800 65400 10000
rect 69000 9800 72200 10000
rect 75800 9800 79000 10000
rect 82600 9800 100000 10000
rect 0 10000 17400 10200
rect 21000 10000 24200 10200
rect 27800 10000 31200 10200
rect 34800 10000 38000 10200
rect 41600 10000 44800 10200
rect 48400 10000 51600 10200
rect 55200 10000 58600 10200
rect 62000 10000 65400 10200
rect 69000 10000 72200 10200
rect 75800 10000 79000 10200
rect 82600 10000 100000 10200
rect 0 10200 17400 10400
rect 21000 10200 24200 10400
rect 27800 10200 31200 10400
rect 34800 10200 38000 10400
rect 41600 10200 44800 10400
rect 48400 10200 51600 10400
rect 55200 10200 58600 10400
rect 62000 10200 65400 10400
rect 69000 10200 72200 10400
rect 75800 10200 79000 10400
rect 82600 10200 100000 10400
rect 0 10400 17400 10600
rect 21000 10400 24200 10600
rect 27800 10400 31200 10600
rect 34800 10400 38000 10600
rect 41600 10400 44800 10600
rect 48400 10400 51600 10600
rect 55200 10400 58600 10600
rect 62000 10400 65400 10600
rect 69000 10400 72200 10600
rect 75800 10400 79000 10600
rect 82600 10400 100000 10600
rect 0 10600 17400 10800
rect 21000 10600 24200 10800
rect 27800 10600 31200 10800
rect 34800 10600 38000 10800
rect 41600 10600 44800 10800
rect 48400 10600 51600 10800
rect 55200 10600 58600 10800
rect 62000 10600 65400 10800
rect 69000 10600 72200 10800
rect 75800 10600 79000 10800
rect 82600 10600 100000 10800
rect 0 10800 17400 11000
rect 21000 10800 24200 11000
rect 27800 10800 31200 11000
rect 34800 10800 38000 11000
rect 41600 10800 44800 11000
rect 48400 10800 51600 11000
rect 55200 10800 58600 11000
rect 62000 10800 65400 11000
rect 69000 10800 72200 11000
rect 75800 10800 79000 11000
rect 82600 10800 100000 11000
rect 0 11000 17400 11200
rect 21000 11000 24200 11200
rect 27800 11000 31200 11200
rect 34800 11000 38000 11200
rect 41600 11000 44800 11200
rect 48400 11000 51600 11200
rect 55200 11000 58600 11200
rect 62000 11000 65400 11200
rect 69000 11000 72200 11200
rect 75800 11000 79000 11200
rect 82600 11000 100000 11200
rect 0 11200 17400 11400
rect 21000 11200 24200 11400
rect 27800 11200 31200 11400
rect 34800 11200 38000 11400
rect 41600 11200 44800 11400
rect 48400 11200 51600 11400
rect 55200 11200 58600 11400
rect 62000 11200 65400 11400
rect 69000 11200 72200 11400
rect 75800 11200 79000 11400
rect 82600 11200 100000 11400
rect 0 11400 17400 11600
rect 21000 11400 24200 11600
rect 27800 11400 31200 11600
rect 34800 11400 38000 11600
rect 41600 11400 44800 11600
rect 48400 11400 51600 11600
rect 55200 11400 58600 11600
rect 62000 11400 65400 11600
rect 69000 11400 72200 11600
rect 75800 11400 79000 11600
rect 82600 11400 100000 11600
rect 0 11600 17400 11800
rect 21000 11600 24200 11800
rect 27800 11600 31200 11800
rect 34800 11600 38000 11800
rect 41600 11600 44800 11800
rect 48400 11600 51600 11800
rect 55200 11600 58600 11800
rect 62000 11600 65400 11800
rect 69000 11600 72200 11800
rect 75800 11600 79000 11800
rect 82600 11600 100000 11800
rect 0 11800 17400 12000
rect 21000 11800 24200 12000
rect 27800 11800 31200 12000
rect 34800 11800 38000 12000
rect 41600 11800 44800 12000
rect 48400 11800 51600 12000
rect 55200 11800 58600 12000
rect 62000 11800 65400 12000
rect 69000 11800 72200 12000
rect 75800 11800 79000 12000
rect 82600 11800 100000 12000
rect 0 12000 17400 12200
rect 21000 12000 24200 12200
rect 27800 12000 31200 12200
rect 34800 12000 38000 12200
rect 41600 12000 44800 12200
rect 48400 12000 51600 12200
rect 55200 12000 58600 12200
rect 62000 12000 65400 12200
rect 69000 12000 72200 12200
rect 75800 12000 79000 12200
rect 82600 12000 100000 12200
rect 0 12200 17400 12400
rect 21000 12200 24200 12400
rect 27800 12200 31200 12400
rect 34800 12200 38000 12400
rect 41600 12200 44800 12400
rect 48400 12200 51600 12400
rect 55200 12200 58600 12400
rect 62000 12200 65400 12400
rect 69000 12200 72200 12400
rect 75800 12200 79000 12400
rect 82600 12200 100000 12400
rect 0 12400 17400 12600
rect 21000 12400 24200 12600
rect 27800 12400 31200 12600
rect 34800 12400 38000 12600
rect 41600 12400 44800 12600
rect 48400 12400 51600 12600
rect 55200 12400 58600 12600
rect 62000 12400 65400 12600
rect 69000 12400 72200 12600
rect 75800 12400 79000 12600
rect 82600 12400 100000 12600
rect 0 12600 17400 12800
rect 21000 12600 24200 12800
rect 27800 12600 31200 12800
rect 34800 12600 38000 12800
rect 41600 12600 44800 12800
rect 48400 12600 51600 12800
rect 55200 12600 58600 12800
rect 62000 12600 65400 12800
rect 69000 12600 72200 12800
rect 75800 12600 79000 12800
rect 82600 12600 100000 12800
rect 0 12800 17400 13000
rect 21000 12800 24200 13000
rect 27800 12800 31200 13000
rect 34800 12800 38000 13000
rect 41600 12800 44800 13000
rect 48400 12800 51600 13000
rect 55200 12800 58600 13000
rect 62000 12800 65400 13000
rect 69000 12800 72200 13000
rect 75800 12800 79000 13000
rect 82600 12800 100000 13000
rect 0 13000 17400 13200
rect 21000 13000 24200 13200
rect 27800 13000 31200 13200
rect 34800 13000 38000 13200
rect 41600 13000 44800 13200
rect 48400 13000 51600 13200
rect 55200 13000 58600 13200
rect 62000 13000 65400 13200
rect 69000 13000 72200 13200
rect 75800 13000 79000 13200
rect 82600 13000 100000 13200
rect 0 13200 17400 13400
rect 21000 13200 24200 13400
rect 27800 13200 31200 13400
rect 34800 13200 38000 13400
rect 41600 13200 44800 13400
rect 48400 13200 51600 13400
rect 55200 13200 58600 13400
rect 62000 13200 65400 13400
rect 69000 13200 72200 13400
rect 75800 13200 79000 13400
rect 82600 13200 100000 13400
rect 0 13400 17400 13600
rect 21000 13400 24200 13600
rect 27800 13400 31200 13600
rect 34800 13400 38000 13600
rect 41600 13400 44800 13600
rect 48400 13400 51600 13600
rect 55200 13400 58600 13600
rect 62000 13400 65400 13600
rect 69000 13400 72200 13600
rect 75800 13400 79000 13600
rect 82600 13400 100000 13600
rect 0 13600 17400 13800
rect 21000 13600 24200 13800
rect 27800 13600 31200 13800
rect 34800 13600 38000 13800
rect 41600 13600 44800 13800
rect 48400 13600 51600 13800
rect 55200 13600 58600 13800
rect 62000 13600 65400 13800
rect 69000 13600 72200 13800
rect 75800 13600 79000 13800
rect 82600 13600 100000 13800
rect 0 13800 17400 14000
rect 21000 13800 24200 14000
rect 27800 13800 31200 14000
rect 34800 13800 38000 14000
rect 41600 13800 44800 14000
rect 48400 13800 51600 14000
rect 55200 13800 58600 14000
rect 62000 13800 65400 14000
rect 69000 13800 72200 14000
rect 75800 13800 79000 14000
rect 82600 13800 100000 14000
rect 0 14000 17400 14200
rect 21000 14000 24200 14200
rect 27800 14000 31200 14200
rect 34800 14000 38000 14200
rect 41600 14000 44800 14200
rect 48400 14000 51600 14200
rect 55200 14000 58600 14200
rect 62000 14000 65400 14200
rect 69000 14000 72200 14200
rect 75800 14000 79000 14200
rect 82600 14000 100000 14200
rect 0 14200 15400 14400
rect 84600 14200 100000 14400
rect 0 14400 15000 14600
rect 85200 14400 100000 14600
rect 0 14600 14600 14800
rect 85400 14600 100000 14800
rect 0 14800 14400 15000
rect 85600 14800 100000 15000
rect 0 15000 14400 15200
rect 85800 15000 100000 15200
rect 0 15200 14200 15400
rect 85800 15200 100000 15400
rect 0 15400 14200 15600
rect 86000 15400 100000 15600
rect 0 15600 14000 15800
rect 86000 15600 100000 15800
rect 0 15800 14000 16000
rect 86000 15800 100000 16000
rect 0 16000 14000 16200
rect 86000 16000 100000 16200
rect 0 16200 14000 16400
rect 86000 16200 100000 16400
rect 0 16400 14000 16600
rect 86000 16400 100000 16600
rect 0 16600 14000 16800
rect 86000 16600 100000 16800
rect 0 16800 14000 17000
rect 86000 16800 100000 17000
rect 0 17000 14000 17200
rect 86000 17000 100000 17200
rect 0 17200 14000 17400
rect 86000 17200 100000 17400
rect 0 17400 14000 17600
rect 86000 17400 100000 17600
rect 0 17600 3400 17800
rect 96600 17600 100000 17800
rect 0 17800 3000 18000
rect 97000 17800 100000 18000
rect 0 18000 2600 18200
rect 97400 18000 100000 18200
rect 0 18200 2400 18400
rect 97600 18200 100000 18400
rect 0 18400 2400 18600
rect 97800 18400 100000 18600
rect 0 18600 2200 18800
rect 97800 18600 100000 18800
rect 0 18800 2200 19000
rect 97800 18800 100000 19000
rect 0 19000 2200 19200
rect 98000 19000 100000 19200
rect 0 19200 2000 19400
rect 18800 19200 43000 19400
rect 51600 19200 81200 19400
rect 98000 19200 100000 19400
rect 0 19400 2000 19600
rect 18800 19400 44200 19600
rect 51600 19400 81200 19600
rect 98000 19400 100000 19600
rect 0 19600 2000 19800
rect 18800 19600 44800 19800
rect 51600 19600 81200 19800
rect 98000 19600 100000 19800
rect 0 19800 2200 20000
rect 18800 19800 45200 20000
rect 51600 19800 81200 20000
rect 98000 19800 100000 20000
rect 0 20000 2200 20200
rect 18800 20000 45600 20200
rect 51600 20000 81200 20200
rect 97800 20000 100000 20200
rect 0 20200 2200 20400
rect 18800 20200 45800 20400
rect 51600 20200 81200 20400
rect 97800 20200 100000 20400
rect 0 20400 2400 20600
rect 18800 20400 46200 20600
rect 51600 20400 81200 20600
rect 97600 20400 100000 20600
rect 0 20600 2600 20800
rect 18800 20600 46400 20800
rect 51600 20600 81200 20800
rect 97400 20600 100000 20800
rect 0 20800 2800 21000
rect 18800 20800 46600 21000
rect 51600 20800 81200 21000
rect 97200 20800 100000 21000
rect 0 21000 3200 21200
rect 18800 21000 46800 21200
rect 51600 21000 81200 21200
rect 96800 21000 100000 21200
rect 0 21200 14000 21400
rect 18800 21200 47000 21400
rect 51600 21200 81200 21400
rect 86000 21200 100000 21400
rect 0 21400 14000 21600
rect 18800 21400 47200 21600
rect 51600 21400 81200 21600
rect 86000 21400 100000 21600
rect 0 21600 14000 21800
rect 18800 21600 47400 21800
rect 51600 21600 81200 21800
rect 86000 21600 100000 21800
rect 0 21800 14000 22000
rect 18800 21800 47400 22000
rect 51600 21800 81200 22000
rect 86000 21800 100000 22000
rect 0 22000 14000 22200
rect 18800 22000 47600 22200
rect 51600 22000 81200 22200
rect 86000 22000 100000 22200
rect 0 22200 14000 22400
rect 18800 22200 47600 22400
rect 51600 22200 81200 22400
rect 86000 22200 100000 22400
rect 0 22400 14000 22600
rect 18800 22400 47800 22600
rect 51600 22400 81200 22600
rect 86000 22400 100000 22600
rect 0 22600 14000 22800
rect 18800 22600 48000 22800
rect 51600 22600 81200 22800
rect 86000 22600 100000 22800
rect 0 22800 14000 23000
rect 18800 22800 48000 23000
rect 51600 22800 81200 23000
rect 86000 22800 100000 23000
rect 0 23000 14000 23200
rect 18800 23000 48000 23200
rect 51600 23000 81200 23200
rect 86000 23000 100000 23200
rect 0 23200 14000 23400
rect 18800 23200 48200 23400
rect 51600 23200 81200 23400
rect 86000 23200 100000 23400
rect 0 23400 14000 23600
rect 18800 23400 48200 23600
rect 51600 23400 81200 23600
rect 86000 23400 100000 23600
rect 0 23600 14000 23800
rect 18800 23600 48200 23800
rect 51600 23600 81200 23800
rect 86000 23600 100000 23800
rect 0 23800 14000 24000
rect 18800 23800 48400 24000
rect 51600 23800 81200 24000
rect 86000 23800 100000 24000
rect 0 24000 14000 24200
rect 18800 24000 48400 24200
rect 51600 24000 81200 24200
rect 86000 24000 100000 24200
rect 0 24200 14000 24400
rect 18800 24200 48400 24400
rect 51600 24200 81200 24400
rect 86000 24200 100000 24400
rect 0 24400 14000 24600
rect 18800 24400 48400 24600
rect 51600 24400 81200 24600
rect 86000 24400 100000 24600
rect 0 24600 3000 24800
rect 18800 24600 48400 24800
rect 51600 24600 81200 24800
rect 97000 24600 100000 24800
rect 0 24800 2800 25000
rect 18800 24800 48400 25000
rect 51600 24800 81200 25000
rect 97200 24800 100000 25000
rect 0 25000 2600 25200
rect 42600 25000 48400 25200
rect 51600 25000 57400 25200
rect 97600 25000 100000 25200
rect 0 25200 2400 25400
rect 42600 25200 48400 25400
rect 51600 25200 57400 25400
rect 97600 25200 100000 25400
rect 0 25400 2200 25600
rect 42600 25400 48400 25600
rect 51600 25400 57400 25600
rect 97800 25400 100000 25600
rect 0 25600 2200 25800
rect 42600 25600 48400 25800
rect 51600 25600 57400 25800
rect 97800 25600 100000 25800
rect 0 25800 2200 26000
rect 42600 25800 48400 26000
rect 51600 25800 57400 26000
rect 98000 25800 100000 26000
rect 0 26000 2000 26200
rect 42600 26000 48400 26200
rect 51600 26000 57400 26200
rect 98000 26000 100000 26200
rect 0 26200 2000 26400
rect 42600 26200 48400 26400
rect 51600 26200 57400 26400
rect 98000 26200 100000 26400
rect 0 26400 2000 26600
rect 42600 26400 48400 26600
rect 51600 26400 57400 26600
rect 98000 26400 100000 26600
rect 0 26600 2200 26800
rect 42600 26600 48400 26800
rect 51600 26600 57400 26800
rect 98000 26600 100000 26800
rect 0 26800 2200 27000
rect 42600 26800 48400 27000
rect 51600 26800 57400 27000
rect 97800 26800 100000 27000
rect 0 27000 2200 27200
rect 42600 27000 48400 27200
rect 51600 27000 57400 27200
rect 97800 27000 100000 27200
rect 0 27200 2400 27400
rect 42600 27200 48400 27400
rect 51600 27200 57400 27400
rect 97600 27200 100000 27400
rect 0 27400 2600 27600
rect 42600 27400 48400 27600
rect 51600 27400 57400 27600
rect 97600 27400 100000 27600
rect 0 27600 2800 27800
rect 42600 27600 48400 27800
rect 51600 27600 57400 27800
rect 97200 27600 100000 27800
rect 0 27800 3200 28000
rect 42600 27800 48400 28000
rect 51600 27800 57400 28000
rect 97000 27800 100000 28000
rect 0 28000 14000 28200
rect 42600 28000 48400 28200
rect 51600 28000 57400 28200
rect 86000 28000 100000 28200
rect 0 28200 14000 28400
rect 42600 28200 48400 28400
rect 51600 28200 57400 28400
rect 86000 28200 100000 28400
rect 0 28400 14000 28600
rect 42600 28400 48400 28600
rect 51600 28400 57400 28600
rect 86000 28400 100000 28600
rect 0 28600 14000 28800
rect 42600 28600 48400 28800
rect 51600 28600 57400 28800
rect 86000 28600 100000 28800
rect 0 28800 14000 29000
rect 42600 28800 48400 29000
rect 51600 28800 57400 29000
rect 86000 28800 100000 29000
rect 0 29000 14000 29200
rect 42600 29000 48400 29200
rect 51600 29000 57400 29200
rect 86000 29000 100000 29200
rect 0 29200 14000 29400
rect 42600 29200 48400 29400
rect 51600 29200 57400 29400
rect 86000 29200 100000 29400
rect 0 29400 14000 29600
rect 42600 29400 48400 29600
rect 51600 29400 57400 29600
rect 86000 29400 100000 29600
rect 0 29600 14000 29800
rect 42600 29600 48400 29800
rect 51600 29600 57400 29800
rect 86000 29600 100000 29800
rect 0 29800 14000 30000
rect 42600 29800 48400 30000
rect 51600 29800 57400 30000
rect 86000 29800 100000 30000
rect 0 30000 14000 30200
rect 42600 30000 48400 30200
rect 51600 30000 57400 30200
rect 86000 30000 100000 30200
rect 0 30200 14000 30400
rect 42600 30200 48400 30400
rect 51600 30200 57400 30400
rect 86000 30200 100000 30400
rect 0 30400 14000 30600
rect 42600 30400 48400 30600
rect 51600 30400 57400 30600
rect 86000 30400 100000 30600
rect 0 30600 14000 30800
rect 42600 30600 48400 30800
rect 51600 30600 57400 30800
rect 86000 30600 100000 30800
rect 0 30800 14000 31000
rect 42600 30800 48400 31000
rect 51600 30800 57400 31000
rect 86000 30800 100000 31000
rect 0 31000 14000 31200
rect 42600 31000 48400 31200
rect 51600 31000 57400 31200
rect 86000 31000 100000 31200
rect 0 31200 14000 31400
rect 23600 31200 48400 31400
rect 51600 31200 76400 31400
rect 86000 31200 100000 31400
rect 0 31400 3200 31600
rect 22800 31400 48400 31600
rect 51600 31400 77200 31600
rect 97000 31400 100000 31600
rect 0 31600 2800 31800
rect 22400 31600 48400 31800
rect 51600 31600 77600 31800
rect 97200 31600 100000 31800
rect 0 31800 2600 32000
rect 22000 31800 48400 32000
rect 51600 31800 78000 32000
rect 97400 31800 100000 32000
rect 0 32000 2400 32200
rect 21600 32000 48400 32200
rect 51600 32000 78400 32200
rect 97600 32000 100000 32200
rect 0 32200 2200 32400
rect 21400 32200 48400 32400
rect 51600 32200 78800 32400
rect 97800 32200 100000 32400
rect 0 32400 2200 32600
rect 21000 32400 48200 32600
rect 51800 32400 79000 32600
rect 97800 32400 100000 32600
rect 0 32600 2200 32800
rect 20800 32600 48200 32800
rect 51800 32600 79200 32800
rect 98000 32600 100000 32800
rect 0 32800 2000 33000
rect 20600 32800 48200 33000
rect 51800 32800 79400 33000
rect 98000 32800 100000 33000
rect 0 33000 2000 33200
rect 20400 33000 48200 33200
rect 52000 33000 79600 33200
rect 98000 33000 100000 33200
rect 0 33200 2000 33400
rect 20200 33200 48000 33400
rect 52000 33200 79800 33400
rect 98000 33200 100000 33400
rect 0 33400 2000 33600
rect 20000 33400 48000 33600
rect 52000 33400 80000 33600
rect 98000 33400 100000 33600
rect 0 33600 2200 33800
rect 20000 33600 47800 33800
rect 52200 33600 80200 33800
rect 97800 33600 100000 33800
rect 0 33800 2200 34000
rect 19800 33800 47800 34000
rect 52400 33800 80200 34000
rect 97800 33800 100000 34000
rect 0 34000 2400 34200
rect 19600 34000 47600 34200
rect 52400 34000 80400 34200
rect 97800 34000 100000 34200
rect 0 34200 2400 34400
rect 19600 34200 47600 34400
rect 52600 34200 80400 34400
rect 97600 34200 100000 34400
rect 0 34400 2800 34600
rect 19400 34400 47400 34600
rect 52600 34400 80600 34600
rect 97400 34400 100000 34600
rect 0 34600 3000 34800
rect 19400 34600 47200 34800
rect 52800 34600 80600 34800
rect 97000 34600 100000 34800
rect 0 34800 3600 35000
rect 19200 34800 47000 35000
rect 53000 34800 80800 35000
rect 96400 34800 100000 35000
rect 0 35000 14000 35200
rect 19200 35000 46800 35200
rect 53200 35000 80800 35200
rect 86000 35000 100000 35200
rect 0 35200 14000 35400
rect 19200 35200 46800 35400
rect 53400 35200 81000 35400
rect 86000 35200 100000 35400
rect 0 35400 14000 35600
rect 19000 35400 46400 35600
rect 53600 35400 81000 35600
rect 86000 35400 100000 35600
rect 0 35600 14000 35800
rect 19000 35600 46200 35800
rect 53800 35600 81000 35800
rect 86000 35600 100000 35800
rect 0 35800 14000 36000
rect 19000 35800 46000 36000
rect 54000 35800 81000 36000
rect 86000 35800 100000 36000
rect 0 36000 14000 36200
rect 19000 36000 45600 36200
rect 54400 36000 81200 36200
rect 86000 36000 100000 36200
rect 0 36200 14000 36400
rect 18800 36200 45400 36400
rect 54800 36200 81200 36400
rect 86000 36200 100000 36400
rect 0 36400 14000 36600
rect 18800 36400 45000 36600
rect 55000 36400 81200 36600
rect 86000 36400 100000 36600
rect 0 36600 14000 36800
rect 18800 36600 44400 36800
rect 55600 36600 81200 36800
rect 86000 36600 100000 36800
rect 0 36800 14000 37000
rect 18800 36800 43600 37000
rect 56400 36800 81200 37000
rect 86000 36800 100000 37000
rect 0 37000 14000 37200
rect 18800 37000 24600 37200
rect 75400 37000 81200 37200
rect 86000 37000 100000 37200
rect 0 37200 14000 37400
rect 18800 37200 24600 37400
rect 75400 37200 81200 37400
rect 86000 37200 100000 37400
rect 0 37400 14000 37600
rect 18800 37400 24600 37600
rect 75400 37400 81200 37600
rect 86000 37400 100000 37600
rect 0 37600 14000 37800
rect 18800 37600 24600 37800
rect 75400 37600 81200 37800
rect 86000 37600 100000 37800
rect 0 37800 14000 38000
rect 18800 37800 24600 38000
rect 75400 37800 81200 38000
rect 86000 37800 100000 38000
rect 0 38000 14000 38200
rect 18800 38000 24600 38200
rect 75400 38000 81200 38200
rect 86000 38000 100000 38200
rect 0 38200 3200 38400
rect 18800 38200 24600 38400
rect 75400 38200 81200 38400
rect 96800 38200 100000 38400
rect 0 38400 2800 38600
rect 18800 38400 24600 38600
rect 75400 38400 81200 38600
rect 97200 38400 100000 38600
rect 0 38600 2600 38800
rect 18800 38600 24600 38800
rect 75400 38600 81200 38800
rect 97400 38600 100000 38800
rect 0 38800 2400 39000
rect 18800 38800 24600 39000
rect 75400 38800 81200 39000
rect 97600 38800 100000 39000
rect 0 39000 2400 39200
rect 18800 39000 24600 39200
rect 75400 39000 81200 39200
rect 97800 39000 100000 39200
rect 0 39200 2200 39400
rect 18800 39200 24600 39400
rect 75400 39200 81200 39400
rect 97800 39200 100000 39400
rect 0 39400 2200 39600
rect 18800 39400 24600 39600
rect 75400 39400 81200 39600
rect 98000 39400 100000 39600
rect 0 39600 2000 39800
rect 18800 39600 24600 39800
rect 75400 39600 81200 39800
rect 98000 39600 100000 39800
rect 0 39800 2000 40000
rect 18800 39800 24600 40000
rect 75400 39800 81200 40000
rect 98000 39800 100000 40000
rect 0 40000 2000 40200
rect 18800 40000 24600 40200
rect 75400 40000 81200 40200
rect 98000 40000 100000 40200
rect 0 40200 2000 40400
rect 18800 40200 24600 40400
rect 75400 40200 81200 40400
rect 98000 40200 100000 40400
rect 0 40400 2200 40600
rect 18800 40400 24600 40600
rect 75400 40400 81200 40600
rect 97800 40400 100000 40600
rect 0 40600 2200 40800
rect 18800 40600 24600 40800
rect 75400 40600 81200 40800
rect 97800 40600 100000 40800
rect 0 40800 2400 41000
rect 18800 40800 24600 41000
rect 75400 40800 81200 41000
rect 97800 40800 100000 41000
rect 0 41000 2400 41200
rect 18800 41000 24600 41200
rect 75400 41000 81200 41200
rect 97600 41000 100000 41200
rect 0 41200 2600 41400
rect 18800 41200 24600 41400
rect 75400 41200 81200 41400
rect 97400 41200 100000 41400
rect 0 41400 3000 41600
rect 18800 41400 24600 41600
rect 75400 41400 81200 41600
rect 97200 41400 100000 41600
rect 0 41600 3400 41800
rect 18800 41600 24600 41800
rect 75400 41600 81200 41800
rect 96600 41600 100000 41800
rect 0 41800 14000 42000
rect 18800 41800 24600 42000
rect 75400 41800 81200 42000
rect 86000 41800 100000 42000
rect 0 42000 14000 42200
rect 18800 42000 24600 42200
rect 75400 42000 81200 42200
rect 86000 42000 100000 42200
rect 0 42200 14000 42400
rect 18800 42200 24600 42400
rect 75400 42200 81200 42400
rect 86000 42200 100000 42400
rect 0 42400 14000 42600
rect 18800 42400 24600 42600
rect 75400 42400 81200 42600
rect 86000 42400 100000 42600
rect 0 42600 14000 42800
rect 18800 42600 24600 42800
rect 75400 42600 81200 42800
rect 86000 42600 100000 42800
rect 0 42800 14000 43000
rect 18800 42800 24600 43000
rect 75400 42800 81200 43000
rect 86000 42800 100000 43000
rect 0 43000 14000 43200
rect 18800 43000 24600 43200
rect 75400 43000 81200 43200
rect 86000 43000 100000 43200
rect 0 43200 14000 43400
rect 18800 43200 48400 43400
rect 51600 43200 81200 43400
rect 86000 43200 100000 43400
rect 0 43400 14000 43600
rect 18800 43400 48400 43600
rect 51600 43400 81200 43600
rect 86000 43400 100000 43600
rect 0 43600 14000 43800
rect 18800 43600 48400 43800
rect 51600 43600 81200 43800
rect 86000 43600 100000 43800
rect 0 43800 14000 44000
rect 18800 43800 48400 44000
rect 51600 43800 81200 44000
rect 86000 43800 100000 44000
rect 0 44000 14000 44200
rect 19000 44000 48400 44200
rect 51600 44000 81200 44200
rect 86000 44000 100000 44200
rect 0 44200 14000 44400
rect 19000 44200 48400 44400
rect 51600 44200 81000 44400
rect 86000 44200 100000 44400
rect 0 44400 14000 44600
rect 19000 44400 48400 44600
rect 51600 44400 81000 44600
rect 86000 44400 100000 44600
rect 0 44600 14000 44800
rect 19000 44600 48400 44800
rect 51600 44600 81000 44800
rect 86000 44600 100000 44800
rect 0 44800 14000 45000
rect 19200 44800 48400 45000
rect 51600 44800 81000 45000
rect 86000 44800 100000 45000
rect 0 45000 3400 45200
rect 19200 45000 48400 45200
rect 51600 45000 80800 45200
rect 96600 45000 100000 45200
rect 0 45200 3000 45400
rect 19200 45200 48400 45400
rect 51600 45200 80800 45400
rect 97000 45200 100000 45400
rect 0 45400 2600 45600
rect 19400 45400 48400 45600
rect 51600 45400 80600 45600
rect 97400 45400 100000 45600
rect 0 45600 2400 45800
rect 19400 45600 48400 45800
rect 51600 45600 80600 45800
rect 97600 45600 100000 45800
rect 0 45800 2400 46000
rect 19600 45800 48400 46000
rect 51600 45800 80400 46000
rect 97800 45800 100000 46000
rect 0 46000 2200 46200
rect 19800 46000 48400 46200
rect 51600 46000 80400 46200
rect 97800 46000 100000 46200
rect 0 46200 2200 46400
rect 19800 46200 48400 46400
rect 51600 46200 80200 46400
rect 97800 46200 100000 46400
rect 0 46400 2200 46600
rect 20000 46400 48400 46600
rect 51600 46400 80000 46600
rect 98000 46400 100000 46600
rect 0 46600 2000 46800
rect 20200 46600 48400 46800
rect 51600 46600 79800 46800
rect 98000 46600 100000 46800
rect 0 46800 2000 47000
rect 20400 46800 48400 47000
rect 51600 46800 79800 47000
rect 98000 46800 100000 47000
rect 0 47000 2000 47200
rect 20400 47000 48400 47200
rect 51600 47000 79600 47200
rect 98000 47000 100000 47200
rect 0 47200 2200 47400
rect 20600 47200 48400 47400
rect 51600 47200 79400 47400
rect 98000 47200 100000 47400
rect 0 47400 2200 47600
rect 21000 47400 48400 47600
rect 51600 47400 79200 47600
rect 97800 47400 100000 47600
rect 0 47600 2200 47800
rect 21200 47600 48400 47800
rect 51600 47600 78800 47800
rect 97800 47600 100000 47800
rect 0 47800 2400 48000
rect 21400 47800 48400 48000
rect 51600 47800 78600 48000
rect 97600 47800 100000 48000
rect 0 48000 2600 48200
rect 21800 48000 48400 48200
rect 51600 48000 78200 48200
rect 97400 48000 100000 48200
rect 0 48200 2800 48400
rect 22200 48200 48400 48400
rect 51600 48200 78000 48400
rect 97200 48200 100000 48400
rect 0 48400 3200 48600
rect 22600 48400 48400 48600
rect 51600 48400 77600 48600
rect 96800 48400 100000 48600
rect 0 48600 14000 48800
rect 23200 48600 48400 48800
rect 51600 48600 77000 48800
rect 86000 48600 100000 48800
rect 0 48800 14000 49000
rect 24200 48800 48400 49000
rect 51600 48800 75800 49000
rect 86000 48800 100000 49000
rect 0 49000 14000 49200
rect 86000 49000 100000 49200
rect 0 49200 14000 49400
rect 86000 49200 100000 49400
rect 0 49400 14000 49600
rect 86000 49400 100000 49600
rect 0 49600 14000 49800
rect 86000 49600 100000 49800
rect 0 49800 14000 50000
rect 86000 49800 100000 50000
rect 0 50000 14000 50200
rect 86000 50000 100000 50200
rect 0 50200 14000 50400
rect 86000 50200 100000 50400
rect 0 50400 14000 50600
rect 86000 50400 100000 50600
rect 0 50600 14000 50800
rect 86000 50600 100000 50800
rect 0 50800 14000 51000
rect 24400 50800 48400 51000
rect 51600 50800 81200 51000
rect 86000 50800 100000 51000
rect 0 51000 14000 51200
rect 23200 51000 48400 51200
rect 51600 51000 81200 51200
rect 86000 51000 100000 51200
rect 0 51200 14000 51400
rect 22600 51200 48400 51400
rect 51600 51200 81200 51400
rect 86000 51200 100000 51400
rect 0 51400 14000 51600
rect 22200 51400 48400 51600
rect 51600 51400 81200 51600
rect 86000 51400 100000 51600
rect 0 51600 14000 51800
rect 21800 51600 48400 51800
rect 51600 51600 81200 51800
rect 86000 51600 100000 51800
rect 0 51800 3600 52000
rect 21400 51800 48400 52000
rect 51600 51800 81200 52000
rect 96400 51800 100000 52000
rect 0 52000 3000 52200
rect 21200 52000 48400 52200
rect 51600 52000 81200 52200
rect 97000 52000 100000 52200
rect 0 52200 2800 52400
rect 21000 52200 48400 52400
rect 51600 52200 81200 52400
rect 97200 52200 100000 52400
rect 0 52400 2600 52600
rect 20600 52400 48400 52600
rect 51600 52400 81200 52600
rect 97600 52400 100000 52600
rect 0 52600 2400 52800
rect 20400 52600 48400 52800
rect 51600 52600 81200 52800
rect 97600 52600 100000 52800
rect 0 52800 2200 53000
rect 20400 52800 48400 53000
rect 51600 52800 81200 53000
rect 97800 52800 100000 53000
rect 0 53000 2200 53200
rect 20200 53000 48400 53200
rect 51600 53000 81200 53200
rect 97800 53000 100000 53200
rect 0 53200 2200 53400
rect 20000 53200 48400 53400
rect 51600 53200 81200 53400
rect 98000 53200 100000 53400
rect 0 53400 2000 53600
rect 19800 53400 48400 53600
rect 51600 53400 81200 53600
rect 98000 53400 100000 53600
rect 0 53600 2000 53800
rect 19800 53600 48400 53800
rect 51600 53600 81200 53800
rect 98000 53600 100000 53800
rect 0 53800 2000 54000
rect 19600 53800 48400 54000
rect 51600 53800 81200 54000
rect 98000 53800 100000 54000
rect 0 54000 2200 54200
rect 19400 54000 48400 54200
rect 51600 54000 81200 54200
rect 98000 54000 100000 54200
rect 0 54200 2200 54400
rect 19400 54200 48400 54400
rect 51600 54200 81200 54400
rect 97800 54200 100000 54400
rect 0 54400 2200 54600
rect 19200 54400 48400 54600
rect 51600 54400 81200 54600
rect 97800 54400 100000 54600
rect 0 54600 2400 54800
rect 19200 54600 48400 54800
rect 51600 54600 81200 54800
rect 97600 54600 100000 54800
rect 0 54800 2600 55000
rect 19200 54800 48400 55000
rect 51600 54800 81200 55000
rect 97600 54800 100000 55000
rect 0 55000 2800 55200
rect 19000 55000 48400 55200
rect 51600 55000 81200 55200
rect 97200 55000 100000 55200
rect 0 55200 3200 55400
rect 19000 55200 48400 55400
rect 51600 55200 81200 55400
rect 97000 55200 100000 55400
rect 0 55400 14000 55600
rect 19000 55400 48400 55600
rect 51600 55400 81200 55600
rect 86000 55400 100000 55600
rect 0 55600 14000 55800
rect 19000 55600 48400 55800
rect 51600 55600 81200 55800
rect 86000 55600 100000 55800
rect 0 55800 14000 56000
rect 18800 55800 48400 56000
rect 51600 55800 81200 56000
rect 86000 55800 100000 56000
rect 0 56000 14000 56200
rect 18800 56000 48400 56200
rect 51600 56000 81200 56200
rect 86000 56000 100000 56200
rect 0 56200 14000 56400
rect 18800 56200 48400 56400
rect 51600 56200 81200 56400
rect 86000 56200 100000 56400
rect 0 56400 14000 56600
rect 18800 56400 48400 56600
rect 51600 56400 81200 56600
rect 86000 56400 100000 56600
rect 0 56600 14000 56800
rect 18800 56600 24600 56800
rect 51600 56600 57400 56800
rect 86000 56600 100000 56800
rect 0 56800 14000 57000
rect 18800 56800 24600 57000
rect 51600 56800 57400 57000
rect 86000 56800 100000 57000
rect 0 57000 14000 57200
rect 18800 57000 24600 57200
rect 51600 57000 57400 57200
rect 86000 57000 100000 57200
rect 0 57200 14000 57400
rect 18800 57200 24600 57400
rect 51600 57200 57400 57400
rect 86000 57200 100000 57400
rect 0 57400 14000 57600
rect 18800 57400 24600 57600
rect 51600 57400 57400 57600
rect 86000 57400 100000 57600
rect 0 57600 14000 57800
rect 18800 57600 24600 57800
rect 51600 57600 57400 57800
rect 86000 57600 100000 57800
rect 0 57800 14000 58000
rect 18800 57800 24600 58000
rect 51600 57800 57400 58000
rect 86000 57800 100000 58000
rect 0 58000 14000 58200
rect 18800 58000 24600 58200
rect 51600 58000 57400 58200
rect 86000 58000 100000 58200
rect 0 58200 14000 58400
rect 18800 58200 24600 58400
rect 51600 58200 57400 58400
rect 86000 58200 100000 58400
rect 0 58400 14000 58600
rect 18800 58400 24600 58600
rect 51600 58400 57400 58600
rect 86000 58400 100000 58600
rect 0 58600 14000 58800
rect 18800 58600 24600 58800
rect 51600 58600 57400 58800
rect 86000 58600 100000 58800
rect 0 58800 3200 59000
rect 18800 58800 24600 59000
rect 51600 58800 57400 59000
rect 97000 58800 100000 59000
rect 0 59000 2800 59200
rect 18800 59000 24600 59200
rect 51600 59000 57400 59200
rect 97200 59000 100000 59200
rect 0 59200 2600 59400
rect 18800 59200 24600 59400
rect 51600 59200 57400 59400
rect 97400 59200 100000 59400
rect 0 59400 2400 59600
rect 18800 59400 24600 59600
rect 51600 59400 57400 59600
rect 97600 59400 100000 59600
rect 0 59600 2200 59800
rect 18800 59600 24600 59800
rect 51600 59600 57400 59800
rect 97800 59600 100000 59800
rect 0 59800 2200 60000
rect 18800 59800 24600 60000
rect 51600 59800 57400 60000
rect 97800 59800 100000 60000
rect 0 60000 2200 60200
rect 18800 60000 24600 60200
rect 51600 60000 57400 60200
rect 98000 60000 100000 60200
rect 0 60200 2000 60400
rect 18800 60200 24600 60400
rect 51600 60200 57400 60400
rect 98000 60200 100000 60400
rect 0 60400 2000 60600
rect 18800 60400 24600 60600
rect 51600 60400 57400 60600
rect 98000 60400 100000 60600
rect 0 60600 2000 60800
rect 18800 60600 24600 60800
rect 51600 60600 57400 60800
rect 98000 60600 100000 60800
rect 0 60800 2000 61000
rect 18800 60800 24600 61000
rect 51600 60800 57400 61000
rect 98000 60800 100000 61000
rect 0 61000 2200 61200
rect 18800 61000 24600 61200
rect 51600 61000 57400 61200
rect 97800 61000 100000 61200
rect 0 61200 2200 61400
rect 18800 61200 24600 61400
rect 51600 61200 57400 61400
rect 97800 61200 100000 61400
rect 0 61400 2400 61600
rect 18800 61400 24600 61600
rect 51600 61400 57400 61600
rect 97800 61400 100000 61600
rect 0 61600 2400 61800
rect 18800 61600 24600 61800
rect 51600 61600 57400 61800
rect 97600 61600 100000 61800
rect 0 61800 2800 62000
rect 18800 61800 24600 62000
rect 51600 61800 57400 62000
rect 97400 61800 100000 62000
rect 0 62000 3000 62200
rect 18800 62000 24600 62200
rect 51600 62000 57400 62200
rect 97000 62000 100000 62200
rect 0 62200 3600 62400
rect 18800 62200 24600 62400
rect 51600 62200 57400 62400
rect 96400 62200 100000 62400
rect 0 62400 14000 62600
rect 18800 62400 24600 62600
rect 51600 62400 57400 62600
rect 86000 62400 100000 62600
rect 0 62600 14000 62800
rect 18800 62600 24600 62800
rect 51600 62600 57400 62800
rect 86000 62600 100000 62800
rect 0 62800 14000 63000
rect 18800 62800 24600 63000
rect 51600 62800 76400 63000
rect 86000 62800 100000 63000
rect 0 63000 14000 63200
rect 18800 63000 24600 63200
rect 51600 63000 77200 63200
rect 86000 63000 100000 63200
rect 0 63200 14000 63400
rect 18800 63200 24600 63400
rect 51600 63200 77600 63400
rect 86000 63200 100000 63400
rect 0 63400 14000 63600
rect 18800 63400 24600 63600
rect 51600 63400 78000 63600
rect 86000 63400 100000 63600
rect 0 63600 14000 63800
rect 18800 63600 24600 63800
rect 51600 63600 78400 63800
rect 86000 63600 100000 63800
rect 0 63800 14000 64000
rect 18800 63800 24600 64000
rect 51600 63800 78800 64000
rect 86000 63800 100000 64000
rect 0 64000 14000 64200
rect 18800 64000 24600 64200
rect 51800 64000 79000 64200
rect 86000 64000 100000 64200
rect 0 64200 14000 64400
rect 18800 64200 24600 64400
rect 51800 64200 79200 64400
rect 86000 64200 100000 64400
rect 0 64400 14000 64600
rect 18800 64400 24600 64600
rect 51800 64400 79400 64600
rect 86000 64400 100000 64600
rect 0 64600 14000 64800
rect 18800 64600 24600 64800
rect 52000 64600 79600 64800
rect 86000 64600 100000 64800
rect 0 64800 14000 65000
rect 18800 64800 24600 65000
rect 52000 64800 79800 65000
rect 86000 64800 100000 65000
rect 0 65000 14000 65200
rect 18800 65000 24600 65200
rect 52000 65000 80000 65200
rect 86000 65000 100000 65200
rect 0 65200 14000 65400
rect 18800 65200 24600 65400
rect 52200 65200 80200 65400
rect 86000 65200 100000 65400
rect 0 65400 14000 65600
rect 18800 65400 24600 65600
rect 52400 65400 80200 65600
rect 86000 65400 100000 65600
rect 0 65600 3200 65800
rect 18800 65600 24600 65800
rect 52400 65600 80400 65800
rect 97000 65600 100000 65800
rect 0 65800 2800 66000
rect 18800 65800 24600 66000
rect 52600 65800 80400 66000
rect 97200 65800 100000 66000
rect 0 66000 2600 66200
rect 18800 66000 24600 66200
rect 52600 66000 80600 66200
rect 97400 66000 100000 66200
rect 0 66200 2400 66400
rect 18800 66200 24600 66400
rect 52800 66200 80600 66400
rect 97600 66200 100000 66400
rect 0 66400 2200 66600
rect 18800 66400 24600 66600
rect 53000 66400 80800 66600
rect 97800 66400 100000 66600
rect 0 66600 2200 66800
rect 18800 66600 24600 66800
rect 53200 66600 80800 66800
rect 97800 66600 100000 66800
rect 0 66800 2200 67000
rect 18800 66800 24600 67000
rect 53400 66800 81000 67000
rect 98000 66800 100000 67000
rect 0 67000 2000 67200
rect 18800 67000 24600 67200
rect 53600 67000 81000 67200
rect 98000 67000 100000 67200
rect 0 67200 2000 67400
rect 18800 67200 24600 67400
rect 53800 67200 81000 67400
rect 98000 67200 100000 67400
rect 0 67400 2000 67600
rect 18800 67400 24600 67600
rect 54000 67400 81000 67600
rect 98000 67400 100000 67600
rect 0 67600 2000 67800
rect 18800 67600 24600 67800
rect 54400 67600 81200 67800
rect 98000 67600 100000 67800
rect 0 67800 2200 68000
rect 18800 67800 24600 68000
rect 54800 67800 81200 68000
rect 97800 67800 100000 68000
rect 0 68000 2200 68200
rect 18800 68000 24600 68200
rect 55000 68000 81200 68200
rect 97800 68000 100000 68200
rect 0 68200 2400 68400
rect 18800 68200 24600 68400
rect 55600 68200 81200 68400
rect 97800 68200 100000 68400
rect 0 68400 2400 68600
rect 18800 68400 24600 68600
rect 56400 68400 81200 68600
rect 97600 68400 100000 68600
rect 0 68600 2600 68800
rect 18800 68600 24600 68800
rect 75400 68600 81200 68800
rect 97400 68600 100000 68800
rect 0 68800 3000 69000
rect 18800 68800 24600 69000
rect 75400 68800 81200 69000
rect 97200 68800 100000 69000
rect 0 69000 3400 69200
rect 18800 69000 24600 69200
rect 75400 69000 81200 69200
rect 96600 69000 100000 69200
rect 0 69200 14000 69400
rect 18800 69200 24600 69400
rect 75400 69200 81200 69400
rect 86000 69200 100000 69400
rect 0 69400 14000 69600
rect 18800 69400 24600 69600
rect 75400 69400 81200 69600
rect 86000 69400 100000 69600
rect 0 69600 14000 69800
rect 18800 69600 24600 69800
rect 75400 69600 81200 69800
rect 86000 69600 100000 69800
rect 0 69800 14000 70000
rect 18800 69800 24600 70000
rect 75400 69800 81200 70000
rect 86000 69800 100000 70000
rect 0 70000 14000 70200
rect 18800 70000 24600 70200
rect 75400 70000 81200 70200
rect 86000 70000 100000 70200
rect 0 70200 14000 70400
rect 18800 70200 24600 70400
rect 75400 70200 81200 70400
rect 86000 70200 100000 70400
rect 0 70400 14000 70600
rect 18800 70400 24600 70600
rect 75400 70400 81200 70600
rect 86000 70400 100000 70600
rect 0 70600 14000 70800
rect 18800 70600 24600 70800
rect 75400 70600 81200 70800
rect 86000 70600 100000 70800
rect 0 70800 14000 71000
rect 18800 70800 24600 71000
rect 75400 70800 81200 71000
rect 86000 70800 100000 71000
rect 0 71000 14000 71200
rect 18800 71000 24600 71200
rect 75400 71000 81200 71200
rect 86000 71000 100000 71200
rect 0 71200 14000 71400
rect 18800 71200 24600 71400
rect 75400 71200 81200 71400
rect 86000 71200 100000 71400
rect 0 71400 14000 71600
rect 18800 71400 24600 71600
rect 75400 71400 81200 71600
rect 86000 71400 100000 71600
rect 0 71600 14000 71800
rect 18800 71600 24600 71800
rect 75400 71600 81200 71800
rect 86000 71600 100000 71800
rect 0 71800 14000 72000
rect 18800 71800 24600 72000
rect 75400 71800 81200 72000
rect 86000 71800 100000 72000
rect 0 72000 14000 72200
rect 18800 72000 24600 72200
rect 75400 72000 81200 72200
rect 86000 72000 100000 72200
rect 0 72200 14000 72400
rect 18800 72200 24600 72400
rect 75400 72200 81200 72400
rect 86000 72200 100000 72400
rect 0 72400 3200 72600
rect 18800 72400 24600 72600
rect 75400 72400 81200 72600
rect 96800 72400 100000 72600
rect 0 72600 2800 72800
rect 18800 72600 24600 72800
rect 75400 72600 81200 72800
rect 97200 72600 100000 72800
rect 0 72800 2600 73000
rect 18800 72800 24600 73000
rect 75400 72800 81200 73000
rect 97400 72800 100000 73000
rect 0 73000 2400 73200
rect 18800 73000 24600 73200
rect 75400 73000 81200 73200
rect 97600 73000 100000 73200
rect 0 73200 2400 73400
rect 18800 73200 24600 73400
rect 75400 73200 81200 73400
rect 97800 73200 100000 73400
rect 0 73400 2200 73600
rect 18800 73400 24600 73600
rect 75400 73400 81200 73600
rect 97800 73400 100000 73600
rect 0 73600 2200 73800
rect 18800 73600 24600 73800
rect 75400 73600 81200 73800
rect 98000 73600 100000 73800
rect 0 73800 2000 74000
rect 18800 73800 24600 74000
rect 75400 73800 81200 74000
rect 98000 73800 100000 74000
rect 0 74000 2000 74200
rect 18800 74000 24600 74200
rect 75400 74000 81200 74200
rect 98000 74000 100000 74200
rect 0 74200 2000 74400
rect 18800 74200 24600 74400
rect 75400 74200 81200 74400
rect 98000 74200 100000 74400
rect 0 74400 2000 74600
rect 18800 74400 24600 74600
rect 75400 74400 81200 74600
rect 98000 74400 100000 74600
rect 0 74600 2200 74800
rect 18800 74600 24600 74800
rect 75400 74600 81200 74800
rect 98000 74600 100000 74800
rect 0 74800 2200 75000
rect 18800 74800 48400 75000
rect 51600 74800 81200 75000
rect 97800 74800 100000 75000
rect 0 75000 2200 75200
rect 18800 75000 48400 75200
rect 51600 75000 81200 75200
rect 97800 75000 100000 75200
rect 0 75200 2400 75400
rect 18800 75200 48400 75400
rect 51600 75200 81200 75400
rect 97600 75200 100000 75400
rect 0 75400 2600 75600
rect 18800 75400 48400 75600
rect 51600 75400 81200 75600
rect 97400 75400 100000 75600
rect 0 75600 2800 75800
rect 19000 75600 48400 75800
rect 51600 75600 81200 75800
rect 97200 75600 100000 75800
rect 0 75800 3200 76000
rect 19000 75800 48400 76000
rect 51600 75800 81000 76000
rect 96800 75800 100000 76000
rect 0 76000 14000 76200
rect 19000 76000 48400 76200
rect 51600 76000 81000 76200
rect 86000 76000 100000 76200
rect 0 76200 14000 76400
rect 19000 76200 48400 76400
rect 51600 76200 81000 76400
rect 86000 76200 100000 76400
rect 0 76400 14000 76600
rect 19200 76400 48400 76600
rect 51600 76400 81000 76600
rect 86000 76400 100000 76600
rect 0 76600 14000 76800
rect 19200 76600 48400 76800
rect 51600 76600 80800 76800
rect 86000 76600 100000 76800
rect 0 76800 14000 77000
rect 19200 76800 48400 77000
rect 51600 76800 80800 77000
rect 86000 76800 100000 77000
rect 0 77000 14000 77200
rect 19400 77000 48400 77200
rect 51600 77000 80600 77200
rect 86000 77000 100000 77200
rect 0 77200 14000 77400
rect 19400 77200 48400 77400
rect 51600 77200 80600 77400
rect 86000 77200 100000 77400
rect 0 77400 14000 77600
rect 19600 77400 48400 77600
rect 51600 77400 80400 77600
rect 86000 77400 100000 77600
rect 0 77600 14000 77800
rect 19800 77600 48400 77800
rect 51600 77600 80400 77800
rect 86000 77600 100000 77800
rect 0 77800 14000 78000
rect 19800 77800 48400 78000
rect 51600 77800 80200 78000
rect 86000 77800 100000 78000
rect 0 78000 14000 78200
rect 20000 78000 48400 78200
rect 51600 78000 80000 78200
rect 86000 78000 100000 78200
rect 0 78200 14000 78400
rect 20200 78200 48400 78400
rect 51600 78200 79800 78400
rect 86000 78200 100000 78400
rect 0 78400 14000 78600
rect 20400 78400 48400 78600
rect 51600 78400 79800 78600
rect 86000 78400 100000 78600
rect 0 78600 14000 78800
rect 20400 78600 48400 78800
rect 51600 78600 79600 78800
rect 86000 78600 100000 78800
rect 0 78800 14000 79000
rect 20600 78800 48400 79000
rect 51600 78800 79400 79000
rect 86000 78800 100000 79000
rect 0 79000 14000 79200
rect 21000 79000 48400 79200
rect 51600 79000 79200 79200
rect 86000 79000 100000 79200
rect 0 79200 3400 79400
rect 21200 79200 48400 79400
rect 51600 79200 78800 79400
rect 96600 79200 100000 79400
rect 0 79400 3000 79600
rect 21400 79400 48400 79600
rect 51600 79400 78600 79600
rect 97000 79400 100000 79600
rect 0 79600 2600 79800
rect 21800 79600 48400 79800
rect 51600 79600 78200 79800
rect 97400 79600 100000 79800
rect 0 79800 2400 80000
rect 22200 79800 48400 80000
rect 51600 79800 78000 80000
rect 97600 79800 100000 80000
rect 0 80000 2400 80200
rect 22600 80000 48400 80200
rect 51600 80000 77600 80200
rect 97800 80000 100000 80200
rect 0 80200 2200 80400
rect 23200 80200 48400 80400
rect 51600 80200 77000 80400
rect 97800 80200 100000 80400
rect 0 80400 2200 80600
rect 24200 80400 48400 80600
rect 51600 80400 75800 80600
rect 97800 80400 100000 80600
rect 0 80600 2200 80800
rect 98000 80600 100000 80800
rect 0 80800 2000 81000
rect 98000 80800 100000 81000
rect 0 81000 2000 81200
rect 98000 81000 100000 81200
rect 0 81200 2000 81400
rect 98000 81200 100000 81400
rect 0 81400 2200 81600
rect 98000 81400 100000 81600
rect 0 81600 2200 81800
rect 97800 81600 100000 81800
rect 0 81800 2200 82000
rect 97800 81800 100000 82000
rect 0 82000 2400 82200
rect 97600 82000 100000 82200
rect 0 82200 2600 82400
rect 97600 82200 100000 82400
rect 0 82400 2800 82600
rect 97200 82400 100000 82600
rect 0 82600 3200 82800
rect 97000 82600 100000 82800
rect 0 82800 14000 83000
rect 86000 82800 100000 83000
rect 0 83000 14000 83200
rect 86000 83000 100000 83200
rect 0 83200 14000 83400
rect 86000 83200 100000 83400
rect 0 83400 14000 83600
rect 86000 83400 100000 83600
rect 0 83600 14000 83800
rect 86000 83600 100000 83800
rect 0 83800 14000 84000
rect 86000 83800 100000 84000
rect 0 84000 14000 84200
rect 86000 84000 100000 84200
rect 0 84200 14000 84400
rect 86000 84200 100000 84400
rect 0 84400 14000 84600
rect 86000 84400 100000 84600
rect 0 84600 14000 84800
rect 86000 84600 100000 84800
rect 0 84800 14000 85000
rect 86000 84800 100000 85000
rect 0 85000 14200 85200
rect 86000 85000 100000 85200
rect 0 85200 14200 85400
rect 85800 85200 100000 85400
rect 0 85400 14400 85600
rect 85800 85400 100000 85600
rect 0 85600 14600 85800
rect 85600 85600 100000 85800
rect 0 85800 14800 86000
rect 85400 85800 100000 86000
rect 0 86000 15000 86200
rect 85000 86000 100000 86200
rect 0 86200 17400 86400
rect 21000 86200 24200 86400
rect 27800 86200 31200 86400
rect 34800 86200 38000 86400
rect 41600 86200 44800 86400
rect 48400 86200 51600 86400
rect 55200 86200 58600 86400
rect 62000 86200 65400 86400
rect 69000 86200 72200 86400
rect 75800 86200 79000 86400
rect 82600 86200 100000 86400
rect 0 86400 17400 86600
rect 21000 86400 24200 86600
rect 27800 86400 31200 86600
rect 34800 86400 38000 86600
rect 41600 86400 44800 86600
rect 48400 86400 51600 86600
rect 55200 86400 58600 86600
rect 62000 86400 65400 86600
rect 69000 86400 72200 86600
rect 75800 86400 79000 86600
rect 82600 86400 100000 86600
rect 0 86600 17400 86800
rect 21000 86600 24200 86800
rect 27800 86600 31200 86800
rect 34800 86600 38000 86800
rect 41600 86600 44800 86800
rect 48400 86600 51600 86800
rect 55200 86600 58600 86800
rect 62000 86600 65400 86800
rect 69000 86600 72200 86800
rect 75800 86600 79000 86800
rect 82600 86600 100000 86800
rect 0 86800 17400 87000
rect 21000 86800 24200 87000
rect 27800 86800 31200 87000
rect 34800 86800 38000 87000
rect 41600 86800 44800 87000
rect 48400 86800 51600 87000
rect 55200 86800 58600 87000
rect 62000 86800 65400 87000
rect 69000 86800 72200 87000
rect 75800 86800 79000 87000
rect 82600 86800 100000 87000
rect 0 87000 17400 87200
rect 21000 87000 24200 87200
rect 27800 87000 31200 87200
rect 34800 87000 38000 87200
rect 41600 87000 44800 87200
rect 48400 87000 51600 87200
rect 55200 87000 58600 87200
rect 62000 87000 65400 87200
rect 69000 87000 72200 87200
rect 75800 87000 79000 87200
rect 82600 87000 100000 87200
rect 0 87200 17400 87400
rect 21000 87200 24200 87400
rect 27800 87200 31200 87400
rect 34800 87200 38000 87400
rect 41600 87200 44800 87400
rect 48400 87200 51600 87400
rect 55200 87200 58600 87400
rect 62000 87200 65400 87400
rect 69000 87200 72200 87400
rect 75800 87200 79000 87400
rect 82600 87200 100000 87400
rect 0 87400 17400 87600
rect 21000 87400 24200 87600
rect 27800 87400 31200 87600
rect 34800 87400 38000 87600
rect 41600 87400 44800 87600
rect 48400 87400 51600 87600
rect 55200 87400 58600 87600
rect 62000 87400 65400 87600
rect 69000 87400 72200 87600
rect 75800 87400 79000 87600
rect 82600 87400 100000 87600
rect 0 87600 17400 87800
rect 21000 87600 24200 87800
rect 27800 87600 31200 87800
rect 34800 87600 38000 87800
rect 41600 87600 44800 87800
rect 48400 87600 51600 87800
rect 55200 87600 58600 87800
rect 62000 87600 65400 87800
rect 69000 87600 72200 87800
rect 75800 87600 79000 87800
rect 82600 87600 100000 87800
rect 0 87800 17400 88000
rect 21000 87800 24200 88000
rect 27800 87800 31200 88000
rect 34800 87800 38000 88000
rect 41600 87800 44800 88000
rect 48400 87800 51600 88000
rect 55200 87800 58600 88000
rect 62000 87800 65400 88000
rect 69000 87800 72200 88000
rect 75800 87800 79000 88000
rect 82600 87800 100000 88000
rect 0 88000 17400 88200
rect 21000 88000 24200 88200
rect 27800 88000 31200 88200
rect 34800 88000 38000 88200
rect 41600 88000 44800 88200
rect 48400 88000 51600 88200
rect 55200 88000 58600 88200
rect 62000 88000 65400 88200
rect 69000 88000 72200 88200
rect 75800 88000 79000 88200
rect 82600 88000 100000 88200
rect 0 88200 17400 88400
rect 21000 88200 24200 88400
rect 27800 88200 31200 88400
rect 34800 88200 38000 88400
rect 41600 88200 44800 88400
rect 48400 88200 51600 88400
rect 55200 88200 58600 88400
rect 62000 88200 65400 88400
rect 69000 88200 72200 88400
rect 75800 88200 79000 88400
rect 82600 88200 100000 88400
rect 0 88400 17400 88600
rect 21000 88400 24200 88600
rect 27800 88400 31200 88600
rect 34800 88400 38000 88600
rect 41600 88400 44800 88600
rect 48400 88400 51600 88600
rect 55200 88400 58600 88600
rect 62000 88400 65400 88600
rect 69000 88400 72200 88600
rect 75800 88400 79000 88600
rect 82600 88400 100000 88600
rect 0 88600 17400 88800
rect 21000 88600 24200 88800
rect 27800 88600 31200 88800
rect 34800 88600 38000 88800
rect 41600 88600 44800 88800
rect 48400 88600 51600 88800
rect 55200 88600 58600 88800
rect 62000 88600 65400 88800
rect 69000 88600 72200 88800
rect 75800 88600 79000 88800
rect 82600 88600 100000 88800
rect 0 88800 17400 89000
rect 21000 88800 24200 89000
rect 27800 88800 31200 89000
rect 34800 88800 38000 89000
rect 41600 88800 44800 89000
rect 48400 88800 51600 89000
rect 55200 88800 58600 89000
rect 62000 88800 65400 89000
rect 69000 88800 72200 89000
rect 75800 88800 79000 89000
rect 82600 88800 100000 89000
rect 0 89000 17400 89200
rect 21000 89000 24200 89200
rect 27800 89000 31200 89200
rect 34800 89000 38000 89200
rect 41600 89000 44800 89200
rect 48400 89000 51600 89200
rect 55200 89000 58600 89200
rect 62000 89000 65400 89200
rect 69000 89000 72200 89200
rect 75800 89000 79000 89200
rect 82600 89000 100000 89200
rect 0 89200 17400 89400
rect 21000 89200 24200 89400
rect 27800 89200 31200 89400
rect 34800 89200 38000 89400
rect 41600 89200 44800 89400
rect 48400 89200 51600 89400
rect 55200 89200 58600 89400
rect 62000 89200 65400 89400
rect 69000 89200 72200 89400
rect 75800 89200 79000 89400
rect 82600 89200 100000 89400
rect 0 89400 17400 89600
rect 21000 89400 24200 89600
rect 27800 89400 31200 89600
rect 34800 89400 38000 89600
rect 41600 89400 44800 89600
rect 48400 89400 51600 89600
rect 55200 89400 58600 89600
rect 62000 89400 65400 89600
rect 69000 89400 72200 89600
rect 75800 89400 79000 89600
rect 82600 89400 100000 89600
rect 0 89600 17400 89800
rect 21000 89600 24200 89800
rect 27800 89600 31200 89800
rect 34800 89600 38000 89800
rect 41600 89600 44800 89800
rect 48400 89600 51600 89800
rect 55200 89600 58600 89800
rect 62000 89600 65400 89800
rect 69000 89600 72200 89800
rect 75800 89600 79000 89800
rect 82600 89600 100000 89800
rect 0 89800 17400 90000
rect 21000 89800 24200 90000
rect 27800 89800 31200 90000
rect 34800 89800 38000 90000
rect 41600 89800 44800 90000
rect 48400 89800 51600 90000
rect 55200 89800 58600 90000
rect 62000 89800 65400 90000
rect 69000 89800 72200 90000
rect 75800 89800 79000 90000
rect 82600 89800 100000 90000
rect 0 90000 17400 90200
rect 21000 90000 24200 90200
rect 27800 90000 31200 90200
rect 34800 90000 38000 90200
rect 41600 90000 44800 90200
rect 48400 90000 51600 90200
rect 55200 90000 58600 90200
rect 62000 90000 65400 90200
rect 69000 90000 72200 90200
rect 75800 90000 79000 90200
rect 82600 90000 100000 90200
rect 0 90200 17400 90400
rect 21000 90200 24200 90400
rect 27800 90200 31200 90400
rect 34800 90200 38000 90400
rect 41600 90200 44800 90400
rect 48400 90200 51600 90400
rect 55200 90200 58600 90400
rect 62000 90200 65400 90400
rect 69000 90200 72200 90400
rect 75800 90200 79000 90400
rect 82600 90200 100000 90400
rect 0 90400 17400 90600
rect 21000 90400 24200 90600
rect 27800 90400 31200 90600
rect 34800 90400 38000 90600
rect 41600 90400 44800 90600
rect 48400 90400 51600 90600
rect 55200 90400 58600 90600
rect 62000 90400 65400 90600
rect 69000 90400 72200 90600
rect 75800 90400 79000 90600
rect 82600 90400 100000 90600
rect 0 90600 17400 90800
rect 21000 90600 24200 90800
rect 27800 90600 31200 90800
rect 34800 90600 38000 90800
rect 41600 90600 44800 90800
rect 48400 90600 51600 90800
rect 55200 90600 58600 90800
rect 62000 90600 65400 90800
rect 69000 90600 72200 90800
rect 75800 90600 79000 90800
rect 82600 90600 100000 90800
rect 0 90800 17400 91000
rect 21000 90800 24200 91000
rect 27800 90800 31200 91000
rect 34800 90800 38000 91000
rect 41600 90800 44800 91000
rect 48400 90800 51600 91000
rect 55200 90800 58600 91000
rect 62000 90800 65400 91000
rect 69000 90800 72200 91000
rect 75800 90800 79000 91000
rect 82600 90800 100000 91000
rect 0 91000 17400 91200
rect 21000 91000 24200 91200
rect 27800 91000 31200 91200
rect 34800 91000 38000 91200
rect 41600 91000 44800 91200
rect 48400 91000 51600 91200
rect 55200 91000 58600 91200
rect 62000 91000 65400 91200
rect 69000 91000 72200 91200
rect 75800 91000 79000 91200
rect 82600 91000 100000 91200
rect 0 91200 17400 91400
rect 21000 91200 24200 91400
rect 27800 91200 31200 91400
rect 34800 91200 38000 91400
rect 41600 91200 44800 91400
rect 48400 91200 51600 91400
rect 55200 91200 58600 91400
rect 62000 91200 65400 91400
rect 69000 91200 72200 91400
rect 75800 91200 79000 91400
rect 82600 91200 100000 91400
rect 0 91400 17400 91600
rect 21000 91400 24200 91600
rect 27800 91400 31200 91600
rect 34800 91400 38000 91600
rect 41600 91400 44800 91600
rect 48400 91400 51600 91600
rect 55200 91400 58600 91600
rect 62000 91400 65400 91600
rect 69000 91400 72200 91600
rect 75800 91400 79000 91600
rect 82600 91400 100000 91600
rect 0 91600 17400 91800
rect 21000 91600 24200 91800
rect 27800 91600 31200 91800
rect 34800 91600 38000 91800
rect 41600 91600 44800 91800
rect 48400 91600 51600 91800
rect 55200 91600 58600 91800
rect 62000 91600 65400 91800
rect 69000 91600 72200 91800
rect 75800 91600 79000 91800
rect 82600 91600 100000 91800
rect 0 91800 17400 92000
rect 21000 91800 24200 92000
rect 27800 91800 31200 92000
rect 34800 91800 38000 92000
rect 41600 91800 44800 92000
rect 48400 91800 51600 92000
rect 55200 91800 58600 92000
rect 62000 91800 65400 92000
rect 69000 91800 72200 92000
rect 75800 91800 79000 92000
rect 82600 91800 100000 92000
rect 0 92000 17400 92200
rect 21000 92000 24200 92200
rect 27800 92000 31200 92200
rect 34800 92000 38000 92200
rect 41600 92000 44800 92200
rect 48400 92000 51600 92200
rect 55200 92000 58600 92200
rect 62000 92000 65400 92200
rect 69000 92000 72200 92200
rect 75800 92000 79000 92200
rect 82600 92000 100000 92200
rect 0 92200 17400 92400
rect 21000 92200 24200 92400
rect 27800 92200 31200 92400
rect 34800 92200 38000 92400
rect 41600 92200 44800 92400
rect 48400 92200 51600 92400
rect 55200 92200 58600 92400
rect 62000 92200 65400 92400
rect 69000 92200 72200 92400
rect 75800 92200 79000 92400
rect 82600 92200 100000 92400
rect 0 92400 17400 92600
rect 21000 92400 24200 92600
rect 27800 92400 31200 92600
rect 34800 92400 38000 92600
rect 41600 92400 44800 92600
rect 48400 92400 51600 92600
rect 55200 92400 58600 92600
rect 62000 92400 65400 92600
rect 69000 92400 72200 92600
rect 75800 92400 79000 92600
rect 82600 92400 100000 92600
rect 0 92600 17400 92800
rect 21000 92600 24200 92800
rect 27800 92600 31200 92800
rect 34800 92600 38000 92800
rect 41600 92600 44800 92800
rect 48400 92600 51600 92800
rect 55200 92600 58600 92800
rect 62000 92600 65400 92800
rect 69000 92600 72200 92800
rect 75800 92600 79000 92800
rect 82600 92600 100000 92800
rect 0 92800 17400 93000
rect 21000 92800 24200 93000
rect 27800 92800 31200 93000
rect 34800 92800 38000 93000
rect 41600 92800 44800 93000
rect 48400 92800 51600 93000
rect 55200 92800 58600 93000
rect 62000 92800 65400 93000
rect 69000 92800 72200 93000
rect 75800 92800 79000 93000
rect 82600 92800 100000 93000
rect 0 93000 17400 93200
rect 21000 93000 24200 93200
rect 27800 93000 31200 93200
rect 34800 93000 38000 93200
rect 41600 93000 44800 93200
rect 48400 93000 51600 93200
rect 55200 93000 58600 93200
rect 62000 93000 65400 93200
rect 69000 93000 72200 93200
rect 75800 93000 79000 93200
rect 82600 93000 100000 93200
rect 0 93200 17400 93400
rect 21000 93200 24200 93400
rect 27800 93200 31200 93400
rect 34800 93200 38000 93400
rect 41600 93200 44800 93400
rect 48400 93200 51600 93400
rect 55200 93200 58600 93400
rect 62000 93200 65400 93400
rect 69000 93200 72200 93400
rect 75800 93200 79000 93400
rect 82600 93200 100000 93400
rect 0 93400 17400 93600
rect 21000 93400 24200 93600
rect 27800 93400 31200 93600
rect 34800 93400 38000 93600
rect 41600 93400 44800 93600
rect 48400 93400 51600 93600
rect 55200 93400 58600 93600
rect 62000 93400 65400 93600
rect 69000 93400 72200 93600
rect 75800 93400 79000 93600
rect 82600 93400 100000 93600
rect 0 93600 17400 93800
rect 21000 93600 24200 93800
rect 27800 93600 31200 93800
rect 34800 93600 38000 93800
rect 41600 93600 44800 93800
rect 48400 93600 51600 93800
rect 55200 93600 58600 93800
rect 62000 93600 65400 93800
rect 69000 93600 72200 93800
rect 75800 93600 79000 93800
rect 82600 93600 100000 93800
rect 0 93800 17400 94000
rect 21000 93800 24200 94000
rect 27800 93800 31200 94000
rect 34800 93800 38000 94000
rect 41600 93800 44800 94000
rect 48400 93800 51600 94000
rect 55200 93800 58600 94000
rect 62000 93800 65400 94000
rect 69000 93800 72200 94000
rect 75800 93800 79000 94000
rect 82600 93800 100000 94000
rect 0 94000 17400 94200
rect 21000 94000 24200 94200
rect 27800 94000 31200 94200
rect 34800 94000 38000 94200
rect 41600 94000 44800 94200
rect 48400 94000 51600 94200
rect 55200 94000 58600 94200
rect 62000 94000 65400 94200
rect 69000 94000 72200 94200
rect 75800 94000 79000 94200
rect 82600 94000 100000 94200
rect 0 94200 17400 94400
rect 21000 94200 24200 94400
rect 27800 94200 31200 94400
rect 34800 94200 38000 94400
rect 41600 94200 44800 94400
rect 48400 94200 51600 94400
rect 55200 94200 58600 94400
rect 62000 94200 65400 94400
rect 69000 94200 72200 94400
rect 75800 94200 79000 94400
rect 82600 94200 100000 94400
rect 0 94400 17400 94600
rect 21000 94400 24200 94600
rect 27800 94400 31200 94600
rect 34800 94400 38000 94600
rect 41600 94400 44800 94600
rect 48400 94400 51600 94600
rect 55200 94400 58600 94600
rect 62000 94400 65400 94600
rect 69000 94400 72200 94600
rect 75800 94400 79000 94600
rect 82600 94400 100000 94600
rect 0 94600 17400 94800
rect 21000 94600 24200 94800
rect 27800 94600 31200 94800
rect 34800 94600 38000 94800
rect 41600 94600 44800 94800
rect 48400 94600 51600 94800
rect 55200 94600 58600 94800
rect 62000 94600 65400 94800
rect 69000 94600 72200 94800
rect 75800 94600 79000 94800
rect 82600 94600 100000 94800
rect 0 94800 17400 95000
rect 21000 94800 24200 95000
rect 27800 94800 31200 95000
rect 34800 94800 38000 95000
rect 41600 94800 44800 95000
rect 48400 94800 51600 95000
rect 55200 94800 58600 95000
rect 62000 94800 65400 95000
rect 69000 94800 72200 95000
rect 75800 94800 79000 95000
rect 82600 94800 100000 95000
rect 0 95000 17400 95200
rect 21000 95000 24200 95200
rect 27800 95000 31200 95200
rect 34800 95000 38000 95200
rect 41600 95000 44800 95200
rect 48400 95000 51600 95200
rect 55200 95000 58600 95200
rect 62000 95000 65400 95200
rect 69000 95000 72200 95200
rect 75800 95000 79000 95200
rect 82600 95000 100000 95200
rect 0 95200 17400 95400
rect 21000 95200 24200 95400
rect 27800 95200 31200 95400
rect 34800 95200 38000 95400
rect 41600 95200 44800 95400
rect 48400 95200 51600 95400
rect 55200 95200 58600 95400
rect 62000 95200 65400 95400
rect 69000 95200 72200 95400
rect 75800 95200 79000 95400
rect 82600 95200 100000 95400
rect 0 95400 17400 95600
rect 21000 95400 24200 95600
rect 27800 95400 31200 95600
rect 34800 95400 38000 95600
rect 41600 95400 44800 95600
rect 48400 95400 51600 95600
rect 55200 95400 58600 95600
rect 62000 95400 65400 95600
rect 69000 95400 72200 95600
rect 75800 95400 79000 95600
rect 82600 95400 100000 95600
rect 0 95600 17400 95800
rect 21000 95600 24200 95800
rect 27800 95600 31200 95800
rect 34800 95600 38000 95800
rect 41600 95600 44800 95800
rect 48400 95600 51600 95800
rect 55200 95600 58600 95800
rect 62000 95600 65400 95800
rect 69000 95600 72200 95800
rect 75800 95600 79000 95800
rect 82600 95600 100000 95800
rect 0 95800 17400 96000
rect 21000 95800 24200 96000
rect 27800 95800 31200 96000
rect 34800 95800 38000 96000
rect 41600 95800 44800 96000
rect 48400 95800 51600 96000
rect 55200 95800 58600 96000
rect 62000 95800 65400 96000
rect 69000 95800 72200 96000
rect 75800 95800 79000 96000
rect 82600 95800 100000 96000
rect 0 96000 17400 96200
rect 21000 96000 24200 96200
rect 27800 96000 31200 96200
rect 34800 96000 38000 96200
rect 41600 96000 44800 96200
rect 48400 96000 51600 96200
rect 55200 96000 58600 96200
rect 62000 96000 65400 96200
rect 69000 96000 72200 96200
rect 75800 96000 79000 96200
rect 82600 96000 100000 96200
rect 0 96200 17400 96400
rect 21000 96200 24200 96400
rect 27800 96200 31200 96400
rect 34800 96200 38000 96400
rect 41600 96200 44800 96400
rect 48400 96200 51600 96400
rect 55200 96200 58600 96400
rect 62000 96200 65400 96400
rect 69000 96200 72200 96400
rect 75800 96200 79000 96400
rect 82600 96200 100000 96400
rect 0 96400 17400 96600
rect 21000 96400 24400 96600
rect 27800 96400 31200 96600
rect 34800 96400 38000 96600
rect 41600 96400 44800 96600
rect 48400 96400 51600 96600
rect 55200 96400 58600 96600
rect 62000 96400 65400 96600
rect 69000 96400 72200 96600
rect 75800 96400 79000 96600
rect 82600 96400 100000 96600
rect 0 96600 17400 96800
rect 21000 96600 24400 96800
rect 27800 96600 31200 96800
rect 34600 96600 38000 96800
rect 41600 96600 44800 96800
rect 48400 96600 51600 96800
rect 55200 96600 58600 96800
rect 62000 96600 65400 96800
rect 69000 96600 72200 96800
rect 75800 96600 79000 96800
rect 82600 96600 100000 96800
rect 0 96800 17400 97000
rect 21000 96800 24400 97000
rect 27800 96800 31200 97000
rect 34600 96800 38000 97000
rect 41600 96800 44800 97000
rect 48400 96800 51800 97000
rect 55200 96800 58600 97000
rect 62000 96800 65400 97000
rect 68800 96800 72200 97000
rect 75800 96800 79000 97000
rect 82600 96800 100000 97000
rect 0 97000 17600 97200
rect 21000 97000 24400 97200
rect 27800 97000 31200 97200
rect 34600 97000 38000 97200
rect 41400 97000 45000 97200
rect 48200 97000 51800 97200
rect 55200 97000 58600 97200
rect 62000 97000 65400 97200
rect 68800 97000 72200 97200
rect 75600 97000 79200 97200
rect 82400 97000 100000 97200
rect 0 97200 17600 97400
rect 20800 97200 24400 97400
rect 27600 97200 31400 97400
rect 34600 97200 38200 97400
rect 41400 97200 45000 97400
rect 48200 97200 51800 97400
rect 55000 97200 58800 97400
rect 61800 97200 65600 97400
rect 68800 97200 72400 97400
rect 75600 97200 79200 97400
rect 82400 97200 100000 97400
rect 0 97400 17800 97600
rect 20800 97400 24600 97600
rect 27600 97400 31400 97600
rect 34400 97400 38200 97600
rect 41200 97400 45200 97600
rect 48000 97400 52000 97600
rect 55000 97400 58800 97600
rect 61800 97400 65600 97600
rect 68600 97400 72400 97600
rect 75400 97400 79400 97600
rect 82200 97400 100000 97600
rect 0 97600 18000 97800
rect 20600 97600 24800 97800
rect 27400 97600 31600 97800
rect 34200 97600 38400 97800
rect 41000 97600 45200 97800
rect 48000 97600 52200 97800
rect 54800 97600 59000 97800
rect 61600 97600 65800 97800
rect 68400 97600 72600 97800
rect 75200 97600 79600 97800
rect 82200 97600 100000 97800
rect 0 97800 18200 98000
rect 20400 97800 25000 98000
rect 27200 97800 31800 98000
rect 34000 97800 38600 98000
rect 40800 97800 45600 98000
rect 47600 97800 52400 98000
rect 54600 97800 59200 98000
rect 61400 97800 66000 98000
rect 68200 97800 72800 98000
rect 75000 97800 79800 98000
rect 81800 97800 100000 98000
rect 0 98000 18600 98200
rect 20000 98000 25400 98200
rect 26800 98000 32200 98200
rect 33600 98000 39000 98200
rect 40600 98000 45800 98200
rect 47400 98000 52800 98200
rect 54200 98000 59600 98200
rect 61000 98000 66400 98200
rect 67800 98000 73200 98200
rect 74800 98000 80000 98200
rect 81600 98000 100000 98200
rect 0 98200 100000 98400
rect 0 98400 100000 98600
rect 0 98600 100000 98800
rect 0 98800 100000 99000
rect 0 99000 100000 99200
rect 0 99200 100000 99400
rect 0 99400 100000 99600
rect 0 99600 100000 99800
rect 0 99800 100000 100000
<< labels >>
rlabel metal4 s 100500 0 100600 100000 6 vccd1
port 1 nsew power input
rlabel metal4 s -600 0 -500 100000 6 vssd1
port 2 nsew ground input
<< end >>
