magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< pwell >>
rect -710 -700 710 700
<< nmos >>
rect -524 -500 -424 500
rect -366 -500 -266 500
rect -208 -500 -108 500
rect -50 -500 50 500
rect 108 -500 208 500
rect 266 -500 366 500
rect 424 -500 524 500
<< ndiff >>
rect -582 459 -524 500
rect -582 425 -570 459
rect -536 425 -524 459
rect -582 391 -524 425
rect -582 357 -570 391
rect -536 357 -524 391
rect -582 323 -524 357
rect -582 289 -570 323
rect -536 289 -524 323
rect -582 255 -524 289
rect -582 221 -570 255
rect -536 221 -524 255
rect -582 187 -524 221
rect -582 153 -570 187
rect -536 153 -524 187
rect -582 119 -524 153
rect -582 85 -570 119
rect -536 85 -524 119
rect -582 51 -524 85
rect -582 17 -570 51
rect -536 17 -524 51
rect -582 -17 -524 17
rect -582 -51 -570 -17
rect -536 -51 -524 -17
rect -582 -85 -524 -51
rect -582 -119 -570 -85
rect -536 -119 -524 -85
rect -582 -153 -524 -119
rect -582 -187 -570 -153
rect -536 -187 -524 -153
rect -582 -221 -524 -187
rect -582 -255 -570 -221
rect -536 -255 -524 -221
rect -582 -289 -524 -255
rect -582 -323 -570 -289
rect -536 -323 -524 -289
rect -582 -357 -524 -323
rect -582 -391 -570 -357
rect -536 -391 -524 -357
rect -582 -425 -524 -391
rect -582 -459 -570 -425
rect -536 -459 -524 -425
rect -582 -500 -524 -459
rect -424 459 -366 500
rect -424 425 -412 459
rect -378 425 -366 459
rect -424 391 -366 425
rect -424 357 -412 391
rect -378 357 -366 391
rect -424 323 -366 357
rect -424 289 -412 323
rect -378 289 -366 323
rect -424 255 -366 289
rect -424 221 -412 255
rect -378 221 -366 255
rect -424 187 -366 221
rect -424 153 -412 187
rect -378 153 -366 187
rect -424 119 -366 153
rect -424 85 -412 119
rect -378 85 -366 119
rect -424 51 -366 85
rect -424 17 -412 51
rect -378 17 -366 51
rect -424 -17 -366 17
rect -424 -51 -412 -17
rect -378 -51 -366 -17
rect -424 -85 -366 -51
rect -424 -119 -412 -85
rect -378 -119 -366 -85
rect -424 -153 -366 -119
rect -424 -187 -412 -153
rect -378 -187 -366 -153
rect -424 -221 -366 -187
rect -424 -255 -412 -221
rect -378 -255 -366 -221
rect -424 -289 -366 -255
rect -424 -323 -412 -289
rect -378 -323 -366 -289
rect -424 -357 -366 -323
rect -424 -391 -412 -357
rect -378 -391 -366 -357
rect -424 -425 -366 -391
rect -424 -459 -412 -425
rect -378 -459 -366 -425
rect -424 -500 -366 -459
rect -266 459 -208 500
rect -266 425 -254 459
rect -220 425 -208 459
rect -266 391 -208 425
rect -266 357 -254 391
rect -220 357 -208 391
rect -266 323 -208 357
rect -266 289 -254 323
rect -220 289 -208 323
rect -266 255 -208 289
rect -266 221 -254 255
rect -220 221 -208 255
rect -266 187 -208 221
rect -266 153 -254 187
rect -220 153 -208 187
rect -266 119 -208 153
rect -266 85 -254 119
rect -220 85 -208 119
rect -266 51 -208 85
rect -266 17 -254 51
rect -220 17 -208 51
rect -266 -17 -208 17
rect -266 -51 -254 -17
rect -220 -51 -208 -17
rect -266 -85 -208 -51
rect -266 -119 -254 -85
rect -220 -119 -208 -85
rect -266 -153 -208 -119
rect -266 -187 -254 -153
rect -220 -187 -208 -153
rect -266 -221 -208 -187
rect -266 -255 -254 -221
rect -220 -255 -208 -221
rect -266 -289 -208 -255
rect -266 -323 -254 -289
rect -220 -323 -208 -289
rect -266 -357 -208 -323
rect -266 -391 -254 -357
rect -220 -391 -208 -357
rect -266 -425 -208 -391
rect -266 -459 -254 -425
rect -220 -459 -208 -425
rect -266 -500 -208 -459
rect -108 459 -50 500
rect -108 425 -96 459
rect -62 425 -50 459
rect -108 391 -50 425
rect -108 357 -96 391
rect -62 357 -50 391
rect -108 323 -50 357
rect -108 289 -96 323
rect -62 289 -50 323
rect -108 255 -50 289
rect -108 221 -96 255
rect -62 221 -50 255
rect -108 187 -50 221
rect -108 153 -96 187
rect -62 153 -50 187
rect -108 119 -50 153
rect -108 85 -96 119
rect -62 85 -50 119
rect -108 51 -50 85
rect -108 17 -96 51
rect -62 17 -50 51
rect -108 -17 -50 17
rect -108 -51 -96 -17
rect -62 -51 -50 -17
rect -108 -85 -50 -51
rect -108 -119 -96 -85
rect -62 -119 -50 -85
rect -108 -153 -50 -119
rect -108 -187 -96 -153
rect -62 -187 -50 -153
rect -108 -221 -50 -187
rect -108 -255 -96 -221
rect -62 -255 -50 -221
rect -108 -289 -50 -255
rect -108 -323 -96 -289
rect -62 -323 -50 -289
rect -108 -357 -50 -323
rect -108 -391 -96 -357
rect -62 -391 -50 -357
rect -108 -425 -50 -391
rect -108 -459 -96 -425
rect -62 -459 -50 -425
rect -108 -500 -50 -459
rect 50 459 108 500
rect 50 425 62 459
rect 96 425 108 459
rect 50 391 108 425
rect 50 357 62 391
rect 96 357 108 391
rect 50 323 108 357
rect 50 289 62 323
rect 96 289 108 323
rect 50 255 108 289
rect 50 221 62 255
rect 96 221 108 255
rect 50 187 108 221
rect 50 153 62 187
rect 96 153 108 187
rect 50 119 108 153
rect 50 85 62 119
rect 96 85 108 119
rect 50 51 108 85
rect 50 17 62 51
rect 96 17 108 51
rect 50 -17 108 17
rect 50 -51 62 -17
rect 96 -51 108 -17
rect 50 -85 108 -51
rect 50 -119 62 -85
rect 96 -119 108 -85
rect 50 -153 108 -119
rect 50 -187 62 -153
rect 96 -187 108 -153
rect 50 -221 108 -187
rect 50 -255 62 -221
rect 96 -255 108 -221
rect 50 -289 108 -255
rect 50 -323 62 -289
rect 96 -323 108 -289
rect 50 -357 108 -323
rect 50 -391 62 -357
rect 96 -391 108 -357
rect 50 -425 108 -391
rect 50 -459 62 -425
rect 96 -459 108 -425
rect 50 -500 108 -459
rect 208 459 266 500
rect 208 425 220 459
rect 254 425 266 459
rect 208 391 266 425
rect 208 357 220 391
rect 254 357 266 391
rect 208 323 266 357
rect 208 289 220 323
rect 254 289 266 323
rect 208 255 266 289
rect 208 221 220 255
rect 254 221 266 255
rect 208 187 266 221
rect 208 153 220 187
rect 254 153 266 187
rect 208 119 266 153
rect 208 85 220 119
rect 254 85 266 119
rect 208 51 266 85
rect 208 17 220 51
rect 254 17 266 51
rect 208 -17 266 17
rect 208 -51 220 -17
rect 254 -51 266 -17
rect 208 -85 266 -51
rect 208 -119 220 -85
rect 254 -119 266 -85
rect 208 -153 266 -119
rect 208 -187 220 -153
rect 254 -187 266 -153
rect 208 -221 266 -187
rect 208 -255 220 -221
rect 254 -255 266 -221
rect 208 -289 266 -255
rect 208 -323 220 -289
rect 254 -323 266 -289
rect 208 -357 266 -323
rect 208 -391 220 -357
rect 254 -391 266 -357
rect 208 -425 266 -391
rect 208 -459 220 -425
rect 254 -459 266 -425
rect 208 -500 266 -459
rect 366 459 424 500
rect 366 425 378 459
rect 412 425 424 459
rect 366 391 424 425
rect 366 357 378 391
rect 412 357 424 391
rect 366 323 424 357
rect 366 289 378 323
rect 412 289 424 323
rect 366 255 424 289
rect 366 221 378 255
rect 412 221 424 255
rect 366 187 424 221
rect 366 153 378 187
rect 412 153 424 187
rect 366 119 424 153
rect 366 85 378 119
rect 412 85 424 119
rect 366 51 424 85
rect 366 17 378 51
rect 412 17 424 51
rect 366 -17 424 17
rect 366 -51 378 -17
rect 412 -51 424 -17
rect 366 -85 424 -51
rect 366 -119 378 -85
rect 412 -119 424 -85
rect 366 -153 424 -119
rect 366 -187 378 -153
rect 412 -187 424 -153
rect 366 -221 424 -187
rect 366 -255 378 -221
rect 412 -255 424 -221
rect 366 -289 424 -255
rect 366 -323 378 -289
rect 412 -323 424 -289
rect 366 -357 424 -323
rect 366 -391 378 -357
rect 412 -391 424 -357
rect 366 -425 424 -391
rect 366 -459 378 -425
rect 412 -459 424 -425
rect 366 -500 424 -459
rect 524 459 582 500
rect 524 425 536 459
rect 570 425 582 459
rect 524 391 582 425
rect 524 357 536 391
rect 570 357 582 391
rect 524 323 582 357
rect 524 289 536 323
rect 570 289 582 323
rect 524 255 582 289
rect 524 221 536 255
rect 570 221 582 255
rect 524 187 582 221
rect 524 153 536 187
rect 570 153 582 187
rect 524 119 582 153
rect 524 85 536 119
rect 570 85 582 119
rect 524 51 582 85
rect 524 17 536 51
rect 570 17 582 51
rect 524 -17 582 17
rect 524 -51 536 -17
rect 570 -51 582 -17
rect 524 -85 582 -51
rect 524 -119 536 -85
rect 570 -119 582 -85
rect 524 -153 582 -119
rect 524 -187 536 -153
rect 570 -187 582 -153
rect 524 -221 582 -187
rect 524 -255 536 -221
rect 570 -255 582 -221
rect 524 -289 582 -255
rect 524 -323 536 -289
rect 570 -323 582 -289
rect 524 -357 582 -323
rect 524 -391 536 -357
rect 570 -391 582 -357
rect 524 -425 582 -391
rect 524 -459 536 -425
rect 570 -459 582 -425
rect 524 -500 582 -459
<< ndiffc >>
rect -570 425 -536 459
rect -570 357 -536 391
rect -570 289 -536 323
rect -570 221 -536 255
rect -570 153 -536 187
rect -570 85 -536 119
rect -570 17 -536 51
rect -570 -51 -536 -17
rect -570 -119 -536 -85
rect -570 -187 -536 -153
rect -570 -255 -536 -221
rect -570 -323 -536 -289
rect -570 -391 -536 -357
rect -570 -459 -536 -425
rect -412 425 -378 459
rect -412 357 -378 391
rect -412 289 -378 323
rect -412 221 -378 255
rect -412 153 -378 187
rect -412 85 -378 119
rect -412 17 -378 51
rect -412 -51 -378 -17
rect -412 -119 -378 -85
rect -412 -187 -378 -153
rect -412 -255 -378 -221
rect -412 -323 -378 -289
rect -412 -391 -378 -357
rect -412 -459 -378 -425
rect -254 425 -220 459
rect -254 357 -220 391
rect -254 289 -220 323
rect -254 221 -220 255
rect -254 153 -220 187
rect -254 85 -220 119
rect -254 17 -220 51
rect -254 -51 -220 -17
rect -254 -119 -220 -85
rect -254 -187 -220 -153
rect -254 -255 -220 -221
rect -254 -323 -220 -289
rect -254 -391 -220 -357
rect -254 -459 -220 -425
rect -96 425 -62 459
rect -96 357 -62 391
rect -96 289 -62 323
rect -96 221 -62 255
rect -96 153 -62 187
rect -96 85 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -85
rect -96 -187 -62 -153
rect -96 -255 -62 -221
rect -96 -323 -62 -289
rect -96 -391 -62 -357
rect -96 -459 -62 -425
rect 62 425 96 459
rect 62 357 96 391
rect 62 289 96 323
rect 62 221 96 255
rect 62 153 96 187
rect 62 85 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -85
rect 62 -187 96 -153
rect 62 -255 96 -221
rect 62 -323 96 -289
rect 62 -391 96 -357
rect 62 -459 96 -425
rect 220 425 254 459
rect 220 357 254 391
rect 220 289 254 323
rect 220 221 254 255
rect 220 153 254 187
rect 220 85 254 119
rect 220 17 254 51
rect 220 -51 254 -17
rect 220 -119 254 -85
rect 220 -187 254 -153
rect 220 -255 254 -221
rect 220 -323 254 -289
rect 220 -391 254 -357
rect 220 -459 254 -425
rect 378 425 412 459
rect 378 357 412 391
rect 378 289 412 323
rect 378 221 412 255
rect 378 153 412 187
rect 378 85 412 119
rect 378 17 412 51
rect 378 -51 412 -17
rect 378 -119 412 -85
rect 378 -187 412 -153
rect 378 -255 412 -221
rect 378 -323 412 -289
rect 378 -391 412 -357
rect 378 -459 412 -425
rect 536 425 570 459
rect 536 357 570 391
rect 536 289 570 323
rect 536 221 570 255
rect 536 153 570 187
rect 536 85 570 119
rect 536 17 570 51
rect 536 -51 570 -17
rect 536 -119 570 -85
rect 536 -187 570 -153
rect 536 -255 570 -221
rect 536 -323 570 -289
rect 536 -391 570 -357
rect 536 -459 570 -425
<< psubdiff >>
rect -684 640 -561 674
rect -527 640 -493 674
rect -459 640 -425 674
rect -391 640 -357 674
rect -323 640 -289 674
rect -255 640 -221 674
rect -187 640 -153 674
rect -119 640 -85 674
rect -51 640 -17 674
rect 17 640 51 674
rect 85 640 119 674
rect 153 640 187 674
rect 221 640 255 674
rect 289 640 323 674
rect 357 640 391 674
rect 425 640 459 674
rect 493 640 527 674
rect 561 640 684 674
rect -684 561 -650 640
rect -684 493 -650 527
rect 650 561 684 640
rect -684 425 -650 459
rect -684 357 -650 391
rect -684 289 -650 323
rect -684 221 -650 255
rect -684 153 -650 187
rect -684 85 -650 119
rect -684 17 -650 51
rect -684 -51 -650 -17
rect -684 -119 -650 -85
rect -684 -187 -650 -153
rect -684 -255 -650 -221
rect -684 -323 -650 -289
rect -684 -391 -650 -357
rect -684 -459 -650 -425
rect -684 -527 -650 -493
rect 650 493 684 527
rect 650 425 684 459
rect 650 357 684 391
rect 650 289 684 323
rect 650 221 684 255
rect 650 153 684 187
rect 650 85 684 119
rect 650 17 684 51
rect 650 -51 684 -17
rect 650 -119 684 -85
rect 650 -187 684 -153
rect 650 -255 684 -221
rect 650 -323 684 -289
rect 650 -391 684 -357
rect 650 -459 684 -425
rect -684 -640 -650 -561
rect 650 -527 684 -493
rect 650 -640 684 -561
rect -684 -674 -561 -640
rect -527 -674 -493 -640
rect -459 -674 -425 -640
rect -391 -674 -357 -640
rect -323 -674 -289 -640
rect -255 -674 -221 -640
rect -187 -674 -153 -640
rect -119 -674 -85 -640
rect -51 -674 -17 -640
rect 17 -674 51 -640
rect 85 -674 119 -640
rect 153 -674 187 -640
rect 221 -674 255 -640
rect 289 -674 323 -640
rect 357 -674 391 -640
rect 425 -674 459 -640
rect 493 -674 527 -640
rect 561 -674 684 -640
<< psubdiffcont >>
rect -561 640 -527 674
rect -493 640 -459 674
rect -425 640 -391 674
rect -357 640 -323 674
rect -289 640 -255 674
rect -221 640 -187 674
rect -153 640 -119 674
rect -85 640 -51 674
rect -17 640 17 674
rect 51 640 85 674
rect 119 640 153 674
rect 187 640 221 674
rect 255 640 289 674
rect 323 640 357 674
rect 391 640 425 674
rect 459 640 493 674
rect 527 640 561 674
rect -684 527 -650 561
rect 650 527 684 561
rect -684 459 -650 493
rect -684 391 -650 425
rect -684 323 -650 357
rect -684 255 -650 289
rect -684 187 -650 221
rect -684 119 -650 153
rect -684 51 -650 85
rect -684 -17 -650 17
rect -684 -85 -650 -51
rect -684 -153 -650 -119
rect -684 -221 -650 -187
rect -684 -289 -650 -255
rect -684 -357 -650 -323
rect -684 -425 -650 -391
rect -684 -493 -650 -459
rect 650 459 684 493
rect 650 391 684 425
rect 650 323 684 357
rect 650 255 684 289
rect 650 187 684 221
rect 650 119 684 153
rect 650 51 684 85
rect 650 -17 684 17
rect 650 -85 684 -51
rect 650 -153 684 -119
rect 650 -221 684 -187
rect 650 -289 684 -255
rect 650 -357 684 -323
rect 650 -425 684 -391
rect 650 -493 684 -459
rect -684 -561 -650 -527
rect 650 -561 684 -527
rect -561 -674 -527 -640
rect -493 -674 -459 -640
rect -425 -674 -391 -640
rect -357 -674 -323 -640
rect -289 -674 -255 -640
rect -221 -674 -187 -640
rect -153 -674 -119 -640
rect -85 -674 -51 -640
rect -17 -674 17 -640
rect 51 -674 85 -640
rect 119 -674 153 -640
rect 187 -674 221 -640
rect 255 -674 289 -640
rect 323 -674 357 -640
rect 391 -674 425 -640
rect 459 -674 493 -640
rect 527 -674 561 -640
<< poly >>
rect -524 572 -424 588
rect -524 538 -491 572
rect -457 538 -424 572
rect -524 500 -424 538
rect -366 572 -266 588
rect -366 538 -333 572
rect -299 538 -266 572
rect -366 500 -266 538
rect -208 572 -108 588
rect -208 538 -175 572
rect -141 538 -108 572
rect -208 500 -108 538
rect -50 572 50 588
rect -50 538 -17 572
rect 17 538 50 572
rect -50 500 50 538
rect 108 572 208 588
rect 108 538 141 572
rect 175 538 208 572
rect 108 500 208 538
rect 266 572 366 588
rect 266 538 299 572
rect 333 538 366 572
rect 266 500 366 538
rect 424 572 524 588
rect 424 538 457 572
rect 491 538 524 572
rect 424 500 524 538
rect -524 -538 -424 -500
rect -524 -572 -491 -538
rect -457 -572 -424 -538
rect -524 -588 -424 -572
rect -366 -538 -266 -500
rect -366 -572 -333 -538
rect -299 -572 -266 -538
rect -366 -588 -266 -572
rect -208 -538 -108 -500
rect -208 -572 -175 -538
rect -141 -572 -108 -538
rect -208 -588 -108 -572
rect -50 -538 50 -500
rect -50 -572 -17 -538
rect 17 -572 50 -538
rect -50 -588 50 -572
rect 108 -538 208 -500
rect 108 -572 141 -538
rect 175 -572 208 -538
rect 108 -588 208 -572
rect 266 -538 366 -500
rect 266 -572 299 -538
rect 333 -572 366 -538
rect 266 -588 366 -572
rect 424 -538 524 -500
rect 424 -572 457 -538
rect 491 -572 524 -538
rect 424 -588 524 -572
<< polycont >>
rect -491 538 -457 572
rect -333 538 -299 572
rect -175 538 -141 572
rect -17 538 17 572
rect 141 538 175 572
rect 299 538 333 572
rect 457 538 491 572
rect -491 -572 -457 -538
rect -333 -572 -299 -538
rect -175 -572 -141 -538
rect -17 -572 17 -538
rect 141 -572 175 -538
rect 299 -572 333 -538
rect 457 -572 491 -538
<< locali >>
rect -684 640 -561 674
rect -527 640 -493 674
rect -459 640 -425 674
rect -391 640 -357 674
rect -323 640 -305 674
rect -255 640 -233 674
rect -187 640 -161 674
rect -119 640 -89 674
rect -51 640 -17 674
rect 17 640 51 674
rect 89 640 119 674
rect 161 640 187 674
rect 233 640 255 674
rect 305 640 323 674
rect 357 640 391 674
rect 425 640 459 674
rect 493 640 527 674
rect 561 640 684 674
rect -684 561 -650 640
rect -524 538 -491 572
rect -457 538 -424 572
rect -366 538 -333 572
rect -299 538 -266 572
rect -208 538 -175 572
rect -141 538 -108 572
rect -50 538 -17 572
rect 17 538 50 572
rect 108 538 141 572
rect 175 538 208 572
rect 266 538 299 572
rect 333 538 366 572
rect 424 538 457 572
rect 491 538 524 572
rect 650 561 684 640
rect -684 493 -650 527
rect -684 425 -650 459
rect -684 357 -650 391
rect -684 289 -650 323
rect -684 221 -650 255
rect -684 153 -650 187
rect -684 85 -650 119
rect -684 17 -650 51
rect -684 -51 -650 -17
rect -684 -119 -650 -85
rect -684 -187 -650 -153
rect -684 -255 -650 -221
rect -684 -323 -650 -289
rect -684 -391 -650 -357
rect -684 -459 -650 -425
rect -684 -527 -650 -493
rect -570 485 -536 504
rect -570 413 -536 425
rect -570 341 -536 357
rect -570 269 -536 289
rect -570 197 -536 221
rect -570 125 -536 153
rect -570 53 -536 85
rect -570 -17 -536 17
rect -570 -85 -536 -53
rect -570 -153 -536 -125
rect -570 -221 -536 -197
rect -570 -289 -536 -269
rect -570 -357 -536 -341
rect -570 -425 -536 -413
rect -570 -504 -536 -485
rect -412 485 -378 504
rect -412 413 -378 425
rect -412 341 -378 357
rect -412 269 -378 289
rect -412 197 -378 221
rect -412 125 -378 153
rect -412 53 -378 85
rect -412 -17 -378 17
rect -412 -85 -378 -53
rect -412 -153 -378 -125
rect -412 -221 -378 -197
rect -412 -289 -378 -269
rect -412 -357 -378 -341
rect -412 -425 -378 -413
rect -412 -504 -378 -485
rect -254 485 -220 504
rect -254 413 -220 425
rect -254 341 -220 357
rect -254 269 -220 289
rect -254 197 -220 221
rect -254 125 -220 153
rect -254 53 -220 85
rect -254 -17 -220 17
rect -254 -85 -220 -53
rect -254 -153 -220 -125
rect -254 -221 -220 -197
rect -254 -289 -220 -269
rect -254 -357 -220 -341
rect -254 -425 -220 -413
rect -254 -504 -220 -485
rect -96 485 -62 504
rect -96 413 -62 425
rect -96 341 -62 357
rect -96 269 -62 289
rect -96 197 -62 221
rect -96 125 -62 153
rect -96 53 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -53
rect -96 -153 -62 -125
rect -96 -221 -62 -197
rect -96 -289 -62 -269
rect -96 -357 -62 -341
rect -96 -425 -62 -413
rect -96 -504 -62 -485
rect 62 485 96 504
rect 62 413 96 425
rect 62 341 96 357
rect 62 269 96 289
rect 62 197 96 221
rect 62 125 96 153
rect 62 53 96 85
rect 62 -17 96 17
rect 62 -85 96 -53
rect 62 -153 96 -125
rect 62 -221 96 -197
rect 62 -289 96 -269
rect 62 -357 96 -341
rect 62 -425 96 -413
rect 62 -504 96 -485
rect 220 485 254 504
rect 220 413 254 425
rect 220 341 254 357
rect 220 269 254 289
rect 220 197 254 221
rect 220 125 254 153
rect 220 53 254 85
rect 220 -17 254 17
rect 220 -85 254 -53
rect 220 -153 254 -125
rect 220 -221 254 -197
rect 220 -289 254 -269
rect 220 -357 254 -341
rect 220 -425 254 -413
rect 220 -504 254 -485
rect 378 485 412 504
rect 378 413 412 425
rect 378 341 412 357
rect 378 269 412 289
rect 378 197 412 221
rect 378 125 412 153
rect 378 53 412 85
rect 378 -17 412 17
rect 378 -85 412 -53
rect 378 -153 412 -125
rect 378 -221 412 -197
rect 378 -289 412 -269
rect 378 -357 412 -341
rect 378 -425 412 -413
rect 378 -504 412 -485
rect 536 485 570 504
rect 536 413 570 425
rect 536 341 570 357
rect 536 269 570 289
rect 536 197 570 221
rect 536 125 570 153
rect 536 53 570 85
rect 536 -17 570 17
rect 536 -85 570 -53
rect 536 -153 570 -125
rect 536 -221 570 -197
rect 536 -289 570 -269
rect 536 -357 570 -341
rect 536 -425 570 -413
rect 536 -504 570 -485
rect 650 493 684 527
rect 650 425 684 459
rect 650 357 684 391
rect 650 289 684 323
rect 650 221 684 255
rect 650 153 684 187
rect 650 85 684 119
rect 650 17 684 51
rect 650 -51 684 -17
rect 650 -119 684 -85
rect 650 -187 684 -153
rect 650 -255 684 -221
rect 650 -323 684 -289
rect 650 -391 684 -357
rect 650 -459 684 -425
rect 650 -527 684 -493
rect -684 -640 -650 -561
rect -524 -572 -491 -538
rect -457 -572 -424 -538
rect -366 -572 -333 -538
rect -299 -572 -266 -538
rect -208 -572 -175 -538
rect -141 -572 -108 -538
rect -50 -572 -17 -538
rect 17 -572 50 -538
rect 108 -572 141 -538
rect 175 -572 208 -538
rect 266 -572 299 -538
rect 333 -572 366 -538
rect 424 -572 457 -538
rect 491 -572 524 -538
rect 650 -640 684 -561
rect -684 -674 -561 -640
rect -527 -674 -493 -640
rect -459 -674 -425 -640
rect -391 -674 -357 -640
rect -323 -674 -305 -640
rect -255 -674 -233 -640
rect -187 -674 -161 -640
rect -119 -674 -89 -640
rect -51 -674 -17 -640
rect 17 -674 51 -640
rect 89 -674 119 -640
rect 161 -674 187 -640
rect 233 -674 255 -640
rect 305 -674 323 -640
rect 357 -674 391 -640
rect 425 -674 459 -640
rect 493 -674 527 -640
rect 561 -674 684 -640
<< viali >>
rect -305 640 -289 674
rect -289 640 -271 674
rect -233 640 -221 674
rect -221 640 -199 674
rect -161 640 -153 674
rect -153 640 -127 674
rect -89 640 -85 674
rect -85 640 -55 674
rect -17 640 17 674
rect 55 640 85 674
rect 85 640 89 674
rect 127 640 153 674
rect 153 640 161 674
rect 199 640 221 674
rect 221 640 233 674
rect 271 640 289 674
rect 289 640 305 674
rect -491 538 -457 572
rect -333 538 -299 572
rect -175 538 -141 572
rect -17 538 17 572
rect 141 538 175 572
rect 299 538 333 572
rect 457 538 491 572
rect -570 459 -536 485
rect -570 451 -536 459
rect -570 391 -536 413
rect -570 379 -536 391
rect -570 323 -536 341
rect -570 307 -536 323
rect -570 255 -536 269
rect -570 235 -536 255
rect -570 187 -536 197
rect -570 163 -536 187
rect -570 119 -536 125
rect -570 91 -536 119
rect -570 51 -536 53
rect -570 19 -536 51
rect -570 -51 -536 -19
rect -570 -53 -536 -51
rect -570 -119 -536 -91
rect -570 -125 -536 -119
rect -570 -187 -536 -163
rect -570 -197 -536 -187
rect -570 -255 -536 -235
rect -570 -269 -536 -255
rect -570 -323 -536 -307
rect -570 -341 -536 -323
rect -570 -391 -536 -379
rect -570 -413 -536 -391
rect -570 -459 -536 -451
rect -570 -485 -536 -459
rect -412 459 -378 485
rect -412 451 -378 459
rect -412 391 -378 413
rect -412 379 -378 391
rect -412 323 -378 341
rect -412 307 -378 323
rect -412 255 -378 269
rect -412 235 -378 255
rect -412 187 -378 197
rect -412 163 -378 187
rect -412 119 -378 125
rect -412 91 -378 119
rect -412 51 -378 53
rect -412 19 -378 51
rect -412 -51 -378 -19
rect -412 -53 -378 -51
rect -412 -119 -378 -91
rect -412 -125 -378 -119
rect -412 -187 -378 -163
rect -412 -197 -378 -187
rect -412 -255 -378 -235
rect -412 -269 -378 -255
rect -412 -323 -378 -307
rect -412 -341 -378 -323
rect -412 -391 -378 -379
rect -412 -413 -378 -391
rect -412 -459 -378 -451
rect -412 -485 -378 -459
rect -254 459 -220 485
rect -254 451 -220 459
rect -254 391 -220 413
rect -254 379 -220 391
rect -254 323 -220 341
rect -254 307 -220 323
rect -254 255 -220 269
rect -254 235 -220 255
rect -254 187 -220 197
rect -254 163 -220 187
rect -254 119 -220 125
rect -254 91 -220 119
rect -254 51 -220 53
rect -254 19 -220 51
rect -254 -51 -220 -19
rect -254 -53 -220 -51
rect -254 -119 -220 -91
rect -254 -125 -220 -119
rect -254 -187 -220 -163
rect -254 -197 -220 -187
rect -254 -255 -220 -235
rect -254 -269 -220 -255
rect -254 -323 -220 -307
rect -254 -341 -220 -323
rect -254 -391 -220 -379
rect -254 -413 -220 -391
rect -254 -459 -220 -451
rect -254 -485 -220 -459
rect -96 459 -62 485
rect -96 451 -62 459
rect -96 391 -62 413
rect -96 379 -62 391
rect -96 323 -62 341
rect -96 307 -62 323
rect -96 255 -62 269
rect -96 235 -62 255
rect -96 187 -62 197
rect -96 163 -62 187
rect -96 119 -62 125
rect -96 91 -62 119
rect -96 51 -62 53
rect -96 19 -62 51
rect -96 -51 -62 -19
rect -96 -53 -62 -51
rect -96 -119 -62 -91
rect -96 -125 -62 -119
rect -96 -187 -62 -163
rect -96 -197 -62 -187
rect -96 -255 -62 -235
rect -96 -269 -62 -255
rect -96 -323 -62 -307
rect -96 -341 -62 -323
rect -96 -391 -62 -379
rect -96 -413 -62 -391
rect -96 -459 -62 -451
rect -96 -485 -62 -459
rect 62 459 96 485
rect 62 451 96 459
rect 62 391 96 413
rect 62 379 96 391
rect 62 323 96 341
rect 62 307 96 323
rect 62 255 96 269
rect 62 235 96 255
rect 62 187 96 197
rect 62 163 96 187
rect 62 119 96 125
rect 62 91 96 119
rect 62 51 96 53
rect 62 19 96 51
rect 62 -51 96 -19
rect 62 -53 96 -51
rect 62 -119 96 -91
rect 62 -125 96 -119
rect 62 -187 96 -163
rect 62 -197 96 -187
rect 62 -255 96 -235
rect 62 -269 96 -255
rect 62 -323 96 -307
rect 62 -341 96 -323
rect 62 -391 96 -379
rect 62 -413 96 -391
rect 62 -459 96 -451
rect 62 -485 96 -459
rect 220 459 254 485
rect 220 451 254 459
rect 220 391 254 413
rect 220 379 254 391
rect 220 323 254 341
rect 220 307 254 323
rect 220 255 254 269
rect 220 235 254 255
rect 220 187 254 197
rect 220 163 254 187
rect 220 119 254 125
rect 220 91 254 119
rect 220 51 254 53
rect 220 19 254 51
rect 220 -51 254 -19
rect 220 -53 254 -51
rect 220 -119 254 -91
rect 220 -125 254 -119
rect 220 -187 254 -163
rect 220 -197 254 -187
rect 220 -255 254 -235
rect 220 -269 254 -255
rect 220 -323 254 -307
rect 220 -341 254 -323
rect 220 -391 254 -379
rect 220 -413 254 -391
rect 220 -459 254 -451
rect 220 -485 254 -459
rect 378 459 412 485
rect 378 451 412 459
rect 378 391 412 413
rect 378 379 412 391
rect 378 323 412 341
rect 378 307 412 323
rect 378 255 412 269
rect 378 235 412 255
rect 378 187 412 197
rect 378 163 412 187
rect 378 119 412 125
rect 378 91 412 119
rect 378 51 412 53
rect 378 19 412 51
rect 378 -51 412 -19
rect 378 -53 412 -51
rect 378 -119 412 -91
rect 378 -125 412 -119
rect 378 -187 412 -163
rect 378 -197 412 -187
rect 378 -255 412 -235
rect 378 -269 412 -255
rect 378 -323 412 -307
rect 378 -341 412 -323
rect 378 -391 412 -379
rect 378 -413 412 -391
rect 378 -459 412 -451
rect 378 -485 412 -459
rect 536 459 570 485
rect 536 451 570 459
rect 536 391 570 413
rect 536 379 570 391
rect 536 323 570 341
rect 536 307 570 323
rect 536 255 570 269
rect 536 235 570 255
rect 536 187 570 197
rect 536 163 570 187
rect 536 119 570 125
rect 536 91 570 119
rect 536 51 570 53
rect 536 19 570 51
rect 536 -51 570 -19
rect 536 -53 570 -51
rect 536 -119 570 -91
rect 536 -125 570 -119
rect 536 -187 570 -163
rect 536 -197 570 -187
rect 536 -255 570 -235
rect 536 -269 570 -255
rect 536 -323 570 -307
rect 536 -341 570 -323
rect 536 -391 570 -379
rect 536 -413 570 -391
rect 536 -459 570 -451
rect 536 -485 570 -459
rect -491 -572 -457 -538
rect -333 -572 -299 -538
rect -175 -572 -141 -538
rect -17 -572 17 -538
rect 141 -572 175 -538
rect 299 -572 333 -538
rect 457 -572 491 -538
rect -305 -674 -289 -640
rect -289 -674 -271 -640
rect -233 -674 -221 -640
rect -221 -674 -199 -640
rect -161 -674 -153 -640
rect -153 -674 -127 -640
rect -89 -674 -85 -640
rect -85 -674 -55 -640
rect -17 -674 17 -640
rect 55 -674 85 -640
rect 85 -674 89 -640
rect 127 -674 153 -640
rect 153 -674 161 -640
rect 199 -674 221 -640
rect 221 -674 233 -640
rect 271 -674 289 -640
rect 289 -674 305 -640
<< metal1 >>
rect -337 674 337 680
rect -337 640 -305 674
rect -271 640 -233 674
rect -199 640 -161 674
rect -127 640 -89 674
rect -55 640 -17 674
rect 17 640 55 674
rect 89 640 127 674
rect 161 640 199 674
rect 233 640 271 674
rect 305 640 337 674
rect -337 634 337 640
rect -520 572 -428 578
rect -520 538 -491 572
rect -457 538 -428 572
rect -520 532 -428 538
rect -362 572 -270 578
rect -362 538 -333 572
rect -299 538 -270 572
rect -362 532 -270 538
rect -204 572 -112 578
rect -204 538 -175 572
rect -141 538 -112 572
rect -204 532 -112 538
rect -46 572 46 578
rect -46 538 -17 572
rect 17 538 46 572
rect -46 532 46 538
rect 112 572 204 578
rect 112 538 141 572
rect 175 538 204 572
rect 112 532 204 538
rect 270 572 362 578
rect 270 538 299 572
rect 333 538 362 572
rect 270 532 362 538
rect 428 572 520 578
rect 428 538 457 572
rect 491 538 520 572
rect 428 532 520 538
rect -576 485 -530 500
rect -576 451 -570 485
rect -536 451 -530 485
rect -576 413 -530 451
rect -576 379 -570 413
rect -536 379 -530 413
rect -576 341 -530 379
rect -576 307 -570 341
rect -536 307 -530 341
rect -576 269 -530 307
rect -576 235 -570 269
rect -536 235 -530 269
rect -576 197 -530 235
rect -576 163 -570 197
rect -536 163 -530 197
rect -576 125 -530 163
rect -576 91 -570 125
rect -536 91 -530 125
rect -576 53 -530 91
rect -576 19 -570 53
rect -536 19 -530 53
rect -576 -19 -530 19
rect -576 -53 -570 -19
rect -536 -53 -530 -19
rect -576 -91 -530 -53
rect -576 -125 -570 -91
rect -536 -125 -530 -91
rect -576 -163 -530 -125
rect -576 -197 -570 -163
rect -536 -197 -530 -163
rect -576 -235 -530 -197
rect -576 -269 -570 -235
rect -536 -269 -530 -235
rect -576 -307 -530 -269
rect -576 -341 -570 -307
rect -536 -341 -530 -307
rect -576 -379 -530 -341
rect -576 -413 -570 -379
rect -536 -413 -530 -379
rect -576 -451 -530 -413
rect -576 -485 -570 -451
rect -536 -485 -530 -451
rect -576 -500 -530 -485
rect -418 485 -372 500
rect -418 451 -412 485
rect -378 451 -372 485
rect -418 413 -372 451
rect -418 379 -412 413
rect -378 379 -372 413
rect -418 341 -372 379
rect -418 307 -412 341
rect -378 307 -372 341
rect -418 269 -372 307
rect -418 235 -412 269
rect -378 235 -372 269
rect -418 197 -372 235
rect -418 163 -412 197
rect -378 163 -372 197
rect -418 125 -372 163
rect -418 91 -412 125
rect -378 91 -372 125
rect -418 53 -372 91
rect -418 19 -412 53
rect -378 19 -372 53
rect -418 -19 -372 19
rect -418 -53 -412 -19
rect -378 -53 -372 -19
rect -418 -91 -372 -53
rect -418 -125 -412 -91
rect -378 -125 -372 -91
rect -418 -163 -372 -125
rect -418 -197 -412 -163
rect -378 -197 -372 -163
rect -418 -235 -372 -197
rect -418 -269 -412 -235
rect -378 -269 -372 -235
rect -418 -307 -372 -269
rect -418 -341 -412 -307
rect -378 -341 -372 -307
rect -418 -379 -372 -341
rect -418 -413 -412 -379
rect -378 -413 -372 -379
rect -418 -451 -372 -413
rect -418 -485 -412 -451
rect -378 -485 -372 -451
rect -418 -500 -372 -485
rect -260 485 -214 500
rect -260 451 -254 485
rect -220 451 -214 485
rect -260 413 -214 451
rect -260 379 -254 413
rect -220 379 -214 413
rect -260 341 -214 379
rect -260 307 -254 341
rect -220 307 -214 341
rect -260 269 -214 307
rect -260 235 -254 269
rect -220 235 -214 269
rect -260 197 -214 235
rect -260 163 -254 197
rect -220 163 -214 197
rect -260 125 -214 163
rect -260 91 -254 125
rect -220 91 -214 125
rect -260 53 -214 91
rect -260 19 -254 53
rect -220 19 -214 53
rect -260 -19 -214 19
rect -260 -53 -254 -19
rect -220 -53 -214 -19
rect -260 -91 -214 -53
rect -260 -125 -254 -91
rect -220 -125 -214 -91
rect -260 -163 -214 -125
rect -260 -197 -254 -163
rect -220 -197 -214 -163
rect -260 -235 -214 -197
rect -260 -269 -254 -235
rect -220 -269 -214 -235
rect -260 -307 -214 -269
rect -260 -341 -254 -307
rect -220 -341 -214 -307
rect -260 -379 -214 -341
rect -260 -413 -254 -379
rect -220 -413 -214 -379
rect -260 -451 -214 -413
rect -260 -485 -254 -451
rect -220 -485 -214 -451
rect -260 -500 -214 -485
rect -102 485 -56 500
rect -102 451 -96 485
rect -62 451 -56 485
rect -102 413 -56 451
rect -102 379 -96 413
rect -62 379 -56 413
rect -102 341 -56 379
rect -102 307 -96 341
rect -62 307 -56 341
rect -102 269 -56 307
rect -102 235 -96 269
rect -62 235 -56 269
rect -102 197 -56 235
rect -102 163 -96 197
rect -62 163 -56 197
rect -102 125 -56 163
rect -102 91 -96 125
rect -62 91 -56 125
rect -102 53 -56 91
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -91 -56 -53
rect -102 -125 -96 -91
rect -62 -125 -56 -91
rect -102 -163 -56 -125
rect -102 -197 -96 -163
rect -62 -197 -56 -163
rect -102 -235 -56 -197
rect -102 -269 -96 -235
rect -62 -269 -56 -235
rect -102 -307 -56 -269
rect -102 -341 -96 -307
rect -62 -341 -56 -307
rect -102 -379 -56 -341
rect -102 -413 -96 -379
rect -62 -413 -56 -379
rect -102 -451 -56 -413
rect -102 -485 -96 -451
rect -62 -485 -56 -451
rect -102 -500 -56 -485
rect 56 485 102 500
rect 56 451 62 485
rect 96 451 102 485
rect 56 413 102 451
rect 56 379 62 413
rect 96 379 102 413
rect 56 341 102 379
rect 56 307 62 341
rect 96 307 102 341
rect 56 269 102 307
rect 56 235 62 269
rect 96 235 102 269
rect 56 197 102 235
rect 56 163 62 197
rect 96 163 102 197
rect 56 125 102 163
rect 56 91 62 125
rect 96 91 102 125
rect 56 53 102 91
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -91 102 -53
rect 56 -125 62 -91
rect 96 -125 102 -91
rect 56 -163 102 -125
rect 56 -197 62 -163
rect 96 -197 102 -163
rect 56 -235 102 -197
rect 56 -269 62 -235
rect 96 -269 102 -235
rect 56 -307 102 -269
rect 56 -341 62 -307
rect 96 -341 102 -307
rect 56 -379 102 -341
rect 56 -413 62 -379
rect 96 -413 102 -379
rect 56 -451 102 -413
rect 56 -485 62 -451
rect 96 -485 102 -451
rect 56 -500 102 -485
rect 214 485 260 500
rect 214 451 220 485
rect 254 451 260 485
rect 214 413 260 451
rect 214 379 220 413
rect 254 379 260 413
rect 214 341 260 379
rect 214 307 220 341
rect 254 307 260 341
rect 214 269 260 307
rect 214 235 220 269
rect 254 235 260 269
rect 214 197 260 235
rect 214 163 220 197
rect 254 163 260 197
rect 214 125 260 163
rect 214 91 220 125
rect 254 91 260 125
rect 214 53 260 91
rect 214 19 220 53
rect 254 19 260 53
rect 214 -19 260 19
rect 214 -53 220 -19
rect 254 -53 260 -19
rect 214 -91 260 -53
rect 214 -125 220 -91
rect 254 -125 260 -91
rect 214 -163 260 -125
rect 214 -197 220 -163
rect 254 -197 260 -163
rect 214 -235 260 -197
rect 214 -269 220 -235
rect 254 -269 260 -235
rect 214 -307 260 -269
rect 214 -341 220 -307
rect 254 -341 260 -307
rect 214 -379 260 -341
rect 214 -413 220 -379
rect 254 -413 260 -379
rect 214 -451 260 -413
rect 214 -485 220 -451
rect 254 -485 260 -451
rect 214 -500 260 -485
rect 372 485 418 500
rect 372 451 378 485
rect 412 451 418 485
rect 372 413 418 451
rect 372 379 378 413
rect 412 379 418 413
rect 372 341 418 379
rect 372 307 378 341
rect 412 307 418 341
rect 372 269 418 307
rect 372 235 378 269
rect 412 235 418 269
rect 372 197 418 235
rect 372 163 378 197
rect 412 163 418 197
rect 372 125 418 163
rect 372 91 378 125
rect 412 91 418 125
rect 372 53 418 91
rect 372 19 378 53
rect 412 19 418 53
rect 372 -19 418 19
rect 372 -53 378 -19
rect 412 -53 418 -19
rect 372 -91 418 -53
rect 372 -125 378 -91
rect 412 -125 418 -91
rect 372 -163 418 -125
rect 372 -197 378 -163
rect 412 -197 418 -163
rect 372 -235 418 -197
rect 372 -269 378 -235
rect 412 -269 418 -235
rect 372 -307 418 -269
rect 372 -341 378 -307
rect 412 -341 418 -307
rect 372 -379 418 -341
rect 372 -413 378 -379
rect 412 -413 418 -379
rect 372 -451 418 -413
rect 372 -485 378 -451
rect 412 -485 418 -451
rect 372 -500 418 -485
rect 530 485 576 500
rect 530 451 536 485
rect 570 451 576 485
rect 530 413 576 451
rect 530 379 536 413
rect 570 379 576 413
rect 530 341 576 379
rect 530 307 536 341
rect 570 307 576 341
rect 530 269 576 307
rect 530 235 536 269
rect 570 235 576 269
rect 530 197 576 235
rect 530 163 536 197
rect 570 163 576 197
rect 530 125 576 163
rect 530 91 536 125
rect 570 91 576 125
rect 530 53 576 91
rect 530 19 536 53
rect 570 19 576 53
rect 530 -19 576 19
rect 530 -53 536 -19
rect 570 -53 576 -19
rect 530 -91 576 -53
rect 530 -125 536 -91
rect 570 -125 576 -91
rect 530 -163 576 -125
rect 530 -197 536 -163
rect 570 -197 576 -163
rect 530 -235 576 -197
rect 530 -269 536 -235
rect 570 -269 576 -235
rect 530 -307 576 -269
rect 530 -341 536 -307
rect 570 -341 576 -307
rect 530 -379 576 -341
rect 530 -413 536 -379
rect 570 -413 576 -379
rect 530 -451 576 -413
rect 530 -485 536 -451
rect 570 -485 576 -451
rect 530 -500 576 -485
rect -520 -538 -428 -532
rect -520 -572 -491 -538
rect -457 -572 -428 -538
rect -520 -578 -428 -572
rect -362 -538 -270 -532
rect -362 -572 -333 -538
rect -299 -572 -270 -538
rect -362 -578 -270 -572
rect -204 -538 -112 -532
rect -204 -572 -175 -538
rect -141 -572 -112 -538
rect -204 -578 -112 -572
rect -46 -538 46 -532
rect -46 -572 -17 -538
rect 17 -572 46 -538
rect -46 -578 46 -572
rect 112 -538 204 -532
rect 112 -572 141 -538
rect 175 -572 204 -538
rect 112 -578 204 -572
rect 270 -538 362 -532
rect 270 -572 299 -538
rect 333 -572 362 -538
rect 270 -578 362 -572
rect 428 -538 520 -532
rect 428 -572 457 -538
rect 491 -572 520 -538
rect 428 -578 520 -572
rect -337 -640 337 -634
rect -337 -674 -305 -640
rect -271 -674 -233 -640
rect -199 -674 -161 -640
rect -127 -674 -89 -640
rect -55 -674 -17 -640
rect 17 -674 55 -640
rect 89 -674 127 -640
rect 161 -674 199 -640
rect 233 -674 271 -640
rect 305 -674 337 -640
rect -337 -680 337 -674
<< properties >>
string FIXED_BBOX -667 -657 667 657
<< end >>
