magic
tech sky130A
magscale 1 2
timestamp 1709390584
<< metal3 >>
rect -1786 6892 1786 6920
rect -1786 3668 1702 6892
rect 1766 3668 1786 6892
rect -1786 3640 1786 3668
rect -1786 3372 1786 3400
rect -1786 148 1702 3372
rect 1766 148 1786 3372
rect -1786 120 1786 148
rect -1786 -148 1786 -120
rect -1786 -3372 1702 -148
rect 1766 -3372 1786 -148
rect -1786 -3400 1786 -3372
rect -1786 -3668 1786 -3640
rect -1786 -6892 1702 -3668
rect 1766 -6892 1786 -3668
rect -1786 -6920 1786 -6892
<< via3 >>
rect 1702 3668 1766 6892
rect 1702 148 1766 3372
rect 1702 -3372 1766 -148
rect 1702 -6892 1766 -3668
<< mimcap >>
rect -1746 6840 1454 6880
rect -1746 3720 -1706 6840
rect 1414 3720 1454 6840
rect -1746 3680 1454 3720
rect -1746 3320 1454 3360
rect -1746 200 -1706 3320
rect 1414 200 1454 3320
rect -1746 160 1454 200
rect -1746 -200 1454 -160
rect -1746 -3320 -1706 -200
rect 1414 -3320 1454 -200
rect -1746 -3360 1454 -3320
rect -1746 -3720 1454 -3680
rect -1746 -6840 -1706 -3720
rect 1414 -6840 1454 -3720
rect -1746 -6880 1454 -6840
<< mimcapcontact >>
rect -1706 3720 1414 6840
rect -1706 200 1414 3320
rect -1706 -3320 1414 -200
rect -1706 -6840 1414 -3720
<< metal4 >>
rect -198 6841 -94 7040
rect 1682 6892 1786 7040
rect -1707 6840 1415 6841
rect -1707 3720 -1706 6840
rect 1414 3720 1415 6840
rect -1707 3719 1415 3720
rect -198 3321 -94 3719
rect 1682 3668 1702 6892
rect 1766 3668 1786 6892
rect 1682 3372 1786 3668
rect -1707 3320 1415 3321
rect -1707 200 -1706 3320
rect 1414 200 1415 3320
rect -1707 199 1415 200
rect -198 -199 -94 199
rect 1682 148 1702 3372
rect 1766 148 1786 3372
rect 1682 -148 1786 148
rect -1707 -200 1415 -199
rect -1707 -3320 -1706 -200
rect 1414 -3320 1415 -200
rect -1707 -3321 1415 -3320
rect -198 -3719 -94 -3321
rect 1682 -3372 1702 -148
rect 1766 -3372 1786 -148
rect 1682 -3668 1786 -3372
rect -1707 -3720 1415 -3719
rect -1707 -6840 -1706 -3720
rect 1414 -6840 1415 -3720
rect -1707 -6841 1415 -6840
rect -198 -7040 -94 -6841
rect 1682 -6892 1702 -3668
rect 1766 -6892 1786 -3668
rect 1682 -7040 1786 -6892
<< properties >>
string FIXED_BBOX -1786 3640 1494 6920
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16.0 l 16.0 val 524.159 carea 2.00 cperi 0.19 nx 1 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
