magic
tech sky130A
magscale 1 2
timestamp 1715652275
<< error_p >>
rect -29 281 29 287
rect -29 247 -17 281
rect -29 241 29 247
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect -29 -287 29 -281
<< nwell >>
rect -226 -419 226 419
<< pmos >>
rect -30 -200 30 200
<< pdiff >>
rect -88 188 -30 200
rect -88 -188 -76 188
rect -42 -188 -30 188
rect -88 -200 -30 -188
rect 30 188 88 200
rect 30 -188 42 188
rect 76 -188 88 188
rect 30 -200 88 -188
<< pdiffc >>
rect -76 -188 -42 188
rect 42 -188 76 188
<< nsubdiff >>
rect -190 349 190 383
rect -190 287 -156 349
rect 156 287 190 349
rect -190 -349 -156 -287
rect 156 -349 190 -287
rect -190 -383 -94 -349
rect 94 -383 190 -349
<< nsubdiffcont >>
rect -190 -287 -156 287
rect 156 -287 190 287
rect -94 -383 94 -349
<< poly >>
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect -30 200 30 231
rect -30 -231 30 -200
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
<< polycont >>
rect -17 247 17 281
rect -17 -281 17 -247
<< locali >>
rect -190 349 190 383
rect -190 287 -156 349
rect 156 287 190 349
rect -33 247 -17 281
rect 17 247 33 281
rect -76 188 -42 204
rect -76 -204 -42 -188
rect 42 188 76 204
rect 42 -204 76 -188
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -190 -349 -156 -287
rect 156 -349 190 -287
rect -190 -383 -94 -349
rect 94 -383 190 -349
<< viali >>
rect -17 247 17 281
rect -76 -188 -42 188
rect 42 -188 76 188
rect -17 -281 17 -247
<< metal1 >>
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect -82 188 -36 200
rect -82 -188 -76 188
rect -42 -188 -36 188
rect -82 -200 -36 -188
rect 36 188 82 200
rect 36 -188 42 188
rect 76 -188 82 188
rect 36 -200 82 -188
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
<< properties >>
string FIXED_BBOX -173 -366 173 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2. l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
