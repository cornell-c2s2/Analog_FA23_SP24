magic
tech sky130A
magscale 1 2
timestamp 1712787074
<< nwell >>
rect -1630 -250 2190 180
rect 450 -450 2190 -250
rect 450 -490 590 -450
rect 630 -490 2190 -450
rect 450 -510 2190 -490
rect 450 -1770 2190 -1120
rect 440 -3010 2190 -2360
rect 450 -4020 2190 -3610
rect 450 -4026 1310 -4020
rect 450 -4030 1134 -4026
rect 1160 -4030 1240 -4026
rect 1258 -4030 1310 -4026
rect 1430 -4030 2190 -4020
rect 450 -4170 2190 -4030
rect 450 -4230 1060 -4170
rect 450 -4250 660 -4230
rect 740 -4250 1060 -4230
rect 1130 -4250 2190 -4170
rect 1158 -4251 1540 -4250
rect 440 -5490 2190 -4840
rect 440 -6730 2190 -6070
<< pwell >>
rect -1600 230 170 500
rect 250 -1020 1940 -570
rect 250 -2280 1500 -1830
rect 250 -3550 940 -3070
rect 250 -4310 660 -4300
rect 740 -4310 1150 -4300
rect 1220 -4310 1250 -4300
rect 1390 -4310 1430 -4300
rect 1510 -4310 1690 -4300
rect 250 -4790 1790 -4310
rect 250 -6030 1140 -5530
rect 250 -6970 1970 -6760
<< pdiff >>
rect 630 -460 660 -450
rect 690 -460 730 -450
<< psubdiff >>
rect 20 460 130 480
rect 20 410 50 460
rect 100 410 130 460
rect 20 340 130 410
rect 20 290 50 340
rect 100 290 130 340
rect 20 260 130 290
rect 330 -660 450 -630
rect 330 -720 360 -660
rect 420 -720 450 -660
rect 330 -750 450 -720
rect 330 -860 450 -830
rect 330 -920 360 -860
rect 420 -920 450 -860
rect 330 -950 450 -920
rect 310 -1900 430 -1870
rect 310 -1960 340 -1900
rect 400 -1960 430 -1900
rect 310 -1990 430 -1960
rect 310 -2150 430 -2120
rect 310 -2210 340 -2150
rect 400 -2210 430 -2150
rect 310 -2240 430 -2210
rect 330 -3160 450 -3130
rect 330 -3220 360 -3160
rect 420 -3220 450 -3160
rect 330 -3330 450 -3220
rect 330 -3390 360 -3330
rect 420 -3390 450 -3330
rect 330 -3420 450 -3390
rect 320 -4410 440 -4380
rect 320 -4470 350 -4410
rect 410 -4470 440 -4410
rect 320 -4500 440 -4470
rect 320 -4590 440 -4560
rect 320 -4650 350 -4590
rect 410 -4650 440 -4590
rect 320 -4680 440 -4650
rect 310 -5580 430 -5550
rect 310 -5640 340 -5580
rect 400 -5640 430 -5580
rect 310 -5670 430 -5640
rect 310 -5830 430 -5800
rect 310 -5890 340 -5830
rect 400 -5890 430 -5830
rect 310 -5920 430 -5890
rect 300 -6830 420 -6800
rect 300 -6890 330 -6830
rect 390 -6890 420 -6830
rect 300 -6920 420 -6890
<< nsubdiff >>
rect -160 0 -50 30
rect -160 -50 -130 0
rect -80 -50 -50 0
rect -160 -130 -50 -50
rect -160 -180 -130 -130
rect -80 -180 -50 -130
rect -160 -210 -50 -180
rect 1160 -1420 1270 -1390
rect 1160 -1470 1190 -1420
rect 1240 -1470 1270 -1420
rect 1160 -1500 1270 -1470
rect 1470 -1420 1580 -1390
rect 1470 -1470 1500 -1420
rect 1550 -1470 1580 -1420
rect 1470 -1500 1580 -1470
rect 1710 -1420 1820 -1390
rect 1710 -1470 1740 -1420
rect 1790 -1470 1820 -1420
rect 1710 -1500 1820 -1470
rect 1970 -1420 2080 -1390
rect 1970 -1470 2000 -1420
rect 2050 -1470 2080 -1420
rect 1970 -1500 2080 -1470
rect 1540 -2660 1650 -2630
rect 1540 -2710 1570 -2660
rect 1620 -2710 1650 -2660
rect 1540 -2740 1650 -2710
rect 1760 -2660 1870 -2630
rect 1760 -2710 1790 -2660
rect 1840 -2710 1870 -2660
rect 1760 -2740 1870 -2710
rect 2000 -2660 2110 -2630
rect 2000 -2710 2030 -2660
rect 2080 -2710 2110 -2660
rect 2000 -2740 2110 -2710
rect 1850 -3910 1960 -3880
rect 1850 -3960 1880 -3910
rect 1930 -3960 1960 -3910
rect 1850 -3990 1960 -3960
rect 2040 -3910 2150 -3880
rect 2040 -3960 2070 -3910
rect 2120 -3960 2150 -3910
rect 2040 -3990 2150 -3960
rect 1190 -5140 1300 -5110
rect 1190 -5190 1220 -5140
rect 1270 -5190 1300 -5140
rect 1190 -5220 1300 -5190
rect 1490 -5140 1600 -5110
rect 1490 -5190 1520 -5140
rect 1570 -5190 1600 -5140
rect 1490 -5220 1600 -5190
rect 1790 -5140 1900 -5110
rect 1790 -5190 1820 -5140
rect 1870 -5190 1900 -5140
rect 1790 -5220 1900 -5190
rect 2030 -6380 2140 -6350
rect 2030 -6430 2060 -6380
rect 2110 -6430 2140 -6380
rect 2030 -6460 2140 -6430
<< psubdiffcont >>
rect 50 410 100 460
rect 50 290 100 340
rect 360 -720 420 -660
rect 360 -920 420 -860
rect 340 -1960 400 -1900
rect 340 -2210 400 -2150
rect 360 -3220 420 -3160
rect 360 -3390 420 -3330
rect 350 -4470 410 -4410
rect 350 -4650 410 -4590
rect 340 -5640 400 -5580
rect 340 -5890 400 -5830
rect 330 -6890 390 -6830
<< nsubdiffcont >>
rect -130 -50 -80 0
rect -130 -180 -80 -130
rect 1190 -1470 1240 -1420
rect 1500 -1470 1550 -1420
rect 1740 -1470 1790 -1420
rect 2000 -1470 2050 -1420
rect 1570 -2710 1620 -2660
rect 1790 -2710 1840 -2660
rect 2030 -2710 2080 -2660
rect 1880 -3960 1930 -3910
rect 2070 -3960 2120 -3910
rect 1220 -5190 1270 -5140
rect 1520 -5190 1570 -5140
rect 1820 -5190 1870 -5140
rect 2060 -6430 2110 -6380
<< locali >>
rect 320 -300 690 -290
rect 320 -340 340 -300
rect 430 -340 690 -300
rect 970 -340 1290 -290
rect 320 -350 450 -340
rect 1430 -440 1580 -430
rect 1450 -500 1580 -440
rect 130 -580 570 -510
rect 1450 -540 1500 -500
rect 1540 -510 1580 -500
rect 1940 -510 2080 -280
rect 1540 -540 1570 -510
rect 1450 -550 1570 -540
rect 1480 -560 1520 -550
rect 1940 -570 1990 -510
rect 2050 -570 2080 -510
rect 130 -620 230 -580
rect 130 -660 150 -620
rect 210 -660 230 -620
rect 1940 -620 2080 -570
rect 130 -690 230 -660
rect 1940 -680 1990 -620
rect 2050 -680 2080 -620
rect 1940 -720 2080 -680
rect 60 -960 190 -930
rect 60 -1010 80 -960
rect 170 -1010 190 -960
rect 990 -960 1130 -940
rect 990 -1000 1070 -960
rect 1110 -1000 1130 -960
rect 60 -1120 570 -1010
rect 990 -1070 1130 -1000
rect 990 -1110 1070 -1070
rect 1110 -1110 1130 -1070
rect 990 -1190 1130 -1110
rect 990 -1230 1070 -1190
rect 1110 -1230 1130 -1190
rect 990 -1270 1130 -1230
rect 310 -1290 400 -1270
rect 310 -1340 330 -1290
rect 380 -1340 550 -1290
rect 310 -1360 400 -1340
rect 320 -1720 560 -1690
rect 320 -1770 370 -1720
rect 420 -1750 560 -1720
rect 890 -1700 970 -1540
rect 890 -1740 910 -1700
rect 950 -1740 970 -1700
rect 420 -1770 650 -1750
rect 320 -1800 650 -1770
rect 890 -1790 970 -1740
rect 890 -1830 910 -1790
rect 950 -1830 970 -1790
rect 890 -1870 970 -1830
rect 890 -1910 910 -1870
rect 950 -1910 970 -1870
rect 890 -1960 970 -1910
rect 1450 -2200 1570 -2180
rect 340 -2350 630 -2320
rect 340 -2390 380 -2350
rect 420 -2360 630 -2350
rect 1450 -2270 1480 -2200
rect 1550 -2270 1570 -2200
rect 420 -2390 560 -2360
rect 340 -2430 560 -2390
rect 1450 -2340 1570 -2270
rect 1450 -2410 1480 -2340
rect 1550 -2410 1570 -2340
rect 1450 -2480 1570 -2410
rect 890 -2590 1290 -2530
rect 1450 -2550 1480 -2480
rect 1550 -2550 1570 -2480
rect 1450 -2590 1570 -2550
rect 380 -2960 600 -2930
rect 380 -3010 420 -2960
rect 470 -3010 600 -2960
rect 380 -3040 600 -3010
rect 350 -3600 600 -3570
rect 350 -3650 400 -3600
rect 450 -3650 600 -3600
rect 350 -3680 600 -3650
rect 480 -4110 550 -4100
rect 480 -4160 490 -4110
rect 540 -4160 550 -4110
rect 480 -4360 550 -4160
rect 1080 -4680 1210 -4660
rect 1080 -4730 1110 -4680
rect 1190 -4730 1210 -4680
rect 1080 -4820 1210 -4730
rect 1080 -4870 1110 -4820
rect 1190 -4870 1210 -4820
rect 330 -4940 550 -4870
rect 330 -4990 350 -4940
rect 400 -4990 550 -4940
rect 1080 -4960 1210 -4870
rect 330 -5010 440 -4990
rect 1080 -5010 1110 -4960
rect 1190 -5010 1210 -4960
rect 1080 -5050 1210 -5010
<< viali >>
rect 20 460 130 480
rect 20 410 50 460
rect 50 410 100 460
rect 100 410 130 460
rect 20 340 130 410
rect -1420 279 -1386 313
rect -1148 276 -1114 310
rect -873 277 -839 311
rect -598 277 -564 311
rect -322 275 -288 309
rect 20 290 50 340
rect 50 290 100 340
rect 100 290 130 340
rect 20 260 130 290
rect -1510 180 -1470 220
rect -1420 187 -1386 221
rect -1228 193 -1194 227
rect -1143 187 -1109 221
rect -962 186 -928 220
rect -866 186 -832 220
rect -686 187 -652 221
rect -593 187 -559 221
rect -410 187 -376 221
rect -318 186 -284 220
rect -1420 98 -1386 132
rect -1147 93 -1113 127
rect -875 92 -841 126
rect -598 93 -564 127
rect -322 93 -288 127
rect -872 20 -838 54
rect -160 0 -50 30
rect -160 -50 -130 0
rect -130 -50 -80 0
rect -80 -50 -50 0
rect -160 -130 -50 -50
rect -160 -180 -130 -130
rect -130 -180 -80 -130
rect -80 -180 -50 -130
rect -160 -210 -50 -180
rect 340 -340 430 -300
rect 690 -490 730 -450
rect 810 -560 850 -520
rect 1070 -560 1110 -520
rect 1200 -560 1240 -520
rect 1280 -560 1320 -520
rect 1500 -540 1540 -500
rect 1710 -550 1760 -510
rect 1990 -570 2050 -510
rect 150 -660 210 -620
rect 330 -660 450 -630
rect 330 -720 360 -660
rect 360 -720 420 -660
rect 420 -720 450 -660
rect 1990 -680 2050 -620
rect 330 -750 450 -720
rect 330 -860 450 -830
rect 330 -920 360 -860
rect 360 -920 420 -860
rect 420 -920 450 -860
rect 330 -950 450 -920
rect 80 -1010 170 -960
rect 1070 -1000 1110 -960
rect 810 -1110 850 -1070
rect 1070 -1110 1110 -1070
rect 680 -1170 720 -1130
rect 1070 -1230 1110 -1190
rect 330 -1340 380 -1290
rect 1160 -1420 1270 -1390
rect 1160 -1470 1190 -1420
rect 1190 -1470 1240 -1420
rect 1240 -1470 1270 -1420
rect 1160 -1500 1270 -1470
rect 1470 -1420 1580 -1390
rect 1470 -1470 1500 -1420
rect 1500 -1470 1550 -1420
rect 1550 -1470 1580 -1420
rect 1470 -1500 1580 -1470
rect 1710 -1420 1820 -1390
rect 1710 -1470 1740 -1420
rect 1740 -1470 1790 -1420
rect 1790 -1470 1820 -1420
rect 1710 -1500 1820 -1470
rect 1970 -1420 2080 -1390
rect 1970 -1470 2000 -1420
rect 2000 -1470 2050 -1420
rect 2050 -1470 2080 -1420
rect 1970 -1500 2080 -1470
rect 370 -1770 420 -1720
rect 910 -1740 950 -1700
rect 700 -1800 740 -1760
rect 910 -1830 950 -1790
rect 310 -1900 430 -1870
rect 310 -1960 340 -1900
rect 340 -1960 400 -1900
rect 400 -1960 430 -1900
rect 910 -1910 950 -1870
rect 310 -1990 430 -1960
rect 310 -2150 430 -2120
rect 310 -2210 340 -2150
rect 340 -2210 400 -2150
rect 400 -2210 430 -2150
rect 310 -2240 430 -2210
rect 380 -2390 420 -2350
rect 700 -2360 740 -2320
rect 980 -2350 1020 -2260
rect 1480 -2270 1550 -2200
rect 1100 -2400 1190 -2310
rect 1270 -2350 1310 -2310
rect 1480 -2410 1550 -2340
rect 1480 -2550 1550 -2480
rect 1540 -2660 1650 -2630
rect 1540 -2710 1570 -2660
rect 1570 -2710 1620 -2660
rect 1620 -2710 1650 -2660
rect 1540 -2740 1650 -2710
rect 1760 -2660 1870 -2630
rect 1760 -2710 1790 -2660
rect 1790 -2710 1840 -2660
rect 1840 -2710 1870 -2660
rect 1760 -2740 1870 -2710
rect 2000 -2660 2110 -2630
rect 2000 -2710 2030 -2660
rect 2030 -2710 2080 -2660
rect 2080 -2710 2110 -2660
rect 2000 -2740 2110 -2710
rect 890 -2950 930 -2910
rect 420 -3010 470 -2960
rect 700 -3040 740 -3000
rect 890 -3070 930 -3030
rect 330 -3160 450 -3130
rect 330 -3220 360 -3160
rect 360 -3220 420 -3160
rect 420 -3220 450 -3160
rect 890 -3170 930 -3130
rect 330 -3330 450 -3220
rect 330 -3390 360 -3330
rect 360 -3390 420 -3330
rect 420 -3390 450 -3330
rect 330 -3420 450 -3390
rect 890 -3550 930 -3510
rect 400 -3650 450 -3600
rect 700 -3610 740 -3570
rect 890 -3630 930 -3590
rect 890 -3730 930 -3690
rect 890 -3810 930 -3770
rect 1850 -3910 1960 -3880
rect 1850 -3960 1880 -3910
rect 1880 -3960 1930 -3910
rect 1930 -3960 1960 -3910
rect 1850 -3990 1960 -3960
rect 2040 -3910 2150 -3880
rect 2040 -3960 2070 -3910
rect 2070 -3960 2120 -3910
rect 2120 -3960 2150 -3910
rect 2040 -3990 2150 -3960
rect 490 -4160 540 -4110
rect 680 -4300 720 -4260
rect 780 -4330 820 -4290
rect 320 -4410 440 -4380
rect 780 -4410 820 -4370
rect 320 -4470 350 -4410
rect 350 -4470 410 -4410
rect 410 -4470 440 -4410
rect 880 -4420 920 -4380
rect 320 -4500 440 -4470
rect 320 -4590 440 -4560
rect 320 -4650 350 -4590
rect 350 -4650 410 -4590
rect 410 -4650 440 -4590
rect 320 -4680 440 -4650
rect 680 -4730 720 -4690
rect 780 -4750 820 -4710
rect 1110 -4730 1190 -4680
rect 680 -4820 720 -4780
rect 780 -4830 820 -4790
rect 880 -4840 920 -4800
rect 1110 -4870 1190 -4820
rect 350 -4990 400 -4940
rect 1110 -5010 1190 -4960
rect 1190 -5140 1300 -5110
rect 1190 -5190 1220 -5140
rect 1220 -5190 1270 -5140
rect 1270 -5190 1300 -5140
rect 1190 -5220 1300 -5190
rect 1490 -5140 1600 -5110
rect 1490 -5190 1520 -5140
rect 1520 -5190 1570 -5140
rect 1570 -5190 1600 -5140
rect 1490 -5220 1600 -5190
rect 1790 -5140 1900 -5110
rect 1790 -5190 1820 -5140
rect 1820 -5190 1870 -5140
rect 1870 -5190 1900 -5140
rect 1790 -5220 1900 -5190
rect 310 -5580 430 -5550
rect 310 -5640 340 -5580
rect 340 -5640 400 -5580
rect 400 -5640 430 -5580
rect 310 -5670 430 -5640
rect 310 -5830 430 -5800
rect 310 -5890 340 -5830
rect 340 -5890 400 -5830
rect 400 -5890 430 -5830
rect 310 -5920 430 -5890
rect 2030 -6380 2140 -6350
rect 2030 -6430 2060 -6380
rect 2060 -6430 2110 -6380
rect 2110 -6430 2140 -6380
rect 2030 -6460 2140 -6430
rect 300 -6830 420 -6800
rect 300 -6890 330 -6830
rect 330 -6890 390 -6830
rect 390 -6890 420 -6830
rect 300 -6920 420 -6890
<< metal1 >>
rect -3910 470 -3710 690
rect -3910 280 -3870 470
rect -3750 280 -3710 470
rect -3910 270 -3710 280
rect -3660 470 -3460 690
rect -3660 280 -3620 470
rect -3500 280 -3460 470
rect -3660 270 -3460 280
rect -3410 470 -3210 690
rect -3410 280 -3370 470
rect -3250 280 -3210 470
rect -3410 270 -3210 280
rect -3160 470 -2960 690
rect -3160 280 -3120 470
rect -3000 280 -2960 470
rect -3160 270 -2960 280
rect -2910 470 -2710 690
rect -2910 280 -2870 470
rect -2750 280 -2710 470
rect -2910 270 -2710 280
rect -2660 470 -2460 690
rect -2660 280 -2620 470
rect -2500 280 -2460 470
rect -2660 270 -2460 280
rect -2410 470 -2210 690
rect -2410 280 -2370 470
rect -2250 280 -2210 470
rect -2410 270 -2210 280
rect -2160 470 -1960 690
rect -2160 280 -2120 470
rect -2000 280 -1960 470
rect -2160 270 -1960 280
rect -1910 680 -1530 690
rect -1910 560 -1700 680
rect -1540 560 -1530 680
rect -1910 550 -1530 560
rect -1910 470 -1710 550
rect -210 490 170 494
rect -1910 280 -1870 470
rect -1750 280 -1710 470
rect -1590 480 170 490
rect -1590 420 20 480
rect -1590 390 -170 420
rect -1429 330 -1362 336
rect -1910 270 -1710 280
rect -1430 313 -1362 330
rect -1430 279 -1420 313
rect -1386 279 -1362 313
rect -1430 260 -1362 279
rect -1157 310 -1079 338
rect -325 332 -273 338
rect -1157 276 -1148 310
rect -1114 276 -1079 310
rect -1157 260 -1079 276
rect -886 311 -822 327
rect -886 277 -873 311
rect -839 277 -822 311
rect -886 260 -822 277
rect -607 311 -541 324
rect -607 277 -598 311
rect -564 277 -541 311
rect -1690 240 -1610 250
rect -1430 247 -1326 260
rect -1700 234 -1680 240
rect -3380 182 -3367 234
rect -3250 182 -1680 234
rect -1690 180 -1680 182
rect -1620 234 -1600 240
rect -1530 234 -1460 240
rect -1620 220 -1460 234
rect -1620 182 -1510 220
rect -1620 180 -1610 182
rect -1690 170 -1610 180
rect -1530 180 -1510 182
rect -1470 180 -1460 220
rect -1530 160 -1460 180
rect -1430 221 -1417 247
rect -1430 187 -1420 221
rect -1430 169 -1417 187
rect -1339 169 -1326 247
rect -1430 156 -1326 169
rect -1250 248 -1190 249
rect -1250 227 -1188 248
rect -1250 193 -1228 227
rect -1194 193 -1188 227
rect -1250 167 -1188 193
rect -1157 247 -1053 260
rect -1157 169 -1144 247
rect -1066 169 -1053 247
rect -1430 132 -1360 156
rect -1430 98 -1420 132
rect -1386 98 -1360 132
rect -2880 70 -1650 80
rect -1430 70 -1360 98
rect -2880 -10 -2870 70
rect -2750 40 -1650 70
rect -1250 40 -1190 167
rect -1157 156 -1053 169
rect -988 247 -923 260
rect -886 247 -767 260
rect -607 247 -541 277
rect -331 309 -273 332
rect -331 275 -322 309
rect -288 275 -273 309
rect -331 247 -273 275
rect -208 300 -170 390
rect -30 300 20 420
rect -208 260 20 300
rect 130 260 170 480
rect -208 250 170 260
rect -923 169 -922 234
rect -886 220 -858 247
rect -886 186 -866 220
rect -886 169 -858 186
rect -780 169 -767 247
rect -988 156 -923 169
rect -886 156 -767 169
rect -728 236 -637 247
rect -728 230 -635 236
rect -728 170 -710 230
rect -650 170 -635 230
rect -728 167 -635 170
rect -607 234 -494 247
rect -607 221 -585 234
rect -607 187 -593 221
rect -607 169 -585 187
rect -507 169 -494 234
rect -728 156 -637 167
rect -607 156 -494 169
rect -455 234 -364 247
rect -455 156 -442 234
rect -1157 127 -1079 156
rect -1157 93 -1147 127
rect -1113 93 -1079 127
rect -1157 52 -1079 93
rect -886 126 -822 156
rect -720 150 -640 156
rect -886 92 -875 126
rect -841 92 -822 126
rect -886 54 -822 92
rect -607 127 -541 156
rect -455 143 -364 156
rect -331 234 -247 247
rect -331 220 -299 234
rect -331 186 -318 220
rect -331 156 -299 186
rect -331 143 -247 156
rect -607 93 -598 127
rect -564 93 -541 127
rect -607 76 -541 93
rect -331 127 -273 143
rect -331 93 -322 127
rect -288 93 -273 127
rect -331 74 -273 93
rect -2750 0 -1190 40
rect -886 20 -872 54
rect -838 20 -822 54
rect -886 7 -822 20
rect -325 0 -273 74
rect -240 40 1960 70
rect -240 30 80 40
rect -2750 -10 -1650 0
rect -2880 -20 -1650 -10
rect -240 -50 -160 30
rect -1590 -150 -160 -50
rect -240 -210 -160 -150
rect -50 -210 80 30
rect 340 -210 1960 40
rect -240 -250 1960 -210
rect -3630 -350 -3610 -290
rect -3510 -300 450 -290
rect -3510 -340 340 -300
rect 430 -340 450 -300
rect 1510 -310 1960 -250
rect -3510 -350 450 -340
rect -3380 -460 -3360 -400
rect -3260 -440 600 -400
rect 2960 -440 3370 -410
rect -3260 -450 750 -440
rect -3260 -460 690 -450
rect 490 -490 690 -460
rect 730 -490 750 -450
rect 490 -500 750 -490
rect 1480 -490 1560 -480
rect -3880 -510 420 -500
rect -3880 -570 -3860 -510
rect -3760 -530 420 -510
rect 780 -520 880 -500
rect 770 -530 810 -520
rect -3760 -560 810 -530
rect 850 -560 880 -520
rect -3760 -570 880 -560
rect -3880 -580 880 -570
rect 1050 -510 1130 -500
rect 1180 -510 1260 -500
rect 1050 -570 1060 -510
rect 1120 -570 1130 -510
rect 1050 -580 1130 -570
rect 1160 -570 1190 -510
rect 1250 -520 1340 -510
rect 1250 -560 1280 -520
rect 1320 -560 1340 -520
rect 1480 -550 1490 -490
rect 1550 -550 1560 -490
rect 1480 -560 1560 -550
rect 1700 -500 1770 -490
rect 1700 -560 1710 -500
rect 1250 -570 1340 -560
rect 1700 -570 1770 -560
rect 1970 -510 2180 -500
rect 1160 -573 1320 -570
rect 1180 -580 1260 -573
rect 130 -670 140 -610
rect 220 -670 230 -610
rect 130 -680 230 -670
rect 310 -630 470 -610
rect 310 -720 330 -630
rect -190 -740 330 -720
rect -190 -890 -170 -740
rect -30 -750 330 -740
rect 450 -720 470 -630
rect 1970 -680 1990 -510
rect 2050 -520 2180 -510
rect 2160 -680 2180 -520
rect 1970 -690 2180 -680
rect 450 -750 1960 -720
rect -30 -830 1960 -750
rect 2960 -750 2990 -440
rect 3340 -500 3370 -440
rect 3340 -700 3570 -500
rect 3340 -750 3370 -700
rect 2960 -780 3370 -750
rect -30 -890 330 -830
rect -190 -910 330 -890
rect 70 -950 180 -940
rect 70 -1020 80 -950
rect 170 -1020 180 -950
rect 310 -950 330 -910
rect 450 -910 1960 -830
rect 2960 -850 3370 -820
rect 450 -950 470 -910
rect 310 -970 470 -950
rect 1050 -960 1130 -940
rect 70 -1030 180 -1020
rect 600 -1060 870 -1050
rect -2880 -1120 -2860 -1060
rect -2760 -1070 870 -1060
rect -2760 -1090 810 -1070
rect -2760 -1120 610 -1090
rect 770 -1110 810 -1090
rect 850 -1110 870 -1070
rect 770 -1120 870 -1110
rect 660 -1130 740 -1120
rect 660 -1150 680 -1130
rect -2380 -1210 -2360 -1150
rect -2260 -1170 680 -1150
rect 720 -1170 740 -1130
rect -2260 -1210 740 -1170
rect 1050 -1250 1060 -960
rect 1120 -1250 1130 -960
rect 1050 -1270 1130 -1250
rect 2960 -1230 2990 -850
rect 3340 -950 3370 -850
rect 3340 -1150 3570 -950
rect 3340 -1230 3370 -1150
rect 2960 -1260 3370 -1230
rect 310 -1280 400 -1270
rect 310 -1350 320 -1280
rect 390 -1350 400 -1280
rect 2290 -1320 2620 -1290
rect 2290 -1350 2320 -1320
rect 310 -1360 400 -1350
rect 480 -1390 2320 -1350
rect 480 -1500 1160 -1390
rect 1270 -1500 1470 -1390
rect 1580 -1500 1710 -1390
rect 1820 -1500 1970 -1390
rect 2080 -1500 2320 -1390
rect 480 -1530 2320 -1500
rect 2290 -1560 2320 -1530
rect 2590 -1560 2620 -1320
rect 2290 -1580 2620 -1560
rect 890 -1700 1330 -1680
rect 350 -1710 440 -1700
rect 350 -1780 360 -1710
rect 430 -1780 440 -1710
rect 890 -1740 910 -1700
rect 950 -1740 1330 -1700
rect 350 -1790 440 -1780
rect 680 -1800 690 -1740
rect 750 -1800 760 -1740
rect 680 -1810 760 -1800
rect 890 -1790 1330 -1740
rect 890 -1830 910 -1790
rect 950 -1820 1330 -1790
rect 950 -1830 1220 -1820
rect 290 -1870 450 -1850
rect 290 -1970 310 -1870
rect -190 -1990 310 -1970
rect 430 -1970 450 -1870
rect 890 -1870 1220 -1830
rect 890 -1910 910 -1870
rect 950 -1910 1220 -1870
rect 890 -1930 1220 -1910
rect 1320 -1930 1330 -1820
rect 890 -1940 1330 -1930
rect 430 -1990 1500 -1970
rect -190 -2130 -170 -1990
rect -30 -2120 1500 -1990
rect -30 -2130 310 -2120
rect -190 -2150 310 -2130
rect 290 -2240 310 -2150
rect 430 -2150 1500 -2120
rect 2960 -2080 3370 -2050
rect 430 -2240 450 -2150
rect 290 -2260 450 -2240
rect 1460 -2200 1700 -2190
rect 960 -2260 1040 -2250
rect 680 -2310 760 -2300
rect 350 -2330 450 -2320
rect 350 -2410 360 -2330
rect 440 -2410 450 -2330
rect 680 -2370 690 -2310
rect 750 -2370 760 -2310
rect 960 -2350 970 -2260
rect 1030 -2350 1040 -2260
rect 1460 -2270 1480 -2200
rect 1550 -2270 1580 -2200
rect 1260 -2300 1320 -2290
rect 960 -2360 1040 -2350
rect 1080 -2310 1210 -2300
rect 680 -2380 760 -2370
rect 350 -2420 450 -2410
rect 1080 -2410 1090 -2310
rect 1200 -2410 1210 -2310
rect 1260 -2370 1320 -2360
rect 1460 -2340 1580 -2270
rect 1080 -2420 1210 -2410
rect 1460 -2410 1480 -2340
rect 1550 -2410 1580 -2340
rect 1460 -2480 1580 -2410
rect 1460 -2550 1480 -2480
rect 1550 -2550 1580 -2480
rect 1690 -2550 1700 -2200
rect 2960 -2460 2990 -2080
rect 3340 -2170 3370 -2080
rect 3340 -2370 3570 -2170
rect 3340 -2460 3370 -2370
rect 2960 -2490 3370 -2460
rect 1460 -2560 1700 -2550
rect 2290 -2550 2620 -2520
rect 2290 -2590 2320 -2550
rect 480 -2630 2320 -2590
rect 480 -2740 1540 -2630
rect 1650 -2740 1760 -2630
rect 1870 -2740 2000 -2630
rect 2110 -2740 2320 -2630
rect 480 -2770 2320 -2740
rect 2290 -2790 2320 -2770
rect 2590 -2790 2620 -2550
rect 2290 -2820 2620 -2790
rect 870 -2900 1510 -2890
rect 870 -2910 1080 -2900
rect 390 -2940 500 -2930
rect 390 -3030 400 -2940
rect 490 -3030 500 -2940
rect 870 -2950 890 -2910
rect 930 -2950 1080 -2910
rect 390 -3040 500 -3030
rect 680 -3040 690 -2980
rect 750 -3040 760 -2980
rect 680 -3050 760 -3040
rect 870 -3030 1080 -2950
rect 870 -3070 890 -3030
rect 930 -3070 1080 -3030
rect 310 -3130 470 -3110
rect 310 -3210 330 -3130
rect -190 -3230 330 -3210
rect -190 -3390 -170 -3230
rect -30 -3390 330 -3230
rect -190 -3410 330 -3390
rect 310 -3420 330 -3410
rect 450 -3210 470 -3130
rect 870 -3130 1080 -3070
rect 870 -3170 890 -3130
rect 930 -3170 1080 -3130
rect 1200 -3170 1440 -2900
rect 1500 -3170 1510 -2900
rect 870 -3180 1510 -3170
rect 450 -3410 950 -3210
rect 450 -3420 470 -3410
rect 310 -3440 470 -3420
rect 870 -3510 1400 -3500
rect 870 -3550 890 -3510
rect 930 -3550 970 -3510
rect 370 -3580 480 -3570
rect 370 -3670 380 -3580
rect 470 -3670 480 -3580
rect 680 -3610 690 -3550
rect 750 -3610 760 -3550
rect 680 -3620 760 -3610
rect 870 -3590 970 -3550
rect 370 -3680 480 -3670
rect 870 -3630 890 -3590
rect 930 -3630 970 -3590
rect 870 -3690 970 -3630
rect 870 -3730 890 -3690
rect 930 -3730 970 -3690
rect 870 -3770 970 -3730
rect 870 -3810 890 -3770
rect 930 -3810 970 -3770
rect 1030 -3810 1400 -3510
rect 870 -3820 1400 -3810
rect 2290 -3810 2620 -3780
rect 2290 -3850 2320 -3810
rect 480 -3880 2320 -3850
rect 480 -3990 1850 -3880
rect 1960 -3990 2040 -3880
rect 2150 -3990 2320 -3880
rect 480 -4007 2320 -3990
rect 480 -4010 1276 -4007
rect 480 -4020 1120 -4010
rect 1487 -4020 2320 -4007
rect 2290 -4050 2320 -4020
rect 2590 -4050 2620 -3810
rect 2290 -4080 2620 -4050
rect 370 -4100 550 -4090
rect 370 -4170 380 -4100
rect 450 -4110 550 -4100
rect 450 -4160 490 -4110
rect 540 -4160 550 -4110
rect 450 -4170 550 -4160
rect 370 -4180 550 -4170
rect 3010 -4190 3210 -3990
rect 770 -4220 830 -4210
rect 100 -4250 180 -4240
rect -1170 -4310 -1150 -4250
rect -1040 -4310 110 -4250
rect 170 -4260 740 -4250
rect 170 -4300 680 -4260
rect 720 -4300 740 -4260
rect 170 -4310 740 -4300
rect 770 -4290 830 -4280
rect 100 -4320 180 -4310
rect 770 -4330 780 -4290
rect 820 -4330 830 -4290
rect 300 -4380 460 -4360
rect 300 -4460 320 -4380
rect -190 -4480 320 -4460
rect -190 -4620 -170 -4480
rect -30 -4500 320 -4480
rect 440 -4460 460 -4380
rect 770 -4370 830 -4330
rect 770 -4410 780 -4370
rect 820 -4410 830 -4370
rect 770 -4430 830 -4410
rect 860 -4360 940 -4350
rect 860 -4420 870 -4360
rect 930 -4420 940 -4360
rect 860 -4430 940 -4420
rect 440 -4500 1790 -4460
rect -30 -4560 1790 -4500
rect -30 -4620 320 -4560
rect -190 -4640 320 -4620
rect 300 -4680 320 -4640
rect 440 -4640 1790 -4560
rect 440 -4680 460 -4640
rect 100 -4700 180 -4690
rect 300 -4700 460 -4680
rect 670 -4690 730 -4670
rect 100 -4760 110 -4700
rect 170 -4730 180 -4700
rect 670 -4730 680 -4690
rect 720 -4730 730 -4690
rect 170 -4760 730 -4730
rect 100 -4770 730 -4760
rect 670 -4780 730 -4770
rect 670 -4820 680 -4780
rect 720 -4820 730 -4780
rect 670 -4840 730 -4820
rect 760 -4840 770 -4670
rect 830 -4840 840 -4670
rect 1080 -4680 1150 -4670
rect 1080 -4730 1110 -4680
rect 760 -4850 840 -4840
rect 870 -4790 940 -4780
rect 870 -4850 880 -4790
rect 870 -4860 940 -4850
rect 1080 -4820 1150 -4730
rect 1080 -4870 1110 -4820
rect 330 -4930 420 -4920
rect 330 -5000 340 -4930
rect 410 -5000 420 -4930
rect 330 -5010 420 -5000
rect 1080 -4960 1150 -4870
rect 1080 -5010 1110 -4960
rect 1080 -5040 1150 -5010
rect 1210 -5040 1220 -4670
rect 1140 -5050 1220 -5040
rect 2290 -5030 2620 -5000
rect 2290 -5080 2320 -5030
rect 480 -5110 2320 -5080
rect 480 -5220 1190 -5110
rect 1300 -5220 1490 -5110
rect 1600 -5220 1790 -5110
rect 1900 -5220 2320 -5110
rect 480 -5250 2320 -5220
rect 2290 -5270 2320 -5250
rect 2590 -5270 2620 -5030
rect 2290 -5300 2620 -5270
rect 290 -5550 450 -5530
rect 290 -5670 310 -5550
rect 430 -5670 450 -5550
rect -190 -5690 450 -5670
rect -190 -5780 -170 -5690
rect -30 -5780 1140 -5690
rect -190 -5800 1140 -5780
rect 290 -5920 310 -5800
rect 430 -5870 1140 -5800
rect 430 -5920 450 -5870
rect 290 -5940 450 -5920
rect 2290 -6290 2620 -6260
rect 2290 -6310 2320 -6290
rect 480 -6350 2320 -6310
rect 480 -6460 2030 -6350
rect 2140 -6460 2320 -6350
rect 480 -6490 2320 -6460
rect 2290 -6530 2320 -6490
rect 2590 -6530 2620 -6290
rect 2290 -6560 2620 -6530
rect 290 -6790 430 -6780
rect -190 -6800 430 -6790
rect -190 -6810 300 -6800
rect -190 -6910 -170 -6810
rect -30 -6910 300 -6810
rect -190 -6920 300 -6910
rect 420 -6920 430 -6800
rect -190 -6930 430 -6920
rect 290 -7050 1970 -6930
<< via1 >>
rect -3870 280 -3750 470
rect -3620 280 -3500 470
rect -3370 280 -3250 470
rect -3120 280 -3000 470
rect -2870 280 -2750 470
rect -2620 280 -2500 470
rect -2370 280 -2250 470
rect -2120 280 -2000 470
rect -1700 560 -1540 680
rect -1870 280 -1750 470
rect -3367 182 -3250 234
rect -1680 180 -1620 240
rect -1417 221 -1339 247
rect -1417 187 -1386 221
rect -1386 187 -1339 221
rect -1417 169 -1339 187
rect -1144 221 -1066 247
rect -1144 187 -1143 221
rect -1143 187 -1109 221
rect -1109 187 -1066 221
rect -1144 169 -1066 187
rect -2870 -10 -2750 70
rect -988 220 -923 247
rect -170 300 -30 420
rect -988 186 -962 220
rect -962 186 -928 220
rect -928 186 -923 220
rect -988 169 -923 186
rect -858 220 -780 247
rect -858 186 -832 220
rect -832 186 -780 220
rect -858 169 -780 186
rect -710 221 -650 230
rect -710 187 -686 221
rect -686 187 -652 221
rect -652 187 -650 221
rect -710 170 -650 187
rect -585 221 -507 234
rect -585 187 -559 221
rect -559 187 -507 221
rect -585 169 -507 187
rect -442 221 -364 234
rect -442 187 -410 221
rect -410 187 -376 221
rect -376 187 -364 221
rect -442 156 -364 187
rect -299 220 -247 234
rect -299 186 -284 220
rect -284 186 -247 220
rect -299 156 -247 186
rect 80 -210 340 40
rect -3610 -350 -3510 -290
rect -3360 -460 -3260 -400
rect -3860 -570 -3760 -510
rect 1060 -520 1120 -510
rect 1060 -560 1070 -520
rect 1070 -560 1110 -520
rect 1110 -560 1120 -520
rect 1060 -570 1120 -560
rect 1190 -520 1250 -510
rect 1190 -560 1200 -520
rect 1200 -560 1240 -520
rect 1240 -560 1250 -520
rect 1490 -500 1550 -490
rect 1490 -540 1500 -500
rect 1500 -540 1540 -500
rect 1540 -540 1550 -500
rect 1490 -550 1550 -540
rect 1710 -510 1770 -500
rect 1710 -550 1760 -510
rect 1760 -550 1770 -510
rect 1710 -560 1770 -550
rect 1190 -570 1250 -560
rect 140 -620 220 -610
rect 140 -660 150 -620
rect 150 -660 210 -620
rect 210 -660 220 -620
rect 140 -670 220 -660
rect -170 -890 -30 -740
rect 1990 -570 2050 -520
rect 2050 -570 2160 -520
rect 1990 -620 2160 -570
rect 1990 -680 2050 -620
rect 2050 -680 2160 -620
rect 2990 -750 3340 -440
rect 80 -960 170 -950
rect 80 -1010 170 -960
rect 80 -1020 170 -1010
rect -2860 -1120 -2760 -1060
rect -2360 -1210 -2260 -1150
rect 1060 -1000 1070 -960
rect 1070 -1000 1110 -960
rect 1110 -1000 1120 -960
rect 1060 -1070 1120 -1000
rect 1060 -1110 1070 -1070
rect 1070 -1110 1110 -1070
rect 1110 -1110 1120 -1070
rect 1060 -1190 1120 -1110
rect 1060 -1230 1070 -1190
rect 1070 -1230 1110 -1190
rect 1110 -1230 1120 -1190
rect 1060 -1250 1120 -1230
rect 2990 -1230 3340 -850
rect 320 -1290 390 -1280
rect 320 -1340 330 -1290
rect 330 -1340 380 -1290
rect 380 -1340 390 -1290
rect 320 -1350 390 -1340
rect 2320 -1560 2590 -1320
rect 360 -1720 430 -1710
rect 360 -1770 370 -1720
rect 370 -1770 420 -1720
rect 420 -1770 430 -1720
rect 360 -1780 430 -1770
rect 690 -1760 750 -1740
rect 690 -1800 700 -1760
rect 700 -1800 740 -1760
rect 740 -1800 750 -1760
rect 1220 -1930 1320 -1820
rect -170 -2130 -30 -1990
rect 360 -2350 440 -2330
rect 360 -2390 380 -2350
rect 380 -2390 420 -2350
rect 420 -2390 440 -2350
rect 360 -2410 440 -2390
rect 690 -2320 750 -2310
rect 690 -2360 700 -2320
rect 700 -2360 740 -2320
rect 740 -2360 750 -2320
rect 690 -2370 750 -2360
rect 970 -2350 980 -2260
rect 980 -2350 1020 -2260
rect 1020 -2350 1030 -2260
rect 1090 -2400 1100 -2310
rect 1100 -2400 1190 -2310
rect 1190 -2400 1200 -2310
rect 1090 -2410 1200 -2400
rect 1260 -2310 1320 -2300
rect 1260 -2350 1270 -2310
rect 1270 -2350 1310 -2310
rect 1310 -2350 1320 -2310
rect 1260 -2360 1320 -2350
rect 1580 -2550 1690 -2200
rect 2990 -2460 3340 -2080
rect 2320 -2790 2590 -2550
rect 400 -2960 490 -2940
rect 400 -3010 420 -2960
rect 420 -3010 470 -2960
rect 470 -3010 490 -2960
rect 400 -3030 490 -3010
rect 690 -3000 750 -2980
rect 690 -3040 700 -3000
rect 700 -3040 740 -3000
rect 740 -3040 750 -3000
rect -170 -3390 -30 -3230
rect 1080 -3170 1200 -2900
rect 1440 -3170 1500 -2900
rect 380 -3600 470 -3580
rect 380 -3650 400 -3600
rect 400 -3650 450 -3600
rect 450 -3650 470 -3600
rect 380 -3670 470 -3650
rect 690 -3570 750 -3550
rect 690 -3610 700 -3570
rect 700 -3610 740 -3570
rect 740 -3610 750 -3570
rect 970 -3810 1030 -3510
rect 2320 -4050 2590 -3810
rect 380 -4170 450 -4100
rect -1150 -4310 -1040 -4250
rect 110 -4310 170 -4250
rect 770 -4280 830 -4220
rect -170 -4620 -30 -4480
rect 870 -4380 930 -4360
rect 870 -4420 880 -4380
rect 880 -4420 920 -4380
rect 920 -4420 930 -4380
rect 110 -4760 170 -4700
rect 770 -4710 830 -4670
rect 770 -4750 780 -4710
rect 780 -4750 820 -4710
rect 820 -4750 830 -4710
rect 770 -4790 830 -4750
rect 770 -4830 780 -4790
rect 780 -4830 820 -4790
rect 820 -4830 830 -4790
rect 770 -4840 830 -4830
rect 1150 -4680 1210 -4670
rect 1150 -4730 1190 -4680
rect 1190 -4730 1210 -4680
rect 880 -4800 940 -4790
rect 880 -4840 920 -4800
rect 920 -4840 940 -4800
rect 880 -4850 940 -4840
rect 1150 -4820 1210 -4730
rect 1150 -4870 1190 -4820
rect 1190 -4870 1210 -4820
rect 340 -4940 410 -4930
rect 340 -4990 350 -4940
rect 350 -4990 400 -4940
rect 400 -4990 410 -4940
rect 340 -5000 410 -4990
rect 1150 -4960 1210 -4870
rect 1150 -5010 1190 -4960
rect 1190 -5010 1210 -4960
rect 1150 -5040 1210 -5010
rect 2320 -5270 2590 -5030
rect -170 -5780 -30 -5690
rect 2320 -6530 2590 -6290
rect -170 -6910 -30 -6810
<< metal2 >>
rect -1710 680 -1530 690
rect -1710 560 -1700 680
rect -1540 560 -1530 680
rect -1710 550 -1530 560
rect 1670 680 1810 690
rect 1670 560 1680 680
rect 1800 560 1810 680
rect 1670 550 1810 560
rect -3880 470 -3740 480
rect -3880 280 -3870 470
rect -3750 280 -3740 470
rect -3880 -510 -3740 280
rect -3880 -570 -3860 -510
rect -3760 -570 -3740 -510
rect -3880 -7030 -3740 -570
rect -3630 470 -3490 480
rect -3630 280 -3620 470
rect -3500 280 -3490 470
rect -3630 -290 -3490 280
rect -3630 -350 -3610 -290
rect -3510 -350 -3490 -290
rect -3630 -7030 -3490 -350
rect -3380 470 -3240 480
rect -3380 280 -3370 470
rect -3250 280 -3240 470
rect -3380 234 -3240 280
rect -3380 182 -3367 234
rect -3250 182 -3240 234
rect -3380 -400 -3240 182
rect -3380 -460 -3360 -400
rect -3260 -460 -3240 -400
rect -3380 -4100 -3240 -460
rect -3380 -4170 -3370 -4100
rect -3250 -4170 -3240 -4100
rect -3380 -7030 -3240 -4170
rect -3130 470 -2990 480
rect -3130 280 -3120 470
rect -3000 280 -2990 470
rect -3130 -600 -2990 280
rect -3130 -660 -3120 -600
rect -3000 -660 -2990 -600
rect -3130 -4930 -2990 -660
rect -3130 -5000 -3120 -4930
rect -3000 -5000 -2990 -4930
rect -3130 -7030 -2990 -5000
rect -2880 470 -2740 480
rect -2880 280 -2870 470
rect -2750 280 -2740 470
rect -2880 70 -2740 280
rect -2880 -10 -2870 70
rect -2750 -10 -2740 70
rect -2880 -1060 -2740 -10
rect -2880 -1120 -2860 -1060
rect -2760 -1120 -2740 -1060
rect -2880 -1560 -2740 -1120
rect -2880 -1620 -2870 -1560
rect -2750 -1620 -2740 -1560
rect -2880 -7030 -2740 -1620
rect -2630 470 -2490 480
rect -2630 280 -2620 470
rect -2500 280 -2490 470
rect -2630 260 -2490 280
rect -2630 156 -2613 260
rect -2496 156 -2490 260
rect -2630 -1280 -2490 156
rect -2630 -1350 -2620 -1280
rect -2500 -1350 -2490 -1280
rect -2630 -2490 -2490 -1350
rect -2630 -2550 -2620 -2490
rect -2500 -2550 -2490 -2490
rect -2630 -7030 -2490 -2550
rect -2380 470 -2240 480
rect -2380 280 -2370 470
rect -2250 280 -2240 470
rect -2380 78 -2240 280
rect -2380 0 -2366 78
rect -2249 0 -2240 78
rect -2380 -1150 -2240 0
rect -2380 -1210 -2360 -1150
rect -2260 -1210 -2240 -1150
rect -2380 -2800 -2240 -1210
rect -2380 -2860 -2370 -2800
rect -2250 -2860 -2240 -2800
rect -2380 -7030 -2240 -2860
rect -2130 470 -1990 480
rect -2130 280 -2120 470
rect -2000 280 -1990 470
rect -2130 -950 -1990 280
rect -2130 -1020 -2110 -950
rect -2010 -1020 -1990 -950
rect -2130 -3440 -1990 -1020
rect -2130 -3500 -2120 -3440
rect -2000 -3500 -1990 -3440
rect -2130 -7030 -1990 -3500
rect -1880 470 -1740 480
rect -1880 280 -1870 470
rect -1750 280 -1740 470
rect -180 420 -20 430
rect -1880 -1710 -1740 280
rect -455 390 -351 403
rect -455 325 -442 390
rect -364 325 -351 390
rect -1690 240 -1610 250
rect -1690 180 -1680 240
rect -1620 180 -1610 240
rect -1690 170 -1610 180
rect -1443 247 -1313 260
rect -1690 169 -1612 170
rect -1443 169 -1417 247
rect -1339 169 -1313 247
rect -1443 -260 -1313 169
rect -1157 247 -1027 260
rect -1157 169 -1144 247
rect -1066 169 -1027 247
rect -1157 -110 -1027 169
rect -988 247 -897 260
rect -910 169 -897 247
rect -988 156 -897 169
rect -860 247 -767 260
rect -860 169 -858 247
rect -780 169 -767 247
rect -860 160 -767 169
rect -858 -52 -767 160
rect -730 230 -630 250
rect -730 170 -710 230
rect -650 170 -630 230
rect -730 150 -630 170
rect -598 234 -494 247
rect -598 169 -585 234
rect -507 169 -494 234
rect -598 156 -494 169
rect -728 104 -637 150
rect -728 26 -715 104
rect -650 26 -637 104
rect -728 13 -637 26
rect -1880 -1780 -1870 -1710
rect -1750 -1780 -1740 -1710
rect -1880 -2330 -1740 -1780
rect -1880 -2410 -1870 -2330
rect -1750 -2410 -1740 -2330
rect -1880 -2940 -1740 -2410
rect -1880 -3030 -1870 -2940
rect -1750 -3030 -1740 -2940
rect -1880 -3580 -1740 -3030
rect -1880 -3670 -1870 -3580
rect -1750 -3670 -1740 -3580
rect -1880 -4360 -1740 -3670
rect -1880 -4420 -1870 -4360
rect -1750 -4420 -1740 -4360
rect -1880 -4790 -1740 -4420
rect -1880 -4850 -1870 -4790
rect -1750 -4850 -1740 -4790
rect -1880 -7030 -1740 -4850
rect -1450 -7030 -1310 -260
rect -1170 -4250 -1020 -110
rect -871 -250 -767 -52
rect -585 -180 -494 156
rect -455 234 -351 325
rect -180 300 -170 420
rect -30 300 -20 420
rect -180 290 -20 300
rect -455 156 -442 234
rect -364 156 -351 234
rect -455 143 -351 156
rect -320 234 -220 250
rect -320 200 -299 234
rect -247 200 -220 234
rect -320 130 -310 200
rect -230 130 -220 200
rect -320 110 -220 130
rect 1180 200 1270 210
rect 1180 130 1190 200
rect 1260 130 1270 200
rect 70 40 350 50
rect -1170 -4310 -1150 -4250
rect -1040 -4310 -1020 -4250
rect -1170 -7030 -1020 -4310
rect -890 -4240 -740 -250
rect -890 -4300 -880 -4240
rect -750 -4300 -740 -4240
rect -890 -7030 -740 -4300
rect -610 -7030 -470 -180
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect 1050 -510 1130 -500
rect 1050 -570 1060 -510
rect 1120 -570 1130 -510
rect 130 -610 230 -600
rect 130 -670 140 -610
rect 220 -670 230 -610
rect 130 -680 230 -670
rect -180 -740 -20 -730
rect -180 -890 -170 -740
rect -30 -890 -20 -740
rect -180 -900 -20 -890
rect 70 -950 180 -940
rect 70 -1020 80 -950
rect 170 -1020 180 -950
rect 70 -1030 180 -1020
rect 1050 -960 1130 -570
rect 1180 -510 1270 130
rect 1180 -570 1190 -510
rect 1250 -570 1270 -510
rect 1180 -580 1270 -570
rect 1480 -490 1560 -480
rect 1480 -550 1490 -490
rect 1550 -550 1560 -490
rect 1050 -1250 1060 -960
rect 1120 -1250 1130 -960
rect 1480 -1010 1560 -550
rect 1700 -500 1780 550
rect 2960 -440 3370 -410
rect 1700 -560 1710 -500
rect 1770 -560 1780 -500
rect 1700 -570 1780 -560
rect 1970 -520 2180 -500
rect 1970 -680 1990 -520
rect 2160 -680 2180 -520
rect 1970 -690 2180 -680
rect 2960 -750 2990 -440
rect 3340 -750 3370 -440
rect 2960 -780 3370 -750
rect 1480 -1070 1490 -1010
rect 1550 -1070 1560 -1010
rect 1480 -1090 1560 -1070
rect 2960 -850 3370 -820
rect 1050 -1270 1130 -1250
rect 2960 -1230 2990 -850
rect 3340 -1230 3370 -850
rect 2960 -1260 3370 -1230
rect 310 -1280 400 -1270
rect 310 -1350 320 -1280
rect 390 -1350 400 -1280
rect 310 -1360 400 -1350
rect 2310 -1320 2600 -1310
rect 680 -1560 760 -1550
rect 680 -1620 690 -1560
rect 750 -1620 760 -1560
rect 2310 -1560 2320 -1320
rect 2590 -1560 2600 -1320
rect 2310 -1570 2600 -1560
rect 350 -1710 440 -1700
rect 350 -1780 360 -1710
rect 430 -1780 440 -1710
rect 350 -1790 440 -1780
rect 680 -1740 760 -1620
rect 680 -1800 690 -1740
rect 750 -1800 760 -1740
rect 680 -1810 760 -1800
rect 1210 -1820 1330 -1810
rect 1210 -1930 1220 -1820
rect 1320 -1930 1330 -1820
rect 1210 -1940 1330 -1930
rect -180 -1990 -20 -1980
rect -180 -2130 -170 -1990
rect -30 -2130 -20 -1990
rect -180 -2140 -20 -2130
rect 960 -2260 1040 -2250
rect 680 -2310 760 -2300
rect 350 -2330 450 -2320
rect 350 -2410 360 -2330
rect 440 -2410 450 -2330
rect 350 -2420 450 -2410
rect 680 -2370 690 -2310
rect 750 -2370 760 -2310
rect 680 -2490 760 -2370
rect 680 -2550 690 -2490
rect 750 -2550 760 -2490
rect 680 -2560 760 -2550
rect 960 -2350 970 -2260
rect 1030 -2350 1040 -2260
rect 1250 -2300 1330 -1940
rect 2960 -2080 3370 -2050
rect 680 -2800 760 -2790
rect 680 -2860 690 -2800
rect 750 -2860 760 -2800
rect 390 -2940 500 -2930
rect 390 -3030 400 -2940
rect 490 -3030 500 -2940
rect 390 -3040 500 -3030
rect 680 -2980 760 -2860
rect 680 -3040 690 -2980
rect 750 -3040 760 -2980
rect 680 -3050 760 -3040
rect -180 -3230 -20 -3220
rect -180 -3390 -170 -3230
rect -30 -3390 -20 -3230
rect -180 -3400 -20 -3390
rect 680 -3440 760 -3430
rect 680 -3500 690 -3440
rect 750 -3500 760 -3440
rect 680 -3550 760 -3500
rect 370 -3580 480 -3570
rect 370 -3670 380 -3580
rect 470 -3670 480 -3580
rect 680 -3610 690 -3550
rect 750 -3610 760 -3550
rect 680 -3620 760 -3610
rect 960 -3510 1040 -2350
rect 1070 -2310 1210 -2300
rect 1070 -2410 1090 -2310
rect 1200 -2410 1210 -2310
rect 1250 -2360 1260 -2300
rect 1320 -2360 1330 -2300
rect 1250 -2370 1330 -2360
rect 1570 -2200 1700 -2190
rect 1070 -2430 1210 -2410
rect 1110 -2890 1210 -2430
rect 1570 -2550 1580 -2200
rect 1690 -2550 1700 -2200
rect 2960 -2460 2990 -2080
rect 3340 -2460 3370 -2080
rect 2960 -2490 3370 -2460
rect 1570 -2560 1700 -2550
rect 2310 -2550 2600 -2540
rect 2310 -2790 2320 -2550
rect 2590 -2790 2600 -2550
rect 2310 -2800 2600 -2790
rect 1070 -2900 1210 -2890
rect 1070 -3170 1080 -2900
rect 1200 -3170 1210 -2900
rect 1070 -3180 1210 -3170
rect 1430 -2900 1510 -2890
rect 1430 -3170 1440 -2900
rect 1500 -3170 1510 -2900
rect 370 -3680 480 -3670
rect 960 -3810 970 -3510
rect 1030 -3810 1040 -3510
rect 960 -3820 1040 -3810
rect 1430 -3500 1510 -3170
rect 1430 -3820 1570 -3500
rect 2310 -3810 2600 -3800
rect 2310 -4050 2320 -3810
rect 2590 -4050 2600 -3810
rect 2310 -4060 2600 -4050
rect 370 -4100 460 -4090
rect 370 -4170 380 -4100
rect 450 -4170 460 -4100
rect 370 -4180 460 -4170
rect 760 -4220 840 -4210
rect 100 -4250 180 -4240
rect 100 -4310 110 -4250
rect 170 -4310 180 -4250
rect 760 -4280 770 -4220
rect 830 -4280 840 -4220
rect 760 -4290 840 -4280
rect -180 -4480 -20 -4470
rect -180 -4620 -170 -4480
rect -30 -4620 -20 -4480
rect -180 -4630 -20 -4620
rect 100 -4700 180 -4310
rect 100 -4760 110 -4700
rect 170 -4760 180 -4700
rect 100 -4770 180 -4760
rect 770 -4670 830 -4290
rect 860 -4360 940 -4350
rect 860 -4420 870 -4360
rect 930 -4420 940 -4360
rect 860 -4430 940 -4420
rect 1150 -4670 1300 -4650
rect 770 -4850 830 -4840
rect 870 -4790 950 -4780
rect 870 -4850 880 -4790
rect 940 -4850 950 -4790
rect 870 -4860 950 -4850
rect 330 -4930 420 -4920
rect 330 -5000 340 -4930
rect 410 -5000 420 -4930
rect 330 -5010 420 -5000
rect 1210 -5040 1300 -4670
rect 1150 -5050 1300 -5040
rect 2310 -5030 2600 -5020
rect 2310 -5270 2320 -5030
rect 2590 -5270 2600 -5030
rect 2310 -5280 2600 -5270
rect -180 -5690 -20 -5680
rect -180 -5780 -170 -5690
rect -30 -5780 -20 -5690
rect -180 -5790 -20 -5780
rect 2310 -6290 2600 -6280
rect 2310 -6530 2320 -6290
rect 2590 -6530 2600 -6290
rect 2310 -6540 2600 -6530
rect -180 -6810 -20 -6800
rect -180 -6910 -170 -6810
rect -30 -6910 -20 -6810
rect -180 -6920 -20 -6910
<< via2 >>
rect -1700 560 -1540 680
rect 1680 560 1800 680
rect -3370 -4170 -3250 -4100
rect -3120 -660 -3000 -600
rect -3120 -5000 -3000 -4930
rect -2870 -1620 -2750 -1560
rect -2613 156 -2496 260
rect -2620 -1350 -2500 -1280
rect -2620 -2550 -2500 -2490
rect -2366 0 -2249 78
rect -2370 -2860 -2250 -2800
rect -2110 -1020 -2010 -950
rect -2120 -3500 -2000 -3440
rect -1859 338 -1768 403
rect -442 325 -364 390
rect -988 169 -923 247
rect -923 169 -910 247
rect -715 26 -650 104
rect -1870 -1780 -1750 -1710
rect -1870 -2410 -1750 -2330
rect -1870 -3030 -1750 -2940
rect -1870 -3670 -1750 -3580
rect -1870 -4420 -1750 -4360
rect -1870 -4850 -1750 -4790
rect -170 300 -30 420
rect -310 156 -299 200
rect -299 156 -247 200
rect -247 156 -230 200
rect -310 130 -230 156
rect 1190 130 1260 200
rect -880 -4300 -750 -4240
rect 80 -210 340 40
rect 140 -670 220 -610
rect -170 -890 -30 -740
rect 80 -1020 170 -950
rect 1990 -680 2160 -520
rect 2990 -750 3340 -440
rect 1490 -1070 1550 -1010
rect 2990 -1230 3340 -850
rect 320 -1350 390 -1280
rect 690 -1620 750 -1560
rect 2320 -1560 2590 -1320
rect 360 -1780 430 -1710
rect -170 -2130 -30 -1990
rect 360 -2410 440 -2330
rect 690 -2550 750 -2490
rect 690 -2860 750 -2800
rect 400 -3030 490 -2940
rect -170 -3380 -30 -3230
rect 690 -3500 750 -3440
rect 380 -3670 470 -3580
rect 1580 -2350 1690 -2200
rect 2990 -2460 3340 -2080
rect 2320 -2790 2590 -2550
rect 2320 -4050 2590 -3810
rect 380 -4160 450 -4100
rect 770 -4280 830 -4220
rect -170 -4620 -30 -4480
rect 870 -4420 930 -4360
rect 880 -4850 940 -4790
rect 340 -5000 410 -4930
rect 2320 -5270 2590 -5030
rect -170 -5780 -30 -5690
rect 2320 -6530 2590 -6290
rect -170 -6910 -30 -6810
<< metal3 >>
rect -1710 680 1810 690
rect -1710 560 -1700 680
rect -1540 560 1680 680
rect 1800 560 1810 680
rect -1710 550 1810 560
rect -190 430 -10 440
rect -1890 403 -1710 420
rect -1890 338 -1859 403
rect -1768 390 -1710 403
rect -455 390 -351 403
rect -1768 338 -442 390
rect -1890 325 -442 338
rect -364 325 -351 390
rect -1890 320 -351 325
rect -455 312 -351 320
rect -190 290 -180 430
rect -20 290 -10 430
rect -190 280 -10 290
rect -2639 260 -2470 273
rect -2639 156 -2613 260
rect -2496 247 -897 260
rect -2496 169 -988 247
rect -910 169 -897 247
rect -2496 156 -897 169
rect -320 200 1270 210
rect -2639 143 -2470 156
rect -320 130 -310 200
rect -230 130 1190 200
rect 1260 130 1270 200
rect -320 120 1270 130
rect -728 104 -637 117
rect -728 91 -715 104
rect -2379 78 -715 91
rect -2379 0 -2366 78
rect -2249 26 -715 78
rect -650 26 -637 104
rect -2249 13 -637 26
rect 70 40 350 50
rect -2249 0 -2236 13
rect -2379 -13 -2236 0
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect 2960 -440 3370 -410
rect 2960 -500 2990 -440
rect 1970 -520 2990 -500
rect -3130 -600 240 -590
rect -3130 -660 -3120 -600
rect -3000 -610 240 -600
rect -3000 -660 140 -610
rect -3130 -670 140 -660
rect 220 -670 240 -610
rect 110 -690 240 -670
rect 1970 -680 1990 -520
rect 2160 -680 2990 -520
rect 1970 -690 2990 -680
rect -180 -740 -20 -730
rect -180 -890 -170 -740
rect -30 -890 -20 -740
rect 2960 -750 2990 -690
rect 3340 -750 3370 -440
rect 2960 -760 3370 -750
rect -180 -900 -20 -890
rect 2960 -850 3370 -820
rect -2130 -950 -470 -940
rect -2130 -1020 -2110 -950
rect -2010 -960 -470 -950
rect 40 -950 180 -940
rect 40 -960 80 -950
rect -2010 -1020 80 -960
rect 170 -1020 180 -950
rect 2960 -990 2990 -850
rect -2130 -1030 180 -1020
rect 1480 -1010 2990 -990
rect 1480 -1070 1490 -1010
rect 1550 -1070 2990 -1010
rect 1480 -1090 2990 -1070
rect 2960 -1230 2990 -1090
rect 3340 -1230 3370 -850
rect 2960 -1260 3370 -1230
rect -2630 -1280 400 -1270
rect -2630 -1350 -2620 -1280
rect -2500 -1350 320 -1280
rect 390 -1350 400 -1280
rect -2630 -1360 400 -1350
rect 2310 -1320 2600 -1310
rect -2880 -1560 760 -1550
rect -2880 -1620 -2870 -1560
rect -2750 -1620 690 -1560
rect 750 -1620 760 -1560
rect 2310 -1560 2320 -1320
rect 2590 -1560 2600 -1320
rect 2310 -1570 2600 -1560
rect -2880 -1630 760 -1620
rect -1880 -1710 440 -1700
rect -1880 -1780 -1870 -1710
rect -1750 -1780 360 -1710
rect 430 -1780 440 -1710
rect -1880 -1790 440 -1780
rect -180 -1990 -20 -1980
rect -180 -2130 -170 -1990
rect -30 -2130 -20 -1990
rect -180 -2140 -20 -2130
rect 2960 -2080 3370 -2050
rect 2960 -2190 2990 -2080
rect 1570 -2200 2990 -2190
rect -1880 -2330 450 -2320
rect -1880 -2410 -1870 -2330
rect -1750 -2410 360 -2330
rect 440 -2410 450 -2330
rect 1570 -2350 1580 -2200
rect 1690 -2350 2990 -2200
rect 1570 -2360 2990 -2350
rect -1880 -2420 450 -2410
rect 2960 -2460 2990 -2360
rect 3340 -2460 3370 -2080
rect -2630 -2490 760 -2480
rect 2960 -2490 3370 -2460
rect -2630 -2550 -2620 -2490
rect -2500 -2550 690 -2490
rect 750 -2550 760 -2490
rect -2630 -2560 760 -2550
rect 2310 -2550 2600 -2540
rect 2310 -2790 2320 -2550
rect 2590 -2790 2600 -2550
rect -2380 -2800 760 -2790
rect 2310 -2800 2600 -2790
rect -2380 -2860 -2370 -2800
rect -2250 -2860 690 -2800
rect 750 -2860 760 -2800
rect -2380 -2870 760 -2860
rect -1880 -2940 500 -2930
rect -1880 -3030 -1870 -2940
rect -1750 -3030 400 -2940
rect 490 -3030 500 -2940
rect -1880 -3040 500 -3030
rect -180 -3230 -20 -3220
rect -180 -3390 -170 -3230
rect -30 -3390 -20 -3230
rect -2130 -3440 -240 -3430
rect -2130 -3500 -2120 -3440
rect -2000 -3450 -240 -3440
rect 40 -3440 760 -3430
rect 40 -3450 690 -3440
rect -2000 -3500 690 -3450
rect 750 -3500 760 -3440
rect -2130 -3510 760 -3500
rect -240 -3520 40 -3510
rect -1880 -3580 -300 -3570
rect 100 -3580 480 -3570
rect -1880 -3670 -1870 -3580
rect -1750 -3670 380 -3580
rect 470 -3670 480 -3580
rect -1880 -3680 480 -3670
rect 2310 -3810 2600 -3800
rect 2310 -4050 2320 -3810
rect 2590 -4050 2600 -3810
rect 2310 -4060 2600 -4050
rect -3380 -4100 460 -4090
rect -3380 -4170 -3370 -4100
rect -3250 -4160 380 -4100
rect 450 -4160 460 -4100
rect -3250 -4170 460 -4160
rect -3380 -4180 -3240 -4170
rect 650 -4220 840 -4210
rect 650 -4230 770 -4220
rect -890 -4240 770 -4230
rect -890 -4300 -880 -4240
rect -750 -4280 770 -4240
rect 830 -4280 840 -4220
rect -750 -4290 840 -4280
rect -750 -4300 -740 -4290
rect -890 -4310 -740 -4300
rect -1880 -4360 -950 -4350
rect -1880 -4420 -1870 -4360
rect -1750 -4370 -950 -4360
rect -680 -4360 940 -4350
rect -680 -4370 870 -4360
rect -1750 -4410 870 -4370
rect -1750 -4420 -250 -4410
rect -1880 -4430 -250 -4420
rect 30 -4420 870 -4410
rect 930 -4420 940 -4360
rect 30 -4430 940 -4420
rect -180 -4480 -20 -4470
rect -180 -4620 -170 -4480
rect -30 -4620 -20 -4480
rect -180 -4630 -20 -4620
rect -1880 -4790 950 -4780
rect -1880 -4850 -1870 -4790
rect -1750 -4850 880 -4790
rect 940 -4850 950 -4790
rect -1880 -4860 950 -4850
rect -3130 -4930 420 -4920
rect -3130 -5000 -3120 -4930
rect -3000 -5000 340 -4930
rect 410 -5000 420 -4930
rect -3130 -5010 420 -5000
rect 2310 -5030 2600 -5020
rect 2310 -5270 2320 -5030
rect 2590 -5270 2600 -5030
rect 2310 -5280 2600 -5270
rect -180 -5690 -20 -5680
rect -180 -5780 -170 -5690
rect -30 -5780 -20 -5690
rect -180 -5790 -20 -5780
rect 2310 -6290 2600 -6280
rect 2310 -6530 2320 -6290
rect 2590 -6530 2600 -6290
rect 2310 -6540 2600 -6530
rect -180 -6810 -20 -6800
rect -180 -6910 -170 -6810
rect -30 -6910 -20 -6810
rect -180 -6920 -20 -6910
<< via3 >>
rect -180 420 -20 430
rect -180 300 -170 420
rect -170 300 -30 420
rect -30 300 -20 420
rect -180 290 -20 300
rect 80 -210 340 40
rect -170 -890 -30 -740
rect 2320 -1560 2590 -1320
rect -170 -2130 -30 -1990
rect 2320 -2790 2590 -2550
rect -170 -3380 -30 -3230
rect -170 -3390 -30 -3380
rect 2320 -4050 2590 -3810
rect -170 -4620 -30 -4480
rect 2320 -5270 2590 -5030
rect -170 -5780 -30 -5690
rect 2320 -6530 2590 -6290
rect -170 -6910 -30 -6810
<< metal4 >>
rect -190 430 -10 700
rect -190 290 -180 430
rect -20 290 -10 430
rect -190 -740 -10 290
rect 70 40 350 50
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect -190 -890 -170 -740
rect -30 -890 -10 -740
rect -190 -1990 -10 -890
rect 2310 -1320 2600 -1310
rect 2310 -1560 2320 -1320
rect 2590 -1560 2600 -1320
rect 2310 -1570 2600 -1560
rect -190 -2130 -170 -1990
rect -30 -2130 -10 -1990
rect -190 -3230 -10 -2130
rect 2310 -2550 2600 -2540
rect 2310 -2790 2320 -2550
rect 2590 -2790 2600 -2550
rect 2310 -2800 2600 -2790
rect -190 -3390 -170 -3230
rect -30 -3390 -10 -3230
rect -190 -4480 -10 -3390
rect 2310 -3810 2600 -3800
rect 2310 -4050 2320 -3810
rect 2590 -4050 2600 -3810
rect 2310 -4060 2600 -4050
rect -190 -4620 -170 -4480
rect -30 -4620 -10 -4480
rect -190 -5690 -10 -4620
rect 2310 -5030 2600 -5020
rect 2310 -5270 2320 -5030
rect 2590 -5270 2600 -5030
rect 2310 -5280 2600 -5270
rect -190 -5780 -170 -5690
rect -30 -5780 -10 -5690
rect -190 -6810 -10 -5780
rect 2310 -6290 2600 -6280
rect 2310 -6530 2320 -6290
rect 2590 -6530 2600 -6290
rect 2310 -6540 2600 -6530
rect -190 -6910 -170 -6810
rect -30 -6910 -10 -6810
rect -190 -7030 -10 -6910
<< via4 >>
rect 80 -210 340 40
rect 2320 -1560 2590 -1320
rect 2320 -2790 2590 -2550
rect 2320 -4050 2590 -3810
rect 2320 -5270 2590 -5030
rect 2320 -6530 2590 -6290
<< metal5 >>
rect 2290 70 2620 700
rect -1590 40 2620 70
rect -1590 -210 80 40
rect 340 -210 2620 40
rect -1590 -250 2620 -210
rect 2290 -1320 2620 -250
rect 2290 -1560 2320 -1320
rect 2590 -1560 2620 -1320
rect 2290 -2550 2620 -1560
rect 2290 -2790 2320 -2550
rect 2590 -2790 2620 -2550
rect 2290 -3810 2620 -2790
rect 2290 -4050 2320 -3810
rect 2590 -4050 2620 -3810
rect 2290 -5030 2620 -4050
rect 2290 -5270 2320 -5030
rect 2590 -5270 2620 -5030
rect 2290 -6290 2620 -5270
rect 2290 -6530 2320 -6290
rect 2590 -6530 2620 -6290
rect 2290 -6560 2620 -6530
use sky130_fd_sc_hd__or4_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 488 0 1 -772
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  x2
timestamp 1701704242
transform 1 0 488 0 -1 -858
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 -758 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1040 0 1 -772
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1701704242
transform 1 0 -1034 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1701704242
transform 1 0 -1308 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1701704242
transform 1 0 -1584 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1500 0 1 -772
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1701704242
transform 1 0 -482 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x10
timestamp 1701704242
transform 1 0 488 0 1 -2022
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x11
timestamp 1701704242
transform 1 0 488 0 -1 -2098
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x12
timestamp 1701704242
transform 1 0 488 0 1 -3262
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x13
timestamp 1701704242
transform 1 0 490 0 -1 -3352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x14
timestamp 1701704242
transform 1 0 948 0 -1 -2098
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 488 0 1 -4512
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x16
timestamp 1701704242
transform 1 0 488 0 -1 -4584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  x17
timestamp 1701704242
transform 1 0 1232 0 1 -4512
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x18
timestamp 1701704242
transform 1 0 488 0 1 -5744
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x19
timestamp 1701704242
transform 1 0 488 0 -1 -5818
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 488 0 1 -6982
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x21
timestamp 1701704242
transform 1 0 948 0 1 -6982
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x22
timestamp 1701704242
transform -1 0 1960 0 1 -6982
box -38 -48 590 592
<< labels >>
flabel metal1 -3910 490 -3710 690 0 FreeSans 256 0 0 0 I0
port 3 nsew
flabel metal1 -3660 490 -3460 690 0 FreeSans 256 0 0 0 I1
port 0 nsew
flabel metal1 -3410 490 -3210 690 0 FreeSans 256 0 0 0 I2
port 4 nsew
flabel metal1 -3160 490 -2960 690 0 FreeSans 256 0 0 0 I3
port 2 nsew
flabel metal1 -2910 490 -2710 690 0 FreeSans 256 0 0 0 I4
port 7 nsew
flabel metal1 -2660 490 -2460 690 0 FreeSans 256 0 0 0 I5
port 1 nsew
flabel metal1 -2410 490 -2210 690 0 FreeSans 256 0 0 0 I6
port 5 nsew
flabel metal1 -2160 490 -1960 690 0 FreeSans 256 0 0 0 I7
port 6 nsew
flabel metal1 -1910 490 -1710 690 0 FreeSans 256 0 0 0 EI
port 13 nsew
flabel metal1 3010 -4190 3210 -3990 0 FreeSans 256 0 0 0 A1
port 11 nsew
flabel metal1 3370 -1150 3570 -950 0 FreeSans 256 0 0 0 EO
port 8 nsew
flabel metal1 3370 -700 3570 -500 0 FreeSans 256 0 0 0 GS
port 9 nsew
flabel metal1 3370 -2370 3570 -2170 0 FreeSans 256 0 0 0 A2
port 10 nsew
<< end >>
