magic
tech sky130A
timestamp 1714793356
<< metal1 >>
rect -2200 16045 2920 16265
rect -2205 15020 2915 15515
rect -2200 13995 2920 14490
rect -2200 12975 2920 13470
rect -2200 11950 2920 12445
rect -2200 10930 2920 11425
rect -2200 10385 2920 10405
rect -2200 9910 2925 10385
rect -2195 9890 2925 9910
rect -2195 9360 2925 9380
rect -2195 8885 2930 9360
rect -2190 8865 2930 8885
rect -2195 8340 2925 8360
rect -2195 7865 2930 8340
rect -2190 7845 2930 7865
rect -2205 6840 2915 7335
rect -2200 5815 2920 6310
rect -2200 4795 2920 5290
rect -2200 3770 2920 4265
rect -2200 2750 2920 3245
rect -2195 1710 2920 2225
rect -2190 685 2925 1200
rect -2190 -335 2925 180
rect -2200 -1345 2915 -830
rect -2205 -2085 2915 -1865
use sky130_fd_pr__res_xhigh_po_5p73_2GP8TG  XR1
timestamp 1714792946
transform 1 0 261 0 1 7090
box -2543 -9255 2543 9255
<< end >>
