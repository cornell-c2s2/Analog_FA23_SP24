magic
tech sky130A
magscale 1 2
timestamp 1709390584
<< error_p >>
rect -797 581 -739 587
rect -605 581 -547 587
rect -413 581 -355 587
rect -221 581 -163 587
rect -29 581 29 587
rect 163 581 221 587
rect 355 581 413 587
rect 547 581 605 587
rect 739 581 797 587
rect -797 547 -785 581
rect -605 547 -593 581
rect -413 547 -401 581
rect -221 547 -209 581
rect -29 547 -17 581
rect 163 547 175 581
rect 355 547 367 581
rect 547 547 559 581
rect 739 547 751 581
rect -797 541 -739 547
rect -605 541 -547 547
rect -413 541 -355 547
rect -221 541 -163 547
rect -29 541 29 547
rect 163 541 221 547
rect 355 541 413 547
rect 547 541 605 547
rect 739 541 797 547
rect -893 -547 -835 -541
rect -701 -547 -643 -541
rect -509 -547 -451 -541
rect -317 -547 -259 -541
rect -125 -547 -67 -541
rect 67 -547 125 -541
rect 259 -547 317 -541
rect 451 -547 509 -541
rect 643 -547 701 -541
rect 835 -547 893 -541
rect -893 -581 -881 -547
rect -701 -581 -689 -547
rect -509 -581 -497 -547
rect -317 -581 -305 -547
rect -125 -581 -113 -547
rect 67 -581 79 -547
rect 259 -581 271 -547
rect 451 -581 463 -547
rect 643 -581 655 -547
rect 835 -581 847 -547
rect -893 -587 -835 -581
rect -701 -587 -643 -581
rect -509 -587 -451 -581
rect -317 -587 -259 -581
rect -125 -587 -67 -581
rect 67 -587 125 -581
rect 259 -587 317 -581
rect 451 -587 509 -581
rect 643 -587 701 -581
rect 835 -587 893 -581
<< nwell >>
rect -1079 -719 1079 719
<< pmos >>
rect -879 -500 -849 500
rect -783 -500 -753 500
rect -687 -500 -657 500
rect -591 -500 -561 500
rect -495 -500 -465 500
rect -399 -500 -369 500
rect -303 -500 -273 500
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
rect 273 -500 303 500
rect 369 -500 399 500
rect 465 -500 495 500
rect 561 -500 591 500
rect 657 -500 687 500
rect 753 -500 783 500
rect 849 -500 879 500
<< pdiff >>
rect -941 488 -879 500
rect -941 -488 -929 488
rect -895 -488 -879 488
rect -941 -500 -879 -488
rect -849 488 -783 500
rect -849 -488 -833 488
rect -799 -488 -783 488
rect -849 -500 -783 -488
rect -753 488 -687 500
rect -753 -488 -737 488
rect -703 -488 -687 488
rect -753 -500 -687 -488
rect -657 488 -591 500
rect -657 -488 -641 488
rect -607 -488 -591 488
rect -657 -500 -591 -488
rect -561 488 -495 500
rect -561 -488 -545 488
rect -511 -488 -495 488
rect -561 -500 -495 -488
rect -465 488 -399 500
rect -465 -488 -449 488
rect -415 -488 -399 488
rect -465 -500 -399 -488
rect -369 488 -303 500
rect -369 -488 -353 488
rect -319 -488 -303 488
rect -369 -500 -303 -488
rect -273 488 -207 500
rect -273 -488 -257 488
rect -223 -488 -207 488
rect -273 -500 -207 -488
rect -177 488 -111 500
rect -177 -488 -161 488
rect -127 -488 -111 488
rect -177 -500 -111 -488
rect -81 488 -15 500
rect -81 -488 -65 488
rect -31 -488 -15 488
rect -81 -500 -15 -488
rect 15 488 81 500
rect 15 -488 31 488
rect 65 -488 81 488
rect 15 -500 81 -488
rect 111 488 177 500
rect 111 -488 127 488
rect 161 -488 177 488
rect 111 -500 177 -488
rect 207 488 273 500
rect 207 -488 223 488
rect 257 -488 273 488
rect 207 -500 273 -488
rect 303 488 369 500
rect 303 -488 319 488
rect 353 -488 369 488
rect 303 -500 369 -488
rect 399 488 465 500
rect 399 -488 415 488
rect 449 -488 465 488
rect 399 -500 465 -488
rect 495 488 561 500
rect 495 -488 511 488
rect 545 -488 561 488
rect 495 -500 561 -488
rect 591 488 657 500
rect 591 -488 607 488
rect 641 -488 657 488
rect 591 -500 657 -488
rect 687 488 753 500
rect 687 -488 703 488
rect 737 -488 753 488
rect 687 -500 753 -488
rect 783 488 849 500
rect 783 -488 799 488
rect 833 -488 849 488
rect 783 -500 849 -488
rect 879 488 941 500
rect 879 -488 895 488
rect 929 -488 941 488
rect 879 -500 941 -488
<< pdiffc >>
rect -929 -488 -895 488
rect -833 -488 -799 488
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
rect 799 -488 833 488
rect 895 -488 929 488
<< nsubdiff >>
rect -1043 649 -947 683
rect 947 649 1043 683
rect -1043 587 -1009 649
rect 1009 587 1043 649
rect -1043 -649 -1009 -587
rect 1009 -649 1043 -587
rect -1043 -683 -947 -649
rect 947 -683 1043 -649
<< nsubdiffcont >>
rect -947 649 947 683
rect -1043 -587 -1009 587
rect 1009 -587 1043 587
rect -947 -683 947 -649
<< poly >>
rect -801 581 -735 597
rect -801 547 -785 581
rect -751 547 -735 581
rect -801 531 -735 547
rect -609 581 -543 597
rect -609 547 -593 581
rect -559 547 -543 581
rect -609 531 -543 547
rect -417 581 -351 597
rect -417 547 -401 581
rect -367 547 -351 581
rect -417 531 -351 547
rect -225 581 -159 597
rect -225 547 -209 581
rect -175 547 -159 581
rect -225 531 -159 547
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect 159 581 225 597
rect 159 547 175 581
rect 209 547 225 581
rect 159 531 225 547
rect 351 581 417 597
rect 351 547 367 581
rect 401 547 417 581
rect 351 531 417 547
rect 543 581 609 597
rect 543 547 559 581
rect 593 547 609 581
rect 543 531 609 547
rect 735 581 801 597
rect 735 547 751 581
rect 785 547 801 581
rect 735 531 801 547
rect -879 500 -849 526
rect -783 500 -753 531
rect -687 500 -657 526
rect -591 500 -561 531
rect -495 500 -465 526
rect -399 500 -369 531
rect -303 500 -273 526
rect -207 500 -177 531
rect -111 500 -81 526
rect -15 500 15 531
rect 81 500 111 526
rect 177 500 207 531
rect 273 500 303 526
rect 369 500 399 531
rect 465 500 495 526
rect 561 500 591 531
rect 657 500 687 526
rect 753 500 783 531
rect 849 500 879 526
rect -879 -531 -849 -500
rect -783 -526 -753 -500
rect -687 -531 -657 -500
rect -591 -526 -561 -500
rect -495 -531 -465 -500
rect -399 -526 -369 -500
rect -303 -531 -273 -500
rect -207 -526 -177 -500
rect -111 -531 -81 -500
rect -15 -526 15 -500
rect 81 -531 111 -500
rect 177 -526 207 -500
rect 273 -531 303 -500
rect 369 -526 399 -500
rect 465 -531 495 -500
rect 561 -526 591 -500
rect 657 -531 687 -500
rect 753 -526 783 -500
rect 849 -531 879 -500
rect -897 -547 -831 -531
rect -897 -581 -881 -547
rect -847 -581 -831 -547
rect -897 -597 -831 -581
rect -705 -547 -639 -531
rect -705 -581 -689 -547
rect -655 -581 -639 -547
rect -705 -597 -639 -581
rect -513 -547 -447 -531
rect -513 -581 -497 -547
rect -463 -581 -447 -547
rect -513 -597 -447 -581
rect -321 -547 -255 -531
rect -321 -581 -305 -547
rect -271 -581 -255 -547
rect -321 -597 -255 -581
rect -129 -547 -63 -531
rect -129 -581 -113 -547
rect -79 -581 -63 -547
rect -129 -597 -63 -581
rect 63 -547 129 -531
rect 63 -581 79 -547
rect 113 -581 129 -547
rect 63 -597 129 -581
rect 255 -547 321 -531
rect 255 -581 271 -547
rect 305 -581 321 -547
rect 255 -597 321 -581
rect 447 -547 513 -531
rect 447 -581 463 -547
rect 497 -581 513 -547
rect 447 -597 513 -581
rect 639 -547 705 -531
rect 639 -581 655 -547
rect 689 -581 705 -547
rect 639 -597 705 -581
rect 831 -547 897 -531
rect 831 -581 847 -547
rect 881 -581 897 -547
rect 831 -597 897 -581
<< polycont >>
rect -785 547 -751 581
rect -593 547 -559 581
rect -401 547 -367 581
rect -209 547 -175 581
rect -17 547 17 581
rect 175 547 209 581
rect 367 547 401 581
rect 559 547 593 581
rect 751 547 785 581
rect -881 -581 -847 -547
rect -689 -581 -655 -547
rect -497 -581 -463 -547
rect -305 -581 -271 -547
rect -113 -581 -79 -547
rect 79 -581 113 -547
rect 271 -581 305 -547
rect 463 -581 497 -547
rect 655 -581 689 -547
rect 847 -581 881 -547
<< locali >>
rect -1043 649 -947 683
rect 947 649 1043 683
rect -1043 587 -1009 649
rect 1009 587 1043 649
rect -801 547 -785 581
rect -751 547 -735 581
rect -609 547 -593 581
rect -559 547 -543 581
rect -417 547 -401 581
rect -367 547 -351 581
rect -225 547 -209 581
rect -175 547 -159 581
rect -33 547 -17 581
rect 17 547 33 581
rect 159 547 175 581
rect 209 547 225 581
rect 351 547 367 581
rect 401 547 417 581
rect 543 547 559 581
rect 593 547 609 581
rect 735 547 751 581
rect 785 547 801 581
rect -929 488 -895 504
rect -929 -504 -895 -488
rect -833 488 -799 504
rect -833 -504 -799 -488
rect -737 488 -703 504
rect -737 -504 -703 -488
rect -641 488 -607 504
rect -641 -504 -607 -488
rect -545 488 -511 504
rect -545 -504 -511 -488
rect -449 488 -415 504
rect -449 -504 -415 -488
rect -353 488 -319 504
rect -353 -504 -319 -488
rect -257 488 -223 504
rect -257 -504 -223 -488
rect -161 488 -127 504
rect -161 -504 -127 -488
rect -65 488 -31 504
rect -65 -504 -31 -488
rect 31 488 65 504
rect 31 -504 65 -488
rect 127 488 161 504
rect 127 -504 161 -488
rect 223 488 257 504
rect 223 -504 257 -488
rect 319 488 353 504
rect 319 -504 353 -488
rect 415 488 449 504
rect 415 -504 449 -488
rect 511 488 545 504
rect 511 -504 545 -488
rect 607 488 641 504
rect 607 -504 641 -488
rect 703 488 737 504
rect 703 -504 737 -488
rect 799 488 833 504
rect 799 -504 833 -488
rect 895 488 929 504
rect 895 -504 929 -488
rect -897 -581 -881 -547
rect -847 -581 -831 -547
rect -705 -581 -689 -547
rect -655 -581 -639 -547
rect -513 -581 -497 -547
rect -463 -581 -447 -547
rect -321 -581 -305 -547
rect -271 -581 -255 -547
rect -129 -581 -113 -547
rect -79 -581 -63 -547
rect 63 -581 79 -547
rect 113 -581 129 -547
rect 255 -581 271 -547
rect 305 -581 321 -547
rect 447 -581 463 -547
rect 497 -581 513 -547
rect 639 -581 655 -547
rect 689 -581 705 -547
rect 831 -581 847 -547
rect 881 -581 897 -547
rect -1043 -649 -1009 -587
rect 1009 -649 1043 -587
rect -1043 -683 -947 -649
rect 947 -683 1043 -649
<< viali >>
rect -785 547 -751 581
rect -593 547 -559 581
rect -401 547 -367 581
rect -209 547 -175 581
rect -17 547 17 581
rect 175 547 209 581
rect 367 547 401 581
rect 559 547 593 581
rect 751 547 785 581
rect -929 -488 -895 488
rect -833 -488 -799 488
rect -737 -488 -703 488
rect -641 -488 -607 488
rect -545 -488 -511 488
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect 511 -488 545 488
rect 607 -488 641 488
rect 703 -488 737 488
rect 799 -488 833 488
rect 895 -488 929 488
rect -881 -581 -847 -547
rect -689 -581 -655 -547
rect -497 -581 -463 -547
rect -305 -581 -271 -547
rect -113 -581 -79 -547
rect 79 -581 113 -547
rect 271 -581 305 -547
rect 463 -581 497 -547
rect 655 -581 689 -547
rect 847 -581 881 -547
<< metal1 >>
rect -797 581 -739 587
rect -797 547 -785 581
rect -751 547 -739 581
rect -797 541 -739 547
rect -605 581 -547 587
rect -605 547 -593 581
rect -559 547 -547 581
rect -605 541 -547 547
rect -413 581 -355 587
rect -413 547 -401 581
rect -367 547 -355 581
rect -413 541 -355 547
rect -221 581 -163 587
rect -221 547 -209 581
rect -175 547 -163 581
rect -221 541 -163 547
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect 163 581 221 587
rect 163 547 175 581
rect 209 547 221 581
rect 163 541 221 547
rect 355 581 413 587
rect 355 547 367 581
rect 401 547 413 581
rect 355 541 413 547
rect 547 581 605 587
rect 547 547 559 581
rect 593 547 605 581
rect 547 541 605 547
rect 739 581 797 587
rect 739 547 751 581
rect 785 547 797 581
rect 739 541 797 547
rect -935 488 -889 500
rect -935 -488 -929 488
rect -895 -488 -889 488
rect -935 -500 -889 -488
rect -839 488 -793 500
rect -839 -488 -833 488
rect -799 -488 -793 488
rect -839 -500 -793 -488
rect -743 488 -697 500
rect -743 -488 -737 488
rect -703 -488 -697 488
rect -743 -500 -697 -488
rect -647 488 -601 500
rect -647 -488 -641 488
rect -607 -488 -601 488
rect -647 -500 -601 -488
rect -551 488 -505 500
rect -551 -488 -545 488
rect -511 -488 -505 488
rect -551 -500 -505 -488
rect -455 488 -409 500
rect -455 -488 -449 488
rect -415 -488 -409 488
rect -455 -500 -409 -488
rect -359 488 -313 500
rect -359 -488 -353 488
rect -319 -488 -313 488
rect -359 -500 -313 -488
rect -263 488 -217 500
rect -263 -488 -257 488
rect -223 -488 -217 488
rect -263 -500 -217 -488
rect -167 488 -121 500
rect -167 -488 -161 488
rect -127 -488 -121 488
rect -167 -500 -121 -488
rect -71 488 -25 500
rect -71 -488 -65 488
rect -31 -488 -25 488
rect -71 -500 -25 -488
rect 25 488 71 500
rect 25 -488 31 488
rect 65 -488 71 488
rect 25 -500 71 -488
rect 121 488 167 500
rect 121 -488 127 488
rect 161 -488 167 488
rect 121 -500 167 -488
rect 217 488 263 500
rect 217 -488 223 488
rect 257 -488 263 488
rect 217 -500 263 -488
rect 313 488 359 500
rect 313 -488 319 488
rect 353 -488 359 488
rect 313 -500 359 -488
rect 409 488 455 500
rect 409 -488 415 488
rect 449 -488 455 488
rect 409 -500 455 -488
rect 505 488 551 500
rect 505 -488 511 488
rect 545 -488 551 488
rect 505 -500 551 -488
rect 601 488 647 500
rect 601 -488 607 488
rect 641 -488 647 488
rect 601 -500 647 -488
rect 697 488 743 500
rect 697 -488 703 488
rect 737 -488 743 488
rect 697 -500 743 -488
rect 793 488 839 500
rect 793 -488 799 488
rect 833 -488 839 488
rect 793 -500 839 -488
rect 889 488 935 500
rect 889 -488 895 488
rect 929 -488 935 488
rect 889 -500 935 -488
rect -893 -547 -835 -541
rect -893 -581 -881 -547
rect -847 -581 -835 -547
rect -893 -587 -835 -581
rect -701 -547 -643 -541
rect -701 -581 -689 -547
rect -655 -581 -643 -547
rect -701 -587 -643 -581
rect -509 -547 -451 -541
rect -509 -581 -497 -547
rect -463 -581 -451 -547
rect -509 -587 -451 -581
rect -317 -547 -259 -541
rect -317 -581 -305 -547
rect -271 -581 -259 -547
rect -317 -587 -259 -581
rect -125 -547 -67 -541
rect -125 -581 -113 -547
rect -79 -581 -67 -547
rect -125 -587 -67 -581
rect 67 -547 125 -541
rect 67 -581 79 -547
rect 113 -581 125 -547
rect 67 -587 125 -581
rect 259 -547 317 -541
rect 259 -581 271 -547
rect 305 -581 317 -547
rect 259 -587 317 -581
rect 451 -547 509 -541
rect 451 -581 463 -547
rect 497 -581 509 -547
rect 451 -587 509 -581
rect 643 -547 701 -541
rect 643 -581 655 -547
rect 689 -581 701 -547
rect 643 -587 701 -581
rect 835 -547 893 -541
rect 835 -581 847 -547
rect 881 -581 893 -547
rect 835 -587 893 -581
<< properties >>
string FIXED_BBOX -1026 -666 1026 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 19 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
