magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< nwell >>
rect -941 -719 941 719
<< pmos >>
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
<< pdiff >>
rect -803 459 -745 500
rect -803 425 -791 459
rect -757 425 -745 459
rect -803 391 -745 425
rect -803 357 -791 391
rect -757 357 -745 391
rect -803 323 -745 357
rect -803 289 -791 323
rect -757 289 -745 323
rect -803 255 -745 289
rect -803 221 -791 255
rect -757 221 -745 255
rect -803 187 -745 221
rect -803 153 -791 187
rect -757 153 -745 187
rect -803 119 -745 153
rect -803 85 -791 119
rect -757 85 -745 119
rect -803 51 -745 85
rect -803 17 -791 51
rect -757 17 -745 51
rect -803 -17 -745 17
rect -803 -51 -791 -17
rect -757 -51 -745 -17
rect -803 -85 -745 -51
rect -803 -119 -791 -85
rect -757 -119 -745 -85
rect -803 -153 -745 -119
rect -803 -187 -791 -153
rect -757 -187 -745 -153
rect -803 -221 -745 -187
rect -803 -255 -791 -221
rect -757 -255 -745 -221
rect -803 -289 -745 -255
rect -803 -323 -791 -289
rect -757 -323 -745 -289
rect -803 -357 -745 -323
rect -803 -391 -791 -357
rect -757 -391 -745 -357
rect -803 -425 -745 -391
rect -803 -459 -791 -425
rect -757 -459 -745 -425
rect -803 -500 -745 -459
rect -545 459 -487 500
rect -545 425 -533 459
rect -499 425 -487 459
rect -545 391 -487 425
rect -545 357 -533 391
rect -499 357 -487 391
rect -545 323 -487 357
rect -545 289 -533 323
rect -499 289 -487 323
rect -545 255 -487 289
rect -545 221 -533 255
rect -499 221 -487 255
rect -545 187 -487 221
rect -545 153 -533 187
rect -499 153 -487 187
rect -545 119 -487 153
rect -545 85 -533 119
rect -499 85 -487 119
rect -545 51 -487 85
rect -545 17 -533 51
rect -499 17 -487 51
rect -545 -17 -487 17
rect -545 -51 -533 -17
rect -499 -51 -487 -17
rect -545 -85 -487 -51
rect -545 -119 -533 -85
rect -499 -119 -487 -85
rect -545 -153 -487 -119
rect -545 -187 -533 -153
rect -499 -187 -487 -153
rect -545 -221 -487 -187
rect -545 -255 -533 -221
rect -499 -255 -487 -221
rect -545 -289 -487 -255
rect -545 -323 -533 -289
rect -499 -323 -487 -289
rect -545 -357 -487 -323
rect -545 -391 -533 -357
rect -499 -391 -487 -357
rect -545 -425 -487 -391
rect -545 -459 -533 -425
rect -499 -459 -487 -425
rect -545 -500 -487 -459
rect -287 459 -229 500
rect -287 425 -275 459
rect -241 425 -229 459
rect -287 391 -229 425
rect -287 357 -275 391
rect -241 357 -229 391
rect -287 323 -229 357
rect -287 289 -275 323
rect -241 289 -229 323
rect -287 255 -229 289
rect -287 221 -275 255
rect -241 221 -229 255
rect -287 187 -229 221
rect -287 153 -275 187
rect -241 153 -229 187
rect -287 119 -229 153
rect -287 85 -275 119
rect -241 85 -229 119
rect -287 51 -229 85
rect -287 17 -275 51
rect -241 17 -229 51
rect -287 -17 -229 17
rect -287 -51 -275 -17
rect -241 -51 -229 -17
rect -287 -85 -229 -51
rect -287 -119 -275 -85
rect -241 -119 -229 -85
rect -287 -153 -229 -119
rect -287 -187 -275 -153
rect -241 -187 -229 -153
rect -287 -221 -229 -187
rect -287 -255 -275 -221
rect -241 -255 -229 -221
rect -287 -289 -229 -255
rect -287 -323 -275 -289
rect -241 -323 -229 -289
rect -287 -357 -229 -323
rect -287 -391 -275 -357
rect -241 -391 -229 -357
rect -287 -425 -229 -391
rect -287 -459 -275 -425
rect -241 -459 -229 -425
rect -287 -500 -229 -459
rect -29 459 29 500
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -500 29 -459
rect 229 459 287 500
rect 229 425 241 459
rect 275 425 287 459
rect 229 391 287 425
rect 229 357 241 391
rect 275 357 287 391
rect 229 323 287 357
rect 229 289 241 323
rect 275 289 287 323
rect 229 255 287 289
rect 229 221 241 255
rect 275 221 287 255
rect 229 187 287 221
rect 229 153 241 187
rect 275 153 287 187
rect 229 119 287 153
rect 229 85 241 119
rect 275 85 287 119
rect 229 51 287 85
rect 229 17 241 51
rect 275 17 287 51
rect 229 -17 287 17
rect 229 -51 241 -17
rect 275 -51 287 -17
rect 229 -85 287 -51
rect 229 -119 241 -85
rect 275 -119 287 -85
rect 229 -153 287 -119
rect 229 -187 241 -153
rect 275 -187 287 -153
rect 229 -221 287 -187
rect 229 -255 241 -221
rect 275 -255 287 -221
rect 229 -289 287 -255
rect 229 -323 241 -289
rect 275 -323 287 -289
rect 229 -357 287 -323
rect 229 -391 241 -357
rect 275 -391 287 -357
rect 229 -425 287 -391
rect 229 -459 241 -425
rect 275 -459 287 -425
rect 229 -500 287 -459
rect 487 459 545 500
rect 487 425 499 459
rect 533 425 545 459
rect 487 391 545 425
rect 487 357 499 391
rect 533 357 545 391
rect 487 323 545 357
rect 487 289 499 323
rect 533 289 545 323
rect 487 255 545 289
rect 487 221 499 255
rect 533 221 545 255
rect 487 187 545 221
rect 487 153 499 187
rect 533 153 545 187
rect 487 119 545 153
rect 487 85 499 119
rect 533 85 545 119
rect 487 51 545 85
rect 487 17 499 51
rect 533 17 545 51
rect 487 -17 545 17
rect 487 -51 499 -17
rect 533 -51 545 -17
rect 487 -85 545 -51
rect 487 -119 499 -85
rect 533 -119 545 -85
rect 487 -153 545 -119
rect 487 -187 499 -153
rect 533 -187 545 -153
rect 487 -221 545 -187
rect 487 -255 499 -221
rect 533 -255 545 -221
rect 487 -289 545 -255
rect 487 -323 499 -289
rect 533 -323 545 -289
rect 487 -357 545 -323
rect 487 -391 499 -357
rect 533 -391 545 -357
rect 487 -425 545 -391
rect 487 -459 499 -425
rect 533 -459 545 -425
rect 487 -500 545 -459
rect 745 459 803 500
rect 745 425 757 459
rect 791 425 803 459
rect 745 391 803 425
rect 745 357 757 391
rect 791 357 803 391
rect 745 323 803 357
rect 745 289 757 323
rect 791 289 803 323
rect 745 255 803 289
rect 745 221 757 255
rect 791 221 803 255
rect 745 187 803 221
rect 745 153 757 187
rect 791 153 803 187
rect 745 119 803 153
rect 745 85 757 119
rect 791 85 803 119
rect 745 51 803 85
rect 745 17 757 51
rect 791 17 803 51
rect 745 -17 803 17
rect 745 -51 757 -17
rect 791 -51 803 -17
rect 745 -85 803 -51
rect 745 -119 757 -85
rect 791 -119 803 -85
rect 745 -153 803 -119
rect 745 -187 757 -153
rect 791 -187 803 -153
rect 745 -221 803 -187
rect 745 -255 757 -221
rect 791 -255 803 -221
rect 745 -289 803 -255
rect 745 -323 757 -289
rect 791 -323 803 -289
rect 745 -357 803 -323
rect 745 -391 757 -357
rect 791 -391 803 -357
rect 745 -425 803 -391
rect 745 -459 757 -425
rect 791 -459 803 -425
rect 745 -500 803 -459
<< pdiffc >>
rect -791 425 -757 459
rect -791 357 -757 391
rect -791 289 -757 323
rect -791 221 -757 255
rect -791 153 -757 187
rect -791 85 -757 119
rect -791 17 -757 51
rect -791 -51 -757 -17
rect -791 -119 -757 -85
rect -791 -187 -757 -153
rect -791 -255 -757 -221
rect -791 -323 -757 -289
rect -791 -391 -757 -357
rect -791 -459 -757 -425
rect -533 425 -499 459
rect -533 357 -499 391
rect -533 289 -499 323
rect -533 221 -499 255
rect -533 153 -499 187
rect -533 85 -499 119
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -119 -499 -85
rect -533 -187 -499 -153
rect -533 -255 -499 -221
rect -533 -323 -499 -289
rect -533 -391 -499 -357
rect -533 -459 -499 -425
rect -275 425 -241 459
rect -275 357 -241 391
rect -275 289 -241 323
rect -275 221 -241 255
rect -275 153 -241 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -275 -187 -241 -153
rect -275 -255 -241 -221
rect -275 -323 -241 -289
rect -275 -391 -241 -357
rect -275 -459 -241 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 241 425 275 459
rect 241 357 275 391
rect 241 289 275 323
rect 241 221 275 255
rect 241 153 275 187
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect 241 -187 275 -153
rect 241 -255 275 -221
rect 241 -323 275 -289
rect 241 -391 275 -357
rect 241 -459 275 -425
rect 499 425 533 459
rect 499 357 533 391
rect 499 289 533 323
rect 499 221 533 255
rect 499 153 533 187
rect 499 85 533 119
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -119 533 -85
rect 499 -187 533 -153
rect 499 -255 533 -221
rect 499 -323 533 -289
rect 499 -391 533 -357
rect 499 -459 533 -425
rect 757 425 791 459
rect 757 357 791 391
rect 757 289 791 323
rect 757 221 791 255
rect 757 153 791 187
rect 757 85 791 119
rect 757 17 791 51
rect 757 -51 791 -17
rect 757 -119 791 -85
rect 757 -187 791 -153
rect 757 -255 791 -221
rect 757 -323 791 -289
rect 757 -391 791 -357
rect 757 -459 791 -425
<< nsubdiff >>
rect -905 649 -799 683
rect -765 649 -731 683
rect -697 649 -663 683
rect -629 649 -595 683
rect -561 649 -527 683
rect -493 649 -459 683
rect -425 649 -391 683
rect -357 649 -323 683
rect -289 649 -255 683
rect -221 649 -187 683
rect -153 649 -119 683
rect -85 649 -51 683
rect -17 649 17 683
rect 51 649 85 683
rect 119 649 153 683
rect 187 649 221 683
rect 255 649 289 683
rect 323 649 357 683
rect 391 649 425 683
rect 459 649 493 683
rect 527 649 561 683
rect 595 649 629 683
rect 663 649 697 683
rect 731 649 765 683
rect 799 649 905 683
rect -905 561 -871 649
rect -905 493 -871 527
rect 871 561 905 649
rect -905 425 -871 459
rect -905 357 -871 391
rect -905 289 -871 323
rect -905 221 -871 255
rect -905 153 -871 187
rect -905 85 -871 119
rect -905 17 -871 51
rect -905 -51 -871 -17
rect -905 -119 -871 -85
rect -905 -187 -871 -153
rect -905 -255 -871 -221
rect -905 -323 -871 -289
rect -905 -391 -871 -357
rect -905 -459 -871 -425
rect -905 -527 -871 -493
rect 871 493 905 527
rect 871 425 905 459
rect 871 357 905 391
rect 871 289 905 323
rect 871 221 905 255
rect 871 153 905 187
rect 871 85 905 119
rect 871 17 905 51
rect 871 -51 905 -17
rect 871 -119 905 -85
rect 871 -187 905 -153
rect 871 -255 905 -221
rect 871 -323 905 -289
rect 871 -391 905 -357
rect 871 -459 905 -425
rect -905 -649 -871 -561
rect 871 -527 905 -493
rect 871 -649 905 -561
rect -905 -683 -799 -649
rect -765 -683 -731 -649
rect -697 -683 -663 -649
rect -629 -683 -595 -649
rect -561 -683 -527 -649
rect -493 -683 -459 -649
rect -425 -683 -391 -649
rect -357 -683 -323 -649
rect -289 -683 -255 -649
rect -221 -683 -187 -649
rect -153 -683 -119 -649
rect -85 -683 -51 -649
rect -17 -683 17 -649
rect 51 -683 85 -649
rect 119 -683 153 -649
rect 187 -683 221 -649
rect 255 -683 289 -649
rect 323 -683 357 -649
rect 391 -683 425 -649
rect 459 -683 493 -649
rect 527 -683 561 -649
rect 595 -683 629 -649
rect 663 -683 697 -649
rect 731 -683 765 -649
rect 799 -683 905 -649
<< nsubdiffcont >>
rect -799 649 -765 683
rect -731 649 -697 683
rect -663 649 -629 683
rect -595 649 -561 683
rect -527 649 -493 683
rect -459 649 -425 683
rect -391 649 -357 683
rect -323 649 -289 683
rect -255 649 -221 683
rect -187 649 -153 683
rect -119 649 -85 683
rect -51 649 -17 683
rect 17 649 51 683
rect 85 649 119 683
rect 153 649 187 683
rect 221 649 255 683
rect 289 649 323 683
rect 357 649 391 683
rect 425 649 459 683
rect 493 649 527 683
rect 561 649 595 683
rect 629 649 663 683
rect 697 649 731 683
rect 765 649 799 683
rect -905 527 -871 561
rect 871 527 905 561
rect -905 459 -871 493
rect -905 391 -871 425
rect -905 323 -871 357
rect -905 255 -871 289
rect -905 187 -871 221
rect -905 119 -871 153
rect -905 51 -871 85
rect -905 -17 -871 17
rect -905 -85 -871 -51
rect -905 -153 -871 -119
rect -905 -221 -871 -187
rect -905 -289 -871 -255
rect -905 -357 -871 -323
rect -905 -425 -871 -391
rect -905 -493 -871 -459
rect 871 459 905 493
rect 871 391 905 425
rect 871 323 905 357
rect 871 255 905 289
rect 871 187 905 221
rect 871 119 905 153
rect 871 51 905 85
rect 871 -17 905 17
rect 871 -85 905 -51
rect 871 -153 905 -119
rect 871 -221 905 -187
rect 871 -289 905 -255
rect 871 -357 905 -323
rect 871 -425 905 -391
rect 871 -493 905 -459
rect -905 -561 -871 -527
rect 871 -561 905 -527
rect -799 -683 -765 -649
rect -731 -683 -697 -649
rect -663 -683 -629 -649
rect -595 -683 -561 -649
rect -527 -683 -493 -649
rect -459 -683 -425 -649
rect -391 -683 -357 -649
rect -323 -683 -289 -649
rect -255 -683 -221 -649
rect -187 -683 -153 -649
rect -119 -683 -85 -649
rect -51 -683 -17 -649
rect 17 -683 51 -649
rect 85 -683 119 -649
rect 153 -683 187 -649
rect 221 -683 255 -649
rect 289 -683 323 -649
rect 357 -683 391 -649
rect 425 -683 459 -649
rect 493 -683 527 -649
rect 561 -683 595 -649
rect 629 -683 663 -649
rect 697 -683 731 -649
rect 765 -683 799 -649
<< poly >>
rect -745 581 -545 597
rect -745 547 -696 581
rect -662 547 -628 581
rect -594 547 -545 581
rect -745 500 -545 547
rect -487 581 -287 597
rect -487 547 -438 581
rect -404 547 -370 581
rect -336 547 -287 581
rect -487 500 -287 547
rect -229 581 -29 597
rect -229 547 -180 581
rect -146 547 -112 581
rect -78 547 -29 581
rect -229 500 -29 547
rect 29 581 229 597
rect 29 547 78 581
rect 112 547 146 581
rect 180 547 229 581
rect 29 500 229 547
rect 287 581 487 597
rect 287 547 336 581
rect 370 547 404 581
rect 438 547 487 581
rect 287 500 487 547
rect 545 581 745 597
rect 545 547 594 581
rect 628 547 662 581
rect 696 547 745 581
rect 545 500 745 547
rect -745 -547 -545 -500
rect -745 -581 -696 -547
rect -662 -581 -628 -547
rect -594 -581 -545 -547
rect -745 -597 -545 -581
rect -487 -547 -287 -500
rect -487 -581 -438 -547
rect -404 -581 -370 -547
rect -336 -581 -287 -547
rect -487 -597 -287 -581
rect -229 -547 -29 -500
rect -229 -581 -180 -547
rect -146 -581 -112 -547
rect -78 -581 -29 -547
rect -229 -597 -29 -581
rect 29 -547 229 -500
rect 29 -581 78 -547
rect 112 -581 146 -547
rect 180 -581 229 -547
rect 29 -597 229 -581
rect 287 -547 487 -500
rect 287 -581 336 -547
rect 370 -581 404 -547
rect 438 -581 487 -547
rect 287 -597 487 -581
rect 545 -547 745 -500
rect 545 -581 594 -547
rect 628 -581 662 -547
rect 696 -581 745 -547
rect 545 -597 745 -581
<< polycont >>
rect -696 547 -662 581
rect -628 547 -594 581
rect -438 547 -404 581
rect -370 547 -336 581
rect -180 547 -146 581
rect -112 547 -78 581
rect 78 547 112 581
rect 146 547 180 581
rect 336 547 370 581
rect 404 547 438 581
rect 594 547 628 581
rect 662 547 696 581
rect -696 -581 -662 -547
rect -628 -581 -594 -547
rect -438 -581 -404 -547
rect -370 -581 -336 -547
rect -180 -581 -146 -547
rect -112 -581 -78 -547
rect 78 -581 112 -547
rect 146 -581 180 -547
rect 336 -581 370 -547
rect 404 -581 438 -547
rect 594 -581 628 -547
rect 662 -581 696 -547
<< locali >>
rect -905 649 -799 683
rect -765 649 -731 683
rect -697 649 -663 683
rect -629 649 -595 683
rect -561 649 -527 683
rect -493 649 -459 683
rect -425 649 -391 683
rect -357 649 -323 683
rect -289 649 -255 683
rect -221 649 -187 683
rect -153 649 -119 683
rect -85 649 -51 683
rect -17 649 17 683
rect 51 649 85 683
rect 119 649 153 683
rect 187 649 221 683
rect 255 649 289 683
rect 323 649 357 683
rect 391 649 425 683
rect 459 649 493 683
rect 527 649 561 683
rect 595 649 629 683
rect 663 649 697 683
rect 731 649 765 683
rect 799 649 905 683
rect -905 561 -871 649
rect -745 547 -698 581
rect -662 547 -628 581
rect -592 547 -545 581
rect -487 547 -440 581
rect -404 547 -370 581
rect -334 547 -287 581
rect -229 547 -182 581
rect -146 547 -112 581
rect -76 547 -29 581
rect 29 547 76 581
rect 112 547 146 581
rect 182 547 229 581
rect 287 547 334 581
rect 370 547 404 581
rect 440 547 487 581
rect 545 547 592 581
rect 628 547 662 581
rect 698 547 745 581
rect 871 561 905 649
rect -905 493 -871 527
rect -905 425 -871 459
rect -905 357 -871 391
rect -905 289 -871 323
rect -905 221 -871 255
rect -905 153 -871 187
rect -905 85 -871 119
rect -905 17 -871 51
rect -905 -51 -871 -17
rect -905 -119 -871 -85
rect -905 -187 -871 -153
rect -905 -255 -871 -221
rect -905 -323 -871 -289
rect -905 -391 -871 -357
rect -905 -459 -871 -425
rect -905 -527 -871 -493
rect -791 485 -757 504
rect -791 413 -757 425
rect -791 341 -757 357
rect -791 269 -757 289
rect -791 197 -757 221
rect -791 125 -757 153
rect -791 53 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -53
rect -791 -153 -757 -125
rect -791 -221 -757 -197
rect -791 -289 -757 -269
rect -791 -357 -757 -341
rect -791 -425 -757 -413
rect -791 -504 -757 -485
rect -533 485 -499 504
rect -533 413 -499 425
rect -533 341 -499 357
rect -533 269 -499 289
rect -533 197 -499 221
rect -533 125 -499 153
rect -533 53 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -53
rect -533 -153 -499 -125
rect -533 -221 -499 -197
rect -533 -289 -499 -269
rect -533 -357 -499 -341
rect -533 -425 -499 -413
rect -533 -504 -499 -485
rect -275 485 -241 504
rect -275 413 -241 425
rect -275 341 -241 357
rect -275 269 -241 289
rect -275 197 -241 221
rect -275 125 -241 153
rect -275 53 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -53
rect -275 -153 -241 -125
rect -275 -221 -241 -197
rect -275 -289 -241 -269
rect -275 -357 -241 -341
rect -275 -425 -241 -413
rect -275 -504 -241 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -504 17 -485
rect 241 485 275 504
rect 241 413 275 425
rect 241 341 275 357
rect 241 269 275 289
rect 241 197 275 221
rect 241 125 275 153
rect 241 53 275 85
rect 241 -17 275 17
rect 241 -85 275 -53
rect 241 -153 275 -125
rect 241 -221 275 -197
rect 241 -289 275 -269
rect 241 -357 275 -341
rect 241 -425 275 -413
rect 241 -504 275 -485
rect 499 485 533 504
rect 499 413 533 425
rect 499 341 533 357
rect 499 269 533 289
rect 499 197 533 221
rect 499 125 533 153
rect 499 53 533 85
rect 499 -17 533 17
rect 499 -85 533 -53
rect 499 -153 533 -125
rect 499 -221 533 -197
rect 499 -289 533 -269
rect 499 -357 533 -341
rect 499 -425 533 -413
rect 499 -504 533 -485
rect 757 485 791 504
rect 757 413 791 425
rect 757 341 791 357
rect 757 269 791 289
rect 757 197 791 221
rect 757 125 791 153
rect 757 53 791 85
rect 757 -17 791 17
rect 757 -85 791 -53
rect 757 -153 791 -125
rect 757 -221 791 -197
rect 757 -289 791 -269
rect 757 -357 791 -341
rect 757 -425 791 -413
rect 757 -504 791 -485
rect 871 493 905 527
rect 871 425 905 459
rect 871 357 905 391
rect 871 289 905 323
rect 871 221 905 255
rect 871 153 905 187
rect 871 85 905 119
rect 871 17 905 51
rect 871 -51 905 -17
rect 871 -119 905 -85
rect 871 -187 905 -153
rect 871 -255 905 -221
rect 871 -323 905 -289
rect 871 -391 905 -357
rect 871 -459 905 -425
rect 871 -527 905 -493
rect -905 -649 -871 -561
rect -745 -581 -698 -547
rect -662 -581 -628 -547
rect -592 -581 -545 -547
rect -487 -581 -440 -547
rect -404 -581 -370 -547
rect -334 -581 -287 -547
rect -229 -581 -182 -547
rect -146 -581 -112 -547
rect -76 -581 -29 -547
rect 29 -581 76 -547
rect 112 -581 146 -547
rect 182 -581 229 -547
rect 287 -581 334 -547
rect 370 -581 404 -547
rect 440 -581 487 -547
rect 545 -581 592 -547
rect 628 -581 662 -547
rect 698 -581 745 -547
rect 871 -649 905 -561
rect -905 -683 -799 -649
rect -765 -683 -731 -649
rect -697 -683 -663 -649
rect -629 -683 -595 -649
rect -561 -683 -527 -649
rect -493 -683 -459 -649
rect -425 -683 -391 -649
rect -357 -683 -323 -649
rect -289 -683 -255 -649
rect -221 -683 -187 -649
rect -153 -683 -119 -649
rect -85 -683 -51 -649
rect -17 -683 17 -649
rect 51 -683 85 -649
rect 119 -683 153 -649
rect 187 -683 221 -649
rect 255 -683 289 -649
rect 323 -683 357 -649
rect 391 -683 425 -649
rect 459 -683 493 -649
rect 527 -683 561 -649
rect 595 -683 629 -649
rect 663 -683 697 -649
rect 731 -683 765 -649
rect 799 -683 905 -649
<< viali >>
rect -698 547 -696 581
rect -696 547 -664 581
rect -626 547 -594 581
rect -594 547 -592 581
rect -440 547 -438 581
rect -438 547 -406 581
rect -368 547 -336 581
rect -336 547 -334 581
rect -182 547 -180 581
rect -180 547 -148 581
rect -110 547 -78 581
rect -78 547 -76 581
rect 76 547 78 581
rect 78 547 110 581
rect 148 547 180 581
rect 180 547 182 581
rect 334 547 336 581
rect 336 547 368 581
rect 406 547 438 581
rect 438 547 440 581
rect 592 547 594 581
rect 594 547 626 581
rect 664 547 696 581
rect 696 547 698 581
rect -791 459 -757 485
rect -791 451 -757 459
rect -791 391 -757 413
rect -791 379 -757 391
rect -791 323 -757 341
rect -791 307 -757 323
rect -791 255 -757 269
rect -791 235 -757 255
rect -791 187 -757 197
rect -791 163 -757 187
rect -791 119 -757 125
rect -791 91 -757 119
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -791 -119 -757 -91
rect -791 -125 -757 -119
rect -791 -187 -757 -163
rect -791 -197 -757 -187
rect -791 -255 -757 -235
rect -791 -269 -757 -255
rect -791 -323 -757 -307
rect -791 -341 -757 -323
rect -791 -391 -757 -379
rect -791 -413 -757 -391
rect -791 -459 -757 -451
rect -791 -485 -757 -459
rect -533 459 -499 485
rect -533 451 -499 459
rect -533 391 -499 413
rect -533 379 -499 391
rect -533 323 -499 341
rect -533 307 -499 323
rect -533 255 -499 269
rect -533 235 -499 255
rect -533 187 -499 197
rect -533 163 -499 187
rect -533 119 -499 125
rect -533 91 -499 119
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -533 -119 -499 -91
rect -533 -125 -499 -119
rect -533 -187 -499 -163
rect -533 -197 -499 -187
rect -533 -255 -499 -235
rect -533 -269 -499 -255
rect -533 -323 -499 -307
rect -533 -341 -499 -323
rect -533 -391 -499 -379
rect -533 -413 -499 -391
rect -533 -459 -499 -451
rect -533 -485 -499 -459
rect -275 459 -241 485
rect -275 451 -241 459
rect -275 391 -241 413
rect -275 379 -241 391
rect -275 323 -241 341
rect -275 307 -241 323
rect -275 255 -241 269
rect -275 235 -241 255
rect -275 187 -241 197
rect -275 163 -241 187
rect -275 119 -241 125
rect -275 91 -241 119
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -275 -119 -241 -91
rect -275 -125 -241 -119
rect -275 -187 -241 -163
rect -275 -197 -241 -187
rect -275 -255 -241 -235
rect -275 -269 -241 -255
rect -275 -323 -241 -307
rect -275 -341 -241 -323
rect -275 -391 -241 -379
rect -275 -413 -241 -391
rect -275 -459 -241 -451
rect -275 -485 -241 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 241 459 275 485
rect 241 451 275 459
rect 241 391 275 413
rect 241 379 275 391
rect 241 323 275 341
rect 241 307 275 323
rect 241 255 275 269
rect 241 235 275 255
rect 241 187 275 197
rect 241 163 275 187
rect 241 119 275 125
rect 241 91 275 119
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 241 -119 275 -91
rect 241 -125 275 -119
rect 241 -187 275 -163
rect 241 -197 275 -187
rect 241 -255 275 -235
rect 241 -269 275 -255
rect 241 -323 275 -307
rect 241 -341 275 -323
rect 241 -391 275 -379
rect 241 -413 275 -391
rect 241 -459 275 -451
rect 241 -485 275 -459
rect 499 459 533 485
rect 499 451 533 459
rect 499 391 533 413
rect 499 379 533 391
rect 499 323 533 341
rect 499 307 533 323
rect 499 255 533 269
rect 499 235 533 255
rect 499 187 533 197
rect 499 163 533 187
rect 499 119 533 125
rect 499 91 533 119
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 499 -119 533 -91
rect 499 -125 533 -119
rect 499 -187 533 -163
rect 499 -197 533 -187
rect 499 -255 533 -235
rect 499 -269 533 -255
rect 499 -323 533 -307
rect 499 -341 533 -323
rect 499 -391 533 -379
rect 499 -413 533 -391
rect 499 -459 533 -451
rect 499 -485 533 -459
rect 757 459 791 485
rect 757 451 791 459
rect 757 391 791 413
rect 757 379 791 391
rect 757 323 791 341
rect 757 307 791 323
rect 757 255 791 269
rect 757 235 791 255
rect 757 187 791 197
rect 757 163 791 187
rect 757 119 791 125
rect 757 91 791 119
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect 757 -119 791 -91
rect 757 -125 791 -119
rect 757 -187 791 -163
rect 757 -197 791 -187
rect 757 -255 791 -235
rect 757 -269 791 -255
rect 757 -323 791 -307
rect 757 -341 791 -323
rect 757 -391 791 -379
rect 757 -413 791 -391
rect 757 -459 791 -451
rect 757 -485 791 -459
rect -698 -581 -696 -547
rect -696 -581 -664 -547
rect -626 -581 -594 -547
rect -594 -581 -592 -547
rect -440 -581 -438 -547
rect -438 -581 -406 -547
rect -368 -581 -336 -547
rect -336 -581 -334 -547
rect -182 -581 -180 -547
rect -180 -581 -148 -547
rect -110 -581 -78 -547
rect -78 -581 -76 -547
rect 76 -581 78 -547
rect 78 -581 110 -547
rect 148 -581 180 -547
rect 180 -581 182 -547
rect 334 -581 336 -547
rect 336 -581 368 -547
rect 406 -581 438 -547
rect 438 -581 440 -547
rect 592 -581 594 -547
rect 594 -581 626 -547
rect 664 -581 696 -547
rect 696 -581 698 -547
<< metal1 >>
rect -741 581 -549 587
rect -741 547 -698 581
rect -664 547 -626 581
rect -592 547 -549 581
rect -741 541 -549 547
rect -483 581 -291 587
rect -483 547 -440 581
rect -406 547 -368 581
rect -334 547 -291 581
rect -483 541 -291 547
rect -225 581 -33 587
rect -225 547 -182 581
rect -148 547 -110 581
rect -76 547 -33 581
rect -225 541 -33 547
rect 33 581 225 587
rect 33 547 76 581
rect 110 547 148 581
rect 182 547 225 581
rect 33 541 225 547
rect 291 581 483 587
rect 291 547 334 581
rect 368 547 406 581
rect 440 547 483 581
rect 291 541 483 547
rect 549 581 741 587
rect 549 547 592 581
rect 626 547 664 581
rect 698 547 741 581
rect 549 541 741 547
rect -797 485 -751 500
rect -797 451 -791 485
rect -757 451 -751 485
rect -797 413 -751 451
rect -797 379 -791 413
rect -757 379 -751 413
rect -797 341 -751 379
rect -797 307 -791 341
rect -757 307 -751 341
rect -797 269 -751 307
rect -797 235 -791 269
rect -757 235 -751 269
rect -797 197 -751 235
rect -797 163 -791 197
rect -757 163 -751 197
rect -797 125 -751 163
rect -797 91 -791 125
rect -757 91 -751 125
rect -797 53 -751 91
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -91 -751 -53
rect -797 -125 -791 -91
rect -757 -125 -751 -91
rect -797 -163 -751 -125
rect -797 -197 -791 -163
rect -757 -197 -751 -163
rect -797 -235 -751 -197
rect -797 -269 -791 -235
rect -757 -269 -751 -235
rect -797 -307 -751 -269
rect -797 -341 -791 -307
rect -757 -341 -751 -307
rect -797 -379 -751 -341
rect -797 -413 -791 -379
rect -757 -413 -751 -379
rect -797 -451 -751 -413
rect -797 -485 -791 -451
rect -757 -485 -751 -451
rect -797 -500 -751 -485
rect -539 485 -493 500
rect -539 451 -533 485
rect -499 451 -493 485
rect -539 413 -493 451
rect -539 379 -533 413
rect -499 379 -493 413
rect -539 341 -493 379
rect -539 307 -533 341
rect -499 307 -493 341
rect -539 269 -493 307
rect -539 235 -533 269
rect -499 235 -493 269
rect -539 197 -493 235
rect -539 163 -533 197
rect -499 163 -493 197
rect -539 125 -493 163
rect -539 91 -533 125
rect -499 91 -493 125
rect -539 53 -493 91
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -91 -493 -53
rect -539 -125 -533 -91
rect -499 -125 -493 -91
rect -539 -163 -493 -125
rect -539 -197 -533 -163
rect -499 -197 -493 -163
rect -539 -235 -493 -197
rect -539 -269 -533 -235
rect -499 -269 -493 -235
rect -539 -307 -493 -269
rect -539 -341 -533 -307
rect -499 -341 -493 -307
rect -539 -379 -493 -341
rect -539 -413 -533 -379
rect -499 -413 -493 -379
rect -539 -451 -493 -413
rect -539 -485 -533 -451
rect -499 -485 -493 -451
rect -539 -500 -493 -485
rect -281 485 -235 500
rect -281 451 -275 485
rect -241 451 -235 485
rect -281 413 -235 451
rect -281 379 -275 413
rect -241 379 -235 413
rect -281 341 -235 379
rect -281 307 -275 341
rect -241 307 -235 341
rect -281 269 -235 307
rect -281 235 -275 269
rect -241 235 -235 269
rect -281 197 -235 235
rect -281 163 -275 197
rect -241 163 -235 197
rect -281 125 -235 163
rect -281 91 -275 125
rect -241 91 -235 125
rect -281 53 -235 91
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -91 -235 -53
rect -281 -125 -275 -91
rect -241 -125 -235 -91
rect -281 -163 -235 -125
rect -281 -197 -275 -163
rect -241 -197 -235 -163
rect -281 -235 -235 -197
rect -281 -269 -275 -235
rect -241 -269 -235 -235
rect -281 -307 -235 -269
rect -281 -341 -275 -307
rect -241 -341 -235 -307
rect -281 -379 -235 -341
rect -281 -413 -275 -379
rect -241 -413 -235 -379
rect -281 -451 -235 -413
rect -281 -485 -275 -451
rect -241 -485 -235 -451
rect -281 -500 -235 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 235 485 281 500
rect 235 451 241 485
rect 275 451 281 485
rect 235 413 281 451
rect 235 379 241 413
rect 275 379 281 413
rect 235 341 281 379
rect 235 307 241 341
rect 275 307 281 341
rect 235 269 281 307
rect 235 235 241 269
rect 275 235 281 269
rect 235 197 281 235
rect 235 163 241 197
rect 275 163 281 197
rect 235 125 281 163
rect 235 91 241 125
rect 275 91 281 125
rect 235 53 281 91
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -91 281 -53
rect 235 -125 241 -91
rect 275 -125 281 -91
rect 235 -163 281 -125
rect 235 -197 241 -163
rect 275 -197 281 -163
rect 235 -235 281 -197
rect 235 -269 241 -235
rect 275 -269 281 -235
rect 235 -307 281 -269
rect 235 -341 241 -307
rect 275 -341 281 -307
rect 235 -379 281 -341
rect 235 -413 241 -379
rect 275 -413 281 -379
rect 235 -451 281 -413
rect 235 -485 241 -451
rect 275 -485 281 -451
rect 235 -500 281 -485
rect 493 485 539 500
rect 493 451 499 485
rect 533 451 539 485
rect 493 413 539 451
rect 493 379 499 413
rect 533 379 539 413
rect 493 341 539 379
rect 493 307 499 341
rect 533 307 539 341
rect 493 269 539 307
rect 493 235 499 269
rect 533 235 539 269
rect 493 197 539 235
rect 493 163 499 197
rect 533 163 539 197
rect 493 125 539 163
rect 493 91 499 125
rect 533 91 539 125
rect 493 53 539 91
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -91 539 -53
rect 493 -125 499 -91
rect 533 -125 539 -91
rect 493 -163 539 -125
rect 493 -197 499 -163
rect 533 -197 539 -163
rect 493 -235 539 -197
rect 493 -269 499 -235
rect 533 -269 539 -235
rect 493 -307 539 -269
rect 493 -341 499 -307
rect 533 -341 539 -307
rect 493 -379 539 -341
rect 493 -413 499 -379
rect 533 -413 539 -379
rect 493 -451 539 -413
rect 493 -485 499 -451
rect 533 -485 539 -451
rect 493 -500 539 -485
rect 751 485 797 500
rect 751 451 757 485
rect 791 451 797 485
rect 751 413 797 451
rect 751 379 757 413
rect 791 379 797 413
rect 751 341 797 379
rect 751 307 757 341
rect 791 307 797 341
rect 751 269 797 307
rect 751 235 757 269
rect 791 235 797 269
rect 751 197 797 235
rect 751 163 757 197
rect 791 163 797 197
rect 751 125 797 163
rect 751 91 757 125
rect 791 91 797 125
rect 751 53 797 91
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -91 797 -53
rect 751 -125 757 -91
rect 791 -125 797 -91
rect 751 -163 797 -125
rect 751 -197 757 -163
rect 791 -197 797 -163
rect 751 -235 797 -197
rect 751 -269 757 -235
rect 791 -269 797 -235
rect 751 -307 797 -269
rect 751 -341 757 -307
rect 791 -341 797 -307
rect 751 -379 797 -341
rect 751 -413 757 -379
rect 791 -413 797 -379
rect 751 -451 797 -413
rect 751 -485 757 -451
rect 791 -485 797 -451
rect 751 -500 797 -485
rect -741 -547 -549 -541
rect -741 -581 -698 -547
rect -664 -581 -626 -547
rect -592 -581 -549 -547
rect -741 -587 -549 -581
rect -483 -547 -291 -541
rect -483 -581 -440 -547
rect -406 -581 -368 -547
rect -334 -581 -291 -547
rect -483 -587 -291 -581
rect -225 -547 -33 -541
rect -225 -581 -182 -547
rect -148 -581 -110 -547
rect -76 -581 -33 -547
rect -225 -587 -33 -581
rect 33 -547 225 -541
rect 33 -581 76 -547
rect 110 -581 148 -547
rect 182 -581 225 -547
rect 33 -587 225 -581
rect 291 -547 483 -541
rect 291 -581 334 -547
rect 368 -581 406 -547
rect 440 -581 483 -547
rect 291 -587 483 -581
rect 549 -547 741 -541
rect 549 -581 592 -547
rect 626 -581 664 -547
rect 698 -581 741 -547
rect 549 -587 741 -581
<< properties >>
string FIXED_BBOX -888 -666 888 666
<< end >>
