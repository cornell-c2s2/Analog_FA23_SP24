* NGSPICE file created from 16to4_PriorityEncoder_v0p0p1_flat.ext - technology: sky130A

.subckt 16to4_PriorityEncoder_v0p0p1_flat I15 I14 I11 I10 I4 I0 A3 I8 I6 I3 I1 A2
+ I9 I2 I12 I5 A1 A0 I13 I7 EI GND VDD
X0 x36.Y x36.A VDD.t427 VDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 A2.t120 x36.Y VDD.t387 VDD.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VDD.t250 x22.A x22.Y VDD.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 A2.t119 x36.Y VDD.t385 VDD.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_6111_n9215# x3.x2.X a_6029_n9459# VDD.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VDD.t425 x36.A x36.Y VDD.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VDD.t383 x36.Y A2.t118 VDD.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 x3.x18.C I2.t0 VDD.t457 VDD.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 a_5751_n6397# x5.x18.C a_5645_n6397# GND.t84 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 x29.A x28.A VDD.t781 VDD.t780 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 A0.t127 x22.Y VDD.t218 VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 GND.t219 x22.Y A0.t63 GND.t218 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VDD.t216 x22.Y A0.t126 VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VDD.t88 I12.t0 a_5507_n2647# VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 x5.x19.C I12.t1 GND.t456 GND.t455 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X15 x5.x22.A a_5509_n4211# VDD.t555 VDD.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X16 VDD.t929 x29.Y A1.t127 VDD.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VDD.t927 x29.Y A1.t126 VDD.t926 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VDD.t796 I12.t2 a_5725_n1939# VDD.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X19 GND.t61 I15.t0 a_5595_n4211# GND.t60 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 A1.t125 x29.Y VDD.t925 VDD.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 A1.t124 x29.Y VDD.t923 VDD.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 GND.t217 x22.Y A0.t62 GND.t216 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 GND.t499 x5.x17.A a_5935_n3179# GND.t498 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X24 A0.t61 x22.Y GND.t215 GND.t214 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VDD.t214 x22.Y A0.t125 VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 GND.t766 x5.x21.B a_6053_n7607# GND.t765 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X27 a_5935_n3179# x5.x22.A GND.t401 GND.t400 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X28 GND.t908 x29.Y A1.t63 GND.t907 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 GND.t391 x36.Y A2.t30 GND.t390 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 x3.x19.X a_5475_n14689# GND.t579 GND.t578 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X31 VDD.t474 EI.t0 a_5475_n7635# VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X32 VDD.t212 x22.Y A0.t124 VDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 A0.t123 x22.Y VDD.t210 VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 GND.t906 x29.Y A1.t62 GND.t905 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 A2.t15 x36.Y GND.t389 GND.t388 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 x29.Y x29.A GND.t36 GND.t35 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 a_5645_n5165# x5.x19.C a_5557_n5165# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X38 a_10858_n5725# x3.A2 a_10776_n5725# VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X39 VDD.t381 x36.Y A2.t117 VDD.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X40 a_5557_n13455# I3.t0 a_5475_n13455# GND.t576 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X41 GND.t433 x36.A x36.Y GND.t432 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X42 a_5725_n9215# I1.t0 a_5653_n9215# VDD.t562 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X43 VDD.t597 I3.t1 a_5475_n14689# VDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X44 A3.t63 x43.Y GND.t730 GND.t729 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X45 a_6183_n9215# x3.x1.X a_6111_n9215# VDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X46 a_6469_n12955# x3.x22.A a_6397_n12955# VDD.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X47 x3.GS a_6519_n9437# GND.t558 GND.t557 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X48 GND.t904 x29.Y A1.t61 GND.t903 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X49 A1.t60 x29.Y GND.t902 GND.t901 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X50 A2.t116 x36.Y VDD.t379 VDD.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X51 VDD.t423 x36.A x36.Y VDD.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X52 GND.t543 x3.x4.A a_6029_n9459# GND.t542 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X53 A3.t127 x43.Y VDD.t749 VDD.t748 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X54 A3.t62 x43.Y GND.t728 GND.t727 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X55 A3.t61 x43.Y GND.t726 GND.t725 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X56 x3.GS a_6519_n9437# VDD.t571 VDD.t570 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X57 A0.t60 x22.Y GND.t213 GND.t212 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X58 A1.t59 x29.Y GND.t900 GND.t899 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X59 VDD.t779 x28.A x29.A VDD.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X60 GND.t577 x3.EI a_5751_n13455# GND.t576 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X61 x3.x11.X a_5507_n10997# VDD.t488 VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X62 a_5475_n14689# x3.EI VDD.t589 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X63 a_5967_n15647# x3.EI VDD.t588 VDD.t587 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X64 A3.t126 x43.Y VDD.t747 VDD.t746 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X65 A3.t125 x43.Y VDD.t745 VDD.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X66 x5.A2 a_5935_n3179# VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X67 GND.t898 x29.Y A1.t58 GND.t897 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X68 A0.t122 x22.Y VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X69 GND.t444 I14.t0 a_5475_n1939# GND.t68 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X70 A0.t59 x22.Y GND.t211 GND.t210 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 a_6301_n4915# x5.x16.X a_6219_n4915# VDD.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X72 GND.t209 x22.Y A0.t58 GND.t208 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X73 GND.t259 I4.t0 a_5593_n10687# GND.t255 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X74 GND.t896 x29.Y A1.t57 GND.t895 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X75 GND.t468 EI.t1 a_5629_n7635# GND.t467 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X76 A1.t123 x29.Y VDD.t921 VDD.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X77 a_6219_n4915# x5.x22.A GND.t399 GND.t398 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X78 VDD.t75 x3.x19.D a_5475_n14689# VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X79 A3.t60 x43.Y GND.t724 GND.t723 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X80 A3.t59 x43.Y GND.t722 GND.t721 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X81 x35.A x34.A GND.t458 GND.t457 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X82 a_5653_n1175# I10.t0 a_5557_n1175# VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X83 x1.A a_6219_n4915# VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X84 A0.t121 x22.Y VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X85 GND.t397 x5.x22.A a_6395_n7385# GND.t396 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X86 x3.x19.C I4.t1 GND.t261 GND.t260 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X87 GND.t207 x22.Y A0.t57 GND.t206 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X88 VDD.t204 x22.Y A0.t120 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X89 GND.t720 x43.Y A3.t58 GND.t719 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X90 GND.t718 x43.Y A3.t57 GND.t717 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X91 a_5509_n4211# EI.t2 VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X92 A2.t14 x36.Y GND.t387 GND.t386 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X93 GND.t205 x22.Y A0.t56 GND.t204 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X94 A3.t124 x43.Y VDD.t743 VDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 A3.t123 x43.Y VDD.t741 VDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X96 a_5557_n1939# I15.t1 a_5475_n1939# VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X97 x35.A x34.A VDD.t453 VDD.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X98 A3.t56 x43.Y GND.t716 GND.t715 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X99 VDD.t504 I1.t1 a_5475_n14437# VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X100 A0.t55 x22.Y GND.t203 GND.t202 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X101 VDD.t202 x22.Y A0.t119 VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X102 VDD.t739 x43.Y A3.t122 VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X103 VDD.t737 x43.Y A3.t121 VDD.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X104 GND.t754 x3.x22.A a_6395_n15425# GND.t753 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X105 GND.t34 x29.A x29.Y GND.t33 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X106 A2.t115 x36.Y VDD.t377 VDD.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X107 x5.x17.A a_5507_n3887# GND.t585 GND.t584 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X108 x5.x20.X a_5475_n7635# GND.t470 GND.t469 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X109 VDD.t200 x22.Y A0.t118 VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 A0.t54 x22.Y GND.t201 GND.t200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X111 A0.t117 x22.Y VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X112 A3.t120 x43.Y VDD.t735 VDD.t734 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X113 A1.t122 x29.Y VDD.t919 VDD.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X114 GND.t199 x22.Y A0.t53 GND.t198 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X115 x5.x18.C I10.t1 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X116 VDD.t917 x29.Y A1.t121 VDD.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X117 VDD.t915 x29.Y A1.t120 VDD.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X118 a_5475_n14437# x3.x19.C VDD.t605 VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X119 x1.A a_6219_n4915# GND.t59 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X120 GND.t556 I4.t2 a_5475_n9979# GND.t257 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X121 A0.t116 x22.Y VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X122 VDD.t440 I14.t1 a_5507_n3887# VDD.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 GND.t487 EI.t3 a_6605_n1397# GND.t486 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X124 A3.t55 x43.Y GND.t714 GND.t713 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X125 x36.Y x36.A GND.t431 GND.t430 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X126 A2.t2 x36.Y GND.t385 GND.t384 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X127 VDD.t196 x22.Y A0.t115 VDD.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X128 A2.t1 x36.Y GND.t383 GND.t382 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X129 a_6519_n1397# x5.EO VDD.t787 VDD.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X130 A0.t52 x22.Y GND.t197 GND.t196 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X131 a_5593_n2957# EI.t4 a_5507_n2957# GND.t57 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X132 GND.t429 x36.A x36.Y GND.t428 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X133 GND.t381 x36.Y A2.t0 GND.t380 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X134 GND.t379 x36.Y A2.t32 GND.t378 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X135 GND.t195 x22.Y A0.t51 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X136 GND.t537 x5.x15.X a_6219_n4915# GND.t398 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X137 VDD.t913 x29.Y A1.t119 VDD.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 GND.t712 x43.Y A3.t54 GND.t711 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X139 a_5475_n5165# x5.x16.C VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X140 x22.Y x22.A GND.t251 GND.t250 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X141 A3.t119 x43.Y VDD.t733 VDD.t732 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X142 a_5645_n6397# I9.t0 a_5557_n6397# GND.t84 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X143 x29.Y x29.A VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X144 x36.Y x36.A VDD.t421 VDD.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X145 A2.t114 x36.Y VDD.t375 VDD.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X146 A2.t113 x36.Y VDD.t373 VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X147 a_6395_n7385# x5.x21.X GND.t501 GND.t500 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X148 VDD.t553 I0.t0 a_5725_n9215# VDD.t552 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X149 VDD.t50 x1.A a_10858_n9865# VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X150 A0.t50 x22.Y GND.t193 GND.t192 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X151 A0.t114 x22.Y VDD.t194 VDD.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X152 VDD.t419 x36.A x36.Y VDD.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X153 VDD.t371 x36.Y A2.t112 VDD.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X154 VDD.t369 x36.Y A2.t111 VDD.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X155 GND.t191 x22.Y A0.t49 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X156 VDD.t73 x3.x19.D a_5475_n14437# VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X157 VDD.t481 x5.x4.A a_6183_n1175# VDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X158 GND.t377 x36.Y A2.t31 GND.t376 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X159 VDD.t192 x22.Y A0.t113 VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X160 x3.A2 a_5935_n11219# GND.t466 GND.t465 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X161 VDD.t731 x43.Y A3.t118 VDD.t730 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X162 x22.Y x22.A VDD.t248 VDD.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X163 VDD.t911 x29.Y A1.t118 VDD.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X164 A0.t112 x22.Y VDD.t190 VDD.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X165 A1.t117 x29.Y VDD.t909 VDD.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X166 GND.t910 x5.x14.A a_5935_n3179# GND.t909 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 VDD.t367 x36.Y A2.t110 VDD.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X168 x21.A x2.X GND.t548 GND.t547 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X169 VDD.t188 x22.Y A0.t111 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X170 x5.x19.X a_5475_n6649# GND.t54 GND.t53 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X171 GND.t38 x5.x2.X a_6029_n1419# GND.t37 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X172 GND.t375 x36.Y A2.t10 GND.t374 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X173 x5.x2.X a_5475_n1939# GND.t393 GND.t392 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X174 GND.t373 x36.Y A2.t9 GND.t372 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X175 VDD.t905 x29.Y A1.t116 VDD.t904 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X176 VDD.t907 x29.Y A1.t115 VDD.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X177 x22.Y x22.A GND.t249 GND.t248 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X178 x36.Y x36.A GND.t427 GND.t426 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X179 x29.Y x29.A VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X180 A1.t114 x29.Y VDD.t903 VDD.t902 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X181 A1.t113 x29.Y VDD.t901 VDD.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X182 x21.A x2.X VDD.t561 VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X183 a_6605_n9437# x3.EO a_6519_n9437# GND.t476 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X184 GND.t189 x22.Y A0.t48 GND.t188 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X185 VDD.t365 x36.Y A2.t109 VDD.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 VDD.t363 x36.Y A2.t108 VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X187 GND.t425 x36.A x36.Y GND.t424 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X188 GND.t371 x36.Y A2.t8 GND.t370 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X189 A0.t47 x22.Y GND.t187 GND.t186 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X190 x36.Y x36.A VDD.t417 VDD.t416 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X191 x2.A a_6395_n7385# GND.t460 GND.t459 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X192 x22.Y x22.A VDD.t246 VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X193 a_5475_n9215# I1.t2 GND.t743 GND.t71 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X194 a_5557_n13205# I2.t1 a_5475_n13205# GND.t564 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X195 x36.Y x36.A GND.t423 GND.t422 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X196 GND.t32 x29.A x29.Y GND.t31 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X197 VDD.t186 x22.Y A0.t110 VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X198 A0.t109 x22.Y VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 VDD.t415 x36.A x36.Y VDD.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X200 VDD.t361 x36.Y A2.t107 VDD.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X201 A3.t53 x43.Y GND.t710 GND.t709 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X202 A1.t56 x29.Y GND.t894 GND.t893 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X203 GND.t536 x43.A x43.Y GND.t535 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X204 x36.Y x36.A VDD.t413 VDD.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X205 VDD.t604 x3.x19.C a_5475_n13455# VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X206 x43.Y x43.A GND.t534 GND.t533 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X207 a_5653_n1939# I14.t2 a_5557_n1939# VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X208 GND.t185 x22.Y A0.t46 GND.t184 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X209 A1.t112 x29.Y VDD.t899 VDD.t898 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X210 A3.t117 x43.Y VDD.t729 VDD.t728 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X211 a_5475_n9979# I7.t0 GND.t586 GND.t257 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X212 GND.t575 x3.EI a_5751_n13205# GND.t564 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X213 VDD.t548 x43.A x43.Y VDD.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X214 a_5935_n3179# x5.x11.X GND.t472 GND.t471 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X215 a_5507_n11927# x3.EI VDD.t586 VDD.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X216 x43.Y x43.A VDD.t546 VDD.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X217 VDD.t180 x22.Y A0.t108 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X218 A1.t55 x29.Y GND.t892 GND.t891 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X219 A0.t45 x22.Y GND.t183 GND.t182 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X220 GND.t30 x29.A x29.Y GND.t29 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X221 GND.t421 x36.A x36.Y GND.t420 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X222 a_5475_n13455# I3.t2 VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X223 A0.t44 x22.Y GND.t181 GND.t180 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X224 x5.x14.A a_5507_n2647# GND.t595 GND.t594 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X225 a_5557_n9215# I3.t3 a_5475_n9215# VDD.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X226 GND.t179 x22.Y A0.t43 GND.t178 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X227 VDD.t82 x5.x19.C a_5475_n5415# VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X228 a_5751_n14689# x3.x19.C a_5645_n14689# GND.t75 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X229 A0.t107 x22.Y VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X230 GND.t706 x43.Y A3.t52 GND.t705 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X231 GND.t708 x43.Y A3.t51 GND.t707 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X232 GND.t704 x43.Y A3.t50 GND.t703 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X233 VDD.t411 x36.A x36.Y VDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 x3.x16.C I5.t0 GND.t435 GND.t434 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X235 x3.x16.X a_5475_n13455# GND.t912 GND.t911 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X236 A0.t106 x22.Y VDD.t176 VDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X237 x5.x14.A a_5507_n2647# VDD.t613 VDD.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X238 GND.t177 x22.Y A0.t42 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X239 VDD.t174 x22.Y A0.t105 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X240 A3.t49 x43.Y GND.t702 GND.t701 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X241 VDD.t725 x43.Y A3.t116 VDD.t724 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X242 VDD.t585 x3.EI a_5475_n13455# VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X243 x3.A1 a_6219_n12955# GND.t744 GND.t73 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X244 VDD.t727 x43.Y A3.t115 VDD.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X245 VDD.t723 x43.Y A3.t114 VDD.t722 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X246 GND.t700 x43.Y A3.t48 GND.t699 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X247 GND.t698 x43.Y A3.t47 GND.t697 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X248 VDD.t1 x3.x21.B a_5967_n15647# VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X249 x43.Y x43.A GND.t532 GND.t531 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X250 a_5475_n15675# x3.x19.D VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X251 x22.Y x22.A GND.t247 GND.t246 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X252 GND.t581 EI.t5 a_5751_n5165# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X253 VDD.t172 x22.Y A0.t104 VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X254 x29.A x28.A GND.t762 GND.t761 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X255 GND.t530 x43.A x43.Y GND.t529 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X256 A3.t113 x43.Y VDD.t721 VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X257 GND.t175 x22.Y A0.t41 GND.t174 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X258 VDD.t719 x43.Y A3.t112 VDD.t718 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X259 VDD.t717 x43.Y A3.t111 VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X260 a_5967_n7607# EI.t6 VDD.t391 VDD.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X261 x43.Y x43.A VDD.t544 VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X262 A0.t40 x22.Y GND.t173 GND.t172 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X263 VDD.t897 x29.Y A1.t111 VDD.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X264 a_5475_n1939# I13.t0 GND.t473 GND.t68 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X265 x22.Y x22.A VDD.t244 VDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X266 VDD.t542 x43.A x43.Y VDD.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X267 GND.t696 x43.Y A3.t46 GND.t695 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X268 GND.t694 x43.Y A3.t45 GND.t693 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X269 A1.t110 x29.Y VDD.t895 VDD.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X270 GND.t245 x22.A x22.Y GND.t244 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X271 GND.t760 x28.A x29.A GND.t759 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X272 x5.x4.A EI.t7 GND.t395 GND.t394 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X273 A1.t109 x29.Y VDD.t893 VDD.t892 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X274 a_6397_n12955# x3.x15.X a_6301_n12955# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X275 VDD.t170 x22.Y A0.t103 VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X276 A0.t39 x22.Y GND.t171 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X277 A0.t102 x22.Y VDD.t168 VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X278 GND.t419 x36.A x36.Y GND.t418 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X279 GND.t169 x22.Y A0.t38 GND.t168 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X280 VDD.t715 x43.Y A3.t110 VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X281 VDD.t713 x43.Y A3.t109 VDD.t712 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X282 VDD.t242 x22.A x22.Y VDD.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X283 GND.t497 x5.x17.A a_6219_n4915# GND.t398 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X284 GND.t692 x43.Y A3.t44 GND.t691 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X285 a_5557_n5165# I10.t2 a_5475_n5165# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X286 a_5507_n10997# x3.EI VDD.t584 VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X287 A3.t43 x43.Y GND.t690 GND.t689 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X288 A2.t34 x36.Y GND.t369 GND.t368 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X289 a_5475_n6649# x5.x19.C VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X290 GND.t167 x22.Y A0.t37 GND.t166 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X291 A0.t101 x22.Y VDD.t166 VDD.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X292 VDD.t409 x36.A x36.Y VDD.t408 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X293 a_5751_n6649# x5.x19.C a_5645_n6649# GND.t85 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X294 x3.x4.A x3.EI VDD.t583 VDD.t582 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X295 VDD.t63 I15.t2 a_5509_n4211# VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X296 VDD.t462 EI.t8 a_5475_n5415# VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X297 GND.t367 x36.Y A2.t33 GND.t366 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X298 GND.t365 x36.Y A2.t26 GND.t364 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X299 x5.x19.X a_5475_n6649# VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X300 a_5629_n7635# x5.x19.D a_5557_n7635# GND.t773 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X301 a_5557_n14437# x3.x19.C a_5475_n14437# GND.t78 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X302 VDD.t164 x22.Y A0.t100 VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X303 GND.t888 x29.Y A1.t54 GND.t887 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X304 VDD.t711 x43.Y A3.t108 VDD.t710 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X305 A1.t53 x29.Y GND.t890 GND.t889 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X306 A2.t106 x36.Y VDD.t359 VDD.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X307 GND.t165 x22.Y A0.t36 GND.t164 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X308 VDD.t162 x22.Y A0.t99 VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X309 A3.t107 x43.Y VDD.t709 VDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X310 A0.t35 x22.Y GND.t163 GND.t162 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X311 A1.t108 x29.Y VDD.t891 VDD.t890 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X312 x5.x11.X a_5507_n2957# GND.t780 GND.t594 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X313 GND.t587 I8.t0 a_5475_n1175# GND.t64 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X314 VDD.t357 x36.Y A2.t105 VDD.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X315 VDD.t355 x36.Y A2.t104 VDD.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X316 A1.t52 x29.Y GND.t886 GND.t885 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X317 GND.t363 x36.Y A2.t25 GND.t362 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X318 x22.Y x22.A GND.t243 GND.t242 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X319 VDD.t160 x22.Y A0.t98 VDD.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X320 VDD.t889 x29.Y A1.t107 VDD.t888 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X321 A0.t34 x22.Y GND.t161 GND.t160 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X322 GND.t79 x3.x19.D a_5751_n14437# GND.t78 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X323 A0.t97 x22.Y VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X324 GND.t775 I6.t0 a_5475_n9979# GND.t257 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X325 x29.Y x29.A VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X326 A1.t106 x29.Y VDD.t885 VDD.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X327 A1.t105 x29.Y VDD.t887 VDD.t886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X328 A1.t51 x29.Y GND.t884 GND.t883 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X329 A3.t42 x43.Y GND.t688 GND.t687 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X330 VDD.t31 x29.A x29.Y VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X331 VDD.t883 x29.Y A1.t104 VDD.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X332 A0.t33 x22.Y GND.t159 GND.t158 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X333 GND.t882 x29.Y A1.t50 GND.t881 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X334 a_5475_n5415# I11.t0 VDD.t487 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X335 VDD.t353 x36.Y A2.t103 VDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X336 x22.Y x22.A VDD.t240 VDD.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X337 GND.t686 x43.Y A3.t41 GND.t685 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X338 GND.t241 x22.A x22.Y GND.t240 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X339 A0.t96 x22.Y VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X340 GND.t361 x36.Y A2.t24 GND.t360 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X341 VDD.t464 EI.t9 a_6519_n1397# VDD.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X342 x5.x19.C I12.t3 VDD.t254 VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X343 GND.t496 I13.t1 a_5593_n2957# GND.t82 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X344 x36.Y x36.A GND.t417 GND.t416 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X345 A2.t53 x36.Y GND.t359 GND.t358 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X346 A2.t52 x36.Y GND.t357 GND.t356 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X347 A3.t106 x43.Y VDD.t707 VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X348 a_5507_n10687# x3.EI VDD.t581 VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X349 GND.t880 x29.Y A1.t49 GND.t879 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X350 a_5653_n9215# I2.t2 a_5557_n9215# VDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X351 A0.t95 x22.Y VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X352 VDD.t705 x43.Y A3.t105 VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X353 VDD.t351 x36.Y A2.t102 VDD.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X354 VDD.t238 x22.A x22.Y VDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X355 GND.t878 x29.Y A1.t48 GND.t877 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X356 A2.t101 x36.Y VDD.t349 VDD.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X357 x36.Y x36.A VDD.t407 VDD.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X358 A2.t100 x36.Y VDD.t347 VDD.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X359 A2.t29 x36.Y GND.t355 GND.t354 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X360 x43.Y x43.A GND.t528 GND.t527 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X361 a_5935_n11219# x3.x22.A GND.t752 GND.t751 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X362 a_5475_n6397# x5.x18.C VDD.t610 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X363 GND.t239 x22.A x22.Y GND.t238 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X364 a_10858_n9865# x3.A1 a_10776_n9865# VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X365 VDD.t881 x29.Y A1.t103 VDD.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X366 A2.t99 x36.Y VDD.t345 VDD.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X367 a_6029_n1419# x5.x1.X GND.t746 GND.t745 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X368 GND.t772 x5.x19.D a_5751_n6397# GND.t84 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X369 A0.t32 x22.Y GND.t157 GND.t156 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X370 x43.Y x43.A VDD.t540 VDD.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X371 x5.x17.A a_5507_n3887# VDD.t599 VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X372 x5.x20.X a_5475_n7635# VDD.t476 VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X373 GND.t155 x22.Y A0.t31 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X374 x36.Y x36.A GND.t415 GND.t414 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X375 A2.t28 x36.Y GND.t353 GND.t352 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X376 VDD.t236 x22.A x22.Y VDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X377 a_6219_n12955# x3.x16.X GND.t749 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X378 a_5593_n2647# EI.t10 a_5507_n2647# GND.t57 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X379 A1.t102 x29.Y VDD.t879 VDD.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X380 GND.t413 x36.A x36.Y GND.t412 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X381 VDD.t29 x29.A x29.Y VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X382 A0.t94 x22.Y VDD.t152 VDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X383 GND.t574 x3.EI a_6605_n9437# GND.t573 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X384 a_5645_n14689# I3.t4 a_5557_n14689# GND.t75 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X385 x5.x16.X a_5475_n5415# GND.t591 GND.t590 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X386 x36.Y x36.A VDD.t405 VDD.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X387 A2.t98 x36.Y VDD.t343 VDD.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X388 VDD.t150 x22.Y A0.t93 VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X389 a_5475_n14689# x3.x19.C VDD.t603 VDD.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X390 a_10858_n13515# x3.A0 a_10776_n13515# VDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X391 VDD.t403 x36.A x36.Y VDD.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X392 x5.x19.D I14.t3 GND.t87 GND.t86 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X393 a_5557_n6397# x5.x19.C a_5475_n6397# GND.t84 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X394 GND.t446 x3.x19.X a_6395_n15425# GND.t445 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X395 a_5725_n9979# I5.t1 a_5653_n9979# VDD.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X396 a_5475_n1175# I11.t1 GND.t580 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X397 GND.t684 x43.Y A3.t40 GND.t683 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X398 GND.t682 x43.Y A3.t39 GND.t681 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X399 VDD.t557 x3.x4.A a_6183_n9215# VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X400 x3.x19.X a_5475_n14689# VDD.t591 VDD.t590 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X401 x43.Y x43.A GND.t526 GND.t525 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X402 A0.t30 x22.Y GND.t153 GND.t152 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X403 x22.Y x22.A GND.t237 GND.t236 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X404 x5.x1.X a_5475_n1175# GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X405 A3.t38 x43.Y GND.t680 GND.t679 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X406 A3.t37 x43.Y GND.t678 GND.t677 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X407 x5.EO a_6029_n1419# GND.t748 GND.t747 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X408 GND.t524 x43.A x43.Y GND.t523 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X409 VDD.t460 I6.t1 a_5507_n11927# VDD.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X410 GND.t151 x22.Y A0.t29 GND.t150 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X411 VDD.t703 x43.Y A3.t104 VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X412 VDD.t701 x43.Y A3.t103 VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X413 x43.Y x43.A VDD.t538 VDD.t537 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X414 A0.t92 x22.Y VDD.t148 VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X415 x3.x19.C I4.t3 VDD.t569 VDD.t568 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X416 x22.Y x22.A VDD.t234 VDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X417 A3.t102 x43.Y VDD.t699 VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X418 A3.t101 x43.Y VDD.t697 VDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X419 A1.t47 x29.Y GND.t876 GND.t875 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X420 VDD.t536 x43.A x43.Y VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X421 A0.t28 x22.Y GND.t149 GND.t148 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X422 VDD.t146 x22.Y A0.t91 VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X423 x28.A x1.X VDD.t566 VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X424 x3.x22.A a_5509_n12251# GND.t452 GND.t451 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X425 a_6477_n7385# x5.x20.X a_6395_n7385# VDD.t461 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X426 a_5645_n6649# I11.t2 a_5557_n6649# GND.t85 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X427 A1.t101 x29.Y VDD.t877 VDD.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X428 A0.t27 x22.Y GND.t147 GND.t146 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X429 A0.t90 x22.Y VDD.t144 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X430 A3.t36 x43.Y GND.t676 GND.t675 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X431 A3.t35 x43.Y GND.t674 GND.t673 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X432 GND.t145 x22.Y A0.t26 GND.t144 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X433 A3.t34 x43.Y GND.t672 GND.t671 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X434 a_6397_n4915# x5.x15.X a_6301_n4915# VDD.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X435 x5.x18.C I10.t3 VDD.t486 VDD.t485 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X436 GND.t522 x43.A x43.Y GND.t521 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X437 x2.A a_6395_n7385# VDD.t455 VDD.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X438 GND.t874 x29.Y A1.t46 GND.t873 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X439 a_10776_n9865# x3.A1 GND.t52 GND.t51 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X440 a_6113_n3179# x5.x17.A a_6017_n3179# VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X441 GND.t351 x36.Y A2.t27 GND.t350 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X442 GND.t349 x36.Y A2.t42 GND.t348 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X443 a_6395_n15425# x3.x20.X GND.t493 GND.t492 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X444 GND.t235 x22.A x22.Y GND.t234 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X445 GND.t555 x3.x14.A a_5935_n11219# GND.t554 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 A2.t41 x36.Y GND.t347 GND.t346 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X447 A0.t89 x22.Y VDD.t142 VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X448 GND.t758 x28.A x29.A GND.t757 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X449 A3.t100 x43.Y VDD.t695 VDD.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X450 GND.t670 x43.Y A3.t33 GND.t669 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X451 a_5475_n14437# x3.x18.C VDD.t458 VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X452 VDD.t140 x22.Y A0.t88 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 x1.X a_10776_n9865# GND.t491 GND.t490 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X454 A3.t99 x43.Y VDD.t693 VDD.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X455 A3.t98 x43.Y VDD.t691 VDD.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 a_6017_n3179# x5.x22.A a_5935_n3179# VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X457 A3.t32 x43.Y GND.t668 GND.t667 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X458 a_5751_n13455# x3.x16.C a_5645_n13455# GND.t576 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X459 GND.t872 x29.Y A1.t45 GND.t871 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X460 VDD.t534 x43.A x43.Y VDD.t533 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X461 VDD.t341 x36.Y A2.t97 VDD.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X462 VDD.t339 x36.Y A2.t96 VDD.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X463 x3.A1 a_6219_n12955# VDD.t766 VDD.t765 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X464 a_5595_n12251# x3.EI a_5509_n12251# GND.t572 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X465 A1.t44 x29.Y GND.t870 GND.t869 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X466 A1.t43 x29.Y GND.t868 GND.t867 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X467 GND.t143 x22.Y A0.t25 GND.t142 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X468 VDD.t772 x3.x22.A a_6645_n15425# VDD.t771 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X469 VDD.t232 x22.A x22.Y VDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X470 VDD.t689 x43.Y A3.t97 VDD.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X471 A2.t95 x36.Y VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X472 x22.Y x22.A GND.t233 GND.t232 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X473 A3.t96 x43.Y VDD.t687 VDD.t686 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X474 VDD.t783 x5.x21.B a_5967_n7607# VDD.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 x29.Y x29.A GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X476 x29.Y x29.A VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X477 A1.t100 x29.Y VDD.t875 VDD.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X478 VDD.t138 x22.Y A0.t87 VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X479 A1.t99 x29.Y VDD.t873 VDD.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X480 VDD.t25 x29.A x29.Y VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X481 VDD.t871 x29.Y A1.t98 VDD.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X482 x22.Y x22.A VDD.t230 VDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X483 VDD.t869 x29.Y A1.t97 VDD.t868 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X484 x3.A2 a_5935_n11219# VDD.t472 VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X485 GND.t345 x36.Y A2.t51 GND.t344 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X486 GND.t464 x2.A a_10776_n13515# GND.t463 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X487 A1.t42 x29.Y GND.t866 GND.t865 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 a_6469_n4915# x5.x22.A a_6397_n4915# VDD.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X489 VDD.t256 I5.t2 a_5507_n10997# VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X490 GND.t26 x29.A x29.Y GND.t25 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X491 A2.t50 x36.Y GND.t343 GND.t342 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X492 A2.t49 x36.Y GND.t341 GND.t340 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X493 A0.t24 x22.Y GND.t141 GND.t140 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X494 x22.A x21.A GND.t740 GND.t739 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X495 a_6185_n3179# x5.x11.X a_6113_n3179# VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X496 GND.t339 x36.Y A2.t55 GND.t338 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X497 VDD.t867 x29.Y A1.t96 VDD.t866 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X498 A1.t41 x29.Y GND.t864 GND.t863 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X499 VDD.t335 x36.Y A2.t94 VDD.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X500 VDD.t466 x2.A a_10858_n13515# VDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X501 a_5593_n3887# EI.t11 a_5507_n3887# GND.t58 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X502 GND.t862 x29.Y A1.t40 GND.t861 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X503 A2.t93 x36.Y VDD.t321 VDD.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X504 A2.t92 x36.Y VDD.t333 VDD.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X505 A0.t86 x22.Y VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X506 x22.A x21.A VDD.t761 VDD.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X507 A2.t54 x36.Y GND.t337 GND.t336 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X508 A2.t37 x36.Y GND.t335 GND.t334 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X509 x5.x16.C I13.t2 GND.t560 GND.t559 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X510 VDD.t331 x36.Y A2.t91 VDD.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X511 GND.t333 x36.Y A2.t36 GND.t332 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X512 GND.t860 x29.Y A1.t39 GND.t859 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X513 GND.t65 I10.t4 a_5475_n1175# GND.t64 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X514 VDD.t468 I4.t4 a_5725_n9979# VDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X515 VDD.t865 x29.Y A1.t95 VDD.t864 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 a_6219_n12955# x3.x22.A GND.t750 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X517 VDD.t863 x29.Y A1.t94 VDD.t862 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X518 A2.t90 x36.Y VDD.t329 VDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X519 A2.t89 x36.Y VDD.t327 VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X520 a_6645_n15425# x3.x21.X a_6573_n15425# VDD.t489 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X521 x3.EI x5.EO GND.t770 GND.t769 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X522 x29.Y x29.A VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X523 GND.t858 x29.Y A1.t38 GND.t857 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X524 a_5751_n5415# x5.x16.C a_5645_n5415# GND.t3 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X525 VDD.t323 x36.Y A2.t88 VDD.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X526 A1.t37 x29.Y GND.t856 GND.t855 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X527 a_5475_n9979# I5.t3 GND.t258 GND.t257 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X528 VDD.t21 x29.A x29.Y VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X529 VDD.t861 x29.Y A1.t93 VDD.t860 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 x29.Y x29.A VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X531 VDD.t470 I4.t5 a_5507_n10687# VDD.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X532 x3.x15.X a_5475_n13205# GND.t74 GND.t73 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X533 x36.A x35.A GND.t443 GND.t442 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X534 GND.t139 x22.Y A0.t23 GND.t138 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X535 x34.A a_10776_n5725# GND.t495 GND.t494 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X536 GND.t441 x35.A x36.A GND.t440 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X537 GND.t331 x36.Y A2.t35 GND.t330 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X538 GND.t329 x36.Y A2.t122 GND.t328 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X539 a_6573_n7385# x5.x19.X a_6477_n7385# VDD.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X540 a_6017_n11219# x3.x22.A a_5935_n11219# VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X541 x36.A x35.A VDD.t438 VDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X542 GND.t129 x22.Y A0.t22 GND.t128 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X543 x5.x2.X a_5475_n1939# VDD.t389 VDD.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X544 GND.t666 x43.Y A3.t31 GND.t665 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X545 GND.t664 x43.Y A3.t30 GND.t663 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X546 x34.A a_10776_n5725# VDD.t501 VDD.t500 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X547 VDD.t325 x36.Y A2.t87 VDD.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X548 x22.Y x22.A GND.t231 GND.t230 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X549 VDD.t134 x22.Y A0.t85 VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 VDD.t436 x35.A x36.A VDD.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X551 VDD.t319 x36.Y A2.t86 VDD.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X552 a_5475_n13455# x3.x16.C VDD.t935 VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X553 A1.t36 x29.Y GND.t854 GND.t853 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X554 GND.t137 x22.Y A0.t21 GND.t136 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X555 A0.t20 x22.Y GND.t135 GND.t134 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X556 VDD.t132 x22.Y A0.t84 VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X557 x5.GS a_6519_n1397# GND.t263 GND.t262 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X558 x22.Y x22.A VDD.t228 VDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X559 VDD.t685 x43.Y A3.t95 VDD.t684 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X560 VDD.t683 x43.Y A3.t94 VDD.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X561 x3.x16.C I5.t4 VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X562 VDD.t17 x29.A x29.Y VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X563 GND.t478 x5.x4.A a_6029_n1419# GND.t477 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X564 x3.x16.X a_5475_n13455# VDD.t940 VDD.t939 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X565 VDD.t130 x22.Y A0.t83 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X566 A0.t19 x22.Y GND.t133 GND.t132 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X567 GND.t83 I12.t4 a_5593_n2647# GND.t82 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X568 x3.A0 a_6395_n15425# GND.t742 GND.t741 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X569 A0.t82 x22.Y VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X570 x3.x20.X a_5475_n15675# GND.t539 GND.t538 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X571 A1.t35 x29.Y GND.t852 GND.t851 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X572 GND.t850 x29.Y A1.t34 GND.t849 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X573 a_6645_n7385# x5.x21.X a_6573_n7385# VDD.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X574 GND.t131 x22.Y A0.t18 GND.t130 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X575 A0.t81 x22.Y VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X576 A3.t29 x43.Y GND.t662 GND.t661 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X577 x3.x20.X a_5475_n15675# VDD.t551 VDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X578 x3.A0 a_6395_n15425# VDD.t763 VDD.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X579 A3.t28 x43.Y GND.t660 GND.t659 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X580 VDD.t503 x5.x17.A a_6469_n4915# VDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X581 x3.x21.X a_5967_n15647# GND.t545 GND.t544 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X582 a_6395_n15425# x3.x21.X GND.t485 GND.t484 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X583 GND.t848 x29.Y A1.t33 GND.t847 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X584 GND.t520 x43.A x43.Y GND.t519 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X585 GND.t658 x43.Y A3.t27 GND.t657 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X586 GND.t656 x43.Y A3.t26 GND.t655 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X587 VDD.t932 x5.x14.A a_6185_n3179# VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X588 GND.t127 x22.Y A0.t17 GND.t126 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X589 VDD.t124 x22.Y A0.t80 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X590 a_5557_n9979# I7.t1 a_5475_n9979# VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X591 a_5645_n13455# x3.x19.C a_5557_n13455# GND.t576 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X592 GND.t846 x29.Y A1.t32 GND.t845 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X593 x5.x4.A EI.t12 VDD.t753 VDD.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X594 A3.t93 x43.Y VDD.t681 VDD.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X595 A3.t92 x43.Y VDD.t679 VDD.t678 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X596 a_5557_n7635# I13.t3 a_5475_n7635# GND.t4 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X597 A3.t25 x43.Y GND.t654 GND.t653 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X598 A3.t24 x43.Y GND.t652 GND.t651 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X599 VDD.t579 x3.EI a_5475_n15675# VDD.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X600 x3.x21.X a_5967_n15647# VDD.t559 VDD.t558 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X601 A1.t31 x29.Y GND.t844 GND.t843 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X602 VDD.t532 x43.A x43.Y VDD.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X603 VDD.t677 x43.Y A3.t91 VDD.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X604 VDD.t675 x43.Y A3.t90 VDD.t674 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X605 VDD.t122 x22.Y A0.t79 VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X606 GND.t650 x43.Y A3.t23 GND.t649 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X607 a_5751_n13205# x3.x16.C a_5645_n13205# GND.t564 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X608 A2.t121 x36.Y GND.t327 GND.t326 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X609 A1.t30 x29.Y GND.t842 GND.t841 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X610 A3.t89 x43.Y VDD.t673 VDD.t672 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X611 A3.t88 x43.Y VDD.t671 VDD.t670 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X612 GND.t840 x29.Y A1.t29 GND.t839 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X613 VDD.t669 x43.Y A3.t87 VDD.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X614 a_5629_n15675# x3.x19.D a_5557_n15675# GND.t77 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X615 x3.x14.A a_5507_n10687# GND.t774 GND.t482 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X616 VDD.t15 x29.A x29.Y VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X617 GND.t229 x22.A x22.Y GND.t228 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X618 A2.t85 x36.Y VDD.t317 VDD.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X619 A2.t13 x36.Y GND.t325 GND.t324 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X620 a_6519_n9437# x3.EO VDD.t479 VDD.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X621 a_6053_n15647# x3.EI a_5967_n15647# GND.t571 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X622 x5.x15.X a_5475_n5165# VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X623 A1.t92 x29.Y VDD.t859 VDD.t858 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X624 VDD.t226 x22.A x22.Y VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X625 A1.t28 x29.Y GND.t838 GND.t837 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X626 GND.t323 x36.Y A2.t12 GND.t322 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X627 GND.t321 x36.Y A2.t11 GND.t320 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X628 VDD.t857 x29.Y A1.t91 VDD.t856 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X629 VDD.t567 x3.x14.A a_6185_n11219# VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X630 VDD.t855 x29.Y A1.t90 VDD.t854 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X631 x3.x21.B a_5475_n14437# GND.t91 GND.t90 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X632 GND.t836 x29.Y A1.t27 GND.t835 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X633 GND.t518 x43.A x43.Y GND.t517 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X634 GND.t648 x43.Y A3.t22 GND.t647 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X635 x29.Y x29.A GND.t24 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X636 GND.t646 x43.Y A3.t21 GND.t645 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X637 A2.t84 x36.Y VDD.t315 VDD.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X638 x43.Y x43.A GND.t516 GND.t515 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X639 A3.t20 x43.Y GND.t644 GND.t643 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X640 A2.t7 x36.Y GND.t319 GND.t318 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X641 A2.t6 x36.Y GND.t317 GND.t316 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X642 A2.t18 x36.Y GND.t315 GND.t314 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X643 A1.t26 x29.Y GND.t834 GND.t833 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X644 VDD.t313 x36.Y A2.t83 VDD.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X645 VDD.t311 x36.Y A2.t82 VDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X646 GND.t46 I7.t2 a_5595_n12251# GND.t45 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X647 GND.t832 x29.Y A1.t25 GND.t831 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X648 GND.t411 x36.A x36.Y GND.t410 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X649 GND.t313 x36.Y A2.t17 GND.t312 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X650 VDD.t530 x43.A x43.Y VDD.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X651 VDD.t667 x43.Y A3.t86 VDD.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X652 VDD.t665 x43.Y A3.t85 VDD.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X653 a_5645_n5415# x5.x19.C a_5557_n5415# GND.t3 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X654 x42.A x5.GS GND.t450 GND.t449 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X655 x3.x19.D I6.t2 GND.t44 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X656 VDD.t853 x29.Y A1.t89 VDD.t852 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X657 VDD.t601 x3.x19.C a_5475_n13205# VDD.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X658 x43.Y x43.A VDD.t528 VDD.t527 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X659 A3.t84 x43.Y VDD.t663 VDD.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X660 A2.t81 x36.Y VDD.t309 VDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X661 GND.t771 x5.x19.D a_5751_n6649# GND.t85 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X662 A2.t80 x36.Y VDD.t307 VDD.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X663 A2.t79 x36.Y VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X664 x5.x1.X a_5475_n1175# VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X665 VDD.t401 x36.A x36.Y VDD.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X666 VDD.t303 x36.Y A2.t78 VDD.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X667 GND.t475 x3.x2.X a_6029_n9459# GND.t474 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X668 x28.A x1.X GND.t553 GND.t552 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X669 x5.EO a_6029_n1419# VDD.t769 VDD.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X670 x3.x2.X a_5475_n9979# GND.t583 GND.t582 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X671 a_5593_n10997# x3.EI a_5507_n10997# GND.t567 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X672 x42.A x5.GS VDD.t447 VDD.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X673 x5.x15.X a_5475_n5165# GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X674 x29.Y x29.A GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X675 VDD.t851 x29.Y A1.t88 VDD.t850 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X676 a_6301_n12955# x3.x16.X a_6219_n12955# VDD.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X677 x29.Y x29.A VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X678 A1.t87 x29.Y VDD.t849 VDD.t848 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X679 A1.t86 x29.Y VDD.t847 VDD.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X680 x36.A x35.A GND.t439 GND.t438 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X681 a_5475_n13205# I2.t3 VDD.t443 VDD.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X682 GND.t830 x29.Y A1.t24 GND.t829 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X683 GND.t311 x36.Y A2.t16 GND.t310 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X684 GND.t309 x36.Y A2.t124 GND.t308 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X685 A1.t23 x29.Y GND.t828 GND.t827 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X686 x5.x11.X a_5507_n2957# VDD.t801 VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X687 a_6185_n11219# x3.x11.X a_6113_n11219# VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X688 VDD.t79 x5.x19.C a_5475_n5165# VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X689 a_5557_n6649# EI.t13 a_5475_n6649# GND.t85 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X690 VDD.t393 x5.x22.A a_6645_n7385# VDD.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X691 A2.t123 x36.Y GND.t307 GND.t306 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X692 A2.t40 x36.Y GND.t305 GND.t304 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X693 x3.x18.C I2.t4 GND.t563 GND.t562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X694 A1.t85 x29.Y VDD.t845 VDD.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X695 x36.A x35.A VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X696 x5.x21.X a_5967_n7607# GND.t589 GND.t588 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X697 GND.t503 I14.t4 a_5593_n3887# GND.t502 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X698 x5.x22.A a_5509_n4211# GND.t541 GND.t540 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X699 VDD.t301 x36.Y A2.t77 VDD.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X700 VDD.t299 x36.Y A2.t76 VDD.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X701 GND.t481 x3.x17.A a_6219_n12955# GND.t88 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X702 x5.A2 a_5935_n3179# GND.t63 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X703 A2.t75 x36.Y VDD.t297 VDD.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X704 A2.t74 x36.Y VDD.t295 VDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X705 a_5475_n5415# x5.x16.C VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X706 VDD.t577 x3.EI a_5475_n13205# VDD.t576 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X707 a_5653_n9979# I6.t3 a_5557_n9979# VDD.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X708 a_5475_n1175# I9.t1 GND.t546 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X709 GND.t227 x22.A x22.Y GND.t226 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X710 GND.t826 x29.Y A1.t22 GND.t825 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X711 x5.x16.X a_5475_n5415# VDD.t609 VDD.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X712 x29.Y x29.A VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X713 A1.t84 x29.Y VDD.t843 VDD.t842 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X714 VDD.t9 x29.A x29.Y VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X715 A3.t19 x43.Y GND.t642 GND.t641 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X716 a_5751_n14437# x3.x18.C a_5645_n14437# GND.t78 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X717 A0.t16 x22.Y GND.t125 GND.t124 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X718 x5.x19.D I14.t5 VDD.t507 VDD.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X719 GND.t640 x43.Y A3.t18 GND.t639 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X720 VDD.t224 x22.A x22.Y VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X721 A1.t21 x29.Y GND.t824 GND.t823 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X722 GND.t570 x3.EI a_5629_n15675# GND.t569 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X723 A0.t78 x22.Y VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X724 A3.t83 x43.Y VDD.t661 VDD.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X725 A1.t20 x29.Y GND.t822 GND.t821 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X726 VDD.t659 x43.Y A3.t82 VDD.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X727 GND.t437 x35.A x36.A GND.t436 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X728 GND.t820 x29.Y A1.t19 GND.t819 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X729 A3.t17 x43.Y GND.t638 GND.t637 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X730 A0.t15 x22.Y GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X731 VDD.t67 I5.t5 a_5475_n15675# VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X732 x3.x15.X a_5475_n13205# VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X733 GND.t480 x3.x17.A a_5935_n11219# GND.t479 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X734 GND.t636 x43.Y A3.t16 GND.t635 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X735 GND.t225 x22.A x22.Y GND.t224 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X736 a_5557_n15675# I5.t6 a_5475_n15675# GND.t254 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X737 a_5509_n12251# x3.EI VDD.t575 VDD.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X738 x3.x17.A a_5507_n11927# GND.t489 GND.t488 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X739 GND.t818 x29.Y A1.t18 GND.t817 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X740 A3.t81 x43.Y VDD.t657 VDD.t656 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X741 VDD.t432 x35.A x36.A VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X742 x3.x11.X a_5507_n10997# GND.t483 GND.t482 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X743 A3.t15 x43.Y GND.t634 GND.t633 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X744 VDD.t937 EI.t14 a_5475_n5165# VDD.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X745 A0.t77 x22.Y VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X746 a_6573_n15425# x3.x19.X a_6477_n15425# VDD.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X747 VDD.t222 x22.A x22.Y VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X748 a_5645_n13205# x3.x19.C a_5557_n13205# GND.t564 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X749 VDD.t655 x43.Y A3.t80 VDD.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X750 GND.t632 x43.Y A3.t14 GND.t631 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X751 GND.t630 x43.Y A3.t13 GND.t629 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X752 x3.x22.A a_5509_n12251# VDD.t449 VDD.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X753 x3.x17.A a_5507_n11927# VDD.t493 VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X754 x43.A x42.A GND.t602 GND.t449 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X755 x29.Y x29.A GND.t20 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X756 A2.t39 x36.Y GND.t303 GND.t302 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X757 A3.t79 x43.Y VDD.t653 VDD.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X758 a_6111_n1175# x5.x2.X a_6029_n1419# VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X759 GND.t816 x29.Y A1.t17 GND.t815 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X760 VDD.t651 x43.Y A3.t78 VDD.t650 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X761 VDD.t649 x43.Y A3.t77 VDD.t648 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X762 x43.A x42.A VDD.t621 VDD.t620 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X763 A1.t16 x29.Y GND.t814 GND.t813 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X764 a_5507_n2957# EI.t15 VDD.t938 VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X765 A2.t73 x36.Y VDD.t293 VDD.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X766 GND.t18 x29.A x29.Y GND.t17 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X767 x22.A x21.A GND.t738 GND.t737 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X768 x5.x21.B a_5475_n6397# GND.t50 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X769 a_5475_n5165# I10.t5 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X770 A1.t15 x29.Y GND.t812 GND.t811 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X771 a_5593_n11927# x3.EI a_5507_n11927# GND.t568 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X772 GND.t810 x29.Y A1.t14 GND.t809 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X773 a_5475_n7635# x5.x19.D VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X774 VDD.t841 x29.Y A1.t83 VDD.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X775 VDD.t839 x29.Y A1.t82 VDD.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X776 x22.A x21.A VDD.t759 VDD.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X777 GND.t628 x43.Y A3.t12 GND.t627 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X778 GND.t626 x43.Y A3.t11 GND.t625 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X779 A1.t81 x29.Y VDD.t837 VDD.t836 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X780 GND.t736 x21.A x22.A GND.t735 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X781 x43.A x42.A GND.t601 GND.t600 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X782 x5.x21.B a_5475_n6397# VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X783 x43.Y x43.A GND.t514 GND.t513 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X784 A3.t10 x43.Y GND.t624 GND.t623 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X785 a_6219_n4915# x5.x16.X GND.t551 GND.t398 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X786 A2.t38 x36.Y GND.t301 GND.t300 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X787 GND.t808 x29.Y A1.t13 GND.t807 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X788 GND.t512 x43.A x43.Y GND.t511 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X789 GND.t299 x36.Y A2.t48 GND.t298 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X790 GND.t297 x36.Y A2.t47 GND.t296 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X791 a_5725_n1175# I9.t2 a_5653_n1175# VDD.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X792 VDD.t641 x43.Y A3.t76 VDD.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X793 a_6477_n15425# x3.x20.X a_6395_n15425# VDD.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X794 a_6183_n1175# x5.x1.X a_6111_n1175# VDD.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X795 x43.A x42.A VDD.t619 VDD.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X796 VDD.t647 x43.Y A3.t75 VDD.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X797 VDD.t757 x21.A x22.A VDD.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X798 GND.t806 x29.Y A1.t12 GND.t805 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X799 x43.Y x43.A VDD.t526 VDD.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X800 A3.t74 x43.Y VDD.t645 VDD.t644 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X801 A3.t9 x43.Y GND.t622 GND.t621 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X802 A3.t8 x43.Y GND.t620 GND.t619 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X803 A2.t72 x36.Y VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X804 GND.t72 I0.t1 a_5475_n9215# GND.t71 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X805 A1.t11 x29.Y GND.t804 GND.t803 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X806 VDD.t524 x43.A x43.Y VDD.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X807 VDD.t289 x36.Y A2.t71 VDD.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X808 VDD.t287 x36.Y A2.t70 VDD.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X809 GND.t295 x36.Y A2.t23 GND.t294 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X810 GND.t121 x22.Y A0.t14 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X811 x36.Y x36.A GND.t409 GND.t408 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X812 x29.Y x29.A GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X813 x5.GS a_6519_n1397# VDD.t258 VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X814 VDD.t835 x29.Y A1.t80 VDD.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X815 A0.t13 x22.Y GND.t119 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X816 A1.t10 x29.Y GND.t802 GND.t801 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X817 A3.t73 x43.Y VDD.t643 VDD.t642 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X818 A3.t72 x43.Y VDD.t639 VDD.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 GND.t1 x3.x21.B a_6053_n15647# GND.t0 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X820 a_5507_n2647# EI.t16 VDD.t512 VDD.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X821 GND.t454 x5.A2 a_10776_n5725# GND.t453 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X822 A1.t79 x29.Y VDD.t833 VDD.t832 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X823 A1.t78 x29.Y VDD.t831 VDD.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X824 x5.x16.C I13.t4 VDD.t593 VDD.t592 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X825 a_5595_n4211# EI.t17 a_5509_n4211# GND.t504 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X826 VDD.t285 x36.Y A2.t69 VDD.t284 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X827 VDD.t829 x29.Y A1.t77 VDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X828 VDD.t116 x22.Y A0.t76 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X829 A1.t9 x29.Y GND.t800 GND.t799 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X830 x36.Y x36.A VDD.t399 VDD.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X831 VDD.t573 x3.EI a_6519_n9437# VDD.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X832 A0.t12 x22.Y GND.t117 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X833 A0.t75 x22.Y VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X834 GND.t14 x29.A x29.Y GND.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X835 GND.t293 x36.Y A2.t22 GND.t292 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X836 a_6053_n7607# EI.t18 a_5967_n7607# GND.t80 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X837 a_5557_n14689# x3.EI a_5475_n14689# GND.t75 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X838 VDD.t451 x5.A2 a_10858_n5725# VDD.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X839 A2.t21 x36.Y GND.t291 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X840 VDD.t931 I11.t3 a_5475_n6649# VDD.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X841 VDD.t495 I13.t5 a_5475_n7635# VDD.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X842 A1.t76 x29.Y VDD.t827 VDD.t826 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 A1.t75 x29.Y VDD.t825 VDD.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X844 A0.t11 x22.Y GND.t115 GND.t114 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X845 x43.Y x43.A GND.t510 GND.t509 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X846 VDD.t823 x29.Y A1.t74 VDD.t822 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X847 GND.t113 x22.Y A0.t10 GND.t112 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X848 A0.t74 x22.Y VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X849 GND.t599 x42.A x43.A GND.t598 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X850 VDD.t283 x36.Y A2.t68 VDD.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X851 GND.t289 x36.Y A2.t44 GND.t288 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X852 GND.t287 x36.Y A2.t43 GND.t286 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X853 A2.t67 x36.Y VDD.t281 VDD.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X854 x36.Y x36.A GND.t407 GND.t406 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X855 A2.t127 x36.Y GND.t285 GND.t284 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X856 A2.t126 x36.Y GND.t283 GND.t282 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X857 a_6395_n7385# x5.x20.X GND.t462 GND.t461 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X858 GND.t111 x22.Y A0.t9 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X859 A0.t73 x22.Y VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X860 x43.Y x43.A VDD.t522 VDD.t521 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 VDD.t108 x22.Y A0.t72 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X862 VDD.t617 x42.A x43.A VDD.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X863 GND.t76 x3.x19.D a_5751_n14689# GND.t75 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X864 VDD.t279 x36.Y A2.t66 VDD.t278 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X865 GND.t256 I5.t7 a_5593_n10997# GND.t255 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X866 GND.t12 x29.A x29.Y GND.t11 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X867 VDD.t277 x36.Y A2.t65 VDD.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X868 a_5645_n14437# I1.t3 a_5557_n14437# GND.t78 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X869 a_6029_n9459# x3.x1.X GND.t593 GND.t592 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X870 GND.t109 x22.Y A0.t8 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X871 x36.Y x36.A VDD.t397 VDD.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X872 A2.t64 x36.Y VDD.t275 VDD.t274 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X873 A2.t63 x36.Y VDD.t273 VDD.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X874 VDD.t106 x22.Y A0.t71 VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X875 A1.t8 x29.Y GND.t798 GND.t797 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X876 GND.t796 x29.Y A1.t7 GND.t795 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X877 x29.A x28.A VDD.t777 VDD.t776 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X878 GND.t81 EI.t19 a_5751_n5415# GND.t3 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X879 a_10776_n5725# x3.A2 GND.t67 GND.t66 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X880 x1.X a_10776_n9865# VDD.t497 VDD.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X881 VDD.t775 x28.A x29.A VDD.t774 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X882 VDD.t821 x29.Y A1.t73 VDD.t820 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X883 VDD.t819 x29.Y A1.t72 VDD.t818 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X884 VDD.t104 x22.Y A0.t70 VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X885 x3.x14.A a_5507_n10687# VDD.t794 VDD.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X886 A2.t125 x36.Y GND.t281 GND.t280 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X887 GND.t69 I12.t5 a_5475_n1939# GND.t68 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X888 x3.EI x5.EO VDD.t785 VDD.t784 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X889 x3.x21.B a_5475_n14437# VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X890 a_5475_n9215# I3.t5 GND.t767 GND.t71 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X891 A2.t62 x36.Y VDD.t271 VDD.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X892 GND.t618 x43.Y A3.t7 GND.t617 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X893 VDD.t790 x5.x19.D a_5475_n6649# VDD.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X894 x3.x1.X a_5475_n9215# GND.t777 GND.t776 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X895 VDD.t800 I9.t3 a_5475_n6397# VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X896 x3.EO a_6029_n9459# GND.t253 GND.t252 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X897 a_5593_n10687# x3.EI a_5507_n10687# GND.t567 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X898 A1.t6 x29.Y GND.t794 GND.t793 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X899 x29.Y x29.A GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X900 A3.t6 x43.Y GND.t616 GND.t615 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X901 A3.t5 x43.Y GND.t614 GND.t613 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X902 VDD.t84 I8.t1 a_5725_n1175# VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X903 a_5557_n5415# I11.t4 a_5475_n5415# GND.t3 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X904 a_5751_n5165# x5.x16.C a_5645_n5165# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X905 GND.t792 x29.Y A1.t5 GND.t791 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X906 VDD.t637 x43.Y A3.t71 VDD.t636 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X907 x3.x1.X a_5475_n9215# VDD.t798 VDD.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X908 x3.EO a_6029_n9459# VDD.t252 VDD.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X909 GND.t612 x43.Y A3.t4 GND.t611 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X910 A3.t70 x43.Y VDD.t631 VDD.t630 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X911 A3.t69 x43.Y VDD.t635 VDD.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X912 a_5725_n1939# I13.t6 a_5653_n1939# VDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X913 A1.t4 x29.Y GND.t790 GND.t789 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X914 a_6113_n11219# x3.x17.A a_6017_n11219# VDD.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X915 x3.x2.X a_5475_n9979# VDD.t595 VDD.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X916 a_5935_n11219# x3.x11.X GND.t764 GND.t763 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X917 VDD.t633 x43.Y A3.t68 VDD.t632 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X918 a_5475_n6649# EI.t20 VDD.t515 VDD.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X919 VDD.t514 I7.t3 a_5509_n12251# VDD.t513 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X920 A0.t7 x22.Y GND.t107 GND.t106 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X921 A1.t3 x29.Y GND.t788 GND.t787 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X922 GND.t786 x29.Y A1.t2 GND.t785 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X923 x43.Y x43.A GND.t508 GND.t507 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X924 a_6605_n1397# x5.EO a_6519_n1397# GND.t768 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X925 a_5507_n3887# EI.t21 VDD.t516 VDD.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X926 GND.t279 x36.Y A2.t46 GND.t278 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X927 GND.t8 x29.A x29.Y GND.t7 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X928 GND.t610 x43.Y A3.t3 GND.t609 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X929 A2.t45 x36.Y GND.t277 GND.t276 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X930 A2.t5 x36.Y GND.t275 GND.t274 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X931 x5.x21.X a_5967_n7607# VDD.t607 VDD.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X932 A0.t69 x22.Y VDD.t102 VDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X933 A1.t71 x29.Y VDD.t817 VDD.t816 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X934 x43.Y x43.A VDD.t520 VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X935 A3.t2 x43.Y GND.t608 GND.t607 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X936 A3.t1 x43.Y GND.t606 GND.t605 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X937 GND.t604 x43.Y A3.t0 GND.t603 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X938 VDD.t269 x36.Y A2.t61 VDD.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X939 GND.t448 x5.x19.X a_6395_n7385# GND.t447 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X940 GND.t105 x22.Y A0.t6 GND.t104 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X941 a_10776_n13515# x3.A0 GND.t550 GND.t549 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X942 GND.t784 x29.Y A1.t1 GND.t783 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X943 VDD.t629 x43.Y A3.t67 VDD.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 A2.t60 x36.Y VDD.t267 VDD.t266 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X945 A2.t59 x36.Y VDD.t265 VDD.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X946 x29.Y x29.A GND.t6 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X947 VDD.t788 x5.x19.D a_5475_n6397# VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X948 GND.t734 x21.A x22.A GND.t733 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X949 x2.X a_10776_n13515# GND.t732 GND.t731 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X950 A3.t66 x43.Y VDD.t627 VDD.t626 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X951 A3.t65 x43.Y VDD.t625 VDD.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X952 A1.t70 x29.Y VDD.t815 VDD.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X953 GND.t103 x22.Y A0.t5 GND.t102 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X954 VDD.t100 x22.Y A0.t68 VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X955 VDD.t623 x43.Y A3.t64 VDD.t622 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X956 VDD.t57 I13.t7 a_5507_n2957# VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X957 A0.t4 x22.Y GND.t101 GND.t100 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X958 A0.t3 x22.Y GND.t99 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X959 GND.t779 I6.t4 a_5593_n11927# GND.t778 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X960 VDD.t813 x29.Y A1.t69 VDD.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X961 VDD.t811 x29.Y A1.t68 VDD.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X962 VDD.t755 x21.A x22.A VDD.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X963 a_5475_n1939# I15.t3 GND.t70 GND.t68 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X964 x2.X a_10776_n13515# VDD.t751 VDD.t750 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X965 GND.t56 x1.A a_10776_n9865# GND.t55 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X966 A2.t4 x36.Y GND.t273 GND.t272 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X967 x3.x4.A x3.EI GND.t566 GND.t565 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X968 x3.x19.D I6.t5 VDD.t429 VDD.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X969 x22.Y x22.A GND.t223 GND.t222 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X970 VDD.t98 x22.Y A0.t67 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X971 A1.t0 x29.Y GND.t782 GND.t781 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X972 x29.A x28.A GND.t756 GND.t755 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X973 A1.t67 x29.Y VDD.t809 VDD.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X974 A1.t66 x29.Y VDD.t807 VDD.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X975 A1.t65 x29.Y VDD.t805 VDD.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X976 A0.t66 x22.Y VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X977 A0.t65 x22.Y VDD.t94 VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X978 VDD.t7 x29.A x29.Y VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X979 VDD.t803 x29.Y A1.t64 VDD.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X980 GND.t597 x42.A x43.A GND.t596 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X981 GND.t89 x3.x15.X a_6219_n12955# GND.t88 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X982 GND.t506 x43.A x43.Y GND.t505 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X983 GND.t271 x36.Y A2.t3 GND.t270 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X984 A0.t2 x22.Y GND.t97 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X985 x22.Y x22.A VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X986 a_5557_n1175# I11.t5 a_5475_n1175# VDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X987 A2.t58 x36.Y VDD.t263 VDD.t262 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X988 a_5475_n6397# x5.x19.C VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X989 GND.t221 x22.A x22.Y GND.t220 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X990 x36.Y x36.A GND.t405 GND.t404 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X991 A2.t20 x36.Y GND.t269 GND.t268 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X992 A2.t19 x36.Y GND.t267 GND.t266 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X993 VDD.t615 x42.A x43.A VDD.t614 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X994 GND.t403 x36.A x36.Y GND.t402 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X995 GND.t265 x36.Y A2.t56 GND.t264 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X996 GND.t561 I2.t5 a_5475_n9215# GND.t71 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X997 VDD.t483 x3.x17.A a_6469_n12955# VDD.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X998 A0.t1 x22.Y GND.t95 GND.t94 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X999 VDD.t518 x43.A x43.Y VDD.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1000 VDD.t261 x36.Y A2.t57 VDD.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1001 A0.t64 x22.Y VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1002 a_5475_n13205# x3.x16.C VDD.t934 VDD.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1003 GND.t93 x22.Y A0.t0 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R0 VDD.n831 VDD 1319.65
R1 VDD.n58 VDD 1319.65
R2 VDD.n672 VDD.t436 584.644
R3 VDD.n1114 VDD.t775 584.644
R4 VDD.n1452 VDD.t757 584.644
R5 VDD.n86 VDD.t615 584.644
R6 VDD.n831 VDD.t582 533.735
R7 VDD.n58 VDD.t752 533.735
R8 VDD.n1557 VDD.n1556 425.228
R9 VDD.n777 VDD.n776 425.228
R10 VDD VDD.t784 421.082
R11 VDD.n1166 VDD.t594 396.079
R12 VDD.n386 VDD.t388 396.079
R13 VDD.n1570 VDD.t588 382.793
R14 VDD.n1209 VDD.t575 382.793
R15 VDD.n1178 VDD.t586 382.793
R16 VDD.n1180 VDD.t584 382.793
R17 VDD.n1157 VDD.t581 382.793
R18 VDD.n790 VDD.t391 382.793
R19 VDD.n429 VDD.t491 382.793
R20 VDD.n398 VDD.t516 382.793
R21 VDD.n400 VDD.t938 382.793
R22 VDD.n377 VDD.t512 382.793
R23 VDD.n812 VDD.t479 382.793
R24 VDD.n6 VDD.t787 382.793
R25 VDD VDD.t428 374.711
R26 VDD VDD.t64 374.711
R27 VDD VDD.t456 374.711
R28 VDD VDD.t506 374.711
R29 VDD VDD.t592 374.711
R30 VDD VDD.t485 374.711
R31 VDD.n1554 VDD.t589 370.341
R32 VDD.n1526 VDD.t509 370.341
R33 VDD.n1522 VDD.t605 370.341
R34 VDD.n1212 VDD.t443 370.341
R35 VDD.n774 VDD.t515 370.341
R36 VDD.n746 VDD.t487 370.341
R37 VDD.n742 VDD.t77 370.341
R38 VDD.n432 VDD.t59 370.341
R39 VDD VDD.t568 370.303
R40 VDD VDD.t253 370.303
R41 VDD VDD.t68 331.981
R42 VDD VDD.t40 331.981
R43 VDD.n365 VDD 323.514
R44 VDD.n1232 VDD.t765 321.801
R45 VDD.n452 VDD.t51 321.801
R46 VDD.n1560 VDD.n1559 318.678
R47 VDD.n780 VDD.n779 318.678
R48 VDD.n1585 VDD.t762 318.108
R49 VDD.n805 VDD.t454 318.108
R50 VDD VDD.t500 313.839
R51 VDD VDD.t496 313.839
R52 VDD VDD.t750 313.839
R53 VDD.n1564 VDD.n1551 307.24
R54 VDD.n1525 VDD.n1524 307.24
R55 VDD.n1530 VDD.n1521 307.24
R56 VDD.n1208 VDD.n1207 307.24
R57 VDD.n784 VDD.n771 307.24
R58 VDD.n745 VDD.n744 307.24
R59 VDD.n750 VDD.n741 307.24
R60 VDD.n428 VDD.n427 307.24
R61 VDD.t68 VDD.t576 246.023
R62 VDD.t40 VDD.t936 246.023
R63 VDD VDD.t558 241.819
R64 VDD VDD.t606 241.819
R65 VDD.t582 VDD 233.643
R66 VDD.t428 VDD 233.643
R67 VDD.t64 VDD 233.643
R68 VDD.t568 VDD 233.643
R69 VDD.t456 VDD 233.643
R70 VDD.t752 VDD 233.643
R71 VDD.t506 VDD 233.643
R72 VDD.t592 VDD 233.643
R73 VDD.t253 VDD 233.643
R74 VDD.t485 VDD 233.643
R75 VDD.t310 VDD 227.321
R76 VDD VDD.t352 227.321
R77 VDD.t380 VDD 227.321
R78 VDD.t402 VDD 227.321
R79 VDD.t810 VDD 227.321
R80 VDD VDD.t852 227.321
R81 VDD.t880 VDD 227.321
R82 VDD VDD.t8 227.321
R83 VDD.t105 VDD 227.321
R84 VDD VDD.t103 227.321
R85 VDD.t179 VDD 227.321
R86 VDD.t237 VDD 227.321
R87 VDD VDD.t435 225.625
R88 VDD VDD.t774 225.625
R89 VDD VDD.t756 225.625
R90 VDD.n510 VDD.t363 204.903
R91 VDD.n907 VDD.t863 204.903
R92 VDD.n1290 VDD.t188 204.903
R93 VDD.n66 VDD.t675 204.9
R94 VDD.n546 VDD.t311 201.012
R95 VDD.n490 VDD.t353 201.012
R96 VDD.n455 VDD.t381 201.012
R97 VDD.n701 VDD.t403 201.012
R98 VDD.n943 VDD.t811 201.012
R99 VDD.n887 VDD.t853 201.012
R100 VDD.n1145 VDD.t881 201.012
R101 VDD.n1078 VDD.t9 201.012
R102 VDD.n1326 VDD.t106 201.012
R103 VDD.n1270 VDD.t104 201.012
R104 VDD.n1235 VDD.t180 201.012
R105 VDD.n1481 VDD.t238 201.012
R106 VDD.n83 VDD.t524 201.012
R107 VDD.n80 VDD.t705 201.012
R108 VDD.n217 VDD.t713 201.012
R109 VDD.n304 VDD.t655 201.012
R110 VDD.n814 VDD.n813 183.363
R111 VDD.n8 VDD.n7 183.363
R112 VDD.t452 VDD 179.821
R113 VDD.t60 VDD 179.821
R114 VDD.n1137 VDD.t565 179.821
R115 VDD.t565 VDD 179.821
R116 VDD.t46 VDD 179.821
R117 VDD.t560 VDD 179.821
R118 VDD.t563 VDD 179.821
R119 VDD.n1545 VDD.n1544 179.131
R120 VDD.n1219 VDD.n1205 179.131
R121 VDD.n1185 VDD.n1173 179.131
R122 VDD.n1177 VDD.n1176 179.131
R123 VDD.n1154 VDD.n1153 179.131
R124 VDD.n765 VDD.n764 179.131
R125 VDD.n439 VDD.n425 179.131
R126 VDD.n405 VDD.n393 179.131
R127 VDD.n397 VDD.n396 179.131
R128 VDD.n374 VDD.n373 179.131
R129 VDD.t251 VDD 174.602
R130 VDD.t768 VDD 174.602
R131 VDD.n674 VDD.n630 174.595
R132 VDD.n527 VDD.n526 174.595
R133 VDD.n553 VDD.n525 174.595
R134 VDD.n523 VDD.n522 174.595
R135 VDD.n560 VDD.n521 174.595
R136 VDD.n519 VDD.n507 174.595
R137 VDD.n509 VDD.n508 174.595
R138 VDD.n512 VDD.n511 174.595
R139 VDD.n493 VDD.n492 174.595
R140 VDD.n579 VDD.n495 174.595
R141 VDD.n497 VDD.n496 174.595
R142 VDD.n572 VDD.n499 174.595
R143 VDD.n537 VDD.n536 174.595
R144 VDD.n540 VDD.n535 174.595
R145 VDD.n534 VDD.n533 174.595
R146 VDD.n606 VDD.n605 174.595
R147 VDD.n612 VDD.n604 174.595
R148 VDD.n602 VDD.n601 174.595
R149 VDD.n619 VDD.n600 174.595
R150 VDD.n598 VDD.n485 174.595
R151 VDD.n487 VDD.n486 174.595
R152 VDD.n591 VDD.n489 174.595
R153 VDD.n473 VDD.n472 174.595
R154 VDD.n708 VDD.n471 174.595
R155 VDD.n470 VDD.n469 174.595
R156 VDD.n715 VDD.n466 174.595
R157 VDD.n464 VDD.n463 174.595
R158 VDD.n459 VDD.n458 174.595
R159 VDD.n726 VDD.n457 174.595
R160 VDD.n666 VDD.n633 174.595
R161 VDD.n635 VDD.n634 174.595
R162 VDD.n660 VDD.n637 174.595
R163 VDD.n654 VDD.n653 174.595
R164 VDD.n651 VDD.n640 174.595
R165 VDD.n646 VDD.n641 174.595
R166 VDD.n643 VDD.n642 174.595
R167 VDD.n1116 VDD.n1024 174.595
R168 VDD.n924 VDD.n923 174.595
R169 VDD.n950 VDD.n922 174.595
R170 VDD.n920 VDD.n919 174.595
R171 VDD.n957 VDD.n918 174.595
R172 VDD.n916 VDD.n904 174.595
R173 VDD.n906 VDD.n905 174.595
R174 VDD.n909 VDD.n908 174.595
R175 VDD.n890 VDD.n889 174.595
R176 VDD.n976 VDD.n892 174.595
R177 VDD.n894 VDD.n893 174.595
R178 VDD.n969 VDD.n896 174.595
R179 VDD.n934 VDD.n933 174.595
R180 VDD.n937 VDD.n932 174.595
R181 VDD.n931 VDD.n930 174.595
R182 VDD.n1003 VDD.n1002 174.595
R183 VDD.n1006 VDD.n1001 174.595
R184 VDD.n999 VDD.n998 174.595
R185 VDD.n1013 VDD.n997 174.595
R186 VDD.n995 VDD.n882 174.595
R187 VDD.n884 VDD.n883 174.595
R188 VDD.n988 VDD.n886 174.595
R189 VDD.n1072 VDD.n1041 174.595
R190 VDD.n1070 VDD.n1042 174.595
R191 VDD.n1064 VDD.n1063 174.595
R192 VDD.n1061 VDD.n1045 174.595
R193 VDD.n1055 VDD.n1054 174.595
R194 VDD.n1051 VDD.n1047 174.595
R195 VDD.n1049 VDD.n1048 174.595
R196 VDD.n1108 VDD.n1027 174.595
R197 VDD.n1029 VDD.n1028 174.595
R198 VDD.n1102 VDD.n1031 174.595
R199 VDD.n1096 VDD.n1095 174.595
R200 VDD.n1093 VDD.n1034 174.595
R201 VDD.n1086 VDD.n1085 174.595
R202 VDD.n1084 VDD.n1037 174.595
R203 VDD.n1454 VDD.n1410 174.595
R204 VDD.n1307 VDD.n1306 174.595
R205 VDD.n1333 VDD.n1305 174.595
R206 VDD.n1303 VDD.n1302 174.595
R207 VDD.n1340 VDD.n1301 174.595
R208 VDD.n1299 VDD.n1287 174.595
R209 VDD.n1289 VDD.n1288 174.595
R210 VDD.n1292 VDD.n1291 174.595
R211 VDD.n1273 VDD.n1272 174.595
R212 VDD.n1359 VDD.n1275 174.595
R213 VDD.n1277 VDD.n1276 174.595
R214 VDD.n1352 VDD.n1279 174.595
R215 VDD.n1317 VDD.n1316 174.595
R216 VDD.n1320 VDD.n1315 174.595
R217 VDD.n1314 VDD.n1313 174.595
R218 VDD.n1386 VDD.n1385 174.595
R219 VDD.n1392 VDD.n1384 174.595
R220 VDD.n1382 VDD.n1381 174.595
R221 VDD.n1399 VDD.n1380 174.595
R222 VDD.n1378 VDD.n1265 174.595
R223 VDD.n1267 VDD.n1266 174.595
R224 VDD.n1371 VDD.n1269 174.595
R225 VDD.n1253 VDD.n1252 174.595
R226 VDD.n1488 VDD.n1251 174.595
R227 VDD.n1250 VDD.n1249 174.595
R228 VDD.n1495 VDD.n1246 174.595
R229 VDD.n1244 VDD.n1243 174.595
R230 VDD.n1239 VDD.n1238 174.595
R231 VDD.n1506 VDD.n1237 174.595
R232 VDD.n1446 VDD.n1413 174.595
R233 VDD.n1415 VDD.n1414 174.595
R234 VDD.n1440 VDD.n1417 174.595
R235 VDD.n1434 VDD.n1433 174.595
R236 VDD.n1431 VDD.n1420 174.595
R237 VDD.n1426 VDD.n1421 174.595
R238 VDD.n1423 VDD.n1422 174.595
R239 VDD.n91 VDD.n90 174.595
R240 VDD.n117 VDD.n116 174.595
R241 VDD.n123 VDD.n122 174.595
R242 VDD.n129 VDD.n128 174.595
R243 VDD.n141 VDD.n140 174.595
R244 VDD.n146 VDD.n145 174.595
R245 VDD.n152 VDD.n151 174.595
R246 VDD.n158 VDD.n157 174.595
R247 VDD.n176 VDD.n175 174.595
R248 VDD.n182 VDD.n181 174.595
R249 VDD.n189 VDD.n188 174.595
R250 VDD.n198 VDD.n197 174.595
R251 VDD.n202 VDD.n201 174.595
R252 VDD.n208 VDD.n207 174.595
R253 VDD.n214 VDD.n213 174.595
R254 VDD.n245 VDD.n244 174.595
R255 VDD.n239 VDD.n238 174.595
R256 VDD.n232 VDD.n231 174.595
R257 VDD.n226 VDD.n225 174.595
R258 VDD.n222 VDD.n221 174.595
R259 VDD.n70 VDD.n69 174.595
R260 VDD.n65 VDD.n64 174.595
R261 VDD.n296 VDD.n295 174.595
R262 VDD.n290 VDD.n289 174.595
R263 VDD.n284 VDD.n283 174.595
R264 VDD.n278 VDD.n277 174.595
R265 VDD.n274 VDD.n273 174.595
R266 VDD.n268 VDD.n267 174.595
R267 VDD.n262 VDD.n261 174.595
R268 VDD.n341 VDD.n340 174.595
R269 VDD.n347 VDD.n346 174.595
R270 VDD.n353 VDD.n352 174.595
R271 VDD.n75 VDD.n74 174.595
R272 VDD.n306 VDD.n305 174.595
R273 VDD.n312 VDD.n311 174.595
R274 VDD.n318 VDD.n317 174.595
R275 VDD.t704 VDD 174.385
R276 VDD.t654 VDD 174.385
R277 VDD VDD.t614 173.083
R278 VDD.n695 VDD.t452 173.036
R279 VDD.n1475 VDD.t560 173.036
R280 VDD.t797 VDD 170.478
R281 VDD.t42 VDD 170.478
R282 VDD.n165 VDD 169.179
R283 VDD.n1583 VDD.n1540 169.107
R284 VDD.n1230 VDD.n1199 169.107
R285 VDD.n1195 VDD.n1169 169.107
R286 VDD.n1164 VDD.n1151 169.107
R287 VDD.n803 VDD.n760 169.107
R288 VDD.n450 VDD.n419 169.107
R289 VDD.n415 VDD.n389 169.107
R290 VDD.n384 VDD.n371 169.107
R291 VDD.n826 VDD.n807 169.107
R292 VDD.n819 VDD.n810 169.107
R293 VDD.n20 VDD.n1 169.107
R294 VDD.n13 VDD.n4 169.107
R295 VDD.n682 VDD.n681 169.017
R296 VDD.n1124 VDD.n1123 169.017
R297 VDD.n1462 VDD.n1461 169.017
R298 VDD.t500 VDD.t450 164.554
R299 VDD.t496 VDD.t49 164.554
R300 VDD.t750 VDD.t465 164.554
R301 VDD.n1550 VDD.n1549 164.215
R302 VDD.n1535 VDD.n1514 164.215
R303 VDD.n1519 VDD.n1518 164.215
R304 VDD.n1224 VDD.n1201 164.215
R305 VDD.n770 VDD.n769 164.215
R306 VDD.n755 VDD.n734 164.215
R307 VDD.n739 VDD.n738 164.215
R308 VDD.n444 VDD.n421 164.215
R309 VDD.n547 VDD.t317 158.117
R310 VDD.n585 VDD.t359 158.117
R311 VDD.n454 VDD.t293 158.117
R312 VDD.n702 VDD.t345 158.117
R313 VDD.n631 VDD.t399 158.117
R314 VDD.n944 VDD.t817 158.117
R315 VDD.n982 VDD.t859 158.117
R316 VDD.n1146 VDD.t921 158.117
R317 VDD.n1077 VDD.t845 158.117
R318 VDD.n1025 VDD.t37 158.117
R319 VDD.n1327 VDD.t178 158.117
R320 VDD.n1365 VDD.t176 158.117
R321 VDD.n1234 VDD.t102 158.117
R322 VDD.n1482 VDD.t120 158.117
R323 VDD.n1411 VDD.t234 158.117
R324 VDD.n85 VDD.t544 158.117
R325 VDD.n82 VDD.t735 158.117
R326 VDD.n79 VDD.t747 158.117
R327 VDD.n251 VDD.t721 158.117
R328 VDD.n302 VDD.t661 158.117
R329 VDD.n679 VDD.t453 158.06
R330 VDD.n1121 VDD.t566 158.06
R331 VDD.n1459 VDD.t561 158.06
R332 VDD.n100 VDD.t447 158.06
R333 VDD.n841 VDD.t457 158.06
R334 VDD.n839 VDD.t569 158.06
R335 VDD.n837 VDD.t65 158.06
R336 VDD.n835 VDD.t429 158.06
R337 VDD.n833 VDD.t583 158.06
R338 VDD.n363 VDD.t785 158.06
R339 VDD.n23 VDD.t753 158.06
R340 VDD.n24 VDD.t507 158.06
R341 VDD.n25 VDD.t593 158.06
R342 VDD.n26 VDD.t254 158.06
R343 VDD.n27 VDD.t486 158.06
R344 VDD.t558 VDD.t0 155.456
R345 VDD.t606 VDD.t782 155.456
R346 VDD.n253 VDD.t712 153.562
R347 VDD VDD.t74 151.137
R348 VDD VDD.t789 151.137
R349 VDD.n678 VDD.t438 151.123
R350 VDD.n1120 VDD.t777 151.123
R351 VDD.n1458 VDD.t759 151.123
R352 VDD.n95 VDD.t621 151.123
R353 VDD.t572 VDD.t570 148.481
R354 VDD.t463 VDD.t257 148.481
R355 VDD.t765 VDD.t482 145.243
R356 VDD.t51 VDD.t502 145.243
R357 VDD.t594 VDD.t467 143.232
R358 VDD.t388 VDD.t795 143.232
R359 VDD.t262 VDD.t362 142.5
R360 VDD.t368 VDD.t262 142.5
R361 VDD.t264 VDD.t368 142.5
R362 VDD.t350 VDD.t264 142.5
R363 VDD.t372 VDD.t350 142.5
R364 VDD.t384 VDD.t268 142.5
R365 VDD.t286 VDD.t384 142.5
R366 VDD.t272 VDD.t286 142.5
R367 VDD.t260 VDD.t272 142.5
R368 VDD.t290 VDD.t260 142.5
R369 VDD.t276 VDD.t290 142.5
R370 VDD.t308 VDD.t276 142.5
R371 VDD.t284 VDD.t308 142.5
R372 VDD.t316 VDD.t284 142.5
R373 VDD.t294 VDD.t310 142.5
R374 VDD.t282 VDD.t294 142.5
R375 VDD.t314 VDD.t282 142.5
R376 VDD.t298 VDD.t314 142.5
R377 VDD.t332 VDD.t318 142.5
R378 VDD.t318 VDD.t348 142.5
R379 VDD.t348 VDD.t334 142.5
R380 VDD.t334 VDD.t304 142.5
R381 VDD.t304 VDD.t338 142.5
R382 VDD.t338 VDD.t326 142.5
R383 VDD.t326 VDD.t354 142.5
R384 VDD.t354 VDD.t376 142.5
R385 VDD.t376 VDD.t366 142.5
R386 VDD.t366 VDD.t358 142.5
R387 VDD.t352 VDD.t342 142.5
R388 VDD.t342 VDD.t364 142.5
R389 VDD.t364 VDD.t346 142.5
R390 VDD.t346 VDD.t370 142.5
R391 VDD.t370 VDD.t266 142.5
R392 VDD.t374 VDD.t382 142.5
R393 VDD.t360 VDD.t374 142.5
R394 VDD.t386 VDD.t360 142.5
R395 VDD.t288 VDD.t386 142.5
R396 VDD.t274 VDD.t288 142.5
R397 VDD.t302 VDD.t274 142.5
R398 VDD.t378 VDD.t302 142.5
R399 VDD.t278 VDD.t378 142.5
R400 VDD.t292 VDD.t278 142.5
R401 VDD.t280 VDD.t380 142.5
R402 VDD.t312 VDD.t280 142.5
R403 VDD.t296 VDD.t312 142.5
R404 VDD.t270 VDD.t330 142.5
R405 VDD.t300 VDD.t270 142.5
R406 VDD.t320 VDD.t300 142.5
R407 VDD.t324 VDD.t320 142.5
R408 VDD.t336 VDD.t324 142.5
R409 VDD.t322 VDD.t336 142.5
R410 VDD.t306 VDD.t322 142.5
R411 VDD.t340 VDD.t306 142.5
R412 VDD.t328 VDD.t340 142.5
R413 VDD.t356 VDD.t328 142.5
R414 VDD.t344 VDD.t356 142.5
R415 VDD.t416 VDD.t402 142.5
R416 VDD.t410 VDD.t404 142.5
R417 VDD.t404 VDD.t408 142.5
R418 VDD.t408 VDD.t406 142.5
R419 VDD.t406 VDD.t418 142.5
R420 VDD.t418 VDD.t412 142.5
R421 VDD.t412 VDD.t424 142.5
R422 VDD.t424 VDD.t420 142.5
R423 VDD.t420 VDD.t414 142.5
R424 VDD.t414 VDD.t426 142.5
R425 VDD.t426 VDD.t422 142.5
R426 VDD.t422 VDD.t396 142.5
R427 VDD.t396 VDD.t400 142.5
R428 VDD.t400 VDD.t398 142.5
R429 VDD.t435 VDD.t433 142.5
R430 VDD.t433 VDD.t431 142.5
R431 VDD.t431 VDD.t437 142.5
R432 VDD.t890 VDD.t862 142.5
R433 VDD.t868 VDD.t890 142.5
R434 VDD.t892 VDD.t868 142.5
R435 VDD.t850 VDD.t892 142.5
R436 VDD.t872 VDD.t850 142.5
R437 VDD.t886 VDD.t896 142.5
R438 VDD.t914 VDD.t886 142.5
R439 VDD.t900 VDD.t914 142.5
R440 VDD.t888 VDD.t900 142.5
R441 VDD.t918 VDD.t888 142.5
R442 VDD.t906 VDD.t918 142.5
R443 VDD.t806 VDD.t906 142.5
R444 VDD.t912 VDD.t806 142.5
R445 VDD.t816 VDD.t912 142.5
R446 VDD.t922 VDD.t810 142.5
R447 VDD.t910 VDD.t922 142.5
R448 VDD.t814 VDD.t910 142.5
R449 VDD.t926 VDD.t814 142.5
R450 VDD.t830 VDD.t818 142.5
R451 VDD.t818 VDD.t846 142.5
R452 VDD.t846 VDD.t834 142.5
R453 VDD.t834 VDD.t804 142.5
R454 VDD.t804 VDD.t838 142.5
R455 VDD.t838 VDD.t824 142.5
R456 VDD.t824 VDD.t854 142.5
R457 VDD.t854 VDD.t876 142.5
R458 VDD.t876 VDD.t866 142.5
R459 VDD.t866 VDD.t858 142.5
R460 VDD.t852 VDD.t842 142.5
R461 VDD.t842 VDD.t864 142.5
R462 VDD.t864 VDD.t848 142.5
R463 VDD.t848 VDD.t870 142.5
R464 VDD.t870 VDD.t894 142.5
R465 VDD.t874 VDD.t882 142.5
R466 VDD.t860 VDD.t874 142.5
R467 VDD.t884 VDD.t860 142.5
R468 VDD.t916 VDD.t884 142.5
R469 VDD.t902 VDD.t916 142.5
R470 VDD.t802 VDD.t902 142.5
R471 VDD.t878 VDD.t802 142.5
R472 VDD.t904 VDD.t878 142.5
R473 VDD.t920 VDD.t904 142.5
R474 VDD.t908 VDD.t880 142.5
R475 VDD.t812 VDD.t908 142.5
R476 VDD.t924 VDD.t812 142.5
R477 VDD.t828 VDD.t898 142.5
R478 VDD.t898 VDD.t928 142.5
R479 VDD.t928 VDD.t832 142.5
R480 VDD.t832 VDD.t820 142.5
R481 VDD.t820 VDD.t836 142.5
R482 VDD.t836 VDD.t822 142.5
R483 VDD.t822 VDD.t808 142.5
R484 VDD.t808 VDD.t840 142.5
R485 VDD.t840 VDD.t826 142.5
R486 VDD.t826 VDD.t856 142.5
R487 VDD.t856 VDD.t844 142.5
R488 VDD.t8 VDD.t22 142.5
R489 VDD.t16 VDD.t10 142.5
R490 VDD.t10 VDD.t14 142.5
R491 VDD.t14 VDD.t12 142.5
R492 VDD.t12 VDD.t24 142.5
R493 VDD.t24 VDD.t18 142.5
R494 VDD.t18 VDD.t30 142.5
R495 VDD.t30 VDD.t26 142.5
R496 VDD.t26 VDD.t20 142.5
R497 VDD.t20 VDD.t32 142.5
R498 VDD.t32 VDD.t28 142.5
R499 VDD.t28 VDD.t34 142.5
R500 VDD.t34 VDD.t6 142.5
R501 VDD.t6 VDD.t36 142.5
R502 VDD.t774 VDD.t780 142.5
R503 VDD.t780 VDD.t778 142.5
R504 VDD.t778 VDD.t776 142.5
R505 VDD.t95 VDD.t187 142.5
R506 VDD.t213 VDD.t95 142.5
R507 VDD.t111 VDD.t213 142.5
R508 VDD.t185 VDD.t111 142.5
R509 VDD.t217 VDD.t185 142.5
R510 VDD.t165 VDD.t115 142.5
R511 VDD.t201 VDD.t165 142.5
R512 VDD.t125 VDD.t201 142.5
R513 VDD.t169 VDD.t125 142.5
R514 VDD.t205 VDD.t169 142.5
R515 VDD.t129 VDD.t205 142.5
R516 VDD.t151 VDD.t129 142.5
R517 VDD.t145 VDD.t151 142.5
R518 VDD.t177 VDD.t145 142.5
R519 VDD.t155 VDD.t105 142.5
R520 VDD.t211 VDD.t155 142.5
R521 VDD.t109 VDD.t211 142.5
R522 VDD.t159 VDD.t109 142.5
R523 VDD.t181 VDD.t121 142.5
R524 VDD.t121 VDD.t147 142.5
R525 VDD.t147 VDD.t199 142.5
R526 VDD.t199 VDD.t189 142.5
R527 VDD.t189 VDD.t97 142.5
R528 VDD.t97 VDD.t141 142.5
R529 VDD.t141 VDD.t171 142.5
R530 VDD.t171 VDD.t207 142.5
R531 VDD.t207 VDD.t133 142.5
R532 VDD.t133 VDD.t175 142.5
R533 VDD.t103 VDD.t153 142.5
R534 VDD.t153 VDD.t191 142.5
R535 VDD.t191 VDD.t183 142.5
R536 VDD.t183 VDD.t215 142.5
R537 VDD.t215 VDD.t113 142.5
R538 VDD.t91 VDD.t163 142.5
R539 VDD.t137 VDD.t91 142.5
R540 VDD.t167 VDD.t137 142.5
R541 VDD.t203 VDD.t167 142.5
R542 VDD.t127 VDD.t203 142.5
R543 VDD.t149 VDD.t127 142.5
R544 VDD.t117 VDD.t149 142.5
R545 VDD.t131 VDD.t117 142.5
R546 VDD.t101 VDD.t131 142.5
R547 VDD.t209 VDD.t179 142.5
R548 VDD.t107 VDD.t209 142.5
R549 VDD.t157 VDD.t107 142.5
R550 VDD.t135 VDD.t195 142.5
R551 VDD.t161 VDD.t135 142.5
R552 VDD.t197 VDD.t161 142.5
R553 VDD.t123 VDD.t197 142.5
R554 VDD.t93 VDD.t123 142.5
R555 VDD.t139 VDD.t93 142.5
R556 VDD.t193 VDD.t139 142.5
R557 VDD.t99 VDD.t193 142.5
R558 VDD.t143 VDD.t99 142.5
R559 VDD.t173 VDD.t143 142.5
R560 VDD.t119 VDD.t173 142.5
R561 VDD.t247 VDD.t237 142.5
R562 VDD.t225 VDD.t239 142.5
R563 VDD.t239 VDD.t223 142.5
R564 VDD.t223 VDD.t245 142.5
R565 VDD.t245 VDD.t249 142.5
R566 VDD.t249 VDD.t229 142.5
R567 VDD.t229 VDD.t241 142.5
R568 VDD.t241 VDD.t219 142.5
R569 VDD.t219 VDD.t231 142.5
R570 VDD.t231 VDD.t243 142.5
R571 VDD.t243 VDD.t221 142.5
R572 VDD.t221 VDD.t227 142.5
R573 VDD.t227 VDD.t235 142.5
R574 VDD.t235 VDD.t233 142.5
R575 VDD.t756 VDD.t760 142.5
R576 VDD.t760 VDD.t754 142.5
R577 VDD.t754 VDD.t758 142.5
R578 VDD.t482 VDD.t773 142.279
R579 VDD.t86 VDD.t770 142.279
R580 VDD.t502 VDD.t394 142.279
R581 VDD.t549 VDD.t564 142.279
R582 VDD.t762 VDD.t771 141.061
R583 VDD.t454 VDD.t392 141.061
R584 VDD.n696 VDD.t416 139.107
R585 VDD.n1139 VDD.t828 139.107
R586 VDD.n1476 VDD.t247 139.107
R587 VDD VDD.t478 138.857
R588 VDD VDD.t786 138.857
R589 VDD.t771 VDD.t489 138.183
R590 VDD.t441 VDD.t499 138.183
R591 VDD.t392 VDD.t505 138.183
R592 VDD.t444 VDD.t461 138.183
R593 VDD.t446 VDD 137.946
R594 VDD.t556 VDD.t251 134.732
R595 VDD.t552 VDD.t797 134.732
R596 VDD.t480 VDD.t768 134.732
R597 VDD.t83 VDD.t42 134.732
R598 VDD.n109 VDD.t446 132.74
R599 VDD VDD.t316 132.321
R600 VDD.t358 VDD 132.321
R601 VDD VDD.t292 132.321
R602 VDD.t330 VDD.n625 132.321
R603 VDD VDD.t344 132.321
R604 VDD.t398 VDD 132.321
R605 VDD VDD.t816 132.321
R606 VDD.t858 VDD 132.321
R607 VDD VDD.t920 132.321
R608 VDD.t844 VDD 132.321
R609 VDD.t22 VDD.n1138 132.321
R610 VDD.t36 VDD 132.321
R611 VDD VDD.t177 132.321
R612 VDD.t175 VDD 132.321
R613 VDD VDD.t101 132.321
R614 VDD.t195 VDD.n1405 132.321
R615 VDD VDD.t119 132.321
R616 VDD.t233 VDD 132.321
R617 VDD.t611 VDD.t556 131.983
R618 VDD.t562 VDD.t552 131.983
R619 VDD.t510 VDD.t259 131.983
R620 VDD.t767 VDD.t480 131.983
R621 VDD.t799 VDD.t83 131.983
R622 VDD.t764 VDD.t39 131.983
R623 VDD VDD.t255 129.228
R624 VDD VDD.t56 129.228
R625 VDD.t437 VDD 127.233
R626 VDD.t776 VDD 127.233
R627 VDD.t758 VDD 127.233
R628 VDD.t450 VDD.t60 122.144
R629 VDD.t49 VDD.t46 122.144
R630 VDD.t465 VDD.t563 122.144
R631 VDD.t933 VDD.t513 121.529
R632 VDD.t4 VDD.t62 121.529
R633 VDD.t0 VDD.t587 120.909
R634 VDD.t70 VDD.t66 120.909
R635 VDD.t782 VDD.t390 120.909
R636 VDD.t791 VDD.t494 120.909
R637 VDD.n1549 VDD.t75 117.451
R638 VDD.n1514 VDD.t585 117.451
R639 VDD.n1518 VDD.t73 117.451
R640 VDD.n1201 VDD.t577 117.451
R641 VDD.n769 VDD.t790 117.451
R642 VDD.n734 VDD.t462 117.451
R643 VDD.n738 VDD.t788 117.451
R644 VDD.n421 VDD.t937 117.451
R645 VDD.n1544 VDD.t1 116.322
R646 VDD.n1205 VDD.t514 116.322
R647 VDD.n1173 VDD.t460 116.322
R648 VDD.n1176 VDD.t256 116.322
R649 VDD.n1153 VDD.t470 116.322
R650 VDD.n764 VDD.t783 116.322
R651 VDD.n425 VDD.t63 116.322
R652 VDD.n393 VDD.t440 116.322
R653 VDD.n396 VDD.t57 116.322
R654 VDD.n373 VDD.t88 116.322
R655 VDD.n813 VDD.t573 116.322
R656 VDD.n7 VDD.t464 116.322
R657 VDD.t478 VDD.t572 115.486
R658 VDD.t786 VDD.t463 115.486
R659 VDD VDD.n695 115.358
R660 VDD.t882 VDD.n1018 115.358
R661 VDD VDD.n1475 115.358
R662 VDD.t578 VDD.t596 110.834
R663 VDD.t473 VDD.t930 110.834
R664 VDD.t718 VDD.t686 109.316
R665 VDD.t746 VDD.t718 109.316
R666 VDD.t732 VDD.t714 109.316
R667 VDD.t714 VDD.t692 109.316
R668 VDD.t692 VDD.t726 109.316
R669 VDD.t738 VDD.t708 109.316
R670 VDD.t630 VDD.t738 109.316
R671 VDD.t622 VDD.t630 109.316
R672 VDD.t730 VDD.t742 109.316
R673 VDD.t626 VDD.t730 109.316
R674 VDD.t650 VDD.t626 109.316
R675 VDD.t642 VDD.t650 109.316
R676 VDD.t658 VDD.t642 109.316
R677 VDD.t734 VDD.t658 109.316
R678 VDD.t523 VDD.t519 109.316
R679 VDD.t519 VDD.t517 109.316
R680 VDD.t517 VDD.t525 109.316
R681 VDD.t527 VDD.t531 109.316
R682 VDD.t533 VDD.t527 109.316
R683 VDD.t521 VDD.t533 109.316
R684 VDD.t529 VDD.t539 109.316
R685 VDD.t539 VDD.t535 109.316
R686 VDD.t535 VDD.t545 109.316
R687 VDD.t537 VDD.t541 109.316
R688 VDD.t547 VDD.t537 109.316
R689 VDD.t614 VDD.t618 109.316
R690 VDD.t618 VDD.t616 109.316
R691 VDD.t616 VDD.t620 109.316
R692 VDD.t656 VDD.t674 109.316
R693 VDD.t646 VDD.t656 109.316
R694 VDD.t678 VDD.t646 109.316
R695 VDD.t664 VDD.t678 109.316
R696 VDD.t690 VDD.t664 109.316
R697 VDD.t724 VDD.t690 109.316
R698 VDD.t696 VDD.t724 109.316
R699 VDD.t682 VDD.t696 109.316
R700 VDD.t670 VDD.t682 109.316
R701 VDD.t700 VDD.t670 109.316
R702 VDD.t728 VDD.t700 109.316
R703 VDD.t716 VDD.t728 109.316
R704 VDD.t744 VDD.t716 109.316
R705 VDD.t688 VDD.t744 109.316
R706 VDD.t720 VDD.t688 109.316
R707 VDD.t712 VDD.t706 109.316
R708 VDD.t706 VDD.t722 109.316
R709 VDD.t722 VDD.t748 109.316
R710 VDD.t748 VDD.t736 109.316
R711 VDD.t736 VDD.t634 109.316
R712 VDD.t634 VDD.t710 109.316
R713 VDD.t710 VDD.t740 109.316
R714 VDD.t624 VDD.t636 109.316
R715 VDD.t648 VDD.t624 109.316
R716 VDD.t638 VDD.t648 109.316
R717 VDD.t628 VDD.t638 109.316
R718 VDD.t652 VDD.t628 109.316
R719 VDD.t632 VDD.t652 109.316
R720 VDD.t660 VDD.t632 109.316
R721 VDD.t644 VDD.t654 109.316
R722 VDD.t382 VDD.n624 108.572
R723 VDD VDD.n1137 108.572
R724 VDD.t163 VDD.n1404 108.572
R725 VDD.t773 VDD.t86 106.709
R726 VDD.t394 VDD.t549 106.709
R727 VDD.t489 VDD.t441 103.636
R728 VDD.t505 VDD.t444 103.636
R729 VDD VDD.t746 101.507
R730 VDD VDD.t734 101.507
R731 VDD.t543 VDD 101.507
R732 VDD VDD.t720 101.507
R733 VDD VDD.t459 99.5409
R734 VDD VDD.t439 99.5409
R735 VDD.t477 VDD.t611 98.9875
R736 VDD.t259 VDD.t562 98.9875
R737 VDD.t38 VDD.t767 98.9875
R738 VDD.t39 VDD.t799 98.9875
R739 VDD.n164 VDD.t622 98.9046
R740 VDD.t550 VDD.t602 97.8793
R741 VDD.t475 VDD.t80 97.8793
R742 VDD.t620 VDD 97.6032
R743 VDD.n1540 VDD.t772 96.1553
R744 VDD.n1199 VDD.t483 96.1553
R745 VDD.n1169 VDD.t567 96.1553
R746 VDD.n1151 VDD.t468 96.1553
R747 VDD.n760 VDD.t393 96.1553
R748 VDD.n419 VDD.t503 96.1553
R749 VDD.n389 VDD.t932 96.1553
R750 VDD.n371 VDD.t796 96.1553
R751 VDD.n807 VDD.t553 96.1553
R752 VDD.n810 VDD.t557 96.1553
R753 VDD.n681 VDD.t451 96.1553
R754 VDD.n1123 VDD.t50 96.1553
R755 VDD.n1461 VDD.t466 96.1553
R756 VDD.n1 VDD.t84 96.1553
R757 VDD.n4 VDD.t481 96.1553
R758 VDD.n566 VDD.t298 95.0005
R759 VDD.n1346 VDD.t159 95.0005
R760 VDD.t770 VDD 94.8523
R761 VDD.t564 VDD 94.8523
R762 VDD.n1556 VDD.t579 93.81
R763 VDD.n776 VDD.t474 93.81
R764 VDD.t66 VDD 93.5611
R765 VDD.t494 VDD 93.5611
R766 VDD.t61 VDD 93.539
R767 VDD.t53 VDD 93.539
R768 VDD VDD.t477 93.4882
R769 VDD VDD.t38 93.4882
R770 VDD.t442 VDD 93.3702
R771 VDD.t58 VDD 93.3702
R772 VDD.t499 VDD 92.1217
R773 VDD.t461 VDD 92.1217
R774 VDD.t600 VDD.t574 91.8882
R775 VDD.t78 VDD.t490 91.8882
R776 VDD.t896 VDD.n962 91.6076
R777 VDD.n110 VDD.t547 91.0964
R778 VDD.t576 VDD.t448 88.9241
R779 VDD.t936 VDD.t554 88.9241
R780 VDD VDD.n109 88.4936
R781 VDD.n963 VDD.t926 88.2148
R782 VDD VDD.t510 87.9889
R783 VDD VDD.t764 87.9889
R784 VDD.t590 VDD 87.8035
R785 VDD.t47 VDD 87.8035
R786 VDD.t793 VDD.t430 87.6928
R787 VDD.t498 VDD.t580 87.6928
R788 VDD.t612 VDD.t445 87.6928
R789 VDD.t85 VDD.t511 87.6928
R790 VDD.n1551 VDD.t603 86.7743
R791 VDD.n1551 VDD.t597 86.7743
R792 VDD.n1524 VDD.t935 86.7743
R793 VDD.n1524 VDD.t604 86.7743
R794 VDD.n1521 VDD.t458 86.7743
R795 VDD.n1521 VDD.t504 86.7743
R796 VDD.n1207 VDD.t934 86.7743
R797 VDD.n1207 VDD.t601 86.7743
R798 VDD.n771 VDD.t81 86.7743
R799 VDD.n771 VDD.t931 86.7743
R800 VDD.n744 VDD.t3 86.7743
R801 VDD.n744 VDD.t82 86.7743
R802 VDD.n741 VDD.t610 86.7743
R803 VDD.n741 VDD.t800 86.7743
R804 VDD.n427 VDD.t5 86.7743
R805 VDD.n427 VDD.t79 86.7743
R806 VDD.t268 VDD.n565 84.8219
R807 VDD.t115 VDD.n1345 84.8219
R808 VDD.n1197 VDD.n1167 83.3098
R809 VDD.n417 VDD.n387 83.3098
R810 VDD.n329 VDD.t660 80.6854
R811 VDD.t676 VDD.t644 78.5727
R812 VDD.n135 VDD.t521 75.48
R813 VDD.t430 VDD.t469 70.1543
R814 VDD.t445 VDD.t87 70.1543
R815 VDD.n1559 VDD.t71 63.3219
R816 VDD.n1559 VDD.t67 63.3219
R817 VDD.n779 VDD.t792 63.3219
R818 VDD.n779 VDD.t495 63.3219
R819 VDD.n330 VDD.t732 59.8635
R820 VDD.n565 VDD.t372 57.6791
R821 VDD.n1345 VDD.t217 57.6791
R822 VDD.t587 VDD.t590 57.5763
R823 VDD.t390 VDD.t47 57.5763
R824 VDD VDD.t508 57.5434
R825 VDD VDD.t2 57.5434
R826 VDD.t574 VDD.t442 56.3188
R827 VDD.t490 VDD.t58 56.3188
R828 VDD.n963 VDD.t830 54.2862
R829 VDD.t467 VDD.t793 52.6159
R830 VDD.t580 VDD.t61 52.6159
R831 VDD.t795 VDD.t612 52.6159
R832 VDD.t511 VDD.t53 52.6159
R833 VDD.n962 VDD.t872 50.8934
R834 VDD.t471 VDD.t484 50.6439
R835 VDD.t54 VDD.t395 50.6439
R836 VDD.n330 VDD.t704 49.4526
R837 VDD.t662 VDD.t676 49.2598
R838 VDD.t640 VDD.t662 49.2598
R839 VDD.t680 VDD.t640 49.2598
R840 VDD.t666 VDD.t680 49.2598
R841 VDD.t694 VDD.t666 49.2598
R842 VDD.t668 VDD.t694 49.2598
R843 VDD.t698 VDD.t668 49.2598
R844 VDD.t684 VDD.t698 49.2598
R845 VDD.t672 VDD.t684 49.2598
R846 VDD.t702 VDD.t672 49.2598
R847 VDD.t686 VDD.t702 47.9846
R848 VDD.n566 VDD.t332 47.5005
R849 VDD.n1346 VDD.t181 47.5005
R850 VDD.n1167 VDD 43.6586
R851 VDD.n387 VDD 43.6586
R852 VDD.n1549 VDD.t591 42.3555
R853 VDD.n1514 VDD.t940 42.3555
R854 VDD.n1518 VDD.t90 42.3555
R855 VDD.n1201 VDD.t69 42.3555
R856 VDD.n769 VDD.t48 42.3555
R857 VDD.n734 VDD.t609 42.3555
R858 VDD.n738 VDD.t45 42.3555
R859 VDD.n421 VDD.t41 42.3555
R860 VDD.n1220 VDD.n1203 39.2858
R861 VDD.n440 VDD.n423 39.2858
R862 VDD.n369 VDD.n368 39.2858
R863 VDD VDD.t72 39.0862
R864 VDD VDD.t76 39.0862
R865 VDD.t602 VDD.t578 38.8641
R866 VDD.t80 VDD.t473 38.8641
R867 VDD.n1159 VDD.n1152 38.7881
R868 VDD.n379 VDD.n372 38.7881
R869 VDD.n1229 VDD.n1228 38.7811
R870 VDD.n449 VDD.n448 38.7811
R871 VDD.t448 VDD.t933 38.534
R872 VDD.t554 VDD.t4 38.534
R873 VDD.t469 VDD.t498 35.0774
R874 VDD.t87 VDD.t85 35.0774
R875 VDD.n1582 VDD.n1581 34.6358
R876 VDD.n1581 VDD.n1541 34.6358
R877 VDD.n1577 VDD.n1541 34.6358
R878 VDD.n1577 VDD.n1576 34.6358
R879 VDD.n1576 VDD.n1542 34.6358
R880 VDD.n1572 VDD.n1571 34.6358
R881 VDD.n1569 VDD.n1546 34.6358
R882 VDD.n1560 VDD.n1558 34.6358
R883 VDD.n1566 VDD.n1565 34.6358
R884 VDD.n1534 VDD.n1516 34.6358
R885 VDD.n1532 VDD.n1531 34.6358
R886 VDD.n1223 VDD.n1202 34.6358
R887 VDD.n1218 VDD.n1206 34.6358
R888 VDD.n1184 VDD.n1174 34.6358
R889 VDD.n1194 VDD.n1193 34.6358
R890 VDD.n1193 VDD.n1170 34.6358
R891 VDD.n1189 VDD.n1170 34.6358
R892 VDD.n1189 VDD.n1188 34.6358
R893 VDD.n1188 VDD.n1171 34.6358
R894 VDD.n1182 VDD.n1181 34.6358
R895 VDD.n1156 VDD.n1155 34.6358
R896 VDD.n1163 VDD.n1152 34.6358
R897 VDD.n802 VDD.n801 34.6358
R898 VDD.n801 VDD.n761 34.6358
R899 VDD.n797 VDD.n761 34.6358
R900 VDD.n797 VDD.n796 34.6358
R901 VDD.n796 VDD.n762 34.6358
R902 VDD.n792 VDD.n791 34.6358
R903 VDD.n789 VDD.n766 34.6358
R904 VDD.n780 VDD.n778 34.6358
R905 VDD.n786 VDD.n785 34.6358
R906 VDD.n754 VDD.n736 34.6358
R907 VDD.n752 VDD.n751 34.6358
R908 VDD.n443 VDD.n422 34.6358
R909 VDD.n438 VDD.n426 34.6358
R910 VDD.n404 VDD.n394 34.6358
R911 VDD.n414 VDD.n413 34.6358
R912 VDD.n413 VDD.n390 34.6358
R913 VDD.n409 VDD.n390 34.6358
R914 VDD.n409 VDD.n408 34.6358
R915 VDD.n408 VDD.n391 34.6358
R916 VDD.n402 VDD.n401 34.6358
R917 VDD.n376 VDD.n375 34.6358
R918 VDD.n383 VDD.n372 34.6358
R919 VDD.n846 VDD.n845 34.6358
R920 VDD.n845 VDD.n840 34.6358
R921 VDD.n850 VDD.n838 34.6358
R922 VDD.n856 VDD.n855 34.6358
R923 VDD.n855 VDD.n836 34.6358
R924 VDD.n861 VDD.n860 34.6358
R925 VDD.n860 VDD.n834 34.6358
R926 VDD.n820 VDD.n808 34.6358
R927 VDD.n824 VDD.n808 34.6358
R928 VDD.n825 VDD.n824 34.6358
R929 VDD.n818 VDD.n811 34.6358
R930 VDD.n518 VDD.n516 34.6358
R931 VDD.n561 VDD.n520 34.6358
R932 VDD.n559 VDD.n558 34.6358
R933 VDD.n555 VDD.n554 34.6358
R934 VDD.n549 VDD.n548 34.6358
R935 VDD.n545 VDD.n531 34.6358
R936 VDD.n539 VDD.n538 34.6358
R937 VDD.n571 VDD.n500 34.6358
R938 VDD.n574 VDD.n573 34.6358
R939 VDD.n578 VDD.n577 34.6358
R940 VDD.n584 VDD.n583 34.6358
R941 VDD.n590 VDD.n589 34.6358
R942 VDD.n597 VDD.n595 34.6358
R943 VDD.n620 VDD.n599 34.6358
R944 VDD.n618 VDD.n617 34.6358
R945 VDD.n614 VDD.n613 34.6358
R946 VDD.n608 VDD.n607 34.6358
R947 VDD.n728 VDD.n727 34.6358
R948 VDD.n721 VDD.n720 34.6358
R949 VDD.n717 VDD.n716 34.6358
R950 VDD.n714 VDD.n467 34.6358
R951 VDD.n710 VDD.n709 34.6358
R952 VDD.n704 VDD.n703 34.6358
R953 VDD.n700 VDD.n477 34.6358
R954 VDD.n650 VDD.n647 34.6358
R955 VDD.n655 VDD.n652 34.6358
R956 VDD.n659 VDD.n638 34.6358
R957 VDD.n662 VDD.n661 34.6358
R958 VDD.n668 VDD.n667 34.6358
R959 VDD.n674 VDD.n673 34.6358
R960 VDD.n674 VDD.n628 34.6358
R961 VDD.n691 VDD.n690 34.6358
R962 VDD.n687 VDD.n686 34.6358
R963 VDD.n686 VDD.n680 34.6358
R964 VDD.n915 VDD.n913 34.6358
R965 VDD.n958 VDD.n917 34.6358
R966 VDD.n956 VDD.n955 34.6358
R967 VDD.n952 VDD.n951 34.6358
R968 VDD.n946 VDD.n945 34.6358
R969 VDD.n942 VDD.n928 34.6358
R970 VDD.n936 VDD.n935 34.6358
R971 VDD.n968 VDD.n897 34.6358
R972 VDD.n971 VDD.n970 34.6358
R973 VDD.n975 VDD.n974 34.6358
R974 VDD.n981 VDD.n980 34.6358
R975 VDD.n987 VDD.n986 34.6358
R976 VDD.n994 VDD.n992 34.6358
R977 VDD.n1014 VDD.n996 34.6358
R978 VDD.n1012 VDD.n1011 34.6358
R979 VDD.n1008 VDD.n1007 34.6358
R980 VDD.n1147 VDD.n872 34.6358
R981 VDD.n1144 VDD.n874 34.6358
R982 VDD.n1056 VDD.n1053 34.6358
R983 VDD.n1060 VDD.n1046 34.6358
R984 VDD.n1065 VDD.n1062 34.6358
R985 VDD.n1069 VDD.n1043 34.6358
R986 VDD.n1073 VDD.n1039 34.6358
R987 VDD.n1083 VDD.n1038 34.6358
R988 VDD.n1092 VDD.n1035 34.6358
R989 VDD.n1097 VDD.n1094 34.6358
R990 VDD.n1101 VDD.n1032 34.6358
R991 VDD.n1104 VDD.n1103 34.6358
R992 VDD.n1110 VDD.n1109 34.6358
R993 VDD.n1116 VDD.n1115 34.6358
R994 VDD.n1116 VDD.n1022 34.6358
R995 VDD.n1133 VDD.n1132 34.6358
R996 VDD.n1129 VDD.n1128 34.6358
R997 VDD.n1128 VDD.n1122 34.6358
R998 VDD.n1298 VDD.n1296 34.6358
R999 VDD.n1341 VDD.n1300 34.6358
R1000 VDD.n1339 VDD.n1338 34.6358
R1001 VDD.n1335 VDD.n1334 34.6358
R1002 VDD.n1329 VDD.n1328 34.6358
R1003 VDD.n1325 VDD.n1311 34.6358
R1004 VDD.n1319 VDD.n1318 34.6358
R1005 VDD.n1351 VDD.n1280 34.6358
R1006 VDD.n1354 VDD.n1353 34.6358
R1007 VDD.n1358 VDD.n1357 34.6358
R1008 VDD.n1364 VDD.n1363 34.6358
R1009 VDD.n1370 VDD.n1369 34.6358
R1010 VDD.n1377 VDD.n1375 34.6358
R1011 VDD.n1400 VDD.n1379 34.6358
R1012 VDD.n1398 VDD.n1397 34.6358
R1013 VDD.n1394 VDD.n1393 34.6358
R1014 VDD.n1388 VDD.n1387 34.6358
R1015 VDD.n1508 VDD.n1507 34.6358
R1016 VDD.n1501 VDD.n1500 34.6358
R1017 VDD.n1497 VDD.n1496 34.6358
R1018 VDD.n1494 VDD.n1247 34.6358
R1019 VDD.n1490 VDD.n1489 34.6358
R1020 VDD.n1484 VDD.n1483 34.6358
R1021 VDD.n1480 VDD.n1257 34.6358
R1022 VDD.n1430 VDD.n1427 34.6358
R1023 VDD.n1435 VDD.n1432 34.6358
R1024 VDD.n1439 VDD.n1418 34.6358
R1025 VDD.n1442 VDD.n1441 34.6358
R1026 VDD.n1448 VDD.n1447 34.6358
R1027 VDD.n1454 VDD.n1453 34.6358
R1028 VDD.n1454 VDD.n1408 34.6358
R1029 VDD.n1471 VDD.n1470 34.6358
R1030 VDD.n1467 VDD.n1466 34.6358
R1031 VDD.n1466 VDD.n1460 34.6358
R1032 VDD.n51 VDD.n50 34.6358
R1033 VDD.n45 VDD.n44 34.6358
R1034 VDD.n33 VDD.n32 34.6358
R1035 VDD.n14 VDD.n2 34.6358
R1036 VDD.n18 VDD.n2 34.6358
R1037 VDD.n19 VDD.n18 34.6358
R1038 VDD.n12 VDD.n5 34.6358
R1039 VDD.n513 VDD.n512 34.2593
R1040 VDD.n541 VDD.n534 34.2593
R1041 VDD.n592 VDD.n591 34.2593
R1042 VDD.n726 VDD.n725 34.2593
R1043 VDD.n645 VDD.n643 34.2593
R1044 VDD.n910 VDD.n909 34.2593
R1045 VDD.n938 VDD.n931 34.2593
R1046 VDD.n989 VDD.n988 34.2593
R1047 VDD.n1050 VDD.n1049 34.2593
R1048 VDD.n1087 VDD.n1084 34.2593
R1049 VDD.n1293 VDD.n1292 34.2593
R1050 VDD.n1321 VDD.n1314 34.2593
R1051 VDD.n1372 VDD.n1371 34.2593
R1052 VDD.n1506 VDD.n1505 34.2593
R1053 VDD.n1425 VDD.n1423 34.2593
R1054 VDD.n624 VDD.t266 33.9291
R1055 VDD.n1404 VDD.t113 33.9291
R1056 VDD.n851 VDD.n850 33.8829
R1057 VDD.n39 VDD.n38 33.8829
R1058 VDD.n135 VDD.t529 33.8361
R1059 VDD.n552 VDD.n527 33.5064
R1060 VDD.n580 VDD.n493 33.5064
R1061 VDD.n611 VDD.n606 33.5064
R1062 VDD.n707 VDD.n473 33.5064
R1063 VDD.n666 VDD.n665 33.5064
R1064 VDD.n949 VDD.n924 33.5064
R1065 VDD.n977 VDD.n890 33.5064
R1066 VDD.n1005 VDD.n1003 33.5064
R1067 VDD.n1072 VDD.n1071 33.5064
R1068 VDD.n1108 VDD.n1107 33.5064
R1069 VDD.n1332 VDD.n1307 33.5064
R1070 VDD.n1360 VDD.n1273 33.5064
R1071 VDD.n1391 VDD.n1386 33.5064
R1072 VDD.n1487 VDD.n1253 33.5064
R1073 VDD.n1446 VDD.n1445 33.5064
R1074 VDD.t513 VDD.t600 32.6058
R1075 VDD.t62 VDD.t78 32.6058
R1076 VDD.n1536 VDD.n1535 32.1329
R1077 VDD.n756 VDD.n755 32.1329
R1078 VDD.t508 VDD.t939 31.4862
R1079 VDD.t72 VDD.t89 31.4862
R1080 VDD.t2 VDD.t608 31.4862
R1081 VDD.t76 VDD.t44 31.4862
R1082 VDD.n553 VDD.n552 29.7417
R1083 VDD.n580 VDD.n579 29.7417
R1084 VDD.n612 VDD.n611 29.7417
R1085 VDD.n708 VDD.n707 29.7417
R1086 VDD.n665 VDD.n635 29.7417
R1087 VDD.n950 VDD.n949 29.7417
R1088 VDD.n977 VDD.n976 29.7417
R1089 VDD.n1006 VDD.n1005 29.7417
R1090 VDD.n1071 VDD.n1070 29.7417
R1091 VDD.n1107 VDD.n1029 29.7417
R1092 VDD.n1333 VDD.n1332 29.7417
R1093 VDD.n1360 VDD.n1359 29.7417
R1094 VDD.n1392 VDD.n1391 29.7417
R1095 VDD.n1488 VDD.n1487 29.7417
R1096 VDD.n1445 VDD.n1415 29.7417
R1097 VDD.n547 VDD.n546 29.3652
R1098 VDD.n585 VDD.n490 29.3652
R1099 VDD.n455 VDD.n454 29.3652
R1100 VDD.n702 VDD.n701 29.3652
R1101 VDD.n944 VDD.n943 29.3652
R1102 VDD.n982 VDD.n887 29.3652
R1103 VDD.n1146 VDD.n1145 29.3652
R1104 VDD.n1078 VDD.n1077 29.3652
R1105 VDD.n1327 VDD.n1326 29.3652
R1106 VDD.n1365 VDD.n1270 29.3652
R1107 VDD.n1235 VDD.n1234 29.3652
R1108 VDD.n1482 VDD.n1481 29.3652
R1109 VDD.n83 VDD.n82 29.3652
R1110 VDD.n80 VDD.n79 29.3652
R1111 VDD.n513 VDD.n509 28.9887
R1112 VDD.n541 VDD.n540 28.9887
R1113 VDD.n592 VDD.n487 28.9887
R1114 VDD.n725 VDD.n459 28.9887
R1115 VDD.n646 VDD.n645 28.9887
R1116 VDD.n672 VDD.n631 28.9887
R1117 VDD.n910 VDD.n906 28.9887
R1118 VDD.n938 VDD.n937 28.9887
R1119 VDD.n989 VDD.n884 28.9887
R1120 VDD.n1051 VDD.n1050 28.9887
R1121 VDD.n1087 VDD.n1086 28.9887
R1122 VDD.n1114 VDD.n1025 28.9887
R1123 VDD.n1293 VDD.n1289 28.9887
R1124 VDD.n1321 VDD.n1320 28.9887
R1125 VDD.n1372 VDD.n1267 28.9887
R1126 VDD.n1505 VDD.n1239 28.9887
R1127 VDD.n1426 VDD.n1425 28.9887
R1128 VDD.n1452 VDD.n1411 28.9887
R1129 VDD.n86 VDD.n85 28.9887
R1130 VDD.n1544 VDD.t559 28.4628
R1131 VDD.n1205 VDD.t449 28.4628
R1132 VDD.n1173 VDD.t493 28.4628
R1133 VDD.n1176 VDD.t488 28.4628
R1134 VDD.n1153 VDD.t794 28.4628
R1135 VDD.n764 VDD.t607 28.4628
R1136 VDD.n425 VDD.t555 28.4628
R1137 VDD.n393 VDD.t599 28.4628
R1138 VDD.n396 VDD.t801 28.4628
R1139 VDD.n373 VDD.t613 28.4628
R1140 VDD.n813 VDD.t571 28.4628
R1141 VDD.n7 VDD.t258 28.4628
R1142 VDD.n1564 VDD.n1563 28.2358
R1143 VDD.n1527 VDD.n1525 28.2358
R1144 VDD.n1530 VDD.n1529 28.2358
R1145 VDD.n1213 VDD.n1208 28.2358
R1146 VDD.n784 VDD.n783 28.2358
R1147 VDD.n747 VDD.n745 28.2358
R1148 VDD.n750 VDD.n749 28.2358
R1149 VDD.n433 VDD.n428 28.2358
R1150 VDD.n1537 VDD 28.2291
R1151 VDD.n757 VDD 28.2291
R1152 VDD.n1558 VDD.n1557 27.4829
R1153 VDD.n778 VDD.n777 27.4829
R1154 VDD.n1018 VDD.t894 27.1434
R1155 VDD.n691 VDD.n678 27.1064
R1156 VDD.n1133 VDD.n1120 27.1064
R1157 VDD.n1471 VDD.n1458 27.1064
R1158 VDD.n1556 VDD.t551 26.9729
R1159 VDD.n776 VDD.t476 26.9729
R1160 VDD.n1540 VDD.t763 26.5955
R1161 VDD.n1199 VDD.t766 26.5955
R1162 VDD.n1169 VDD.t472 26.5955
R1163 VDD.n1151 VDD.t595 26.5955
R1164 VDD.n760 VDD.t455 26.5955
R1165 VDD.n419 VDD.t52 26.5955
R1166 VDD.n389 VDD.t55 26.5955
R1167 VDD.n371 VDD.t389 26.5955
R1168 VDD.n807 VDD.t798 26.5955
R1169 VDD.n810 VDD.t252 26.5955
R1170 VDD.n1 VDD.t43 26.5955
R1171 VDD.n4 VDD.t769 26.5955
R1172 VDD.n630 VDD.t434 26.5955
R1173 VDD.n630 VDD.t432 26.5955
R1174 VDD.n526 VDD.t309 26.5955
R1175 VDD.n526 VDD.t285 26.5955
R1176 VDD.n525 VDD.t291 26.5955
R1177 VDD.n525 VDD.t277 26.5955
R1178 VDD.n522 VDD.t273 26.5955
R1179 VDD.n522 VDD.t261 26.5955
R1180 VDD.n521 VDD.t385 26.5955
R1181 VDD.n521 VDD.t287 26.5955
R1182 VDD.n507 VDD.t373 26.5955
R1183 VDD.n507 VDD.t269 26.5955
R1184 VDD.n508 VDD.t265 26.5955
R1185 VDD.n508 VDD.t351 26.5955
R1186 VDD.n511 VDD.t263 26.5955
R1187 VDD.n511 VDD.t369 26.5955
R1188 VDD.n492 VDD.t377 26.5955
R1189 VDD.n492 VDD.t367 26.5955
R1190 VDD.n495 VDD.t327 26.5955
R1191 VDD.n495 VDD.t355 26.5955
R1192 VDD.n496 VDD.t305 26.5955
R1193 VDD.n496 VDD.t339 26.5955
R1194 VDD.n499 VDD.t349 26.5955
R1195 VDD.n499 VDD.t335 26.5955
R1196 VDD.n536 VDD.t333 26.5955
R1197 VDD.n536 VDD.t319 26.5955
R1198 VDD.n535 VDD.t315 26.5955
R1199 VDD.n535 VDD.t299 26.5955
R1200 VDD.n533 VDD.t295 26.5955
R1201 VDD.n533 VDD.t283 26.5955
R1202 VDD.n605 VDD.t379 26.5955
R1203 VDD.n605 VDD.t279 26.5955
R1204 VDD.n604 VDD.t275 26.5955
R1205 VDD.n604 VDD.t303 26.5955
R1206 VDD.n601 VDD.t387 26.5955
R1207 VDD.n601 VDD.t289 26.5955
R1208 VDD.n600 VDD.t375 26.5955
R1209 VDD.n600 VDD.t361 26.5955
R1210 VDD.n485 VDD.t267 26.5955
R1211 VDD.n485 VDD.t383 26.5955
R1212 VDD.n486 VDD.t347 26.5955
R1213 VDD.n486 VDD.t371 26.5955
R1214 VDD.n489 VDD.t343 26.5955
R1215 VDD.n489 VDD.t365 26.5955
R1216 VDD.n472 VDD.t329 26.5955
R1217 VDD.n472 VDD.t357 26.5955
R1218 VDD.n471 VDD.t307 26.5955
R1219 VDD.n471 VDD.t341 26.5955
R1220 VDD.n469 VDD.t337 26.5955
R1221 VDD.n469 VDD.t323 26.5955
R1222 VDD.n466 VDD.t321 26.5955
R1223 VDD.n466 VDD.t325 26.5955
R1224 VDD.n463 VDD.t271 26.5955
R1225 VDD.n463 VDD.t301 26.5955
R1226 VDD.n458 VDD.t297 26.5955
R1227 VDD.n458 VDD.t331 26.5955
R1228 VDD.n457 VDD.t281 26.5955
R1229 VDD.n457 VDD.t313 26.5955
R1230 VDD.n633 VDD.t397 26.5955
R1231 VDD.n633 VDD.t401 26.5955
R1232 VDD.n634 VDD.t427 26.5955
R1233 VDD.n634 VDD.t423 26.5955
R1234 VDD.n637 VDD.t421 26.5955
R1235 VDD.n637 VDD.t415 26.5955
R1236 VDD.n653 VDD.t413 26.5955
R1237 VDD.n653 VDD.t425 26.5955
R1238 VDD.n640 VDD.t407 26.5955
R1239 VDD.n640 VDD.t419 26.5955
R1240 VDD.n641 VDD.t405 26.5955
R1241 VDD.n641 VDD.t409 26.5955
R1242 VDD.n642 VDD.t417 26.5955
R1243 VDD.n642 VDD.t411 26.5955
R1244 VDD.n1024 VDD.t781 26.5955
R1245 VDD.n1024 VDD.t779 26.5955
R1246 VDD.n923 VDD.t807 26.5955
R1247 VDD.n923 VDD.t913 26.5955
R1248 VDD.n922 VDD.t919 26.5955
R1249 VDD.n922 VDD.t907 26.5955
R1250 VDD.n919 VDD.t901 26.5955
R1251 VDD.n919 VDD.t889 26.5955
R1252 VDD.n918 VDD.t887 26.5955
R1253 VDD.n918 VDD.t915 26.5955
R1254 VDD.n904 VDD.t873 26.5955
R1255 VDD.n904 VDD.t897 26.5955
R1256 VDD.n905 VDD.t893 26.5955
R1257 VDD.n905 VDD.t851 26.5955
R1258 VDD.n908 VDD.t891 26.5955
R1259 VDD.n908 VDD.t869 26.5955
R1260 VDD.n889 VDD.t877 26.5955
R1261 VDD.n889 VDD.t867 26.5955
R1262 VDD.n892 VDD.t825 26.5955
R1263 VDD.n892 VDD.t855 26.5955
R1264 VDD.n893 VDD.t805 26.5955
R1265 VDD.n893 VDD.t839 26.5955
R1266 VDD.n896 VDD.t847 26.5955
R1267 VDD.n896 VDD.t835 26.5955
R1268 VDD.n933 VDD.t831 26.5955
R1269 VDD.n933 VDD.t819 26.5955
R1270 VDD.n932 VDD.t815 26.5955
R1271 VDD.n932 VDD.t927 26.5955
R1272 VDD.n930 VDD.t923 26.5955
R1273 VDD.n930 VDD.t911 26.5955
R1274 VDD.n1002 VDD.t879 26.5955
R1275 VDD.n1002 VDD.t905 26.5955
R1276 VDD.n1001 VDD.t903 26.5955
R1277 VDD.n1001 VDD.t803 26.5955
R1278 VDD.n998 VDD.t885 26.5955
R1279 VDD.n998 VDD.t917 26.5955
R1280 VDD.n997 VDD.t875 26.5955
R1281 VDD.n997 VDD.t861 26.5955
R1282 VDD.n882 VDD.t895 26.5955
R1283 VDD.n882 VDD.t883 26.5955
R1284 VDD.n883 VDD.t849 26.5955
R1285 VDD.n883 VDD.t871 26.5955
R1286 VDD.n886 VDD.t843 26.5955
R1287 VDD.n886 VDD.t865 26.5955
R1288 VDD.n1041 VDD.t827 26.5955
R1289 VDD.n1041 VDD.t857 26.5955
R1290 VDD.n1042 VDD.t809 26.5955
R1291 VDD.n1042 VDD.t841 26.5955
R1292 VDD.n1063 VDD.t837 26.5955
R1293 VDD.n1063 VDD.t823 26.5955
R1294 VDD.n1045 VDD.t833 26.5955
R1295 VDD.n1045 VDD.t821 26.5955
R1296 VDD.n1054 VDD.t899 26.5955
R1297 VDD.n1054 VDD.t929 26.5955
R1298 VDD.n1047 VDD.t925 26.5955
R1299 VDD.n1047 VDD.t829 26.5955
R1300 VDD.n1048 VDD.t909 26.5955
R1301 VDD.n1048 VDD.t813 26.5955
R1302 VDD.n1027 VDD.t35 26.5955
R1303 VDD.n1027 VDD.t7 26.5955
R1304 VDD.n1028 VDD.t33 26.5955
R1305 VDD.n1028 VDD.t29 26.5955
R1306 VDD.n1031 VDD.t27 26.5955
R1307 VDD.n1031 VDD.t21 26.5955
R1308 VDD.n1095 VDD.t19 26.5955
R1309 VDD.n1095 VDD.t31 26.5955
R1310 VDD.n1034 VDD.t13 26.5955
R1311 VDD.n1034 VDD.t25 26.5955
R1312 VDD.n1085 VDD.t11 26.5955
R1313 VDD.n1085 VDD.t15 26.5955
R1314 VDD.n1037 VDD.t23 26.5955
R1315 VDD.n1037 VDD.t17 26.5955
R1316 VDD.n1410 VDD.t761 26.5955
R1317 VDD.n1410 VDD.t755 26.5955
R1318 VDD.n1306 VDD.t152 26.5955
R1319 VDD.n1306 VDD.t146 26.5955
R1320 VDD.n1305 VDD.t206 26.5955
R1321 VDD.n1305 VDD.t130 26.5955
R1322 VDD.n1302 VDD.t126 26.5955
R1323 VDD.n1302 VDD.t170 26.5955
R1324 VDD.n1301 VDD.t166 26.5955
R1325 VDD.n1301 VDD.t202 26.5955
R1326 VDD.n1287 VDD.t218 26.5955
R1327 VDD.n1287 VDD.t116 26.5955
R1328 VDD.n1288 VDD.t112 26.5955
R1329 VDD.n1288 VDD.t186 26.5955
R1330 VDD.n1291 VDD.t96 26.5955
R1331 VDD.n1291 VDD.t214 26.5955
R1332 VDD.n1272 VDD.t208 26.5955
R1333 VDD.n1272 VDD.t134 26.5955
R1334 VDD.n1275 VDD.t142 26.5955
R1335 VDD.n1275 VDD.t172 26.5955
R1336 VDD.n1276 VDD.t190 26.5955
R1337 VDD.n1276 VDD.t98 26.5955
R1338 VDD.n1279 VDD.t148 26.5955
R1339 VDD.n1279 VDD.t200 26.5955
R1340 VDD.n1316 VDD.t182 26.5955
R1341 VDD.n1316 VDD.t122 26.5955
R1342 VDD.n1315 VDD.t110 26.5955
R1343 VDD.n1315 VDD.t160 26.5955
R1344 VDD.n1313 VDD.t156 26.5955
R1345 VDD.n1313 VDD.t212 26.5955
R1346 VDD.n1385 VDD.t118 26.5955
R1347 VDD.n1385 VDD.t132 26.5955
R1348 VDD.n1384 VDD.t128 26.5955
R1349 VDD.n1384 VDD.t150 26.5955
R1350 VDD.n1381 VDD.t168 26.5955
R1351 VDD.n1381 VDD.t204 26.5955
R1352 VDD.n1380 VDD.t92 26.5955
R1353 VDD.n1380 VDD.t138 26.5955
R1354 VDD.n1265 VDD.t114 26.5955
R1355 VDD.n1265 VDD.t164 26.5955
R1356 VDD.n1266 VDD.t184 26.5955
R1357 VDD.n1266 VDD.t216 26.5955
R1358 VDD.n1269 VDD.t154 26.5955
R1359 VDD.n1269 VDD.t192 26.5955
R1360 VDD.n1252 VDD.t144 26.5955
R1361 VDD.n1252 VDD.t174 26.5955
R1362 VDD.n1251 VDD.t194 26.5955
R1363 VDD.n1251 VDD.t100 26.5955
R1364 VDD.n1249 VDD.t94 26.5955
R1365 VDD.n1249 VDD.t140 26.5955
R1366 VDD.n1246 VDD.t198 26.5955
R1367 VDD.n1246 VDD.t124 26.5955
R1368 VDD.n1243 VDD.t136 26.5955
R1369 VDD.n1243 VDD.t162 26.5955
R1370 VDD.n1238 VDD.t158 26.5955
R1371 VDD.n1238 VDD.t196 26.5955
R1372 VDD.n1237 VDD.t210 26.5955
R1373 VDD.n1237 VDD.t108 26.5955
R1374 VDD.n1413 VDD.t228 26.5955
R1375 VDD.n1413 VDD.t236 26.5955
R1376 VDD.n1414 VDD.t244 26.5955
R1377 VDD.n1414 VDD.t222 26.5955
R1378 VDD.n1417 VDD.t220 26.5955
R1379 VDD.n1417 VDD.t232 26.5955
R1380 VDD.n1433 VDD.t230 26.5955
R1381 VDD.n1433 VDD.t242 26.5955
R1382 VDD.n1420 VDD.t246 26.5955
R1383 VDD.n1420 VDD.t250 26.5955
R1384 VDD.n1421 VDD.t240 26.5955
R1385 VDD.n1421 VDD.t224 26.5955
R1386 VDD.n1422 VDD.t248 26.5955
R1387 VDD.n1422 VDD.t226 26.5955
R1388 VDD.n90 VDD.t619 26.5955
R1389 VDD.n90 VDD.t617 26.5955
R1390 VDD.n116 VDD.t538 26.5955
R1391 VDD.n116 VDD.t548 26.5955
R1392 VDD.n122 VDD.t546 26.5955
R1393 VDD.n122 VDD.t542 26.5955
R1394 VDD.n128 VDD.t540 26.5955
R1395 VDD.n128 VDD.t536 26.5955
R1396 VDD.n140 VDD.t522 26.5955
R1397 VDD.n140 VDD.t530 26.5955
R1398 VDD.n145 VDD.t528 26.5955
R1399 VDD.n145 VDD.t534 26.5955
R1400 VDD.n151 VDD.t526 26.5955
R1401 VDD.n151 VDD.t532 26.5955
R1402 VDD.n157 VDD.t520 26.5955
R1403 VDD.n157 VDD.t518 26.5955
R1404 VDD.n175 VDD.t643 26.5955
R1405 VDD.n175 VDD.t659 26.5955
R1406 VDD.n181 VDD.t627 26.5955
R1407 VDD.n181 VDD.t651 26.5955
R1408 VDD.n188 VDD.t743 26.5955
R1409 VDD.n188 VDD.t731 26.5955
R1410 VDD.n197 VDD.t631 26.5955
R1411 VDD.n197 VDD.t623 26.5955
R1412 VDD.n201 VDD.t709 26.5955
R1413 VDD.n201 VDD.t739 26.5955
R1414 VDD.n207 VDD.t693 26.5955
R1415 VDD.n207 VDD.t727 26.5955
R1416 VDD.n213 VDD.t733 26.5955
R1417 VDD.n213 VDD.t715 26.5955
R1418 VDD.n244 VDD.t745 26.5955
R1419 VDD.n244 VDD.t689 26.5955
R1420 VDD.n238 VDD.t729 26.5955
R1421 VDD.n238 VDD.t717 26.5955
R1422 VDD.n231 VDD.t671 26.5955
R1423 VDD.n231 VDD.t701 26.5955
R1424 VDD.n225 VDD.t697 26.5955
R1425 VDD.n225 VDD.t683 26.5955
R1426 VDD.n221 VDD.t691 26.5955
R1427 VDD.n221 VDD.t725 26.5955
R1428 VDD.n69 VDD.t679 26.5955
R1429 VDD.n69 VDD.t665 26.5955
R1430 VDD.n64 VDD.t657 26.5955
R1431 VDD.n64 VDD.t647 26.5955
R1432 VDD.n295 VDD.t653 26.5955
R1433 VDD.n295 VDD.t633 26.5955
R1434 VDD.n289 VDD.t639 26.5955
R1435 VDD.n289 VDD.t629 26.5955
R1436 VDD.n283 VDD.t625 26.5955
R1437 VDD.n283 VDD.t649 26.5955
R1438 VDD.n277 VDD.t741 26.5955
R1439 VDD.n277 VDD.t637 26.5955
R1440 VDD.n273 VDD.t635 26.5955
R1441 VDD.n273 VDD.t711 26.5955
R1442 VDD.n267 VDD.t749 26.5955
R1443 VDD.n267 VDD.t737 26.5955
R1444 VDD.n261 VDD.t707 26.5955
R1445 VDD.n261 VDD.t723 26.5955
R1446 VDD.n340 VDD.t687 26.5955
R1447 VDD.n340 VDD.t719 26.5955
R1448 VDD.n346 VDD.t673 26.5955
R1449 VDD.n346 VDD.t703 26.5955
R1450 VDD.n352 VDD.t699 26.5955
R1451 VDD.n352 VDD.t685 26.5955
R1452 VDD.n74 VDD.t695 26.5955
R1453 VDD.n74 VDD.t669 26.5955
R1454 VDD.n305 VDD.t681 26.5955
R1455 VDD.n305 VDD.t667 26.5955
R1456 VDD.n311 VDD.t663 26.5955
R1457 VDD.n311 VDD.t641 26.5955
R1458 VDD.n317 VDD.t645 26.5955
R1459 VDD.n317 VDD.t677 26.5955
R1460 VDD.n819 VDD.n818 25.977
R1461 VDD.n13 VDD.n12 25.977
R1462 VDD.t74 VDD.t550 25.9096
R1463 VDD.t789 VDD.t475 25.9096
R1464 VDD.n681 VDD.t501 25.6105
R1465 VDD.n1123 VDD.t497 25.6105
R1466 VDD.n1461 VDD.t751 25.6105
R1467 VDD.n826 VDD.n825 25.224
R1468 VDD.n20 VDD.n19 25.224
R1469 VDD.n555 VDD.n523 23.7181
R1470 VDD.n577 VDD.n497 23.7181
R1471 VDD.n614 VDD.n602 23.7181
R1472 VDD.n710 VDD.n470 23.7181
R1473 VDD.n661 VDD.n660 23.7181
R1474 VDD.n952 VDD.n920 23.7181
R1475 VDD.n974 VDD.n894 23.7181
R1476 VDD.n1008 VDD.n999 23.7181
R1477 VDD.n1064 VDD.n1043 23.7181
R1478 VDD.n1103 VDD.n1102 23.7181
R1479 VDD.n1335 VDD.n1303 23.7181
R1480 VDD.n1357 VDD.n1277 23.7181
R1481 VDD.n1394 VDD.n1382 23.7181
R1482 VDD.n1490 VDD.n1250 23.7181
R1483 VDD.n1441 VDD.n1440 23.7181
R1484 VDD.t596 VDD.t70 23.0308
R1485 VDD.t930 VDD.t791 23.0308
R1486 VDD.n1583 VDD.n1582 22.9652
R1487 VDD.n1230 VDD.n1229 22.9652
R1488 VDD.n1195 VDD.n1194 22.9652
R1489 VDD.n1164 VDD.n1163 22.9652
R1490 VDD.n803 VDD.n802 22.9652
R1491 VDD.n450 VDD.n449 22.9652
R1492 VDD.n415 VDD.n414 22.9652
R1493 VDD.n384 VDD.n383 22.9652
R1494 VDD.n519 VDD.n518 22.9652
R1495 VDD.n538 VDD.n537 22.9652
R1496 VDD.n598 VDD.n597 22.9652
R1497 VDD.n720 VDD.n464 22.9652
R1498 VDD.n651 VDD.n650 22.9652
R1499 VDD.n916 VDD.n915 22.9652
R1500 VDD.n935 VDD.n934 22.9652
R1501 VDD.n995 VDD.n994 22.9652
R1502 VDD.n1056 VDD.n1055 22.9652
R1503 VDD.n1093 VDD.n1092 22.9652
R1504 VDD.n1299 VDD.n1298 22.9652
R1505 VDD.n1318 VDD.n1317 22.9652
R1506 VDD.n1378 VDD.n1377 22.9652
R1507 VDD.n1500 VDD.n1244 22.9652
R1508 VDD.n1431 VDD.n1430 22.9652
R1509 VDD.n1167 VDD 22.7027
R1510 VDD.n387 VDD 22.7027
R1511 VDD.n1557 VDD.n1546 22.5887
R1512 VDD.n777 VDD.n766 22.5887
R1513 VDD.n820 VDD.n819 22.2123
R1514 VDD.n673 VDD.n672 22.2123
R1515 VDD.n678 VDD.n628 22.2123
R1516 VDD.n1115 VDD.n1114 22.2123
R1517 VDD.n1120 VDD.n1022 22.2123
R1518 VDD.n1453 VDD.n1452 22.2123
R1519 VDD.n1458 VDD.n1408 22.2123
R1520 VDD.n14 VDD.n13 22.2123
R1521 VDD.n546 VDD.n545 21.8358
R1522 VDD.n589 VDD.n490 21.8358
R1523 VDD.n728 VDD.n455 21.8358
R1524 VDD.n701 VDD.n700 21.8358
R1525 VDD.n943 VDD.n942 21.8358
R1526 VDD.n986 VDD.n887 21.8358
R1527 VDD.n1145 VDD.n1144 21.8358
R1528 VDD.n1078 VDD.n1038 21.8358
R1529 VDD.n1326 VDD.n1325 21.8358
R1530 VDD.n1369 VDD.n1270 21.8358
R1531 VDD.n1508 VDD.n1235 21.8358
R1532 VDD.n1481 VDD.n1480 21.8358
R1533 VDD.n548 VDD.n547 21.0829
R1534 VDD.n585 VDD.n584 21.0829
R1535 VDD.n607 VDD.n454 21.0829
R1536 VDD.n703 VDD.n702 21.0829
R1537 VDD.n668 VDD.n631 21.0829
R1538 VDD.n945 VDD.n944 21.0829
R1539 VDD.n982 VDD.n981 21.0829
R1540 VDD.n1147 VDD.n1146 21.0829
R1541 VDD.n1077 VDD.n1039 21.0829
R1542 VDD.n1110 VDD.n1025 21.0829
R1543 VDD.n1328 VDD.n1327 21.0829
R1544 VDD.n1365 VDD.n1364 21.0829
R1545 VDD.n1387 VDD.n1234 21.0829
R1546 VDD.n1483 VDD.n1482 21.0829
R1547 VDD.n1448 VDD.n1411 21.0829
R1548 VDD.n253 VDD 20.8224
R1549 VDD VDD.n329 20.8224
R1550 VDD.n1563 VDD.n1554 19.9534
R1551 VDD.n1527 VDD.n1526 19.9534
R1552 VDD.n1529 VDD.n1522 19.9534
R1553 VDD.n1213 VDD.n1212 19.9534
R1554 VDD.n783 VDD.n774 19.9534
R1555 VDD.n747 VDD.n746 19.9534
R1556 VDD.n749 VDD.n742 19.9534
R1557 VDD.n433 VDD.n432 19.9534
R1558 VDD.n110 VDD.t543 18.2197
R1559 VDD.n560 VDD.n559 17.6946
R1560 VDD.n573 VDD.n572 17.6946
R1561 VDD.n619 VDD.n618 17.6946
R1562 VDD.n715 VDD.n714 17.6946
R1563 VDD.n654 VDD.n638 17.6946
R1564 VDD.n957 VDD.n956 17.6946
R1565 VDD.n970 VDD.n969 17.6946
R1566 VDD.n1013 VDD.n1012 17.6946
R1567 VDD.n1062 VDD.n1061 17.6946
R1568 VDD.n1096 VDD.n1032 17.6946
R1569 VDD.n1340 VDD.n1339 17.6946
R1570 VDD.n1353 VDD.n1352 17.6946
R1571 VDD.n1399 VDD.n1398 17.6946
R1572 VDD.n1495 VDD.n1494 17.6946
R1573 VDD.n1434 VDD.n1418 17.6946
R1574 VDD.n1566 VDD.n1550 16.9417
R1575 VDD.n1535 VDD.n1534 16.9417
R1576 VDD.n1532 VDD.n1519 16.9417
R1577 VDD.n1224 VDD.n1223 16.9417
R1578 VDD.n786 VDD.n770 16.9417
R1579 VDD.n755 VDD.n754 16.9417
R1580 VDD.n752 VDD.n739 16.9417
R1581 VDD.n444 VDD.n443 16.9417
R1582 VDD.n561 VDD.n560 16.9417
R1583 VDD.n572 VDD.n571 16.9417
R1584 VDD.n620 VDD.n619 16.9417
R1585 VDD.n716 VDD.n715 16.9417
R1586 VDD.n655 VDD.n654 16.9417
R1587 VDD.n958 VDD.n957 16.9417
R1588 VDD.n969 VDD.n968 16.9417
R1589 VDD.n1014 VDD.n1013 16.9417
R1590 VDD.n1061 VDD.n1060 16.9417
R1591 VDD.n1097 VDD.n1096 16.9417
R1592 VDD.n1341 VDD.n1340 16.9417
R1593 VDD.n1352 VDD.n1351 16.9417
R1594 VDD.n1400 VDD.n1399 16.9417
R1595 VDD.n1496 VDD.n1495 16.9417
R1596 VDD.n1435 VDD.n1434 16.9417
R1597 VDD.n142 VDD.n141 16.9417
R1598 VDD.n199 VDD.n198 16.9417
R1599 VDD.n227 VDD.n226 16.9417
R1600 VDD.n279 VDD.n278 16.9417
R1601 VDD.n76 VDD.n75 16.9417
R1602 VDD.n1565 VDD.n1564 16.1887
R1603 VDD.n1525 VDD.n1516 16.1887
R1604 VDD.n1531 VDD.n1530 16.1887
R1605 VDD.n1208 VDD.n1202 16.1887
R1606 VDD.n785 VDD.n784 16.1887
R1607 VDD.n745 VDD.n736 16.1887
R1608 VDD.n751 VDD.n750 16.1887
R1609 VDD.n428 VDD.n422 16.1887
R1610 VDD.n863 VDD.n833 14.6892
R1611 VDD.n366 VDD.n365 14.5711
R1612 VDD.n564 VDD.n503 14.5711
R1613 VDD.n564 VDD.n563 14.5711
R1614 VDD.n568 VDD.n567 14.5711
R1615 VDD.n623 VDD.n481 14.5711
R1616 VDD.n623 VDD.n622 14.5711
R1617 VDD.n461 VDD.n460 14.5711
R1618 VDD.n462 VDD.n461 14.5711
R1619 VDD.n698 VDD.n697 14.5711
R1620 VDD.n697 VDD.n480 14.5711
R1621 VDD.n694 VDD.n626 14.5711
R1622 VDD.n694 VDD.n627 14.5711
R1623 VDD.n961 VDD.n900 14.5711
R1624 VDD.n961 VDD.n960 14.5711
R1625 VDD.n965 VDD.n964 14.5711
R1626 VDD.n1017 VDD.n878 14.5711
R1627 VDD.n1017 VDD.n1016 14.5711
R1628 VDD.n1141 VDD.n1140 14.5711
R1629 VDD.n1140 VDD.n877 14.5711
R1630 VDD.n1081 VDD.n1019 14.5711
R1631 VDD.n1089 VDD.n1019 14.5711
R1632 VDD.n1136 VDD.n1020 14.5711
R1633 VDD.n1136 VDD.n1021 14.5711
R1634 VDD.n1344 VDD.n1283 14.5711
R1635 VDD.n1344 VDD.n1343 14.5711
R1636 VDD.n1348 VDD.n1347 14.5711
R1637 VDD.n1403 VDD.n1261 14.5711
R1638 VDD.n1403 VDD.n1402 14.5711
R1639 VDD.n1241 VDD.n1240 14.5711
R1640 VDD.n1242 VDD.n1241 14.5711
R1641 VDD.n1478 VDD.n1477 14.5711
R1642 VDD.n1477 VDD.n1260 14.5711
R1643 VDD.n1474 VDD.n1406 14.5711
R1644 VDD.n1474 VDD.n1407 14.5711
R1645 VDD.t255 VDD.t471 13.9711
R1646 VDD.t459 VDD.t492 13.9711
R1647 VDD.t56 VDD.t54 13.9711
R1648 VDD.t439 VDD.t598 13.9711
R1649 VDD.n814 VDD.n812 13.3488
R1650 VDD.n8 VDD.n6 13.3488
R1651 VDD.n842 VDD.n841 12.9329
R1652 VDD.n364 VDD.n363 12.9329
R1653 VDD.n28 VDD.n27 12.9329
R1654 VDD.n101 VDD.n100 12.9329
R1655 VDD.n520 VDD.n519 11.6711
R1656 VDD.n537 VDD.n500 11.6711
R1657 VDD.n599 VDD.n598 11.6711
R1658 VDD.n717 VDD.n464 11.6711
R1659 VDD.n652 VDD.n651 11.6711
R1660 VDD.n917 VDD.n916 11.6711
R1661 VDD.n934 VDD.n897 11.6711
R1662 VDD.n996 VDD.n995 11.6711
R1663 VDD.n1055 VDD.n1046 11.6711
R1664 VDD.n1094 VDD.n1093 11.6711
R1665 VDD.n1300 VDD.n1299 11.6711
R1666 VDD.n1317 VDD.n1280 11.6711
R1667 VDD.n1379 VDD.n1378 11.6711
R1668 VDD.n1497 VDD.n1244 11.6711
R1669 VDD.n1432 VDD.n1431 11.6711
R1670 VDD.n147 VDD.n146 11.6711
R1671 VDD.n203 VDD.n202 11.6711
R1672 VDD.n223 VDD.n222 11.6711
R1673 VDD.n275 VDD.n274 11.6711
R1674 VDD.n307 VDD.n306 11.6711
R1675 VDD.n558 VDD.n523 10.9181
R1676 VDD.n574 VDD.n497 10.9181
R1677 VDD.n617 VDD.n602 10.9181
R1678 VDD.n470 VDD.n467 10.9181
R1679 VDD.n660 VDD.n659 10.9181
R1680 VDD.n955 VDD.n920 10.9181
R1681 VDD.n971 VDD.n894 10.9181
R1682 VDD.n1011 VDD.n999 10.9181
R1683 VDD.n1065 VDD.n1064 10.9181
R1684 VDD.n1102 VDD.n1101 10.9181
R1685 VDD.n1338 VDD.n1303 10.9181
R1686 VDD.n1354 VDD.n1277 10.9181
R1687 VDD.n1397 VDD.n1382 10.9181
R1688 VDD.n1250 VDD.n1247 10.9181
R1689 VDD.n1440 VDD.n1439 10.9181
R1690 VDD.n130 VDD.n129 10.9181
R1691 VDD.n190 VDD.n189 10.9181
R1692 VDD.n233 VDD.n232 10.9181
R1693 VDD.n285 VDD.n284 10.9181
R1694 VDD.n354 VDD.n353 10.9181
R1695 VDD.n1537 VDD 10.8576
R1696 VDD.n757 VDD 10.8576
R1697 VDD.n841 VDD.n840 10.5417
R1698 VDD.n839 VDD.n838 10.5417
R1699 VDD.n837 VDD.n836 10.5417
R1700 VDD.n835 VDD.n834 10.5417
R1701 VDD.n368 VDD.n363 10.5417
R1702 VDD.n690 VDD.n679 10.5417
R1703 VDD.n1132 VDD.n1121 10.5417
R1704 VDD.n1470 VDD.n1459 10.5417
R1705 VDD.t742 VDD.n164 10.4115
R1706 VDD.n625 VDD.t296 10.1791
R1707 VDD.n1138 VDD.t16 10.1791
R1708 VDD.n1405 VDD.t157 10.1791
R1709 VDD.n682 VDD.n680 10.1652
R1710 VDD.n1124 VDD.n1122 10.1652
R1711 VDD.n1462 VDD.n1460 10.1652
R1712 VDD.n1571 VDD.n1570 9.41227
R1713 VDD.n1209 VDD.n1206 9.41227
R1714 VDD.n1178 VDD.n1174 9.41227
R1715 VDD.n1181 VDD.n1180 9.41227
R1716 VDD.n1157 VDD.n1156 9.41227
R1717 VDD.n791 VDD.n790 9.41227
R1718 VDD.n429 VDD.n426 9.41227
R1719 VDD.n398 VDD.n394 9.41227
R1720 VDD.n401 VDD.n400 9.41227
R1721 VDD.n377 VDD.n376 9.41227
R1722 VDD.n868 VDD.n828 9.3005
R1723 VDD.n866 VDD.n865 9.3005
R1724 VDD.n865 VDD.n828 9.3005
R1725 VDD.n1210 VDD.n1209 8.79168
R1726 VDD.n1179 VDD.n1178 8.79168
R1727 VDD.n1180 VDD.n1179 8.79168
R1728 VDD.n1158 VDD.n1157 8.79168
R1729 VDD.n430 VDD.n429 8.79168
R1730 VDD.n399 VDD.n398 8.79168
R1731 VDD.n400 VDD.n399 8.79168
R1732 VDD.n378 VDD.n377 8.79168
R1733 VDD.n846 VDD.n839 8.28285
R1734 VDD.n851 VDD.n837 8.28285
R1735 VDD.n856 VDD.n835 8.28285
R1736 VDD.n861 VDD.n833 8.28285
R1737 VDD.n687 VDD.n679 8.28285
R1738 VDD.n1129 VDD.n1121 8.28285
R1739 VDD.n1467 VDD.n1459 8.28285
R1740 VDD.n51 VDD.n23 8.28285
R1741 VDD.n45 VDD.n24 8.28285
R1742 VDD.n39 VDD.n25 8.28285
R1743 VDD.n33 VDD.n26 8.28285
R1744 VDD.n1186 VDD.n1185 7.54105
R1745 VDD.n1154 VDD.n1150 7.54105
R1746 VDD.n406 VDD.n405 7.54105
R1747 VDD.n374 VDD.n370 7.54105
R1748 VDD.n1572 VDD.n1545 6.4005
R1749 VDD.n1219 VDD.n1218 6.4005
R1750 VDD.n1185 VDD.n1184 6.4005
R1751 VDD.n1182 VDD.n1177 6.4005
R1752 VDD.n1155 VDD.n1154 6.4005
R1753 VDD.n792 VDD.n765 6.4005
R1754 VDD.n439 VDD.n438 6.4005
R1755 VDD.n405 VDD.n404 6.4005
R1756 VDD.n402 VDD.n397 6.4005
R1757 VDD.n375 VDD.n374 6.4005
R1758 VDD.n516 VDD.n509 5.64756
R1759 VDD.n540 VDD.n539 5.64756
R1760 VDD.n595 VDD.n487 5.64756
R1761 VDD.n721 VDD.n459 5.64756
R1762 VDD.n647 VDD.n646 5.64756
R1763 VDD.n913 VDD.n906 5.64756
R1764 VDD.n937 VDD.n936 5.64756
R1765 VDD.n992 VDD.n884 5.64756
R1766 VDD.n1053 VDD.n1051 5.64756
R1767 VDD.n1086 VDD.n1035 5.64756
R1768 VDD.n1296 VDD.n1289 5.64756
R1769 VDD.n1320 VDD.n1319 5.64756
R1770 VDD.n1375 VDD.n1267 5.64756
R1771 VDD.n1501 VDD.n1239 5.64756
R1772 VDD.n1427 VDD.n1426 5.64756
R1773 VDD.n153 VDD.n152 5.64756
R1774 VDD.n209 VDD.n208 5.64756
R1775 VDD.n71 VDD.n70 5.64756
R1776 VDD.n269 VDD.n268 5.64756
R1777 VDD.n313 VDD.n312 5.64756
R1778 VDD.n258 VDD.n257 5.27114
R1779 VDD.n98 VDD.n97 5.27114
R1780 VDD.n325 VDD.n324 5.27114
R1781 VDD.n165 VDD.t523 5.20598
R1782 VDD.n866 VDD.n830 4.90677
R1783 VDD.n554 VDD.n553 4.89462
R1784 VDD.n579 VDD.n578 4.89462
R1785 VDD.n613 VDD.n612 4.89462
R1786 VDD.n709 VDD.n708 4.89462
R1787 VDD.n662 VDD.n635 4.89462
R1788 VDD.n951 VDD.n950 4.89462
R1789 VDD.n976 VDD.n975 4.89462
R1790 VDD.n1007 VDD.n1006 4.89462
R1791 VDD.n1070 VDD.n1069 4.89462
R1792 VDD.n1104 VDD.n1029 4.89462
R1793 VDD.n1334 VDD.n1333 4.89462
R1794 VDD.n1359 VDD.n1358 4.89462
R1795 VDD.n1393 VDD.n1392 4.89462
R1796 VDD.n1489 VDD.n1488 4.89462
R1797 VDD.n1442 VDD.n1415 4.89462
R1798 VDD.n124 VDD.n123 4.89462
R1799 VDD.n183 VDD.n182 4.89462
R1800 VDD.n240 VDD.n239 4.89462
R1801 VDD.n291 VDD.n290 4.89462
R1802 VDD.n348 VDD.n347 4.89462
R1803 VDD.n1555 VDD.n1554 4.6505
R1804 VDD.n1564 VDD.n1553 4.6505
R1805 VDD.n1558 VDD.n1553 4.6505
R1806 VDD.n1563 VDD.n1562 4.6505
R1807 VDD.n1557 VDD.n1548 4.6505
R1808 VDD.n1567 VDD.n1546 4.6505
R1809 VDD.n1569 VDD.n1568 4.6505
R1810 VDD.n1571 VDD.n1543 4.6505
R1811 VDD.n1573 VDD.n1572 4.6505
R1812 VDD.n1574 VDD.n1542 4.6505
R1813 VDD.n1576 VDD.n1575 4.6505
R1814 VDD.n1578 VDD.n1577 4.6505
R1815 VDD.n1579 VDD.n1541 4.6505
R1816 VDD.n1581 VDD.n1580 4.6505
R1817 VDD.n1582 VDD.n1539 4.6505
R1818 VDD.n1565 VDD.n1548 4.6505
R1819 VDD.n1567 VDD.n1566 4.6505
R1820 VDD.n1523 VDD.n1522 4.6505
R1821 VDD.n1530 VDD.n1520 4.6505
R1822 VDD.n1529 VDD.n1528 4.6505
R1823 VDD.n1531 VDD.n1517 4.6505
R1824 VDD.n1533 VDD.n1532 4.6505
R1825 VDD.n1526 VDD.n1523 4.6505
R1826 VDD.n1528 VDD.n1527 4.6505
R1827 VDD.n1525 VDD.n1520 4.6505
R1828 VDD.n1517 VDD.n1516 4.6505
R1829 VDD.n1534 VDD.n1533 4.6505
R1830 VDD.n1535 VDD.n1515 4.6505
R1831 VDD.n1212 VDD.n1211 4.6505
R1832 VDD.n1214 VDD.n1213 4.6505
R1833 VDD.n1216 VDD.n1208 4.6505
R1834 VDD.n1204 VDD.n1202 4.6505
R1835 VDD.n1223 VDD.n1222 4.6505
R1836 VDD.n1215 VDD.n1206 4.6505
R1837 VDD.n1218 VDD.n1217 4.6505
R1838 VDD.n1221 VDD.n1220 4.6505
R1839 VDD.n1229 VDD.n1198 4.6505
R1840 VDD.n1175 VDD.n1174 4.6505
R1841 VDD.n1184 VDD.n1183 4.6505
R1842 VDD.n1181 VDD.n1175 4.6505
R1843 VDD.n1183 VDD.n1182 4.6505
R1844 VDD.n1172 VDD.n1171 4.6505
R1845 VDD.n1188 VDD.n1187 4.6505
R1846 VDD.n1190 VDD.n1189 4.6505
R1847 VDD.n1191 VDD.n1170 4.6505
R1848 VDD.n1193 VDD.n1192 4.6505
R1849 VDD.n1194 VDD.n1168 4.6505
R1850 VDD.n1160 VDD.n1156 4.6505
R1851 VDD.n1161 VDD.n1155 4.6505
R1852 VDD.n1161 VDD.n1152 4.6505
R1853 VDD.n1163 VDD.n1162 4.6505
R1854 VDD.n775 VDD.n774 4.6505
R1855 VDD.n784 VDD.n773 4.6505
R1856 VDD.n778 VDD.n773 4.6505
R1857 VDD.n783 VDD.n782 4.6505
R1858 VDD.n777 VDD.n768 4.6505
R1859 VDD.n787 VDD.n766 4.6505
R1860 VDD.n789 VDD.n788 4.6505
R1861 VDD.n791 VDD.n763 4.6505
R1862 VDD.n793 VDD.n792 4.6505
R1863 VDD.n794 VDD.n762 4.6505
R1864 VDD.n796 VDD.n795 4.6505
R1865 VDD.n798 VDD.n797 4.6505
R1866 VDD.n799 VDD.n761 4.6505
R1867 VDD.n801 VDD.n800 4.6505
R1868 VDD.n802 VDD.n759 4.6505
R1869 VDD.n785 VDD.n768 4.6505
R1870 VDD.n787 VDD.n786 4.6505
R1871 VDD.n743 VDD.n742 4.6505
R1872 VDD.n750 VDD.n740 4.6505
R1873 VDD.n749 VDD.n748 4.6505
R1874 VDD.n751 VDD.n737 4.6505
R1875 VDD.n753 VDD.n752 4.6505
R1876 VDD.n746 VDD.n743 4.6505
R1877 VDD.n748 VDD.n747 4.6505
R1878 VDD.n745 VDD.n740 4.6505
R1879 VDD.n737 VDD.n736 4.6505
R1880 VDD.n754 VDD.n753 4.6505
R1881 VDD.n755 VDD.n735 4.6505
R1882 VDD.n432 VDD.n431 4.6505
R1883 VDD.n434 VDD.n433 4.6505
R1884 VDD.n436 VDD.n428 4.6505
R1885 VDD.n424 VDD.n422 4.6505
R1886 VDD.n443 VDD.n442 4.6505
R1887 VDD.n435 VDD.n426 4.6505
R1888 VDD.n438 VDD.n437 4.6505
R1889 VDD.n441 VDD.n440 4.6505
R1890 VDD.n449 VDD.n418 4.6505
R1891 VDD.n395 VDD.n394 4.6505
R1892 VDD.n404 VDD.n403 4.6505
R1893 VDD.n401 VDD.n395 4.6505
R1894 VDD.n403 VDD.n402 4.6505
R1895 VDD.n392 VDD.n391 4.6505
R1896 VDD.n408 VDD.n407 4.6505
R1897 VDD.n410 VDD.n409 4.6505
R1898 VDD.n411 VDD.n390 4.6505
R1899 VDD.n413 VDD.n412 4.6505
R1900 VDD.n414 VDD.n388 4.6505
R1901 VDD.n380 VDD.n376 4.6505
R1902 VDD.n381 VDD.n375 4.6505
R1903 VDD.n381 VDD.n372 4.6505
R1904 VDD.n383 VDD.n382 4.6505
R1905 VDD.n862 VDD.n861 4.6505
R1906 VDD.n860 VDD.n859 4.6505
R1907 VDD.n858 VDD.n834 4.6505
R1908 VDD.n857 VDD.n856 4.6505
R1909 VDD.n855 VDD.n854 4.6505
R1910 VDD.n853 VDD.n836 4.6505
R1911 VDD.n852 VDD.n851 4.6505
R1912 VDD.n850 VDD.n849 4.6505
R1913 VDD.n848 VDD.n838 4.6505
R1914 VDD.n847 VDD.n846 4.6505
R1915 VDD.n845 VDD.n844 4.6505
R1916 VDD.n843 VDD.n840 4.6505
R1917 VDD.n815 VDD.n811 4.6505
R1918 VDD.n819 VDD.n809 4.6505
R1919 VDD.n825 VDD.n806 4.6505
R1920 VDD.n824 VDD.n823 4.6505
R1921 VDD.n822 VDD.n808 4.6505
R1922 VDD.n821 VDD.n820 4.6505
R1923 VDD.n818 VDD.n817 4.6505
R1924 VDD.n368 VDD.n367 4.6505
R1925 VDD.n678 VDD.n677 4.6505
R1926 VDD.n672 VDD.n671 4.6505
R1927 VDD.n670 VDD.n631 4.6505
R1928 VDD.n701 VDD.n476 4.6505
R1929 VDD.n702 VDD.n475 4.6505
R1930 VDD.n730 VDD.n455 4.6505
R1931 VDD.n731 VDD.n454 4.6505
R1932 VDD.n587 VDD.n490 4.6505
R1933 VDD.n586 VDD.n585 4.6505
R1934 VDD.n546 VDD.n530 4.6505
R1935 VDD.n547 VDD.n529 4.6505
R1936 VDD.n684 VDD.n680 4.6505
R1937 VDD.n686 VDD.n685 4.6505
R1938 VDD.n688 VDD.n687 4.6505
R1939 VDD.n690 VDD.n689 4.6505
R1940 VDD.n692 VDD.n691 4.6505
R1941 VDD.n676 VDD.n628 4.6505
R1942 VDD.n675 VDD.n674 4.6505
R1943 VDD.n673 VDD.n629 4.6505
R1944 VDD.n669 VDD.n668 4.6505
R1945 VDD.n667 VDD.n632 4.6505
R1946 VDD.n665 VDD.n664 4.6505
R1947 VDD.n663 VDD.n662 4.6505
R1948 VDD.n661 VDD.n636 4.6505
R1949 VDD.n659 VDD.n658 4.6505
R1950 VDD.n657 VDD.n638 4.6505
R1951 VDD.n656 VDD.n655 4.6505
R1952 VDD.n652 VDD.n639 4.6505
R1953 VDD.n650 VDD.n649 4.6505
R1954 VDD.n648 VDD.n647 4.6505
R1955 VDD.n645 VDD.n644 4.6505
R1956 VDD.n478 VDD.n477 4.6505
R1957 VDD.n700 VDD.n699 4.6505
R1958 VDD.n703 VDD.n474 4.6505
R1959 VDD.n705 VDD.n704 4.6505
R1960 VDD.n707 VDD.n706 4.6505
R1961 VDD.n709 VDD.n468 4.6505
R1962 VDD.n711 VDD.n710 4.6505
R1963 VDD.n712 VDD.n467 4.6505
R1964 VDD.n714 VDD.n713 4.6505
R1965 VDD.n716 VDD.n465 4.6505
R1966 VDD.n718 VDD.n717 4.6505
R1967 VDD.n720 VDD.n719 4.6505
R1968 VDD.n722 VDD.n721 4.6505
R1969 VDD.n725 VDD.n724 4.6505
R1970 VDD.n727 VDD.n456 4.6505
R1971 VDD.n729 VDD.n728 4.6505
R1972 VDD.n607 VDD.n453 4.6505
R1973 VDD.n609 VDD.n608 4.6505
R1974 VDD.n611 VDD.n610 4.6505
R1975 VDD.n613 VDD.n603 4.6505
R1976 VDD.n615 VDD.n614 4.6505
R1977 VDD.n617 VDD.n616 4.6505
R1978 VDD.n618 VDD.n484 4.6505
R1979 VDD.n621 VDD.n620 4.6505
R1980 VDD.n599 VDD.n483 4.6505
R1981 VDD.n597 VDD.n596 4.6505
R1982 VDD.n595 VDD.n594 4.6505
R1983 VDD.n593 VDD.n592 4.6505
R1984 VDD.n590 VDD.n488 4.6505
R1985 VDD.n589 VDD.n588 4.6505
R1986 VDD.n584 VDD.n491 4.6505
R1987 VDD.n583 VDD.n582 4.6505
R1988 VDD.n581 VDD.n580 4.6505
R1989 VDD.n578 VDD.n494 4.6505
R1990 VDD.n577 VDD.n576 4.6505
R1991 VDD.n575 VDD.n574 4.6505
R1992 VDD.n573 VDD.n498 4.6505
R1993 VDD.n571 VDD.n570 4.6505
R1994 VDD.n569 VDD.n500 4.6505
R1995 VDD.n538 VDD.n501 4.6505
R1996 VDD.n539 VDD.n532 4.6505
R1997 VDD.n542 VDD.n541 4.6505
R1998 VDD.n543 VDD.n531 4.6505
R1999 VDD.n545 VDD.n544 4.6505
R2000 VDD.n548 VDD.n528 4.6505
R2001 VDD.n550 VDD.n549 4.6505
R2002 VDD.n552 VDD.n551 4.6505
R2003 VDD.n554 VDD.n524 4.6505
R2004 VDD.n556 VDD.n555 4.6505
R2005 VDD.n558 VDD.n557 4.6505
R2006 VDD.n559 VDD.n506 4.6505
R2007 VDD.n562 VDD.n561 4.6505
R2008 VDD.n520 VDD.n505 4.6505
R2009 VDD.n518 VDD.n517 4.6505
R2010 VDD.n516 VDD.n515 4.6505
R2011 VDD.n514 VDD.n513 4.6505
R2012 VDD.n1120 VDD.n1119 4.6505
R2013 VDD.n1114 VDD.n1113 4.6505
R2014 VDD.n1112 VDD.n1025 4.6505
R2015 VDD.n1079 VDD.n1078 4.6505
R2016 VDD.n1077 VDD.n1076 4.6505
R2017 VDD.n1145 VDD.n873 4.6505
R2018 VDD.n1146 VDD.n871 4.6505
R2019 VDD.n984 VDD.n887 4.6505
R2020 VDD.n983 VDD.n982 4.6505
R2021 VDD.n943 VDD.n927 4.6505
R2022 VDD.n944 VDD.n926 4.6505
R2023 VDD.n1126 VDD.n1122 4.6505
R2024 VDD.n1128 VDD.n1127 4.6505
R2025 VDD.n1130 VDD.n1129 4.6505
R2026 VDD.n1132 VDD.n1131 4.6505
R2027 VDD.n1134 VDD.n1133 4.6505
R2028 VDD.n1118 VDD.n1022 4.6505
R2029 VDD.n1117 VDD.n1116 4.6505
R2030 VDD.n1115 VDD.n1023 4.6505
R2031 VDD.n1111 VDD.n1110 4.6505
R2032 VDD.n1109 VDD.n1026 4.6505
R2033 VDD.n1107 VDD.n1106 4.6505
R2034 VDD.n1105 VDD.n1104 4.6505
R2035 VDD.n1103 VDD.n1030 4.6505
R2036 VDD.n1101 VDD.n1100 4.6505
R2037 VDD.n1099 VDD.n1032 4.6505
R2038 VDD.n1098 VDD.n1097 4.6505
R2039 VDD.n1094 VDD.n1033 4.6505
R2040 VDD.n1092 VDD.n1091 4.6505
R2041 VDD.n1090 VDD.n1035 4.6505
R2042 VDD.n1088 VDD.n1087 4.6505
R2043 VDD.n1083 VDD.n1082 4.6505
R2044 VDD.n1080 VDD.n1038 4.6505
R2045 VDD.n1075 VDD.n1039 4.6505
R2046 VDD.n1074 VDD.n1073 4.6505
R2047 VDD.n1071 VDD.n1040 4.6505
R2048 VDD.n1069 VDD.n1068 4.6505
R2049 VDD.n1067 VDD.n1043 4.6505
R2050 VDD.n1066 VDD.n1065 4.6505
R2051 VDD.n1062 VDD.n1044 4.6505
R2052 VDD.n1060 VDD.n1059 4.6505
R2053 VDD.n1058 VDD.n1046 4.6505
R2054 VDD.n1057 VDD.n1056 4.6505
R2055 VDD.n1053 VDD.n1052 4.6505
R2056 VDD.n1050 VDD.n875 4.6505
R2057 VDD.n1142 VDD.n874 4.6505
R2058 VDD.n1144 VDD.n1143 4.6505
R2059 VDD.n1148 VDD.n1147 4.6505
R2060 VDD.n872 VDD.n870 4.6505
R2061 VDD.n1005 VDD.n1004 4.6505
R2062 VDD.n1007 VDD.n1000 4.6505
R2063 VDD.n1009 VDD.n1008 4.6505
R2064 VDD.n1011 VDD.n1010 4.6505
R2065 VDD.n1012 VDD.n881 4.6505
R2066 VDD.n1015 VDD.n1014 4.6505
R2067 VDD.n996 VDD.n880 4.6505
R2068 VDD.n994 VDD.n993 4.6505
R2069 VDD.n992 VDD.n991 4.6505
R2070 VDD.n990 VDD.n989 4.6505
R2071 VDD.n987 VDD.n885 4.6505
R2072 VDD.n986 VDD.n985 4.6505
R2073 VDD.n981 VDD.n888 4.6505
R2074 VDD.n980 VDD.n979 4.6505
R2075 VDD.n978 VDD.n977 4.6505
R2076 VDD.n975 VDD.n891 4.6505
R2077 VDD.n974 VDD.n973 4.6505
R2078 VDD.n972 VDD.n971 4.6505
R2079 VDD.n970 VDD.n895 4.6505
R2080 VDD.n968 VDD.n967 4.6505
R2081 VDD.n966 VDD.n897 4.6505
R2082 VDD.n935 VDD.n898 4.6505
R2083 VDD.n936 VDD.n929 4.6505
R2084 VDD.n939 VDD.n938 4.6505
R2085 VDD.n940 VDD.n928 4.6505
R2086 VDD.n942 VDD.n941 4.6505
R2087 VDD.n945 VDD.n925 4.6505
R2088 VDD.n947 VDD.n946 4.6505
R2089 VDD.n949 VDD.n948 4.6505
R2090 VDD.n951 VDD.n921 4.6505
R2091 VDD.n953 VDD.n952 4.6505
R2092 VDD.n955 VDD.n954 4.6505
R2093 VDD.n956 VDD.n903 4.6505
R2094 VDD.n959 VDD.n958 4.6505
R2095 VDD.n917 VDD.n902 4.6505
R2096 VDD.n915 VDD.n914 4.6505
R2097 VDD.n913 VDD.n912 4.6505
R2098 VDD.n911 VDD.n910 4.6505
R2099 VDD.n1458 VDD.n1457 4.6505
R2100 VDD.n1452 VDD.n1451 4.6505
R2101 VDD.n1450 VDD.n1411 4.6505
R2102 VDD.n1481 VDD.n1256 4.6505
R2103 VDD.n1482 VDD.n1255 4.6505
R2104 VDD.n1510 VDD.n1235 4.6505
R2105 VDD.n1511 VDD.n1234 4.6505
R2106 VDD.n1367 VDD.n1270 4.6505
R2107 VDD.n1366 VDD.n1365 4.6505
R2108 VDD.n1326 VDD.n1310 4.6505
R2109 VDD.n1327 VDD.n1309 4.6505
R2110 VDD.n1464 VDD.n1460 4.6505
R2111 VDD.n1466 VDD.n1465 4.6505
R2112 VDD.n1468 VDD.n1467 4.6505
R2113 VDD.n1470 VDD.n1469 4.6505
R2114 VDD.n1472 VDD.n1471 4.6505
R2115 VDD.n1456 VDD.n1408 4.6505
R2116 VDD.n1455 VDD.n1454 4.6505
R2117 VDD.n1453 VDD.n1409 4.6505
R2118 VDD.n1449 VDD.n1448 4.6505
R2119 VDD.n1447 VDD.n1412 4.6505
R2120 VDD.n1445 VDD.n1444 4.6505
R2121 VDD.n1443 VDD.n1442 4.6505
R2122 VDD.n1441 VDD.n1416 4.6505
R2123 VDD.n1439 VDD.n1438 4.6505
R2124 VDD.n1437 VDD.n1418 4.6505
R2125 VDD.n1436 VDD.n1435 4.6505
R2126 VDD.n1432 VDD.n1419 4.6505
R2127 VDD.n1430 VDD.n1429 4.6505
R2128 VDD.n1428 VDD.n1427 4.6505
R2129 VDD.n1425 VDD.n1424 4.6505
R2130 VDD.n1258 VDD.n1257 4.6505
R2131 VDD.n1480 VDD.n1479 4.6505
R2132 VDD.n1483 VDD.n1254 4.6505
R2133 VDD.n1485 VDD.n1484 4.6505
R2134 VDD.n1487 VDD.n1486 4.6505
R2135 VDD.n1489 VDD.n1248 4.6505
R2136 VDD.n1491 VDD.n1490 4.6505
R2137 VDD.n1492 VDD.n1247 4.6505
R2138 VDD.n1494 VDD.n1493 4.6505
R2139 VDD.n1496 VDD.n1245 4.6505
R2140 VDD.n1498 VDD.n1497 4.6505
R2141 VDD.n1500 VDD.n1499 4.6505
R2142 VDD.n1502 VDD.n1501 4.6505
R2143 VDD.n1505 VDD.n1504 4.6505
R2144 VDD.n1507 VDD.n1236 4.6505
R2145 VDD.n1509 VDD.n1508 4.6505
R2146 VDD.n1387 VDD.n1233 4.6505
R2147 VDD.n1389 VDD.n1388 4.6505
R2148 VDD.n1391 VDD.n1390 4.6505
R2149 VDD.n1393 VDD.n1383 4.6505
R2150 VDD.n1395 VDD.n1394 4.6505
R2151 VDD.n1397 VDD.n1396 4.6505
R2152 VDD.n1398 VDD.n1264 4.6505
R2153 VDD.n1401 VDD.n1400 4.6505
R2154 VDD.n1379 VDD.n1263 4.6505
R2155 VDD.n1377 VDD.n1376 4.6505
R2156 VDD.n1375 VDD.n1374 4.6505
R2157 VDD.n1373 VDD.n1372 4.6505
R2158 VDD.n1370 VDD.n1268 4.6505
R2159 VDD.n1369 VDD.n1368 4.6505
R2160 VDD.n1364 VDD.n1271 4.6505
R2161 VDD.n1363 VDD.n1362 4.6505
R2162 VDD.n1361 VDD.n1360 4.6505
R2163 VDD.n1358 VDD.n1274 4.6505
R2164 VDD.n1357 VDD.n1356 4.6505
R2165 VDD.n1355 VDD.n1354 4.6505
R2166 VDD.n1353 VDD.n1278 4.6505
R2167 VDD.n1351 VDD.n1350 4.6505
R2168 VDD.n1349 VDD.n1280 4.6505
R2169 VDD.n1318 VDD.n1281 4.6505
R2170 VDD.n1319 VDD.n1312 4.6505
R2171 VDD.n1322 VDD.n1321 4.6505
R2172 VDD.n1323 VDD.n1311 4.6505
R2173 VDD.n1325 VDD.n1324 4.6505
R2174 VDD.n1328 VDD.n1308 4.6505
R2175 VDD.n1330 VDD.n1329 4.6505
R2176 VDD.n1332 VDD.n1331 4.6505
R2177 VDD.n1334 VDD.n1304 4.6505
R2178 VDD.n1336 VDD.n1335 4.6505
R2179 VDD.n1338 VDD.n1337 4.6505
R2180 VDD.n1339 VDD.n1286 4.6505
R2181 VDD.n1342 VDD.n1341 4.6505
R2182 VDD.n1300 VDD.n1285 4.6505
R2183 VDD.n1298 VDD.n1297 4.6505
R2184 VDD.n1296 VDD.n1295 4.6505
R2185 VDD.n1294 VDD.n1293 4.6505
R2186 VDD.n52 VDD.n51 4.6505
R2187 VDD.n50 VDD.n49 4.6505
R2188 VDD.n48 VDD.n47 4.6505
R2189 VDD.n46 VDD.n45 4.6505
R2190 VDD.n44 VDD.n43 4.6505
R2191 VDD.n42 VDD.n41 4.6505
R2192 VDD.n40 VDD.n39 4.6505
R2193 VDD.n38 VDD.n37 4.6505
R2194 VDD.n36 VDD.n35 4.6505
R2195 VDD.n34 VDD.n33 4.6505
R2196 VDD.n32 VDD.n31 4.6505
R2197 VDD.n30 VDD.n29 4.6505
R2198 VDD.n9 VDD.n5 4.6505
R2199 VDD.n13 VDD.n3 4.6505
R2200 VDD.n19 VDD.n0 4.6505
R2201 VDD.n18 VDD.n17 4.6505
R2202 VDD.n16 VDD.n2 4.6505
R2203 VDD.n15 VDD.n14 4.6505
R2204 VDD.n12 VDD.n11 4.6505
R2205 VDD.n345 VDD.n78 4.6505
R2206 VDD.n349 VDD.n348 4.6505
R2207 VDD.n351 VDD.n350 4.6505
R2208 VDD.n355 VDD.n354 4.6505
R2209 VDD.n357 VDD.n356 4.6505
R2210 VDD.n77 VDD.n76 4.6505
R2211 VDD.n308 VDD.n307 4.6505
R2212 VDD.n310 VDD.n309 4.6505
R2213 VDD.n314 VDD.n313 4.6505
R2214 VDD.n316 VDD.n315 4.6505
R2215 VDD.n96 VDD.n95 4.6505
R2216 VDD.n87 VDD.n86 4.6505
R2217 VDD.n85 VDD.n84 4.6505
R2218 VDD.n170 VDD.n83 4.6505
R2219 VDD.n172 VDD.n82 4.6505
R2220 VDD.n336 VDD.n80 4.6505
R2221 VDD.n337 VDD.n79 4.6505
R2222 VDD.n103 VDD.n102 4.6505
R2223 VDD.n106 VDD.n105 4.6505
R2224 VDD.n94 VDD.n93 4.6505
R2225 VDD.n92 VDD.n91 4.6505
R2226 VDD.n89 VDD.n88 4.6505
R2227 VDD.n114 VDD.n113 4.6505
R2228 VDD.n119 VDD.n118 4.6505
R2229 VDD.n121 VDD.n120 4.6505
R2230 VDD.n125 VDD.n124 4.6505
R2231 VDD.n127 VDD.n126 4.6505
R2232 VDD.n131 VDD.n130 4.6505
R2233 VDD.n134 VDD.n133 4.6505
R2234 VDD.n143 VDD.n142 4.6505
R2235 VDD.n148 VDD.n147 4.6505
R2236 VDD.n150 VDD.n149 4.6505
R2237 VDD.n154 VDD.n153 4.6505
R2238 VDD.n156 VDD.n155 4.6505
R2239 VDD.n160 VDD.n159 4.6505
R2240 VDD.n163 VDD.n162 4.6505
R2241 VDD.n174 VDD.n173 4.6505
R2242 VDD.n178 VDD.n177 4.6505
R2243 VDD.n180 VDD.n179 4.6505
R2244 VDD.n184 VDD.n183 4.6505
R2245 VDD.n186 VDD.n185 4.6505
R2246 VDD.n191 VDD.n190 4.6505
R2247 VDD.n196 VDD.n195 4.6505
R2248 VDD.n200 VDD.n199 4.6505
R2249 VDD.n204 VDD.n203 4.6505
R2250 VDD.n206 VDD.n205 4.6505
R2251 VDD.n210 VDD.n209 4.6505
R2252 VDD.n212 VDD.n211 4.6505
R2253 VDD.n216 VDD.n215 4.6505
R2254 VDD.n334 VDD.n333 4.6505
R2255 VDD.n339 VDD.n338 4.6505
R2256 VDD.n343 VDD.n342 4.6505
R2257 VDD.n323 VDD.n304 4.6505
R2258 VDD.n303 VDD.n302 4.6505
R2259 VDD.n218 VDD.n217 4.6505
R2260 VDD.n252 VDD.n251 4.6505
R2261 VDD.n320 VDD.n319 4.6505
R2262 VDD.n322 VDD.n321 4.6505
R2263 VDD.n300 VDD.n299 4.6505
R2264 VDD.n298 VDD.n297 4.6505
R2265 VDD.n294 VDD.n293 4.6505
R2266 VDD.n292 VDD.n291 4.6505
R2267 VDD.n288 VDD.n287 4.6505
R2268 VDD.n286 VDD.n285 4.6505
R2269 VDD.n282 VDD.n281 4.6505
R2270 VDD.n280 VDD.n279 4.6505
R2271 VDD.n276 VDD.n275 4.6505
R2272 VDD.n272 VDD.n271 4.6505
R2273 VDD.n270 VDD.n269 4.6505
R2274 VDD.n266 VDD.n265 4.6505
R2275 VDD.n264 VDD.n263 4.6505
R2276 VDD.n260 VDD.n259 4.6505
R2277 VDD.n249 VDD.n248 4.6505
R2278 VDD.n247 VDD.n246 4.6505
R2279 VDD.n243 VDD.n242 4.6505
R2280 VDD.n241 VDD.n240 4.6505
R2281 VDD.n237 VDD.n236 4.6505
R2282 VDD.n234 VDD.n233 4.6505
R2283 VDD.n230 VDD.n229 4.6505
R2284 VDD.n228 VDD.n227 4.6505
R2285 VDD.n224 VDD.n223 4.6505
R2286 VDD.n220 VDD.n219 4.6505
R2287 VDD.n72 VDD.n71 4.6505
R2288 VDD.n68 VDD.n67 4.6505
R2289 VDD.n66 VDD.n65 4.45149
R2290 VDD.n512 VDD.n510 4.4514
R2291 VDD.n909 VDD.n907 4.4514
R2292 VDD.n1292 VDD.n1290 4.4514
R2293 VDD.n683 VDD.n682 4.14756
R2294 VDD.n1125 VDD.n1124 4.14756
R2295 VDD.n1463 VDD.n1462 4.14756
R2296 VDD.n1570 VDD.n1569 4.14168
R2297 VDD.n790 VDD.n789 4.14168
R2298 VDD.n812 VDD.n811 4.14168
R2299 VDD.n6 VDD.n5 4.14168
R2300 VDD.n1550 VDD.n1547 4.05611
R2301 VDD.n770 VDD.n767 4.05611
R2302 VDD.n1519 VDD.n1513 4.05569
R2303 VDD.n1225 VDD.n1224 4.05569
R2304 VDD.n739 VDD.n733 4.05569
R2305 VDD.n445 VDD.n444 4.05569
R2306 VDD.n1584 VDD.n1583 4.01726
R2307 VDD.n1196 VDD.n1195 4.01726
R2308 VDD.n1165 VDD.n1164 4.01726
R2309 VDD.n804 VDD.n803 4.01726
R2310 VDD.n416 VDD.n415 4.01726
R2311 VDD.n385 VDD.n384 4.01726
R2312 VDD.n1231 VDD.n1230 4.01682
R2313 VDD.n451 VDD.n450 4.01682
R2314 VDD.n827 VDD.n826 3.96556
R2315 VDD.n21 VDD.n20 3.96556
R2316 VDD.n696 VDD.t410 3.39336
R2317 VDD.n1139 VDD.t924 3.39336
R2318 VDD.n1476 VDD.t225 3.39336
R2319 VDD.n1545 VDD.n1542 3.38874
R2320 VDD.n1220 VDD.n1219 3.38874
R2321 VDD.n1177 VDD.n1171 3.38874
R2322 VDD.n765 VDD.n762 3.38874
R2323 VDD.n440 VDD.n439 3.38874
R2324 VDD.n397 VDD.n391 3.38874
R2325 VDD.n1561 VDD.n1560 2.30978
R2326 VDD.n781 VDD.n780 2.30978
R2327 VDD.n549 VDD.n527 1.12991
R2328 VDD.n583 VDD.n493 1.12991
R2329 VDD.n608 VDD.n606 1.12991
R2330 VDD.n704 VDD.n473 1.12991
R2331 VDD.n667 VDD.n666 1.12991
R2332 VDD.n946 VDD.n924 1.12991
R2333 VDD.n980 VDD.n890 1.12991
R2334 VDD.n1003 VDD.n872 1.12991
R2335 VDD.n1073 VDD.n1072 1.12991
R2336 VDD.n1109 VDD.n1108 1.12991
R2337 VDD.n1329 VDD.n1307 1.12991
R2338 VDD.n1363 VDD.n1273 1.12991
R2339 VDD.n1388 VDD.n1386 1.12991
R2340 VDD.n1484 VDD.n1253 1.12991
R2341 VDD.n1447 VDD.n1446 1.12991
R2342 VDD.n118 VDD.n117 1.12991
R2343 VDD.n177 VDD.n176 1.12991
R2344 VDD.n246 VDD.n245 1.12991
R2345 VDD.n297 VDD.n296 1.12991
R2346 VDD.n342 VDD.n341 1.12991
R2347 VDD.n1591 VDD.n1166 0.826983
R2348 VDD.n1599 VDD.n386 0.826983
R2349 VDD.n1590 VDD.n1197 0.557954
R2350 VDD.n1598 VDD.n417 0.557954
R2351 VDD.n1226 VDD 0.476404
R2352 VDD.n446 VDD 0.476404
R2353 VDD VDD.n1226 0.403703
R2354 VDD VDD.n446 0.403703
R2355 VDD.n1587 VDD.n1538 0.399037
R2356 VDD.n1595 VDD.n758 0.399037
R2357 VDD.n534 VDD.n531 0.376971
R2358 VDD.n591 VDD.n590 0.376971
R2359 VDD.n727 VDD.n726 0.376971
R2360 VDD.n643 VDD.n477 0.376971
R2361 VDD.n931 VDD.n928 0.376971
R2362 VDD.n988 VDD.n987 0.376971
R2363 VDD.n1049 VDD.n874 0.376971
R2364 VDD.n1084 VDD.n1083 0.376971
R2365 VDD.n1314 VDD.n1311 0.376971
R2366 VDD.n1371 VDD.n1370 0.376971
R2367 VDD.n1507 VDD.n1506 0.376971
R2368 VDD.n1423 VDD.n1257 0.376971
R2369 VDD.n159 VDD.n158 0.376971
R2370 VDD.n215 VDD.n214 0.376971
R2371 VDD.n263 VDD.n262 0.376971
R2372 VDD.n319 VDD.n318 0.376971
R2373 VDD.n1589 VDD.n1232 0.35558
R2374 VDD.n1597 VDD.n452 0.35558
R2375 VDD.n1200 VDD 0.340206
R2376 VDD.n420 VDD 0.340206
R2377 VDD.n320 VDD 0.330819
R2378 VDD.n1596 VDD.n732 0.303619
R2379 VDD.n1588 VDD.n1512 0.303619
R2380 VDD.n1592 VDD.n1149 0.299064
R2381 VDD.n815 VDD.n814 0.240091
R2382 VDD.n9 VDD.n8 0.240091
R2383 VDD.n1586 VDD.n1585 0.212557
R2384 VDD.n1594 VDD.n805 0.212557
R2385 VDD.n1166 VDD.n1165 0.211096
R2386 VDD.n386 VDD.n385 0.211096
R2387 VDD.n1552 VDD 0.210222
R2388 VDD.n772 VDD 0.210222
R2389 VDD.n1227 VDD 0.196824
R2390 VDD.n447 VDD 0.196824
R2391 VDD.n1232 VDD.n1231 0.183651
R2392 VDD.n452 VDD.n451 0.183651
R2393 VDD.n1593 VDD.n869 0.180844
R2394 VDD.n361 VDD.n63 0.180844
R2395 VDD.n1585 VDD.n1584 0.175873
R2396 VDD.n805 VDD.n804 0.175873
R2397 VDD.n1600 VDD.n369 0.168948
R2398 VDD.n1197 VDD.n1196 0.155541
R2399 VDD.n417 VDD.n416 0.155541
R2400 VDD.n1228 VDD 0.145087
R2401 VDD.n448 VDD 0.145087
R2402 VDD VDD.n827 0.137071
R2403 VDD VDD.n21 0.137071
R2404 VDD.n863 VDD.n862 0.128415
R2405 VDD.n53 VDD.n52 0.12814
R2406 VDD.n1538 VDD.n1536 0.120987
R2407 VDD.n758 VDD.n756 0.120987
R2408 VDD.n864 VDD.n863 0.119283
R2409 VDD.n54 VDD.n53 0.11856
R2410 VDD.n859 VDD.n858 0.1155
R2411 VDD.n858 VDD.n857 0.1155
R2412 VDD.n854 VDD.n853 0.1155
R2413 VDD.n853 VDD.n852 0.1155
R2414 VDD.n849 VDD.n848 0.1155
R2415 VDD.n848 VDD.n847 0.1155
R2416 VDD.n844 VDD.n843 0.1155
R2417 VDD.n843 VDD.n842 0.1155
R2418 VDD.n49 VDD.n48 0.1155
R2419 VDD.n48 VDD.n46 0.1155
R2420 VDD.n43 VDD.n42 0.1155
R2421 VDD.n42 VDD.n40 0.1155
R2422 VDD.n37 VDD.n36 0.1155
R2423 VDD.n36 VDD.n34 0.1155
R2424 VDD.n31 VDD.n30 0.1155
R2425 VDD.n30 VDD.n28 0.1155
R2426 VDD.n869 VDD 0.109094
R2427 VDD.n63 VDD 0.109094
R2428 VDD.n869 VDD.n868 0.107922
R2429 VDD.n63 VDD.n62 0.107922
R2430 VDD.n864 VDD 0.0950313
R2431 VDD.n54 VDD 0.0950313
R2432 VDD.n514 VDD.n510 0.0892839
R2433 VDD.n911 VDD.n907 0.0892839
R2434 VDD.n1294 VDD.n1290 0.0892839
R2435 VDD.n68 VDD.n66 0.088354
R2436 VDD.n1226 VDD.n1225 0.0849867
R2437 VDD.n446 VDD.n445 0.0849867
R2438 VDD.n1231 VDD.n1198 0.0777407
R2439 VDD.n451 VDD.n418 0.0777407
R2440 VDD.n1584 VDD.n1539 0.0734782
R2441 VDD.n1196 VDD.n1168 0.0734782
R2442 VDD.n804 VDD.n759 0.0734782
R2443 VDD.n416 VDD.n388 0.0734782
R2444 VDD.n360 VDD.n73 0.0694387
R2445 VDD.n1533 VDD.n1515 0.0681471
R2446 VDD.n1533 VDD.n1517 0.0681471
R2447 VDD.n1520 VDD.n1517 0.0681471
R2448 VDD.n1528 VDD.n1520 0.0681471
R2449 VDD.n1528 VDD.n1523 0.0681471
R2450 VDD.n753 VDD.n735 0.0681471
R2451 VDD.n753 VDD.n737 0.0681471
R2452 VDD.n740 VDD.n737 0.0681471
R2453 VDD.n748 VDD.n740 0.0681471
R2454 VDD.n748 VDD.n743 0.0681471
R2455 VDD.n1165 VDD.n1150 0.0671334
R2456 VDD.n385 VDD.n370 0.0671334
R2457 VDD.n1222 VDD.n1221 0.065907
R2458 VDD.n1217 VDD.n1204 0.065907
R2459 VDD.n1216 VDD.n1215 0.065907
R2460 VDD.n1214 VDD.n1210 0.065907
R2461 VDD.n442 VDD.n441 0.065907
R2462 VDD.n437 VDD.n424 0.065907
R2463 VDD.n436 VDD.n435 0.065907
R2464 VDD.n434 VDD.n430 0.065907
R2465 VDD.n1562 VDD.n1553 0.0658409
R2466 VDD.n782 VDD.n773 0.0658409
R2467 VDD.n1580 VDD.n1539 0.0643889
R2468 VDD.n1580 VDD.n1579 0.0643889
R2469 VDD.n1579 VDD.n1578 0.0643889
R2470 VDD.n1575 VDD.n1574 0.0643889
R2471 VDD.n1574 VDD.n1573 0.0643889
R2472 VDD.n1573 VDD.n1543 0.0643889
R2473 VDD.n1567 VDD.n1548 0.0643889
R2474 VDD.n1192 VDD.n1168 0.0643889
R2475 VDD.n1192 VDD.n1191 0.0643889
R2476 VDD.n1191 VDD.n1190 0.0643889
R2477 VDD.n1183 VDD.n1172 0.0643889
R2478 VDD.n1183 VDD.n1175 0.0643889
R2479 VDD.n1179 VDD.n1175 0.0643889
R2480 VDD.n1162 VDD.n1161 0.0643889
R2481 VDD.n1161 VDD.n1160 0.0643889
R2482 VDD.n800 VDD.n759 0.0643889
R2483 VDD.n800 VDD.n799 0.0643889
R2484 VDD.n799 VDD.n798 0.0643889
R2485 VDD.n795 VDD.n794 0.0643889
R2486 VDD.n794 VDD.n793 0.0643889
R2487 VDD.n793 VDD.n763 0.0643889
R2488 VDD.n787 VDD.n768 0.0643889
R2489 VDD.n412 VDD.n388 0.0643889
R2490 VDD.n412 VDD.n411 0.0643889
R2491 VDD.n411 VDD.n410 0.0643889
R2492 VDD.n403 VDD.n392 0.0643889
R2493 VDD.n403 VDD.n395 0.0643889
R2494 VDD.n399 VDD.n395 0.0643889
R2495 VDD.n382 VDD.n381 0.0643889
R2496 VDD.n381 VDD.n380 0.0643889
R2497 VDD.n235 VDD 0.0639804
R2498 VDD.n1536 VDD.n1513 0.0599867
R2499 VDD.n756 VDD.n733 0.0599867
R2500 VDD.n1159 VDD.n1158 0.0587674
R2501 VDD.n379 VDD.n378 0.0587674
R2502 VDD.n1187 VDD.n1186 0.0580441
R2503 VDD.n407 VDD.n406 0.0580441
R2504 VDD.n859 VDD 0.058
R2505 VDD.n854 VDD 0.058
R2506 VDD.n844 VDD 0.058
R2507 VDD.n49 VDD 0.058
R2508 VDD.n43 VDD 0.058
R2509 VDD.n31 VDD 0.058
R2510 VDD.n1547 VDD.n1543 0.0567153
R2511 VDD.n767 VDD.n763 0.0567153
R2512 VDD.n849 VDD 0.0555
R2513 VDD.n37 VDD 0.0555
R2514 VDD.n1553 VDD.n1552 0.0516364
R2515 VDD.n773 VDD.n772 0.0516364
R2516 VDD.n1225 VDD.n1200 0.0418891
R2517 VDD.n445 VDD.n420 0.0418891
R2518 VDD.n1227 VDD.n1198 0.0409412
R2519 VDD.n447 VDD.n418 0.0409412
R2520 VDD.n1594 VDD.n1593 0.0407258
R2521 VDD.n827 VDD.n806 0.03976
R2522 VDD.n21 VDD.n0 0.03976
R2523 VDD.n865 VDD.n864 0.0376094
R2524 VDD.n55 VDD.n54 0.0376094
R2525 VDD.n1228 VDD.n1227 0.0371297
R2526 VDD.n448 VDD.n447 0.0371297
R2527 VDD VDD.n1601 0.0351129
R2528 VDD.n1203 VDD.n1200 0.0339302
R2529 VDD.n423 VDD.n420 0.0339302
R2530 VDD.n817 VDD.n809 0.033737
R2531 VDD.n821 VDD.n809 0.033737
R2532 VDD.n822 VDD.n821 0.033737
R2533 VDD.n823 VDD.n822 0.033737
R2534 VDD.n11 VDD.n3 0.033737
R2535 VDD.n15 VDD.n3 0.033737
R2536 VDD.n16 VDD.n15 0.033737
R2537 VDD.n17 VDD.n16 0.033737
R2538 VDD.n1562 VDD.n1561 0.0334425
R2539 VDD.n1561 VDD.n1555 0.0334425
R2540 VDD.n782 VDD.n781 0.0334425
R2541 VDD.n781 VDD.n775 0.0334425
R2542 VDD.n369 VDD.n362 0.0333707
R2543 VDD.n1575 VDD 0.0324444
R2544 VDD VDD.n1567 0.0324444
R2545 VDD.n1187 VDD 0.0324444
R2546 VDD.n795 VDD 0.0324444
R2547 VDD VDD.n787 0.0324444
R2548 VDD.n407 VDD 0.0324444
R2549 VDD.n1598 VDD.n1597 0.0299677
R2550 VDD.n1595 VDD.n1594 0.0299677
R2551 VDD.n1590 VDD.n1589 0.0299677
R2552 VDD.n1587 VDD.n1586 0.0299677
R2553 VDD.n1599 VDD.n1598 0.0292661
R2554 VDD.n1591 VDD.n1590 0.0292661
R2555 VDD.n1588 VDD.n1587 0.0286815
R2556 VDD.n683 VDD 0.0279106
R2557 VDD.n1125 VDD 0.0279106
R2558 VDD.n1463 VDD 0.0279106
R2559 VDD.n344 VDD 0.0260435
R2560 VDD.n336 VDD.n335 0.0254026
R2561 VDD.n343 VDD.n339 0.0249681
R2562 VDD.n339 VDD.n337 0.0249681
R2563 VDD.n216 VDD.n212 0.0249681
R2564 VDD.n212 VDD.n210 0.0249681
R2565 VDD.n210 VDD.n206 0.0249681
R2566 VDD.n206 VDD.n204 0.0249681
R2567 VDD.n204 VDD.n200 0.0249681
R2568 VDD.n200 VDD.n196 0.0249681
R2569 VDD.n186 VDD.n184 0.0249681
R2570 VDD.n184 VDD.n180 0.0249681
R2571 VDD.n180 VDD.n178 0.0249681
R2572 VDD.n178 VDD.n174 0.0249681
R2573 VDD.n174 VDD.n172 0.0249681
R2574 VDD.n160 VDD.n156 0.0249681
R2575 VDD.n156 VDD.n154 0.0249681
R2576 VDD.n154 VDD.n150 0.0249681
R2577 VDD.n150 VDD.n148 0.0249681
R2578 VDD.n131 VDD.n127 0.0249681
R2579 VDD.n127 VDD.n125 0.0249681
R2580 VDD.n125 VDD.n121 0.0249681
R2581 VDD.n121 VDD.n119 0.0249681
R2582 VDD.n89 VDD.n87 0.0249681
R2583 VDD.n92 VDD.n89 0.0249681
R2584 VDD.n94 VDD.n92 0.0249681
R2585 VDD.n96 VDD.n94 0.0249681
R2586 VDD.n103 VDD.n101 0.0249681
R2587 VDD.n241 VDD.n237 0.0249681
R2588 VDD.n243 VDD.n241 0.0249681
R2589 VDD.n247 VDD.n243 0.0249681
R2590 VDD.n249 VDD.n247 0.0249681
R2591 VDD.n264 VDD.n260 0.0249681
R2592 VDD.n266 VDD.n264 0.0249681
R2593 VDD.n270 VDD.n266 0.0249681
R2594 VDD.n272 VDD.n270 0.0249681
R2595 VDD.n276 VDD.n272 0.0249681
R2596 VDD.n280 VDD.n276 0.0249681
R2597 VDD.n282 VDD.n280 0.0249681
R2598 VDD.n286 VDD.n282 0.0249681
R2599 VDD.n288 VDD.n286 0.0249681
R2600 VDD.n292 VDD.n288 0.0249681
R2601 VDD.n294 VDD.n292 0.0249681
R2602 VDD.n298 VDD.n294 0.0249681
R2603 VDD.n300 VDD.n298 0.0249681
R2604 VDD.n323 VDD.n322 0.0249681
R2605 VDD.n322 VDD.n320 0.0249681
R2606 VDD.n1592 VDD 0.0245887
R2607 VDD.n367 VDD.n366 0.0243281
R2608 VDD.n332 VDD.n216 0.0241145
R2609 VDD.n1596 VDD.n1595 0.0228347
R2610 VDD.n112 VDD.n84 0.0218724
R2611 VDD.n862 VDD 0.02175
R2612 VDD.n857 VDD 0.02175
R2613 VDD.n852 VDD 0.02175
R2614 VDD.n847 VDD 0.02175
R2615 VDD.n842 VDD 0.02175
R2616 VDD.n52 VDD 0.02175
R2617 VDD.n46 VDD 0.02175
R2618 VDD.n40 VDD 0.02175
R2619 VDD.n34 VDD 0.02175
R2620 VDD.n28 VDD 0.02175
R2621 VDD.n1601 VDD 0.0213145
R2622 VDD.n148 VDD.n144 0.0212447
R2623 VDD.n260 VDD.n258 0.0207128
R2624 VDD.n196 VDD.n194 0.0198592
R2625 VDD.n303 VDD.n301 0.0188511
R2626 VDD.n106 VDD.n104 0.0172553
R2627 VDD.n817 VDD 0.0171185
R2628 VDD VDD.n806 0.0171185
R2629 VDD.n11 VDD 0.0171185
R2630 VDD VDD.n0 0.0171185
R2631 VDD.n868 VDD.n867 0.0165987
R2632 VDD.n62 VDD.n61 0.0165987
R2633 VDD.n161 VDD.n160 0.0161915
R2634 VDD.n865 VDD.n829 0.016125
R2635 VDD.n56 VDD.n55 0.016125
R2636 VDD.n143 VDD.n139 0.0153936
R2637 VDD.n250 VDD.n249 0.0151277
R2638 VDD.n191 VDD.n187 0.0148617
R2639 VDD.n684 VDD.n683 0.0146339
R2640 VDD.n1126 VDD.n1125 0.0146339
R2641 VDD.n1464 VDD.n1463 0.0146339
R2642 VDD.n132 VDD.n131 0.0145957
R2643 VDD.n115 VDD.n114 0.0145957
R2644 VDD.n1552 VDD.n1548 0.0143889
R2645 VDD.n772 VDD.n768 0.0143889
R2646 VDD.n344 VDD.n343 0.0143298
R2647 VDD.n170 VDD.n169 0.0137979
R2648 VDD.n1523 VDD 0.013
R2649 VDD.n743 VDD 0.013
R2650 VDD VDD.n336 0.012734
R2651 VDD.n87 VDD 0.012734
R2652 VDD VDD.n218 0.012734
R2653 VDD.n366 VDD.n364 0.0126094
R2654 VDD.n515 VDD.n514 0.0126053
R2655 VDD.n562 VDD.n506 0.0126053
R2656 VDD.n557 VDD.n506 0.0126053
R2657 VDD.n557 VDD.n556 0.0126053
R2658 VDD.n556 VDD.n524 0.0126053
R2659 VDD.n551 VDD.n524 0.0126053
R2660 VDD.n551 VDD.n550 0.0126053
R2661 VDD.n550 VDD.n528 0.0126053
R2662 VDD.n529 VDD.n528 0.0126053
R2663 VDD.n544 VDD.n530 0.0126053
R2664 VDD.n544 VDD.n543 0.0126053
R2665 VDD.n543 VDD.n542 0.0126053
R2666 VDD.n542 VDD.n532 0.0126053
R2667 VDD.n570 VDD.n569 0.0126053
R2668 VDD.n570 VDD.n498 0.0126053
R2669 VDD.n575 VDD.n498 0.0126053
R2670 VDD.n576 VDD.n575 0.0126053
R2671 VDD.n576 VDD.n494 0.0126053
R2672 VDD.n581 VDD.n494 0.0126053
R2673 VDD.n582 VDD.n581 0.0126053
R2674 VDD.n582 VDD.n491 0.0126053
R2675 VDD.n586 VDD.n491 0.0126053
R2676 VDD.n588 VDD.n587 0.0126053
R2677 VDD.n588 VDD.n488 0.0126053
R2678 VDD.n593 VDD.n488 0.0126053
R2679 VDD.n594 VDD.n593 0.0126053
R2680 VDD.n621 VDD.n484 0.0126053
R2681 VDD.n616 VDD.n484 0.0126053
R2682 VDD.n616 VDD.n615 0.0126053
R2683 VDD.n615 VDD.n603 0.0126053
R2684 VDD.n610 VDD.n603 0.0126053
R2685 VDD.n610 VDD.n609 0.0126053
R2686 VDD.n609 VDD.n453 0.0126053
R2687 VDD.n730 VDD.n729 0.0126053
R2688 VDD.n729 VDD.n456 0.0126053
R2689 VDD.n719 VDD.n718 0.0126053
R2690 VDD.n718 VDD.n465 0.0126053
R2691 VDD.n713 VDD.n465 0.0126053
R2692 VDD.n713 VDD.n712 0.0126053
R2693 VDD.n712 VDD.n711 0.0126053
R2694 VDD.n711 VDD.n468 0.0126053
R2695 VDD.n706 VDD.n468 0.0126053
R2696 VDD.n706 VDD.n705 0.0126053
R2697 VDD.n705 VDD.n474 0.0126053
R2698 VDD.n475 VDD.n474 0.0126053
R2699 VDD.n699 VDD.n476 0.0126053
R2700 VDD.n649 VDD.n648 0.0126053
R2701 VDD.n649 VDD.n639 0.0126053
R2702 VDD.n656 VDD.n639 0.0126053
R2703 VDD.n657 VDD.n656 0.0126053
R2704 VDD.n658 VDD.n657 0.0126053
R2705 VDD.n658 VDD.n636 0.0126053
R2706 VDD.n663 VDD.n636 0.0126053
R2707 VDD.n664 VDD.n663 0.0126053
R2708 VDD.n664 VDD.n632 0.0126053
R2709 VDD.n669 VDD.n632 0.0126053
R2710 VDD.n670 VDD.n669 0.0126053
R2711 VDD.n671 VDD.n629 0.0126053
R2712 VDD.n675 VDD.n629 0.0126053
R2713 VDD.n676 VDD.n675 0.0126053
R2714 VDD.n677 VDD.n676 0.0126053
R2715 VDD.n689 VDD.n688 0.0126053
R2716 VDD.n685 VDD.n684 0.0126053
R2717 VDD.n912 VDD.n911 0.0126053
R2718 VDD.n959 VDD.n903 0.0126053
R2719 VDD.n954 VDD.n903 0.0126053
R2720 VDD.n954 VDD.n953 0.0126053
R2721 VDD.n953 VDD.n921 0.0126053
R2722 VDD.n948 VDD.n921 0.0126053
R2723 VDD.n948 VDD.n947 0.0126053
R2724 VDD.n947 VDD.n925 0.0126053
R2725 VDD.n926 VDD.n925 0.0126053
R2726 VDD.n941 VDD.n927 0.0126053
R2727 VDD.n941 VDD.n940 0.0126053
R2728 VDD.n940 VDD.n939 0.0126053
R2729 VDD.n939 VDD.n929 0.0126053
R2730 VDD.n967 VDD.n966 0.0126053
R2731 VDD.n967 VDD.n895 0.0126053
R2732 VDD.n972 VDD.n895 0.0126053
R2733 VDD.n973 VDD.n972 0.0126053
R2734 VDD.n973 VDD.n891 0.0126053
R2735 VDD.n978 VDD.n891 0.0126053
R2736 VDD.n979 VDD.n978 0.0126053
R2737 VDD.n979 VDD.n888 0.0126053
R2738 VDD.n983 VDD.n888 0.0126053
R2739 VDD.n985 VDD.n984 0.0126053
R2740 VDD.n985 VDD.n885 0.0126053
R2741 VDD.n990 VDD.n885 0.0126053
R2742 VDD.n991 VDD.n990 0.0126053
R2743 VDD.n1015 VDD.n881 0.0126053
R2744 VDD.n1010 VDD.n881 0.0126053
R2745 VDD.n1010 VDD.n1009 0.0126053
R2746 VDD.n1009 VDD.n1000 0.0126053
R2747 VDD.n1004 VDD.n1000 0.0126053
R2748 VDD.n1004 VDD.n870 0.0126053
R2749 VDD.n1148 VDD.n871 0.0126053
R2750 VDD.n1143 VDD.n873 0.0126053
R2751 VDD.n1143 VDD.n1142 0.0126053
R2752 VDD.n1058 VDD.n1057 0.0126053
R2753 VDD.n1059 VDD.n1058 0.0126053
R2754 VDD.n1059 VDD.n1044 0.0126053
R2755 VDD.n1066 VDD.n1044 0.0126053
R2756 VDD.n1067 VDD.n1066 0.0126053
R2757 VDD.n1068 VDD.n1067 0.0126053
R2758 VDD.n1068 VDD.n1040 0.0126053
R2759 VDD.n1074 VDD.n1040 0.0126053
R2760 VDD.n1075 VDD.n1074 0.0126053
R2761 VDD.n1076 VDD.n1075 0.0126053
R2762 VDD.n1080 VDD.n1079 0.0126053
R2763 VDD.n1091 VDD.n1090 0.0126053
R2764 VDD.n1091 VDD.n1033 0.0126053
R2765 VDD.n1098 VDD.n1033 0.0126053
R2766 VDD.n1099 VDD.n1098 0.0126053
R2767 VDD.n1100 VDD.n1099 0.0126053
R2768 VDD.n1100 VDD.n1030 0.0126053
R2769 VDD.n1105 VDD.n1030 0.0126053
R2770 VDD.n1106 VDD.n1105 0.0126053
R2771 VDD.n1106 VDD.n1026 0.0126053
R2772 VDD.n1111 VDD.n1026 0.0126053
R2773 VDD.n1112 VDD.n1111 0.0126053
R2774 VDD.n1113 VDD.n1023 0.0126053
R2775 VDD.n1117 VDD.n1023 0.0126053
R2776 VDD.n1118 VDD.n1117 0.0126053
R2777 VDD.n1119 VDD.n1118 0.0126053
R2778 VDD.n1131 VDD.n1130 0.0126053
R2779 VDD.n1127 VDD.n1126 0.0126053
R2780 VDD.n1295 VDD.n1294 0.0126053
R2781 VDD.n1342 VDD.n1286 0.0126053
R2782 VDD.n1337 VDD.n1286 0.0126053
R2783 VDD.n1337 VDD.n1336 0.0126053
R2784 VDD.n1336 VDD.n1304 0.0126053
R2785 VDD.n1331 VDD.n1304 0.0126053
R2786 VDD.n1331 VDD.n1330 0.0126053
R2787 VDD.n1330 VDD.n1308 0.0126053
R2788 VDD.n1309 VDD.n1308 0.0126053
R2789 VDD.n1324 VDD.n1310 0.0126053
R2790 VDD.n1324 VDD.n1323 0.0126053
R2791 VDD.n1323 VDD.n1322 0.0126053
R2792 VDD.n1322 VDD.n1312 0.0126053
R2793 VDD.n1350 VDD.n1349 0.0126053
R2794 VDD.n1350 VDD.n1278 0.0126053
R2795 VDD.n1355 VDD.n1278 0.0126053
R2796 VDD.n1356 VDD.n1355 0.0126053
R2797 VDD.n1356 VDD.n1274 0.0126053
R2798 VDD.n1361 VDD.n1274 0.0126053
R2799 VDD.n1362 VDD.n1361 0.0126053
R2800 VDD.n1362 VDD.n1271 0.0126053
R2801 VDD.n1366 VDD.n1271 0.0126053
R2802 VDD.n1368 VDD.n1367 0.0126053
R2803 VDD.n1368 VDD.n1268 0.0126053
R2804 VDD.n1373 VDD.n1268 0.0126053
R2805 VDD.n1374 VDD.n1373 0.0126053
R2806 VDD.n1401 VDD.n1264 0.0126053
R2807 VDD.n1396 VDD.n1264 0.0126053
R2808 VDD.n1396 VDD.n1395 0.0126053
R2809 VDD.n1395 VDD.n1383 0.0126053
R2810 VDD.n1390 VDD.n1383 0.0126053
R2811 VDD.n1390 VDD.n1389 0.0126053
R2812 VDD.n1389 VDD.n1233 0.0126053
R2813 VDD.n1510 VDD.n1509 0.0126053
R2814 VDD.n1509 VDD.n1236 0.0126053
R2815 VDD.n1499 VDD.n1498 0.0126053
R2816 VDD.n1498 VDD.n1245 0.0126053
R2817 VDD.n1493 VDD.n1245 0.0126053
R2818 VDD.n1493 VDD.n1492 0.0126053
R2819 VDD.n1492 VDD.n1491 0.0126053
R2820 VDD.n1491 VDD.n1248 0.0126053
R2821 VDD.n1486 VDD.n1248 0.0126053
R2822 VDD.n1486 VDD.n1485 0.0126053
R2823 VDD.n1485 VDD.n1254 0.0126053
R2824 VDD.n1255 VDD.n1254 0.0126053
R2825 VDD.n1479 VDD.n1256 0.0126053
R2826 VDD.n1429 VDD.n1428 0.0126053
R2827 VDD.n1429 VDD.n1419 0.0126053
R2828 VDD.n1436 VDD.n1419 0.0126053
R2829 VDD.n1437 VDD.n1436 0.0126053
R2830 VDD.n1438 VDD.n1437 0.0126053
R2831 VDD.n1438 VDD.n1416 0.0126053
R2832 VDD.n1443 VDD.n1416 0.0126053
R2833 VDD.n1444 VDD.n1443 0.0126053
R2834 VDD.n1444 VDD.n1412 0.0126053
R2835 VDD.n1449 VDD.n1412 0.0126053
R2836 VDD.n1450 VDD.n1449 0.0126053
R2837 VDD.n1451 VDD.n1409 0.0126053
R2838 VDD.n1455 VDD.n1409 0.0126053
R2839 VDD.n1456 VDD.n1455 0.0126053
R2840 VDD.n1457 VDD.n1456 0.0126053
R2841 VDD.n1469 VDD.n1468 0.0126053
R2842 VDD.n1465 VDD.n1464 0.0126053
R2843 VDD.n1555 VDD 0.0125739
R2844 VDD.n775 VDD 0.0125739
R2845 VDD.n732 VDD.n731 0.0124737
R2846 VDD.n1512 VDD.n1511 0.0124737
R2847 VDD.n1568 VDD 0.0123056
R2848 VDD.n1179 VDD 0.0123056
R2849 VDD.n788 VDD 0.0123056
R2850 VDD.n399 VDD 0.0123056
R2851 VDD.n1149 VDD.n870 0.0122105
R2852 VDD.n532 VDD.n502 0.0119152
R2853 VDD.n1312 VDD.n1282 0.0119152
R2854 VDD.n72 VDD.n68 0.0117745
R2855 VDD.n224 VDD.n220 0.0117745
R2856 VDD.n228 VDD.n224 0.0117745
R2857 VDD.n230 VDD.n228 0.0117745
R2858 VDD.n234 VDD.n230 0.0117745
R2859 VDD.n1578 VDD 0.0116111
R2860 VDD.n1190 VDD 0.0116111
R2861 VDD.n1158 VDD 0.0116111
R2862 VDD.n798 VDD 0.0116111
R2863 VDD.n410 VDD 0.0116111
R2864 VDD.n378 VDD 0.0116111
R2865 VDD.n1211 VDD 0.0114012
R2866 VDD.n431 VDD 0.0114012
R2867 VDD.n929 VDD.n899 0.0113889
R2868 VDD.n1016 VDD.n1015 0.0108947
R2869 VDD.n134 VDD.n132 0.0108723
R2870 VDD.n119 VDD.n115 0.0108723
R2871 VDD.n1057 VDD.n877 0.0106316
R2872 VDD.n1090 VDD.n1089 0.0106316
R2873 VDD.n187 VDD.n186 0.0106064
R2874 VDD.n515 VDD.n503 0.0103684
R2875 VDD.n622 VDD.n621 0.0103684
R2876 VDD.n1295 VDD.n1283 0.0103684
R2877 VDD.n1402 VDD.n1401 0.0103684
R2878 VDD.n167 VDD.n163 0.0103404
R2879 VDD.n252 VDD.n250 0.0103404
R2880 VDD.n235 VDD.n234 0.0103039
R2881 VDD.n719 VDD.n462 0.0101053
R2882 VDD.n648 VDD.n480 0.0101053
R2883 VDD.n1499 VDD.n1242 0.0101053
R2884 VDD.n1428 VDD.n1260 0.0101053
R2885 VDD.n912 VDD.n900 0.00984211
R2886 VDD.n99 VDD 0.00954255
R2887 VDD.n1515 VDD.n1513 0.0095362
R2888 VDD.n735 VDD.n733 0.0095362
R2889 VDD.n163 VDD.n161 0.0092766
R2890 VDD.n1568 VDD.n1547 0.00906279
R2891 VDD.n788 VDD.n767 0.00906279
R2892 VDD.n960 VDD.n959 0.00905263
R2893 VDD.n320 VDD.n316 0.00883333
R2894 VDD.n316 VDD.n314 0.00883333
R2895 VDD.n314 VDD.n310 0.00883333
R2896 VDD.n310 VDD.n308 0.00883333
R2897 VDD.n308 VDD.n77 0.00883333
R2898 VDD.n357 VDD.n355 0.00883333
R2899 VDD.n355 VDD.n351 0.00883333
R2900 VDD.n351 VDD.n349 0.00883333
R2901 VDD.n349 VDD.n345 0.00883333
R2902 VDD.n460 VDD.n456 0.00878947
R2903 VDD.n699 VDD.n698 0.00878947
R2904 VDD.n692 VDD.n627 0.00878947
R2905 VDD.n1240 VDD.n1236 0.00878947
R2906 VDD.n1479 VDD.n1478 0.00878947
R2907 VDD.n1472 VDD.n1407 0.00878947
R2908 VDD.n137 VDD.n134 0.00874468
R2909 VDD.n563 VDD.n562 0.00852632
R2910 VDD.n568 VDD.n501 0.00852632
R2911 VDD.n594 VDD.n481 0.00852632
R2912 VDD.n1343 VDD.n1342 0.00852632
R2913 VDD.n1348 VDD.n1281 0.00852632
R2914 VDD.n1374 VDD.n1261 0.00852632
R2915 VDD.n324 VDD 0.00847872
R2916 VDD.n1142 VDD.n1141 0.00826316
R2917 VDD.n1081 VDD.n1080 0.00826316
R2918 VDD.n1134 VDD.n1021 0.00826316
R2919 VDD.n104 VDD.n103 0.00821277
R2920 VDD.n1160 VDD.n1159 0.00802802
R2921 VDD.n380 VDD.n379 0.00802802
R2922 VDD.n965 VDD.n898 0.008
R2923 VDD.n991 VDD.n878 0.008
R2924 VDD.n880 VDD.n879 0.008
R2925 VDD.n1186 VDD.n1172 0.00775202
R2926 VDD.n1162 VDD.n1150 0.00775202
R2927 VDD.n406 VDD.n392 0.00775202
R2928 VDD.n382 VDD.n370 0.00775202
R2929 VDD.n1052 VDD.n876 0.00773684
R2930 VDD.n1088 VDD.n1036 0.00773684
R2931 VDD.n517 VDD.n504 0.00747368
R2932 VDD.n483 VDD.n482 0.00747368
R2933 VDD.n1297 VDD.n1284 0.00747368
R2934 VDD.n1263 VDD.n1262 0.00747368
R2935 VDD VDD.n171 0.00741489
R2936 VDD.n723 VDD.n722 0.00721053
R2937 VDD.n644 VDD.n479 0.00721053
R2938 VDD.n1503 VDD.n1502 0.00721053
R2939 VDD.n1424 VDD.n1259 0.00721053
R2940 VDD.n364 VDD 0.00714063
R2941 VDD.n358 VDD.n357 0.00702174
R2942 VDD.n823 VDD 0.00700289
R2943 VDD.n17 VDD 0.00700289
R2944 VDD.n914 VDD.n901 0.00694737
R2945 VDD.n816 VDD 0.00675
R2946 VDD.n10 VDD 0.00675
R2947 VDD.n1597 VDD.n1596 0.00669758
R2948 VDD.n73 VDD.n72 0.00662745
R2949 VDD.n301 VDD.n300 0.00661702
R2950 VDD.n530 VDD 0.00655263
R2951 VDD.n587 VDD 0.00655263
R2952 VDD VDD.n730 0.00655263
R2953 VDD.n476 VDD 0.00655263
R2954 VDD.n671 VDD 0.00655263
R2955 VDD.n685 VDD 0.00655263
R2956 VDD.n927 VDD 0.00655263
R2957 VDD.n984 VDD 0.00655263
R2958 VDD.n873 VDD 0.00655263
R2959 VDD.n1079 VDD 0.00655263
R2960 VDD.n1113 VDD 0.00655263
R2961 VDD.n1127 VDD 0.00655263
R2962 VDD.n1310 VDD 0.00655263
R2963 VDD.n1367 VDD 0.00655263
R2964 VDD VDD.n1510 0.00655263
R2965 VDD.n1256 VDD 0.00655263
R2966 VDD.n1451 VDD 0.00655263
R2967 VDD.n1465 VDD 0.00655263
R2968 VDD.n902 VDD.n901 0.00615789
R2969 VDD VDD.n815 0.00609211
R2970 VDD VDD.n9 0.00609211
R2971 VDD.n724 VDD.n723 0.00589474
R2972 VDD.n479 VDD.n478 0.00589474
R2973 VDD.n1504 VDD.n1503 0.00589474
R2974 VDD.n1259 VDD.n1258 0.00589474
R2975 VDD.n171 VDD.n170 0.00581915
R2976 VDD.n220 VDD.n73 0.00564706
R2977 VDD.n505 VDD.n504 0.00563158
R2978 VDD.n596 VDD.n482 0.00563158
R2979 VDD.n693 VDD 0.00563158
R2980 VDD.n1285 VDD.n1284 0.00563158
R2981 VDD.n1376 VDD.n1262 0.00563158
R2982 VDD.n1473 VDD 0.00563158
R2983 VDD.n114 VDD.n112 0.00552129
R2984 VDD.n876 VDD.n875 0.00536842
R2985 VDD.n1082 VDD.n1036 0.00536842
R2986 VDD.n1593 VDD.n1592 0.00517742
R2987 VDD.n966 VDD.n965 0.00510526
R2988 VDD.n993 VDD.n878 0.00510526
R2989 VDD.n993 VDD.n879 0.00510526
R2990 VDD.n1135 VDD 0.00510526
R2991 VDD.n337 VDD 0.00502128
R2992 VDD.n172 VDD 0.00502128
R2993 VDD VDD.n84 0.00502128
R2994 VDD.n101 VDD 0.00502128
R2995 VDD VDD.n252 0.00502128
R2996 VDD.n1141 VDD.n875 0.00484211
R2997 VDD.n1082 VDD.n1081 0.00484211
R2998 VDD.n1131 VDD.n1021 0.00484211
R2999 VDD.n193 VDD.n191 0.00475532
R3000 VDD.n255 VDD 0.00475532
R3001 VDD.n258 VDD.n218 0.00475532
R3002 VDD.n324 VDD.n323 0.00475532
R3003 VDD.n563 VDD.n505 0.00457895
R3004 VDD.n569 VDD.n568 0.00457895
R3005 VDD.n596 VDD.n481 0.00457895
R3006 VDD.n1343 VDD.n1285 0.00457895
R3007 VDD.n1349 VDD.n1348 0.00457895
R3008 VDD.n1376 VDD.n1261 0.00457895
R3009 VDD.n1601 VDD 0.00455181
R3010 VDD.n367 VDD.n362 0.00451563
R3011 VDD.n724 VDD.n460 0.00431579
R3012 VDD.n698 VDD.n478 0.00431579
R3013 VDD.n689 VDD.n627 0.00431579
R3014 VDD.n1504 VDD.n1240 0.00431579
R3015 VDD.n1478 VDD.n1258 0.00431579
R3016 VDD.n1469 VDD.n1407 0.00431579
R3017 VDD.n144 VDD.n143 0.0042234
R3018 VDD.n345 VDD.n344 0.00412319
R3019 VDD VDD.n816 0.00411272
R3020 VDD VDD.n10 0.00411272
R3021 VDD.n960 VDD.n902 0.00405263
R3022 VDD.n1586 VDD 0.00400806
R3023 VDD.n816 VDD 0.00378947
R3024 VDD.n10 VDD 0.00378947
R3025 VDD.n237 VDD.n235 0.00369149
R3026 VDD.n326 VDD 0.00342553
R3027 VDD VDD.n1591 0.00330645
R3028 VDD.n914 VDD.n900 0.00326316
R3029 VDD.n97 VDD.n96 0.00315957
R3030 VDD.n722 VDD.n462 0.003
R3031 VDD.n644 VDD.n480 0.003
R3032 VDD.n1502 VDD.n1242 0.003
R3033 VDD.n1424 VDD.n1260 0.003
R3034 VDD.n517 VDD.n503 0.00273684
R3035 VDD VDD.n529 0.00273684
R3036 VDD VDD.n586 0.00273684
R3037 VDD.n622 VDD.n483 0.00273684
R3038 VDD.n731 VDD 0.00273684
R3039 VDD VDD.n475 0.00273684
R3040 VDD VDD.n670 0.00273684
R3041 VDD.n688 VDD 0.00273684
R3042 VDD VDD.n926 0.00273684
R3043 VDD VDD.n983 0.00273684
R3044 VDD VDD.n871 0.00273684
R3045 VDD.n1076 VDD 0.00273684
R3046 VDD VDD.n1112 0.00273684
R3047 VDD.n1130 VDD 0.00273684
R3048 VDD.n1297 VDD.n1283 0.00273684
R3049 VDD VDD.n1309 0.00273684
R3050 VDD VDD.n1366 0.00273684
R3051 VDD.n1402 VDD.n1263 0.00273684
R3052 VDD.n1511 VDD 0.00273684
R3053 VDD VDD.n1255 0.00273684
R3054 VDD VDD.n1450 0.00273684
R3055 VDD.n1468 VDD 0.00273684
R3056 VDD.n899 VDD.n898 0.00271053
R3057 VDD.n359 VDD 0.00270801
R3058 VDD.n256 VDD 0.00262766
R3059 VDD.n830 VDD.n828 0.00257829
R3060 VDD.n677 VDD.n626 0.00247368
R3061 VDD.n1052 VDD.n877 0.00247368
R3062 VDD.n1089 VDD.n1088 0.00247368
R3063 VDD.n1457 VDD.n1406 0.00247368
R3064 VDD.n360 VDD.n359 0.00243485
R3065 VDD.n97 VDD 0.0023617
R3066 VDD.n107 VDD.n106 0.0023617
R3067 VDD.n334 VDD.n332 0.00232979
R3068 VDD.n194 VDD.n193 0.00232979
R3069 VDD.n358 VDD.n77 0.00231159
R3070 VDD.n1016 VDD.n880 0.00221053
R3071 VDD.n502 VDD.n501 0.00218421
R3072 VDD.n1282 VDD.n1281 0.00218421
R3073 VDD.n1601 VDD.n361 0.00204788
R3074 VDD VDD.n1600 0.00202016
R3075 VDD.n1222 VDD.n1203 0.00195349
R3076 VDD.n1221 VDD.n1204 0.00195349
R3077 VDD.n1217 VDD.n1216 0.00195349
R3078 VDD.n1215 VDD.n1214 0.00195349
R3079 VDD.n1211 VDD.n1210 0.00195349
R3080 VDD.n442 VDD.n423 0.00195349
R3081 VDD.n441 VDD.n424 0.00195349
R3082 VDD.n437 VDD.n436 0.00195349
R3083 VDD.n435 VDD.n434 0.00195349
R3084 VDD.n431 VDD.n430 0.00195349
R3085 VDD.n1119 VDD.n1020 0.00194737
R3086 VDD.n1135 VDD.n1134 0.00194737
R3087 VDD.n169 VDD.n167 0.00182979
R3088 VDD.n139 VDD.n137 0.00182979
R3089 VDD.n107 VDD.n99 0.00182979
R3090 VDD.n256 VDD.n255 0.00182979
R3091 VDD.n327 VDD.n326 0.00182979
R3092 VDD.n1600 VDD.n1599 0.00178629
R3093 VDD.n361 VDD.n360 0.0015471
R3094 VDD.n693 VDD.n692 0.00142105
R3095 VDD.n1473 VDD.n1472 0.00142105
R3096 VDD VDD.n1020 0.00128947
R3097 VDD.n830 VDD.n829 0.00116652
R3098 VDD.n56 VDD.n22 0.00116652
R3099 VDD.n866 VDD.n832 0.00114708
R3100 VDD.n832 VDD.n828 0.00114708
R3101 VDD.n60 VDD.n59 0.00114708
R3102 VDD.n59 VDD.n57 0.00114708
R3103 VDD.n867 VDD.n866 0.00107711
R3104 VDD.n61 VDD.n60 0.00107711
R3105 VDD.n332 VDD.n331 0.00100344
R3106 VDD.n194 VDD.n81 0.00100344
R3107 VDD.n112 VDD.n111 0.00100342
R3108 VDD.n1538 VDD.n1537 0.00100258
R3109 VDD.n758 VDD.n757 0.00100258
R3110 VDD.n567 VDD.n502 0.00100097
R3111 VDD.n964 VDD.n899 0.00100097
R3112 VDD.n1347 VDD.n1282 0.00100097
R3113 VDD.n365 VDD.n362 0.00100097
R3114 VDD.n867 VDD.n829 0.00100013
R3115 VDD.n61 VDD.n56 0.00100013
R3116 VDD.n335 VDD.n334 0.001
R3117 VDD.n832 VDD.n831 0.001
R3118 VDD.n59 VDD.n58 0.001
R3119 VDD.n1149 VDD.n1148 0.000894737
R3120 VDD.n1589 VDD.n1588 0.000850806
R3121 VDD.n327 VDD.n303 0.000765957
R3122 VDD VDD.n626 0.000763158
R3123 VDD VDD.n1406 0.000763158
R3124 VDD.n732 VDD.n453 0.000631579
R3125 VDD.n1512 VDD.n1233 0.000631579
R3126 VDD.n697 VDD.n696 0.000506553
R3127 VDD.n625 VDD.n461 0.000506553
R3128 VDD.n624 VDD.n623 0.000506553
R3129 VDD.n567 VDD.n566 0.000506553
R3130 VDD.n565 VDD.n564 0.000506553
R3131 VDD.n695 VDD.n694 0.000506553
R3132 VDD.n1138 VDD.n1019 0.000506553
R3133 VDD.n1140 VDD.n1139 0.000506553
R3134 VDD.n1018 VDD.n1017 0.000506553
R3135 VDD.n964 VDD.n963 0.000506553
R3136 VDD.n962 VDD.n961 0.000506553
R3137 VDD.n1137 VDD.n1136 0.000506553
R3138 VDD.n1477 VDD.n1476 0.000506553
R3139 VDD.n1405 VDD.n1241 0.000506553
R3140 VDD.n1404 VDD.n1403 0.000506553
R3141 VDD.n1347 VDD.n1346 0.000506553
R3142 VDD.n1345 VDD.n1344 0.000506553
R3143 VDD.n1475 VDD.n1474 0.000506553
R3144 VDD.n166 VDD.n165 0.000506553
R3145 VDD.n331 VDD.n330 0.000506553
R3146 VDD.n164 VDD.n81 0.000506553
R3147 VDD.n136 VDD.n135 0.000506553
R3148 VDD.n111 VDD.n110 0.000506553
R3149 VDD.n109 VDD.n108 0.000506553
R3150 VDD.n254 VDD.n253 0.000506553
R3151 VDD.n329 VDD.n328 0.000506553
R3152 VDD.n167 VDD.n166 0.000503441
R3153 VDD.n137 VDD.n136 0.000503441
R3154 VDD.n108 VDD.n107 0.000503441
R3155 VDD.n328 VDD.n327 0.000503441
R3156 VDD.n255 VDD.n254 0.000503441
R3157 VDD.n193 VDD.n192 0.000501258
R3158 VDD.n139 VDD.n138 0.000501258
R3159 VDD.n99 VDD.n98 0.000501258
R3160 VDD.n169 VDD.n168 0.000501258
R3161 VDD.n326 VDD.n325 0.000501258
R3162 VDD.n257 VDD.n256 0.000501258
R3163 VDD.n697 VDD.n479 0.00050097
R3164 VDD.n723 VDD.n461 0.00050097
R3165 VDD.n623 VDD.n482 0.00050097
R3166 VDD.n564 VDD.n504 0.00050097
R3167 VDD.n1036 VDD.n1019 0.00050097
R3168 VDD.n1140 VDD.n876 0.00050097
R3169 VDD.n1017 VDD.n879 0.00050097
R3170 VDD.n961 VDD.n901 0.00050097
R3171 VDD.n1477 VDD.n1259 0.00050097
R3172 VDD.n1503 VDD.n1241 0.00050097
R3173 VDD.n1403 VDD.n1262 0.00050097
R3174 VDD.n1344 VDD.n1284 0.00050097
R3175 VDD.n694 VDD.n693 0.00050097
R3176 VDD.n1136 VDD.n1135 0.00050097
R3177 VDD.n1474 VDD.n1473 0.00050097
R3178 VDD.n359 VDD.n358 0.000500071
R3179 A2.n82 A2.n80 145.809
R3180 A2.n25 A2.n23 145.809
R3181 A2.n124 A2.n122 145.809
R3182 A2.n62 A2.n60 145.808
R3183 A2.n25 A2.n24 107.409
R3184 A2.n27 A2.n26 107.409
R3185 A2.n29 A2.n28 107.409
R3186 A2.n31 A2.n30 107.409
R3187 A2.n33 A2.n32 107.409
R3188 A2.n35 A2.n34 107.409
R3189 A2.n124 A2.n123 107.409
R3190 A2.n126 A2.n125 107.409
R3191 A2.n128 A2.n127 107.409
R3192 A2.n130 A2.n129 107.409
R3193 A2.n132 A2.n131 107.409
R3194 A2.n134 A2.n133 107.409
R3195 A2.n82 A2.n81 107.407
R3196 A2.n84 A2.n83 107.407
R3197 A2.n86 A2.n85 107.407
R3198 A2.n88 A2.n87 107.407
R3199 A2.n90 A2.n89 107.407
R3200 A2.n92 A2.n91 107.407
R3201 A2.n62 A2.n61 107.407
R3202 A2.n64 A2.n63 107.407
R3203 A2.n66 A2.n65 107.407
R3204 A2.n68 A2.n67 107.407
R3205 A2.n70 A2.n69 107.407
R3206 A2.n72 A2.n71 107.407
R3207 A2.n98 A2.n96 87.1779
R3208 A2.n43 A2.n41 87.1779
R3209 A2.n4 A2.n2 87.1779
R3210 A2.n142 A2.n140 87.1779
R3211 A2.n14 A2.n13 52.82
R3212 A2.n152 A2.n151 52.82
R3213 A2.n98 A2.n97 52.82
R3214 A2.n100 A2.n99 52.82
R3215 A2.n102 A2.n101 52.82
R3216 A2.n104 A2.n103 52.82
R3217 A2.n106 A2.n105 52.82
R3218 A2.n108 A2.n107 52.82
R3219 A2.n43 A2.n42 52.82
R3220 A2.n45 A2.n44 52.82
R3221 A2.n47 A2.n46 52.82
R3222 A2.n49 A2.n48 52.82
R3223 A2.n51 A2.n50 52.82
R3224 A2.n53 A2.n52 52.82
R3225 A2.n4 A2.n3 52.82
R3226 A2.n6 A2.n5 52.82
R3227 A2.n8 A2.n7 52.82
R3228 A2.n10 A2.n9 52.82
R3229 A2.n12 A2.n11 52.82
R3230 A2.n142 A2.n141 52.82
R3231 A2.n144 A2.n143 52.82
R3232 A2.n146 A2.n145 52.82
R3233 A2.n148 A2.n147 52.82
R3234 A2.n150 A2.n149 52.82
R3235 A2 A2.n109 51.0745
R3236 A2 A2.n54 51.0745
R3237 A2.n84 A2.n82 38.4005
R3238 A2.n86 A2.n84 38.4005
R3239 A2.n88 A2.n86 38.4005
R3240 A2.n90 A2.n88 38.4005
R3241 A2.n92 A2.n90 38.4005
R3242 A2.n93 A2.n92 38.4005
R3243 A2.n64 A2.n62 38.4005
R3244 A2.n66 A2.n64 38.4005
R3245 A2.n68 A2.n66 38.4005
R3246 A2.n70 A2.n68 38.4005
R3247 A2.n72 A2.n70 38.4005
R3248 A2.n73 A2.n72 38.4005
R3249 A2.n27 A2.n25 38.4005
R3250 A2.n29 A2.n27 38.4005
R3251 A2.n31 A2.n29 38.4005
R3252 A2.n33 A2.n31 38.4005
R3253 A2.n35 A2.n33 38.4005
R3254 A2.n36 A2.n35 38.4005
R3255 A2.n126 A2.n124 38.4005
R3256 A2.n128 A2.n126 38.4005
R3257 A2.n130 A2.n128 38.4005
R3258 A2.n132 A2.n130 38.4005
R3259 A2.n134 A2.n132 38.4005
R3260 A2.n135 A2.n134 38.4005
R3261 A2.n100 A2.n98 34.3584
R3262 A2.n102 A2.n100 34.3584
R3263 A2.n104 A2.n102 34.3584
R3264 A2.n106 A2.n104 34.3584
R3265 A2.n108 A2.n106 34.3584
R3266 A2.n110 A2.n108 34.3584
R3267 A2.n45 A2.n43 34.3584
R3268 A2.n47 A2.n45 34.3584
R3269 A2.n49 A2.n47 34.3584
R3270 A2.n51 A2.n49 34.3584
R3271 A2.n53 A2.n51 34.3584
R3272 A2.n55 A2.n53 34.3584
R3273 A2.n6 A2.n4 34.3584
R3274 A2.n8 A2.n6 34.3584
R3275 A2.n10 A2.n8 34.3584
R3276 A2.n12 A2.n10 34.3584
R3277 A2.n14 A2.n12 34.3584
R3278 A2.n18 A2.n14 34.3584
R3279 A2.n144 A2.n142 34.3584
R3280 A2.n146 A2.n144 34.3584
R3281 A2.n148 A2.n146 34.3584
R3282 A2.n150 A2.n148 34.3584
R3283 A2.n152 A2.n150 34.3584
R3284 A2.n153 A2.n152 34.3584
R3285 A2.n78 A2.t117 26.5955
R3286 A2.n78 A2.t67 26.5955
R3287 A2.n80 A2.t105 26.5955
R3288 A2.n80 A2.t99 26.5955
R3289 A2.n81 A2.t97 26.5955
R3290 A2.n81 A2.t90 26.5955
R3291 A2.n83 A2.t88 26.5955
R3292 A2.n83 A2.t80 26.5955
R3293 A2.n85 A2.t87 26.5955
R3294 A2.n85 A2.t95 26.5955
R3295 A2.n87 A2.t77 26.5955
R3296 A2.n87 A2.t93 26.5955
R3297 A2.n89 A2.t91 26.5955
R3298 A2.n89 A2.t62 26.5955
R3299 A2.n91 A2.t83 26.5955
R3300 A2.n91 A2.t75 26.5955
R3301 A2.n59 A2.t103 26.5955
R3302 A2.n59 A2.t98 26.5955
R3303 A2.n60 A2.t66 26.5955
R3304 A2.n60 A2.t73 26.5955
R3305 A2.n61 A2.t78 26.5955
R3306 A2.n61 A2.t116 26.5955
R3307 A2.n63 A2.t71 26.5955
R3308 A2.n63 A2.t64 26.5955
R3309 A2.n65 A2.t107 26.5955
R3310 A2.n65 A2.t120 26.5955
R3311 A2.n67 A2.t118 26.5955
R3312 A2.n67 A2.t114 26.5955
R3313 A2.n69 A2.t112 26.5955
R3314 A2.n69 A2.t60 26.5955
R3315 A2.n71 A2.t109 26.5955
R3316 A2.n71 A2.t100 26.5955
R3317 A2.n22 A2.t82 26.5955
R3318 A2.n22 A2.t74 26.5955
R3319 A2.n23 A2.t110 26.5955
R3320 A2.n23 A2.t106 26.5955
R3321 A2.n24 A2.t104 26.5955
R3322 A2.n24 A2.t115 26.5955
R3323 A2.n26 A2.t96 26.5955
R3324 A2.n26 A2.t89 26.5955
R3325 A2.n28 A2.t94 26.5955
R3326 A2.n28 A2.t79 26.5955
R3327 A2.n30 A2.t86 26.5955
R3328 A2.n30 A2.t101 26.5955
R3329 A2.n32 A2.t76 26.5955
R3330 A2.n32 A2.t92 26.5955
R3331 A2.n34 A2.t68 26.5955
R3332 A2.n34 A2.t84 26.5955
R3333 A2.n121 A2.t108 26.5955
R3334 A2.n121 A2.t58 26.5955
R3335 A2.n122 A2.t69 26.5955
R3336 A2.n122 A2.t85 26.5955
R3337 A2.n123 A2.t65 26.5955
R3338 A2.n123 A2.t81 26.5955
R3339 A2.n125 A2.t57 26.5955
R3340 A2.n125 A2.t72 26.5955
R3341 A2.n127 A2.t70 26.5955
R3342 A2.n127 A2.t63 26.5955
R3343 A2.n129 A2.t61 26.5955
R3344 A2.n129 A2.t119 26.5955
R3345 A2.n131 A2.t102 26.5955
R3346 A2.n131 A2.t113 26.5955
R3347 A2.n133 A2.t111 26.5955
R3348 A2.n133 A2.t59 26.5955
R3349 A2.n109 A2.t30 24.9236
R3350 A2.n109 A2.t21 24.9236
R3351 A2.n96 A2.t33 24.9236
R3352 A2.n96 A2.t29 24.9236
R3353 A2.n97 A2.t27 24.9236
R3354 A2.n97 A2.t54 24.9236
R3355 A2.n99 A2.t36 24.9236
R3356 A2.n99 A2.t7 24.9236
R3357 A2.n101 A2.t35 24.9236
R3358 A2.n101 A2.t41 24.9236
R3359 A2.n103 A2.t16 24.9236
R3360 A2.n103 A2.t50 24.9236
R3361 A2.n105 A2.t55 24.9236
R3362 A2.n105 A2.t125 24.9236
R3363 A2.n107 A2.t12 24.9236
R3364 A2.n107 A2.t123 24.9236
R3365 A2.n54 A2.t25 24.9236
R3366 A2.n54 A2.t28 24.9236
R3367 A2.n41 A2.t44 24.9236
R3368 A2.n41 A2.t39 24.9236
R3369 A2.n42 A2.t17 24.9236
R3370 A2.n42 A2.t15 24.9236
R3371 A2.n44 A2.t48 24.9236
R3372 A2.n44 A2.t127 24.9236
R3373 A2.n46 A2.t8 24.9236
R3374 A2.n46 A2.t20 24.9236
R3375 A2.n48 A2.t56 24.9236
R3376 A2.n48 A2.t2 24.9236
R3377 A2.n50 A2.t0 24.9236
R3378 A2.n50 A2.t45 24.9236
R3379 A2.n52 A2.t10 24.9236
R3380 A2.n52 A2.t53 24.9236
R3381 A2.n15 A2.t11 24.9236
R3382 A2.n15 A2.t40 24.9236
R3383 A2.n2 A2.t31 24.9236
R3384 A2.n2 A2.t34 24.9236
R3385 A2.n3 A2.t26 24.9236
R3386 A2.n3 A2.t14 24.9236
R3387 A2.n5 A2.t42 24.9236
R3388 A2.n5 A2.t37 24.9236
R3389 A2.n7 A2.t51 24.9236
R3390 A2.n7 A2.t6 24.9236
R3391 A2.n9 A2.t122 24.9236
R3392 A2.n9 A2.t52 24.9236
R3393 A2.n11 A2.t124 24.9236
R3394 A2.n11 A2.t49 24.9236
R3395 A2.n13 A2.t22 24.9236
R3396 A2.n13 A2.t13 24.9236
R3397 A2.n154 A2.t9 24.9236
R3398 A2.n154 A2.t4 24.9236
R3399 A2.n140 A2.t23 24.9236
R3400 A2.n140 A2.t121 24.9236
R3401 A2.n141 A2.t43 24.9236
R3402 A2.n141 A2.t18 24.9236
R3403 A2.n143 A2.t3 24.9236
R3404 A2.n143 A2.t38 24.9236
R3405 A2.n145 A2.t47 24.9236
R3406 A2.n145 A2.t126 24.9236
R3407 A2.n147 A2.t46 24.9236
R3408 A2.n147 A2.t19 24.9236
R3409 A2.n149 A2.t24 24.9236
R3410 A2.n149 A2.t1 24.9236
R3411 A2.n151 A2.t32 24.9236
R3412 A2.n151 A2.t5 24.9236
R3413 A2 A2.n110 11.4429
R3414 A2 A2.n55 11.4429
R3415 A2 A2.n18 11.4429
R3416 A2.n37 A2.n22 8.55118
R3417 A2.n136 A2.n121 8.55118
R3418 A2.n74 A2.n59 8.55117
R3419 A2.n79 A2.n78 8.47293
R3420 A2.n16 A2.n15 7.80093
R3421 A2.n155 A2.n154 7.80093
R3422 A2.n38 A2.n37 3.20954
R3423 A2.n137 A2.n136 3.20953
R3424 A2.n75 A2.n74 3.20289
R3425 A2.n111 A2 3.10353
R3426 A2.n56 A2 3.10353
R3427 A2.n19 A2 3.10353
R3428 A2 A2.n159 3.10353
R3429 A2.n95 A2.n94 3.1005
R3430 A2.n17 A2.n1 3.1005
R3431 A2.n157 A2.n156 3.1005
R3432 A2.n94 A2.n93 2.71565
R3433 A2.n74 A2.n73 2.13383
R3434 A2.n37 A2.n36 2.13383
R3435 A2.n136 A2.n135 2.13383
R3436 A2.n110 A2 1.74595
R3437 A2.n55 A2 1.74595
R3438 A2.n18 A2.n17 1.16414
R3439 A2.n156 A2.n153 1.16414
R3440 A2.n117 A2.n116 1.07337
R3441 A2.n118 A2.n117 0.69375
R3442 A2.n119 A2.n118 0.68905
R3443 A2.n16 A2 0.488972
R3444 A2.n155 A2 0.488972
R3445 A2.n118 A2.n39 0.414635
R3446 A2.n117 A2.n76 0.382465
R3447 A2.n119 A2 0.380486
R3448 A2.n120 A2.n119 0.368576
R3449 A2.n94 A2.n79 0.196887
R3450 A2.n39 A2.n38 0.157252
R3451 A2.n137 A2.n120 0.139891
R3452 A2.n116 A2.n115 0.139389
R3453 A2.n76 A2.n75 0.132946
R3454 A2.n20 A2.n1 0.113
R3455 A2.n158 A2.n157 0.113
R3456 A2.n114 A2.n95 0.101889
R3457 A2.n17 A2.n16 0.0893205
R3458 A2.n156 A2.n155 0.0893205
R3459 A2.n114 A2.n112 0.0282778
R3460 A2.n95 A2.n77 0.0268889
R3461 A2.n58 A2.n57 0.0213333
R3462 A2.n21 A2.n20 0.0143889
R3463 A2.n158 A2.n139 0.0143889
R3464 A2.n75 A2.n58 0.00100004
R3465 A2.n139 A2.n137 0.00100004
R3466 A2.n38 A2.n21 0.00100004
R3467 A2.n112 A2.n111 0.000513335
R3468 A2.n57 A2.n56 0.000513335
R3469 A2.n20 A2.n19 0.000513218
R3470 A2.n159 A2.n158 0.000513218
R3471 A2.n58 A2.n40 0.00050517
R3472 A2.n114 A2.n113 0.000504838
R3473 A2.n21 A2.n0 0.000504838
R3474 A2.n139 A2.n138 0.000504838
R3475 A2.n115 A2.n114 0.000501713
R3476 I2.n4 I2.t3 323.342
R3477 I2.n0 I2.t0 228.927
R3478 I2.n2 I2.t5 196.549
R3479 I2.n4 I2.t1 194.809
R3480 I2.n0 I2.t4 159.391
R3481 I2.n2 I2.t2 148.35
R3482 I2.n5 I2.n4 76.0005
R3483 I2.n3 I2.n2 76.0005
R3484 I2.n6 I2.n5 29.2624
R3485 I2.n7 I2 9.11
R3486 I2.n1 I2.n0 8.68501
R3487 I2.n3 I2 5.78114
R3488 I2.n8 I2.n1 4.26764
R3489 I2 I2.n3 3.71663
R3490 I2.n1 I2 1.99697
R3491 I2.n5 I2 1.92927
R3492 I2.n7 I2.n6 1.79514
R3493 I2.n8 I2.n7 0.570143
R3494 I2.n6 I2 0.449389
R3495 I2 I2.n8 0.221483
R3496 GND.n1547 GND 2.276e+06
R3497 GND.n1547 GND 2.00869e+06
R3498 GND GND.n542 334900
R3499 GND.n367 GND 334900
R3500 GND GND.n1543 271091
R3501 GND.n461 GND 271091
R3502 GND.n542 GND.n123 215600
R3503 GND.n368 GND.n367 215600
R3504 GND.n537 GND.n536 18654.2
R3505 GND.n1544 GND.t451 10105.3
R3506 GND.t540 GND.n460 10105.3
R3507 GND.n121 GND.n120 7236.84
R3508 GND.n1545 GND.t465 5863.39
R3509 GND.t62 GND.n364 5863.39
R3510 GND.n536 GND 5222.01
R3511 GND.t741 GND.n1534 4783.15
R3512 GND.n369 GND.t262 3113.6
R3513 GND.n367 GND.n366 3003.29
R3514 GND.n371 GND.n370 2817.54
R3515 GND.n493 GND.n492 2786.18
R3516 GND.n1532 GND.n1531 2744.41
R3517 GND.n100 GND.n99 2744.41
R3518 GND.n1546 GND.t557 2656.51
R3519 GND.n1550 GND.n1549 2243.42
R3520 GND.t394 GND.n535 2135.29
R3521 GND.n1548 GND.n122 1899.15
R3522 GND.t544 GND 1848
R3523 GND.n1548 GND.n1547 1742.45
R3524 GND.n1546 GND.n1545 1566.95
R3525 GND.n1545 GND.n1544 1560.68
R3526 GND.n122 GND.n100 1548.15
R3527 GND.n1533 GND.n1532 1548.15
R3528 GND.t569 GND.t538 1408
R3529 GND.t538 GND 1353
R3530 GND.t459 GND.n1548 1269.38
R3531 GND GND.t482 1255.01
R3532 GND.t594 GND 1255.01
R3533 GND.t0 GND.t544 1188
R3534 GND GND.t769 1129.73
R3535 GND GND.t571 1111
R3536 GND.t753 GND.t741 1078
R3537 GND.t492 GND.t445 1056
R3538 GND.n493 GND.n461 940.789
R3539 GND.t484 GND.t753 924
R3540 GND.t445 GND.t484 924
R3541 GND.t571 GND.t0 924
R3542 GND.t252 GND 917.571
R3543 GND GND.t747 917.571
R3544 GND.n1535 GND 909.476
R3545 GND.n1535 GND.n672 892.495
R3546 GND.t831 GND.n834 869.471
R3547 GND.n536 GND 867.972
R3548 GND.t86 GND 860.76
R3549 GND.t559 GND 860.76
R3550 GND.t39 GND 860.76
R3551 GND.t455 GND 850.634
R3552 GND.t482 GND.t255 806.792
R3553 GND.t82 GND.t594 806.792
R3554 GND.t77 GND.t569 792
R3555 GND.t254 GND.t77 792
R3556 GND GND.t71 784.713
R3557 GND GND.t64 784.713
R3558 GND.t573 GND.t557 780.297
R3559 GND.t262 GND.t486 780.297
R3560 GND.t488 GND.t45 777.333
R3561 GND.t60 GND.t584 777.333
R3562 GND.t567 GND 754.5
R3563 GND GND.t57 754.5
R3564 GND.t372 GND.n1119 751.37
R3565 GND.t465 GND.t554 732.088
R3566 GND.t909 GND.t62 732.088
R3567 GND GND.t476 729.721
R3568 GND.t768 GND 729.721
R3569 GND.t568 GND 726
R3570 GND GND.t58 726
R3571 GND.t479 GND.t751 717.149
R3572 GND.t400 GND.t498 717.149
R3573 GND GND.t254 715
R3574 GND.t542 GND.t252 708.047
R3575 GND.t747 GND.t477 708.047
R3576 GND GND.t492 704
R3577 GND.t588 GND 654.159
R3578 GND.n370 GND.n369 654.136
R3579 GND.n371 GND 654.054
R3580 GND.t554 GND.t763 627.505
R3581 GND.t763 GND.t479 627.505
R3582 GND.t255 GND.t567 627.505
R3583 GND.t471 GND.t909 627.505
R3584 GND.t498 GND.t471 627.505
R3585 GND.t57 GND.t82 627.505
R3586 GND.t476 GND.t573 606.898
R3587 GND.t592 GND.t542 606.898
R3588 GND.t474 GND.t592 606.898
R3589 GND.t486 GND.t768 606.898
R3590 GND.t477 GND.t745 606.898
R3591 GND.t745 GND.t37 606.898
R3592 GND.t778 GND.t572 601.333
R3593 GND.t504 GND.t502 601.333
R3594 GND.n122 GND.n121 578.947
R3595 GND GND.t257 546.497
R3596 GND GND.t68 546.497
R3597 GND GND.t394 536.71
R3598 GND GND.t86 536.71
R3599 GND GND.t559 536.71
R3600 GND GND.t455 536.71
R3601 GND GND.t39 536.71
R3602 GND GND.t596 513.333
R3603 GND.t467 GND.t469 498.408
R3604 GND.t469 GND 478.938
R3605 GND.t751 GND 478.099
R3606 GND GND.t400 478.099
R3607 GND.n1543 GND.n1542 459.635
R3608 GND.n370 GND.n364 445.014
R3609 GND.t765 GND.t588 420.531
R3610 GND.n123 GND 420.382
R3611 GND.n368 GND 420.382
R3612 GND.n123 GND.t474 419.048
R3613 GND.t37 GND.n368 419.048
R3614 GND GND.t80 393.274
R3615 GND.t396 GND.t459 381.594
R3616 GND.t461 GND.t447 373.805
R3617 GND.n542 GND.n541 370.385
R3618 GND.t731 GND 352.382
R3619 GND GND.t564 339.942
R3620 GND GND.t2 339.942
R3621 GND.t500 GND.t396 327.08
R3622 GND.t447 GND.t500 327.08
R3623 GND.t80 GND.t765 327.08
R3624 GND.t505 GND.t507 324.212
R3625 GND.t513 GND.t505 324.212
R3626 GND.t519 GND.t515 324.212
R3627 GND.t515 GND.t521 324.212
R3628 GND.t521 GND.t509 324.212
R3629 GND.t509 GND.t517 324.212
R3630 GND.t523 GND.t527 324.212
R3631 GND.t533 GND.t529 324.212
R3632 GND.t529 GND.t525 324.212
R3633 GND.t535 GND.t531 324.212
R3634 GND.t596 GND.t600 324.212
R3635 GND.t600 GND.t598 324.212
R3636 GND.t598 GND.t449 324.212
R3637 GND.t531 GND 301.053
R3638 GND.n1549 GND 299.824
R3639 GND.n373 GND.t525 285.615
R3640 GND.t773 GND.t467 280.354
R3641 GND.t4 GND.t773 280.354
R3642 GND.n410 GND.t519 270.175
R3643 GND GND.t78 266.514
R3644 GND GND.t84 266.514
R3645 GND GND.t490 263.26
R3646 GND GND.t110 255.238
R3647 GND.t108 GND 255.238
R3648 GND GND.t184 255.238
R3649 GND.t240 GND 255.238
R3650 GND GND.t735 253.333
R3651 GND GND.t4 253.097
R3652 GND.t547 GND.n1530 251.429
R3653 GND.n460 GND.n459 250.713
R3654 GND GND.t461 249.204
R3655 GND.n1534 GND.n1533 244.445
R3656 GND GND.t576 230.905
R3657 GND GND.t3 230.905
R3658 GND GND.t494 227.501
R3659 GND.n1547 GND.n1546 213.106
R3660 GND.n372 GND 211.114
R3661 GND GND.t547 201.905
R3662 GND.n370 GND.t523 196.843
R3663 GND.n1353 GND.t443 193.933
R3664 GND.n1066 GND.t762 193.933
R3665 GND.n1506 GND.t738 193.933
R3666 GND.n338 GND.t602 193.933
R3667 GND.n1090 GND.t552 193.532
R3668 GND.n1343 GND.t441 192.982
R3669 GND.n1056 GND.t760 192.982
R3670 GND.n1496 GND.t736 192.982
R3671 GND.n357 GND.t597 192.982
R3672 GND.t879 GND 190.686
R3673 GND GND.t877 190.686
R3674 GND.t825 GND 190.686
R3675 GND GND.t13 190.686
R3676 GND GND.t759 189.263
R3677 GND.t463 GND.t731 184.762
R3678 GND.n123 GND 182.167
R3679 GND.n368 GND 182.167
R3680 GND GND.t75 181.03
R3681 GND GND.t85 181.03
R3682 GND GND.t549 179.048
R3683 GND.n1531 GND 176.386
R3684 GND.n99 GND 176.386
R3685 GND.t320 GND 164.786
R3686 GND GND.t362 164.786
R3687 GND.t390 GND 164.786
R3688 GND GND.t412 164.786
R3689 GND GND.t440 163.555
R3690 GND.n1377 GND.t457 162.326
R3691 GND.t100 GND.t190 160
R3692 GND.t218 GND.t100 160
R3693 GND.t116 GND.t218 160
R3694 GND.t188 GND.t116 160
R3695 GND.t94 GND.t188 160
R3696 GND.t120 GND.t170 160
R3697 GND.t170 GND.t206 160
R3698 GND.t206 GND.t132 160
R3699 GND.t132 GND.t174 160
R3700 GND.t174 GND.t210 160
R3701 GND.t210 GND.t136 160
R3702 GND.t136 GND.t156 160
R3703 GND.t156 GND.t150 160
R3704 GND.t150 GND.t182 160
R3705 GND.t110 GND.t160 160
R3706 GND.t160 GND.t216 160
R3707 GND.t216 GND.t114 160
R3708 GND.t200 GND.t164 160
R3709 GND.t126 GND.t200 160
R3710 GND.t152 GND.t126 160
R3711 GND.t204 GND.t152 160
R3712 GND.t192 GND.t204 160
R3713 GND.t102 GND.t192 160
R3714 GND.t146 GND.t102 160
R3715 GND.t176 GND.t146 160
R3716 GND.t212 GND.t176 160
R3717 GND.t138 GND.t212 160
R3718 GND.t180 GND.t138 160
R3719 GND.t158 GND.t108 160
R3720 GND.t194 GND.t158 160
R3721 GND.t186 GND.t194 160
R3722 GND.t92 GND.t186 160
R3723 GND.t118 GND.t168 160
R3724 GND.t168 GND.t96 160
R3725 GND.t96 GND.t142 160
R3726 GND.t142 GND.t172 160
R3727 GND.t172 GND.t208 160
R3728 GND.t208 GND.t134 160
R3729 GND.t134 GND.t154 160
R3730 GND.t154 GND.t122 160
R3731 GND.t122 GND.t128 160
R3732 GND.t128 GND.t106 160
R3733 GND.t184 GND.t214 160
R3734 GND.t214 GND.t112 160
R3735 GND.t112 GND.t162 160
R3736 GND.t140 GND.t198 160
R3737 GND.t166 GND.t140 160
R3738 GND.t202 GND.t166 160
R3739 GND.t130 GND.t202 160
R3740 GND.t98 GND.t130 160
R3741 GND.t144 GND.t98 160
R3742 GND.t196 GND.t144 160
R3743 GND.t104 GND.t196 160
R3744 GND.t148 GND.t104 160
R3745 GND.t178 GND.t148 160
R3746 GND.t124 GND.t178 160
R3747 GND.t250 GND.t240 160
R3748 GND.t228 GND.t250 160
R3749 GND.t242 GND.t226 160
R3750 GND.t226 GND.t248 160
R3751 GND.t248 GND.t220 160
R3752 GND.t220 GND.t232 160
R3753 GND.t232 GND.t244 160
R3754 GND.t244 GND.t222 160
R3755 GND.t222 GND.t234 160
R3756 GND.t234 GND.t246 160
R3757 GND.t246 GND.t224 160
R3758 GND.t224 GND.t230 160
R3759 GND.t230 GND.t238 160
R3760 GND.t238 GND.t236 160
R3761 GND.t735 GND.t739 160
R3762 GND.t739 GND.t733 160
R3763 GND.t733 GND.t737 160
R3764 GND.t549 GND.t463 160
R3765 GND.n1356 GND.t67 154.006
R3766 GND.n1069 GND.t52 154.006
R3767 GND.n1509 GND.t550 154.006
R3768 GND.t552 GND 150.841
R3769 GND.n75 GND.t462 150.465
R3770 GND.n475 GND.t551 150.465
R3771 GND.n53 GND.t401 150.465
R3772 GND.n3 GND.t70 150.465
R3773 GND.n36 GND.t580 150.465
R3774 GND.n631 GND.t493 150.465
R3775 GND.n556 GND.t749 150.465
R3776 GND.n586 GND.t752 150.465
R3777 GND.n125 GND.t586 150.465
R3778 GND.n158 GND.t767 150.465
R3779 GND GND.t693 149.645
R3780 GND GND.t635 149.645
R3781 GND GND.t685 149.645
R3782 GND.t511 GND 149.645
R3783 GND.t182 GND 148.571
R3784 GND GND.t180 148.571
R3785 GND.t106 GND 148.571
R3786 GND.t198 GND.n1453 148.571
R3787 GND GND.t124 148.571
R3788 GND.t236 GND 148.571
R3789 GND.n1534 GND 146.667
R3790 GND.t737 GND 142.857
R3791 GND.n1533 GND 138.286
R3792 GND.n122 GND 138.286
R3793 GND.t490 GND.t55 138.035
R3794 GND.t51 GND 133.766
R3795 GND.n788 GND.t118 133.333
R3796 GND.t457 GND 130.352
R3797 GND.n459 GND.t507 127.368
R3798 GND.n370 GND.t533 127.368
R3799 GND.t869 GND.t831 119.534
R3800 GND.t859 GND.t869 119.534
R3801 GND.t885 GND.t859 119.534
R3802 GND.t829 GND.t885 119.534
R3803 GND.t863 GND.t829 119.534
R3804 GND.t811 GND.t887 119.534
R3805 GND.t847 GND.t811 119.534
R3806 GND.t899 GND.t847 119.534
R3807 GND.t815 GND.t899 119.534
R3808 GND.t851 GND.t815 119.534
R3809 GND.t903 GND.t851 119.534
R3810 GND.t797 GND.t903 119.534
R3811 GND.t791 GND.t797 119.534
R3812 GND.t823 GND.t791 119.534
R3813 GND.t801 GND.t879 119.534
R3814 GND.t857 GND.t801 119.534
R3815 GND.t883 GND.t857 119.534
R3816 GND.t805 GND.t841 119.534
R3817 GND.t841 GND.t895 119.534
R3818 GND.t895 GND.t793 119.534
R3819 GND.t793 GND.t845 119.534
R3820 GND.t845 GND.t833 119.534
R3821 GND.t833 GND.t871 119.534
R3822 GND.t871 GND.t787 119.534
R3823 GND.t787 GND.t817 119.534
R3824 GND.t817 GND.t853 119.534
R3825 GND.t853 GND.t907 119.534
R3826 GND.t907 GND.t821 119.534
R3827 GND.t877 GND.t799 119.534
R3828 GND.t799 GND.t835 119.534
R3829 GND.t835 GND.t827 119.534
R3830 GND.t827 GND.t861 119.534
R3831 GND.t809 GND.t889 119.534
R3832 GND.t865 GND.t809 119.534
R3833 GND.t783 GND.t865 119.534
R3834 GND.t813 GND.t783 119.534
R3835 GND.t849 GND.t813 119.534
R3836 GND.t901 GND.t849 119.534
R3837 GND.t795 GND.t901 119.534
R3838 GND.t891 GND.t795 119.534
R3839 GND.t905 GND.t891 119.534
R3840 GND.t875 GND.t905 119.534
R3841 GND.t855 GND.t825 119.534
R3842 GND.t881 GND.t855 119.534
R3843 GND.t803 GND.t881 119.534
R3844 GND.t839 GND.t781 119.534
R3845 GND.t781 GND.t807 119.534
R3846 GND.t807 GND.t843 119.534
R3847 GND.t843 GND.t897 119.534
R3848 GND.t897 GND.t867 119.534
R3849 GND.t867 GND.t785 119.534
R3850 GND.t785 GND.t837 119.534
R3851 GND.t837 GND.t873 119.534
R3852 GND.t873 GND.t789 119.534
R3853 GND.t789 GND.t819 119.534
R3854 GND.t819 GND.t893 119.534
R3855 GND.t13 GND.t23 119.534
R3856 GND.t23 GND.t33 119.534
R3857 GND.t15 GND.t31 119.534
R3858 GND.t31 GND.t21 119.534
R3859 GND.t21 GND.t25 119.534
R3860 GND.t25 GND.t5 119.534
R3861 GND.t5 GND.t17 119.534
R3862 GND.t17 GND.t27 119.534
R3863 GND.t27 GND.t7 119.534
R3864 GND.t7 GND.t19 119.534
R3865 GND.t19 GND.t29 119.534
R3866 GND.t29 GND.t35 119.534
R3867 GND.t35 GND.t11 119.534
R3868 GND.t11 GND.t9 119.534
R3869 GND.t759 GND.t755 119.534
R3870 GND.t755 GND.t757 119.534
R3871 GND.t757 GND.t761 119.534
R3872 GND.t55 GND.t51 119.534
R3873 GND.t494 GND.t453 119.285
R3874 GND.t71 GND.t776 119.109
R3875 GND.t257 GND.t582 119.109
R3876 GND.t64 GND.t47 119.109
R3877 GND.t68 GND.t392 119.109
R3878 GND.n1361 GND.n1360 118.1
R3879 GND.n1074 GND.n1073 118.1
R3880 GND.n1514 GND.n1513 118.1
R3881 GND.n14 GND.n13 117.984
R3882 GND.n136 GND.n135 117.984
R3883 GND.n1122 GND.t373 117.626
R3884 GND.n837 GND.t832 117.626
R3885 GND.n683 GND.t191 117.626
R3886 GND.n165 GND.t656 117.007
R3887 GND.n1092 GND.t839 116.689
R3888 GND.n95 GND.n94 116.052
R3889 GND.n651 GND.n650 116.052
R3890 GND.t66 GND 115.596
R3891 GND.n1348 GND.n1347 114.713
R3892 GND.n1300 GND.n1299 114.713
R3893 GND.n1308 GND.n1307 114.713
R3894 GND.n1314 GND.n1313 114.713
R3895 GND.n1318 GND.n1317 114.713
R3896 GND.n1324 GND.n1323 114.713
R3897 GND.n1330 GND.n1329 114.713
R3898 GND.n1336 GND.n1335 114.713
R3899 GND.n1386 GND.n1385 114.713
R3900 GND.n1114 GND.n1113 114.713
R3901 GND.n1266 GND.n1265 114.713
R3902 GND.n1270 GND.n1269 114.713
R3903 GND.n1276 GND.n1275 114.713
R3904 GND.n1282 GND.n1281 114.713
R3905 GND.n1288 GND.n1287 114.713
R3906 GND.n1219 GND.n1218 114.713
R3907 GND.n1226 GND.n1225 114.713
R3908 GND.n1252 GND.n1251 114.713
R3909 GND.n1248 GND.n1247 114.713
R3910 GND.n1242 GND.n1241 114.713
R3911 GND.n1236 GND.n1235 114.713
R3912 GND.n1230 GND.n1229 114.713
R3913 GND.n1135 GND.n1134 114.713
R3914 GND.n1178 GND.n1177 114.713
R3915 GND.n1185 GND.n1184 114.713
R3916 GND.n1189 GND.n1188 114.713
R3917 GND.n1195 GND.n1194 114.713
R3918 GND.n1201 GND.n1200 114.713
R3919 GND.n1207 GND.n1206 114.713
R3920 GND.n1121 GND.n1120 114.713
R3921 GND.n1126 GND.n1125 114.713
R3922 GND.n1168 GND.n1167 114.713
R3923 GND.n1163 GND.n1162 114.713
R3924 GND.n1157 GND.n1156 114.713
R3925 GND.n1151 GND.n1150 114.713
R3926 GND.n1145 GND.n1144 114.713
R3927 GND.n1061 GND.n1060 114.713
R3928 GND.n1013 GND.n1012 114.713
R3929 GND.n1021 GND.n1020 114.713
R3930 GND.n1027 GND.n1026 114.713
R3931 GND.n1031 GND.n1030 114.713
R3932 GND.n1037 GND.n1036 114.713
R3933 GND.n1043 GND.n1042 114.713
R3934 GND.n1049 GND.n1048 114.713
R3935 GND.n1099 GND.n1098 114.713
R3936 GND.n829 GND.n828 114.713
R3937 GND.n978 GND.n977 114.713
R3938 GND.n982 GND.n981 114.713
R3939 GND.n988 GND.n987 114.713
R3940 GND.n994 GND.n993 114.713
R3941 GND.n1000 GND.n999 114.713
R3942 GND.n935 GND.n934 114.713
R3943 GND.n942 GND.n941 114.713
R3944 GND.n964 GND.n963 114.713
R3945 GND.n960 GND.n959 114.713
R3946 GND.n954 GND.n953 114.713
R3947 GND.n948 GND.n947 114.713
R3948 GND.n823 GND.n822 114.713
R3949 GND.n851 GND.n850 114.713
R3950 GND.n894 GND.n893 114.713
R3951 GND.n901 GND.n900 114.713
R3952 GND.n905 GND.n904 114.713
R3953 GND.n911 GND.n910 114.713
R3954 GND.n917 GND.n916 114.713
R3955 GND.n923 GND.n922 114.713
R3956 GND.n836 GND.n835 114.713
R3957 GND.n841 GND.n840 114.713
R3958 GND.n884 GND.n883 114.713
R3959 GND.n879 GND.n878 114.713
R3960 GND.n873 GND.n872 114.713
R3961 GND.n867 GND.n866 114.713
R3962 GND.n861 GND.n860 114.713
R3963 GND.n1501 GND.n1500 114.713
R3964 GND.n674 GND.n673 114.713
R3965 GND.n1461 GND.n1460 114.713
R3966 GND.n1467 GND.n1466 114.713
R3967 GND.n1471 GND.n1470 114.713
R3968 GND.n1477 GND.n1476 114.713
R3969 GND.n1483 GND.n1482 114.713
R3970 GND.n1489 GND.n1488 114.713
R3971 GND.n1404 GND.n1403 114.713
R3972 GND.n1448 GND.n1447 114.713
R3973 GND.n1441 GND.n1440 114.713
R3974 GND.n1437 GND.n1436 114.713
R3975 GND.n1431 GND.n1430 114.713
R3976 GND.n1425 GND.n1424 114.713
R3977 GND.n1419 GND.n1418 114.713
R3978 GND.n743 GND.n742 114.713
R3979 GND.n678 GND.n677 114.713
R3980 GND.n795 GND.n794 114.713
R3981 GND.n799 GND.n798 114.713
R3982 GND.n805 GND.n804 114.713
R3983 GND.n811 GND.n810 114.713
R3984 GND.n817 GND.n816 114.713
R3985 GND.n731 GND.n730 114.713
R3986 GND.n782 GND.n781 114.713
R3987 GND.n775 GND.n774 114.713
R3988 GND.n771 GND.n770 114.713
R3989 GND.n765 GND.n764 114.713
R3990 GND.n759 GND.n758 114.713
R3991 GND.n753 GND.n752 114.713
R3992 GND.n682 GND.n681 114.713
R3993 GND.n687 GND.n686 114.713
R3994 GND.n696 GND.n695 114.713
R3995 GND.n701 GND.n700 114.713
R3996 GND.n707 GND.n706 114.713
R3997 GND.n713 GND.n712 114.713
R3998 GND.n719 GND.n718 114.713
R3999 GND.n354 GND.n353 114.713
R4000 GND.n417 GND.n416 114.713
R4001 GND.n407 GND.n406 114.713
R4002 GND.n400 GND.n399 114.713
R4003 GND.n396 GND.n395 114.713
R4004 GND.n390 GND.n389 114.713
R4005 GND.n384 GND.n383 114.713
R4006 GND.n377 GND.n376 114.713
R4007 GND.n273 GND.n272 114.713
R4008 GND.n267 GND.n266 114.713
R4009 GND.n453 GND.n452 114.713
R4010 GND.n448 GND.n447 114.713
R4011 GND.n441 GND.n440 114.713
R4012 GND.n435 GND.n434 114.713
R4013 GND.n428 GND.n427 114.713
R4014 GND.n248 GND.n247 114.713
R4015 GND.n254 GND.n253 114.713
R4016 GND.n261 GND.n260 114.713
R4017 GND.n302 GND.n301 114.713
R4018 GND.n295 GND.n294 114.713
R4019 GND.n289 GND.n288 114.713
R4020 GND.n283 GND.n282 114.713
R4021 GND.n200 GND.n199 114.713
R4022 GND.n206 GND.n205 114.713
R4023 GND.n212 GND.n211 114.713
R4024 GND.n216 GND.n215 114.713
R4025 GND.n222 GND.n221 114.713
R4026 GND.n230 GND.n229 114.713
R4027 GND.n236 GND.n235 114.713
R4028 GND.n168 GND.n167 114.713
R4029 GND.n176 GND.n175 114.713
R4030 GND.n182 GND.n181 114.713
R4031 GND.n186 GND.n185 114.713
R4032 GND.n329 GND.n328 114.713
R4033 GND.n323 GND.n322 114.713
R4034 GND.n317 GND.n316 114.713
R4035 GND.n1295 GND.t413 113.734
R4036 GND.n1112 GND.t391 113.734
R4037 GND.n1214 GND.t363 113.734
R4038 GND.n1132 GND.t321 113.734
R4039 GND.n1007 GND.t14 113.734
R4040 GND.n827 GND.t826 113.734
R4041 GND.n930 GND.t878 113.734
R4042 GND.n848 GND.t880 113.734
R4043 GND.n1411 GND.t241 113.734
R4044 GND.n1399 GND.t185 113.734
R4045 GND.n738 GND.t109 113.734
R4046 GND.n726 GND.t111 113.734
R4047 GND.n335 GND.t512 113.734
R4048 GND.n265 GND.t686 113.734
R4049 GND.n243 GND.t636 113.734
R4050 GND.n195 GND.t694 113.734
R4051 GND.n87 GND.n86 111.957
R4052 GND.n1605 GND.n1604 111.957
R4053 GND.n1607 GND.n1606 111.957
R4054 GND.n55 GND.n54 111.957
R4055 GND.n60 GND.n45 111.957
R4056 GND.n643 GND.n642 111.957
R4057 GND.n611 GND.n610 111.957
R4058 GND.n613 GND.n612 111.957
R4059 GND.n588 GND.n587 111.957
R4060 GND.n593 GND.n578 111.957
R4061 GND.n1557 GND.t566 111.924
R4062 GND.n1558 GND.t44 111.924
R4063 GND.n1559 GND.t435 111.924
R4064 GND.n1560 GND.t261 111.924
R4065 GND.n1561 GND.t563 111.924
R4066 GND.n1355 GND.t458 111.924
R4067 GND.n1068 GND.t553 111.924
R4068 GND.n1508 GND.t548 111.924
R4069 GND.n343 GND.t450 111.924
R4070 GND.n340 GND.t770 111.924
R4071 GND.n495 GND.t395 111.924
R4072 GND.n496 GND.t87 111.924
R4073 GND.n497 GND.t560 111.924
R4074 GND.n498 GND.t456 111.924
R4075 GND.n499 GND.t40 111.924
R4076 GND.n1342 GND.t409 111.296
R4077 GND.n1294 GND.t355 111.296
R4078 GND.n1111 GND.t303 111.296
R4079 GND.n1213 GND.t369 111.296
R4080 GND.n1131 GND.t327 111.296
R4081 GND.n1055 GND.t10 111.296
R4082 GND.n1006 GND.t894 111.296
R4083 GND.n826 GND.t876 111.296
R4084 GND.n929 GND.t822 111.296
R4085 GND.n847 GND.t824 111.296
R4086 GND.n1495 GND.t237 111.296
R4087 GND.n1410 GND.t125 111.296
R4088 GND.n1398 GND.t107 111.296
R4089 GND.n737 GND.t181 111.296
R4090 GND.n725 GND.t183 111.296
R4091 GND.n336 GND.t532 111.296
R4092 GND.n334 GND.t716 111.296
R4093 GND.n264 GND.t728 111.296
R4094 GND.n241 GND.t642 111.296
R4095 GND.n194 GND.t702 111.296
R4096 GND GND.t823 110.996
R4097 GND.t821 GND 110.996
R4098 GND GND.t875 110.996
R4099 GND.t893 GND 110.996
R4100 GND.t9 GND 110.996
R4101 GND.n77 GND.n76 109.359
R4102 GND.n633 GND.n632 109.359
R4103 GND.n472 GND.n471 109.314
R4104 GND.n50 GND.n49 109.314
R4105 GND.n553 GND.n552 109.314
R4106 GND.n583 GND.n582 109.314
R4107 GND.n107 GND.t772 108.505
R4108 GND.n104 GND.t771 108.505
R4109 GND.n468 GND.t81 108.505
R4110 GND.n465 GND.t581 108.505
R4111 GND.n659 GND.t79 108.505
R4112 GND.n656 GND.t76 108.505
R4113 GND.n549 GND.t577 108.505
R4114 GND.n546 GND.t575 108.505
R4115 GND.n79 GND.n78 108.016
R4116 GND.n473 GND.n470 108.016
R4117 GND.n48 GND.n47 108.016
R4118 GND.n30 GND.n29 108.016
R4119 GND.n34 GND.n4 108.016
R4120 GND.n10 GND.n9 108.016
R4121 GND.n635 GND.n634 108.016
R4122 GND.n554 GND.n551 108.016
R4123 GND.n581 GND.n580 108.016
R4124 GND.n152 GND.n151 108.016
R4125 GND.n156 GND.n126 108.016
R4126 GND.n132 GND.n131 108.016
R4127 GND.t761 GND 106.728
R4128 GND.n1454 GND.t242 106.668
R4129 GND.n27 GND.n26 105.975
R4130 GND.n7 GND.n6 105.975
R4131 GND.n17 GND.n12 105.975
R4132 GND.n149 GND.n148 105.975
R4133 GND.n129 GND.n128 105.975
R4134 GND.n139 GND.n134 105.975
R4135 GND.t889 GND.n972 105.305
R4136 GND.t565 GND.n493 103.51
R4137 GND.t272 GND.t372 103.299
R4138 GND.t378 GND.t272 103.299
R4139 GND.t274 GND.t378 103.299
R4140 GND.t360 GND.t274 103.299
R4141 GND.t382 GND.t360 103.299
R4142 GND.t266 GND.t278 103.299
R4143 GND.t296 GND.t266 103.299
R4144 GND.t282 GND.t296 103.299
R4145 GND.t270 GND.t282 103.299
R4146 GND.t300 GND.t270 103.299
R4147 GND.t286 GND.t300 103.299
R4148 GND.t314 GND.t286 103.299
R4149 GND.t294 GND.t314 103.299
R4150 GND.t326 GND.t294 103.299
R4151 GND.t304 GND.t320 103.299
R4152 GND.t292 GND.t304 103.299
R4153 GND.t324 GND.t292 103.299
R4154 GND.t308 GND.t340 103.299
R4155 GND.t340 GND.t328 103.299
R4156 GND.t328 GND.t356 103.299
R4157 GND.t356 GND.t344 103.299
R4158 GND.t344 GND.t316 103.299
R4159 GND.t316 GND.t348 103.299
R4160 GND.t348 GND.t334 103.299
R4161 GND.t334 GND.t364 103.299
R4162 GND.t364 GND.t386 103.299
R4163 GND.t386 GND.t376 103.299
R4164 GND.t376 GND.t368 103.299
R4165 GND.t362 GND.t352 103.299
R4166 GND.t352 GND.t374 103.299
R4167 GND.t374 GND.t358 103.299
R4168 GND.t358 GND.t380 103.299
R4169 GND.t264 GND.t276 103.299
R4170 GND.t384 GND.t264 103.299
R4171 GND.t370 GND.t384 103.299
R4172 GND.t268 GND.t370 103.299
R4173 GND.t298 GND.t268 103.299
R4174 GND.t284 GND.t298 103.299
R4175 GND.t312 GND.t284 103.299
R4176 GND.t388 GND.t312 103.299
R4177 GND.t288 GND.t388 103.299
R4178 GND.t302 GND.t288 103.299
R4179 GND.t290 GND.t390 103.299
R4180 GND.t322 GND.t290 103.299
R4181 GND.t306 GND.t322 103.299
R4182 GND.t338 GND.t280 103.299
R4183 GND.t280 GND.t310 103.299
R4184 GND.t310 GND.t342 103.299
R4185 GND.t342 GND.t330 103.299
R4186 GND.t330 GND.t346 103.299
R4187 GND.t346 GND.t332 103.299
R4188 GND.t332 GND.t318 103.299
R4189 GND.t318 GND.t350 103.299
R4190 GND.t350 GND.t336 103.299
R4191 GND.t336 GND.t366 103.299
R4192 GND.t366 GND.t354 103.299
R4193 GND.t412 GND.t426 103.299
R4194 GND.t426 GND.t420 103.299
R4195 GND.t414 GND.t418 103.299
R4196 GND.t418 GND.t416 103.299
R4197 GND.t416 GND.t428 103.299
R4198 GND.t428 GND.t422 103.299
R4199 GND.t422 GND.t402 103.299
R4200 GND.t402 GND.t430 103.299
R4201 GND.t430 GND.t424 103.299
R4202 GND.t424 GND.t404 103.299
R4203 GND.t404 GND.t432 103.299
R4204 GND.t432 GND.t406 103.299
R4205 GND.t406 GND.t410 103.299
R4206 GND.t410 GND.t408 103.299
R4207 GND.t440 GND.t438 103.299
R4208 GND.t438 GND.t436 103.299
R4209 GND.t436 GND.t442 103.299
R4210 GND.t453 GND.t66 103.299
R4211 GND.n692 GND.t94 102.858
R4212 GND.t164 GND.n787 102.858
R4213 GND.n94 GND.t468 101.43
R4214 GND.n650 GND.t570 101.43
R4215 GND.t43 GND 98.3051
R4216 GND.t434 GND 98.3051
R4217 GND.t562 GND 98.3051
R4218 GND.t260 GND 97.1486
R4219 GND GND.t326 95.92
R4220 GND.t368 GND 95.92
R4221 GND GND.t302 95.92
R4222 GND.n1379 GND.t338 95.92
R4223 GND.t354 GND 95.92
R4224 GND.t408 GND 95.92
R4225 GND.t637 GND.t655 93.8076
R4226 GND.t625 GND.t659 93.8076
R4227 GND.t659 GND.t645 93.8076
R4228 GND.t645 GND.t673 93.8076
R4229 GND.t673 GND.t703 93.8076
R4230 GND.t703 GND.t677 93.8076
R4231 GND.t677 GND.t663 93.8076
R4232 GND.t681 GND.t651 93.8076
R4233 GND.t709 GND.t681 93.8076
R4234 GND.t697 GND.t709 93.8076
R4235 GND.t725 GND.t697 93.8076
R4236 GND.t669 GND.t725 93.8076
R4237 GND.t693 GND.t687 93.8076
R4238 GND.t687 GND.t707 93.8076
R4239 GND.t707 GND.t729 93.8076
R4240 GND.t729 GND.t717 93.8076
R4241 GND.t717 GND.t613 93.8076
R4242 GND.t613 GND.t691 93.8076
R4243 GND.t691 GND.t721 93.8076
R4244 GND.t721 GND.t617 93.8076
R4245 GND.t617 GND.t605 93.8076
R4246 GND.t605 GND.t629 93.8076
R4247 GND.t619 GND.t609 93.8076
R4248 GND.t609 GND.t633 93.8076
R4249 GND.t633 GND.t611 93.8076
R4250 GND.t611 GND.t641 93.8076
R4251 GND.t635 GND.t623 93.8076
R4252 GND.t623 GND.t657 93.8076
R4253 GND.t657 GND.t643 93.8076
R4254 GND.t643 GND.t627 93.8076
R4255 GND.t627 GND.t661 93.8076
R4256 GND.t661 GND.t647 93.8076
R4257 GND.t675 GND.t649 93.8076
R4258 GND.t649 GND.t679 93.8076
R4259 GND.t679 GND.t665 93.8076
R4260 GND.t665 GND.t653 93.8076
R4261 GND.t653 GND.t683 93.8076
R4262 GND.t683 GND.t667 93.8076
R4263 GND.t667 GND.t699 93.8076
R4264 GND.t699 GND.t727 93.8076
R4265 GND.t685 GND.t713 93.8076
R4266 GND.t713 GND.t695 93.8076
R4267 GND.t695 GND.t671 93.8076
R4268 GND.t671 GND.t705 93.8076
R4269 GND.t705 GND.t689 93.8076
R4270 GND.t615 GND.t719 93.8076
R4271 GND.t603 GND.t615 93.8076
R4272 GND.t723 GND.t603 93.8076
R4273 GND.t711 GND.t723 93.8076
R4274 GND.t607 GND.t711 93.8076
R4275 GND.t631 GND.t607 93.8076
R4276 GND.t621 GND.t631 93.8076
R4277 GND.t639 GND.t621 93.8076
R4278 GND.t715 GND.t639 93.8076
R4279 GND.t442 GND 92.2308
R4280 GND.n309 GND.t669 87.1071
R4281 GND.t701 GND 87.1071
R4282 GND.t641 GND 87.1071
R4283 GND.t727 GND 87.1071
R4284 GND GND.t715 87.1071
R4285 GND.t276 GND.n1260 86.0821
R4286 GND.n1091 GND.t15 85.3821
R4287 GND.n890 GND.t805 82.5361
R4288 GND.n308 GND.t619 80.4066
R4289 GND.t576 GND.t911 73.7614
R4290 GND.t3 GND.t590 73.7614
R4291 GND.n86 GND.t766 72.8576
R4292 GND.n1604 GND.t61 72.8576
R4293 GND.n1606 GND.t503 72.8576
R4294 GND.n54 GND.t496 72.8576
R4295 GND.n45 GND.t83 72.8576
R4296 GND.n13 GND.t487 72.8576
R4297 GND.n642 GND.t1 72.8576
R4298 GND.n610 GND.t46 72.8576
R4299 GND.n612 GND.t779 72.8576
R4300 GND.n587 GND.t256 72.8576
R4301 GND.n578 GND.t259 72.8576
R4302 GND.n135 GND.t574 72.8576
R4303 GND.n1530 GND 72.3815
R4304 GND.n123 GND 72.2501
R4305 GND.n368 GND 72.2501
R4306 GND.n1533 GND.n672 71.4001
R4307 GND.n889 GND.t863 71.1519
R4308 GND.n1378 GND.t414 68.8658
R4309 GND.n108 GND.n107 67.973
R4310 GND.n105 GND.n104 67.973
R4311 GND.n479 GND.n468 67.973
R4312 GND.n466 GND.n465 67.973
R4313 GND.n660 GND.n659 67.973
R4314 GND.n657 GND.n656 67.973
R4315 GND.n560 GND.n549 67.973
R4316 GND.n547 GND.n546 67.973
R4317 GND.n163 GND.t637 67.0056
R4318 GND.n1173 GND.t382 66.4063
R4319 GND.n1174 GND.t308 66.4063
R4320 GND.n458 GND.t689 64.7721
R4321 GND GND.t565 61.2963
R4322 GND GND.t43 61.2963
R4323 GND GND.t434 61.2963
R4324 GND GND.t260 61.2963
R4325 GND GND.t562 61.2963
R4326 GND.t78 GND.t90 57.8291
R4327 GND.t75 GND.t578 57.8291
R4328 GND.t84 GND.t49 57.8291
R4329 GND.t85 GND.t53 57.8291
R4330 GND.n692 GND.t120 57.1434
R4331 GND.n787 GND.t114 57.1434
R4332 GND.n459 GND.t511 56.9548
R4333 GND.n1360 GND.t454 55.7148
R4334 GND.n1073 GND.t56 55.7148
R4335 GND.n1513 GND.t464 55.7148
R4336 GND.t88 GND.t73 54.5194
R4337 GND.n1531 GND 54.5194
R4338 GND.t398 GND.t41 54.5194
R4339 GND.n99 GND 54.5194
R4340 GND.n410 GND.t513 54.0356
R4341 GND.n307 GND.t675 53.6046
R4342 GND.n1454 GND.t228 53.3338
R4343 GND.n76 GND.t397 52.8576
R4344 GND.n471 GND.t497 52.8576
R4345 GND.n49 GND.t910 52.8576
R4346 GND.n26 GND.t69 52.8576
R4347 GND.n6 GND.t587 52.8576
R4348 GND.n12 GND.t478 52.8576
R4349 GND.n632 GND.t754 52.8576
R4350 GND.n552 GND.t481 52.8576
R4351 GND.n582 GND.t555 52.8576
R4352 GND.n148 GND.t556 52.8576
R4353 GND.n128 GND.t72 52.8576
R4354 GND.n134 GND.t543 52.8576
R4355 GND.t887 GND.n889 48.3834
R4356 GND GND.n1090 48.3834
R4357 GND.n1533 GND 47.7719
R4358 GND.n122 GND 47.7719
R4359 GND GND.n1377 46.7305
R4360 GND.t647 GND.n307 40.2035
R4361 GND.n118 GND.n117 39.2858
R4362 GND.n489 GND.n488 39.2858
R4363 GND.n1611 GND.n1601 39.2858
R4364 GND.n1615 GND.n1614 39.2858
R4365 GND.n65 GND.n64 39.2858
R4366 GND.n670 GND.n669 39.2858
R4367 GND.n570 GND.n569 39.2858
R4368 GND.n617 GND.n607 39.2858
R4369 GND.n621 GND.n620 39.2858
R4370 GND.n598 GND.n597 39.2858
R4371 GND.n349 GND.n339 39.2858
R4372 GND.n114 GND.n101 38.7881
R4373 GND.n485 GND.n462 38.7881
R4374 GND.n61 GND.n42 38.7881
R4375 GND.n666 GND.n653 38.7881
R4376 GND.n566 GND.n543 38.7881
R4377 GND.n594 GND.n575 38.7881
R4378 GND.n107 GND.t50 38.7697
R4379 GND.n104 GND.t54 38.7697
R4380 GND.n468 GND.t591 38.7697
R4381 GND.n465 GND.t42 38.7697
R4382 GND.n659 GND.t91 38.7697
R4383 GND.n656 GND.t579 38.7697
R4384 GND.n549 GND.t912 38.7697
R4385 GND.n546 GND.t74 38.7697
R4386 GND.n16 GND.n14 38.7523
R4387 GND.n138 GND.n136 38.7523
R4388 GND.n373 GND.t535 38.597
R4389 GND.n78 GND.t501 38.5719
R4390 GND.n78 GND.t448 38.5719
R4391 GND.n470 GND.t399 38.5719
R4392 GND.n470 GND.t537 38.5719
R4393 GND.n47 GND.t472 38.5719
R4394 GND.n47 GND.t499 38.5719
R4395 GND.n29 GND.t473 38.5719
R4396 GND.n29 GND.t444 38.5719
R4397 GND.n4 GND.t546 38.5719
R4398 GND.n4 GND.t65 38.5719
R4399 GND.n9 GND.t746 38.5719
R4400 GND.n9 GND.t38 38.5719
R4401 GND.n634 GND.t485 38.5719
R4402 GND.n634 GND.t446 38.5719
R4403 GND.n551 GND.t750 38.5719
R4404 GND.n551 GND.t89 38.5719
R4405 GND.n580 GND.t764 38.5719
R4406 GND.n580 GND.t480 38.5719
R4407 GND.n151 GND.t258 38.5719
R4408 GND.n151 GND.t775 38.5719
R4409 GND.n126 GND.t743 38.5719
R4410 GND.n126 GND.t561 38.5719
R4411 GND.n131 GND.t593 38.5719
R4412 GND.n131 GND.t475 38.5719
R4413 GND.n890 GND.t883 36.9992
R4414 GND.t278 GND.n1173 36.8926
R4415 GND.n1174 GND.t324 36.8926
R4416 GND.n1585 GND.n1584 34.6358
R4417 GND.n1579 GND.n1578 34.6358
R4418 GND.n1567 GND.n1566 34.6358
R4419 GND.n85 GND.n84 34.6358
R4420 GND.n88 GND.n73 34.6358
R4421 GND.n92 GND.n73 34.6358
R4422 GND.n93 GND.n92 34.6358
R4423 GND.n110 GND.n109 34.6358
R4424 GND.n109 GND.n102 34.6358
R4425 GND.n117 GND.n102 34.6358
R4426 GND.n113 GND.n112 34.6358
R4427 GND.n114 GND.n113 34.6358
R4428 GND.n481 GND.n480 34.6358
R4429 GND.n480 GND.n463 34.6358
R4430 GND.n488 GND.n463 34.6358
R4431 GND.n484 GND.n483 34.6358
R4432 GND.n485 GND.n484 34.6358
R4433 GND.n1611 GND.n1610 34.6358
R4434 GND.n1614 GND.n1602 34.6358
R4435 GND.n64 GND.n43 34.6358
R4436 GND.n57 GND.n56 34.6358
R4437 GND.n23 GND.n22 34.6358
R4438 GND.n641 GND.n640 34.6358
R4439 GND.n644 GND.n629 34.6358
R4440 GND.n648 GND.n629 34.6358
R4441 GND.n649 GND.n648 34.6358
R4442 GND.n662 GND.n661 34.6358
R4443 GND.n661 GND.n654 34.6358
R4444 GND.n669 GND.n654 34.6358
R4445 GND.n665 GND.n664 34.6358
R4446 GND.n666 GND.n665 34.6358
R4447 GND.n562 GND.n561 34.6358
R4448 GND.n561 GND.n544 34.6358
R4449 GND.n569 GND.n544 34.6358
R4450 GND.n565 GND.n564 34.6358
R4451 GND.n566 GND.n565 34.6358
R4452 GND.n617 GND.n616 34.6358
R4453 GND.n620 GND.n608 34.6358
R4454 GND.n597 GND.n576 34.6358
R4455 GND.n590 GND.n589 34.6358
R4456 GND.n145 GND.n144 34.6358
R4457 GND.n1368 GND.n1367 34.6358
R4458 GND.n1081 GND.n1080 34.6358
R4459 GND.n1521 GND.n1520 34.6358
R4460 GND.n523 GND.n522 34.6358
R4461 GND.n517 GND.n516 34.6358
R4462 GND.n505 GND.n504 34.6358
R4463 GND.t420 GND.n1378 34.4331
R4464 GND.t33 GND.n1091 34.1532
R4465 GND.n1573 GND.n1572 33.8829
R4466 GND.n511 GND.n510 33.8829
R4467 GND.n479 GND.n478 32.1329
R4468 GND.n560 GND.n559 32.1329
R4469 GND.t719 GND.n458 29.036
R4470 GND.n1295 GND.n1294 27.8593
R4471 GND.n1112 GND.n1111 27.8593
R4472 GND.n1214 GND.n1213 27.8593
R4473 GND.n1132 GND.n1131 27.8593
R4474 GND.n1007 GND.n1006 27.8593
R4475 GND.n827 GND.n826 27.8593
R4476 GND.n930 GND.n929 27.8593
R4477 GND.n848 GND.n847 27.8593
R4478 GND.n1411 GND.n1410 27.8593
R4479 GND.n1399 GND.n1398 27.8593
R4480 GND.n738 GND.n737 27.8593
R4481 GND.n726 GND.n725 27.8593
R4482 GND.n335 GND.n334 27.8593
R4483 GND.n265 GND.n264 27.8593
R4484 GND.n195 GND.n194 27.8593
R4485 GND.n76 GND.t460 27.5691
R4486 GND.n471 GND.t59 27.5691
R4487 GND.n49 GND.t63 27.5691
R4488 GND.n26 GND.t393 27.5691
R4489 GND.n6 GND.t48 27.5691
R4490 GND.n12 GND.t748 27.5691
R4491 GND.n632 GND.t742 27.5691
R4492 GND.n552 GND.t744 27.5691
R4493 GND.n582 GND.t466 27.5691
R4494 GND.n148 GND.t583 27.5691
R4495 GND.n128 GND.t777 27.5691
R4496 GND.n134 GND.t253 27.5691
R4497 GND.n347 GND.n338 27.1064
R4498 GND.n1360 GND.t495 26.8576
R4499 GND.n1073 GND.t491 26.8576
R4500 GND.n1513 GND.t732 26.8576
R4501 GND.n163 GND.t625 26.8025
R4502 GND.n788 GND.t92 26.6672
R4503 GND.t449 GND.n372 26.1036
R4504 GND.n94 GND.t470 25.9346
R4505 GND.n650 GND.t539 25.9346
R4506 GND.n1347 GND.t439 24.9236
R4507 GND.n1347 GND.t437 24.9236
R4508 GND.n1299 GND.t427 24.9236
R4509 GND.n1299 GND.t421 24.9236
R4510 GND.n1307 GND.t415 24.9236
R4511 GND.n1307 GND.t419 24.9236
R4512 GND.n1313 GND.t417 24.9236
R4513 GND.n1313 GND.t429 24.9236
R4514 GND.n1317 GND.t423 24.9236
R4515 GND.n1317 GND.t403 24.9236
R4516 GND.n1323 GND.t431 24.9236
R4517 GND.n1323 GND.t425 24.9236
R4518 GND.n1329 GND.t405 24.9236
R4519 GND.n1329 GND.t433 24.9236
R4520 GND.n1335 GND.t407 24.9236
R4521 GND.n1335 GND.t411 24.9236
R4522 GND.n1385 GND.t291 24.9236
R4523 GND.n1385 GND.t323 24.9236
R4524 GND.n1113 GND.t307 24.9236
R4525 GND.n1113 GND.t339 24.9236
R4526 GND.n1265 GND.t281 24.9236
R4527 GND.n1265 GND.t311 24.9236
R4528 GND.n1269 GND.t343 24.9236
R4529 GND.n1269 GND.t331 24.9236
R4530 GND.n1275 GND.t347 24.9236
R4531 GND.n1275 GND.t333 24.9236
R4532 GND.n1281 GND.t319 24.9236
R4533 GND.n1281 GND.t351 24.9236
R4534 GND.n1287 GND.t337 24.9236
R4535 GND.n1287 GND.t367 24.9236
R4536 GND.n1218 GND.t353 24.9236
R4537 GND.n1218 GND.t375 24.9236
R4538 GND.n1225 GND.t359 24.9236
R4539 GND.n1225 GND.t381 24.9236
R4540 GND.n1251 GND.t277 24.9236
R4541 GND.n1251 GND.t265 24.9236
R4542 GND.n1247 GND.t385 24.9236
R4543 GND.n1247 GND.t371 24.9236
R4544 GND.n1241 GND.t269 24.9236
R4545 GND.n1241 GND.t299 24.9236
R4546 GND.n1235 GND.t285 24.9236
R4547 GND.n1235 GND.t313 24.9236
R4548 GND.n1229 GND.t389 24.9236
R4549 GND.n1229 GND.t289 24.9236
R4550 GND.n1134 GND.t305 24.9236
R4551 GND.n1134 GND.t293 24.9236
R4552 GND.n1177 GND.t325 24.9236
R4553 GND.n1177 GND.t309 24.9236
R4554 GND.n1184 GND.t341 24.9236
R4555 GND.n1184 GND.t329 24.9236
R4556 GND.n1188 GND.t357 24.9236
R4557 GND.n1188 GND.t345 24.9236
R4558 GND.n1194 GND.t317 24.9236
R4559 GND.n1194 GND.t349 24.9236
R4560 GND.n1200 GND.t335 24.9236
R4561 GND.n1200 GND.t365 24.9236
R4562 GND.n1206 GND.t387 24.9236
R4563 GND.n1206 GND.t377 24.9236
R4564 GND.n1120 GND.t273 24.9236
R4565 GND.n1120 GND.t379 24.9236
R4566 GND.n1125 GND.t275 24.9236
R4567 GND.n1125 GND.t361 24.9236
R4568 GND.n1167 GND.t383 24.9236
R4569 GND.n1167 GND.t279 24.9236
R4570 GND.n1162 GND.t267 24.9236
R4571 GND.n1162 GND.t297 24.9236
R4572 GND.n1156 GND.t283 24.9236
R4573 GND.n1156 GND.t271 24.9236
R4574 GND.n1150 GND.t301 24.9236
R4575 GND.n1150 GND.t287 24.9236
R4576 GND.n1144 GND.t315 24.9236
R4577 GND.n1144 GND.t295 24.9236
R4578 GND.n1060 GND.t756 24.9236
R4579 GND.n1060 GND.t758 24.9236
R4580 GND.n1012 GND.t24 24.9236
R4581 GND.n1012 GND.t34 24.9236
R4582 GND.n1020 GND.t16 24.9236
R4583 GND.n1020 GND.t32 24.9236
R4584 GND.n1026 GND.t22 24.9236
R4585 GND.n1026 GND.t26 24.9236
R4586 GND.n1030 GND.t6 24.9236
R4587 GND.n1030 GND.t18 24.9236
R4588 GND.n1036 GND.t28 24.9236
R4589 GND.n1036 GND.t8 24.9236
R4590 GND.n1042 GND.t20 24.9236
R4591 GND.n1042 GND.t30 24.9236
R4592 GND.n1048 GND.t36 24.9236
R4593 GND.n1048 GND.t12 24.9236
R4594 GND.n1098 GND.t856 24.9236
R4595 GND.n1098 GND.t882 24.9236
R4596 GND.n828 GND.t804 24.9236
R4597 GND.n828 GND.t840 24.9236
R4598 GND.n977 GND.t782 24.9236
R4599 GND.n977 GND.t808 24.9236
R4600 GND.n981 GND.t844 24.9236
R4601 GND.n981 GND.t898 24.9236
R4602 GND.n987 GND.t868 24.9236
R4603 GND.n987 GND.t786 24.9236
R4604 GND.n993 GND.t838 24.9236
R4605 GND.n993 GND.t874 24.9236
R4606 GND.n999 GND.t790 24.9236
R4607 GND.n999 GND.t820 24.9236
R4608 GND.n934 GND.t800 24.9236
R4609 GND.n934 GND.t836 24.9236
R4610 GND.n941 GND.t828 24.9236
R4611 GND.n941 GND.t862 24.9236
R4612 GND.n963 GND.t890 24.9236
R4613 GND.n963 GND.t810 24.9236
R4614 GND.n959 GND.t866 24.9236
R4615 GND.n959 GND.t784 24.9236
R4616 GND.n953 GND.t814 24.9236
R4617 GND.n953 GND.t850 24.9236
R4618 GND.n947 GND.t902 24.9236
R4619 GND.n947 GND.t796 24.9236
R4620 GND.n822 GND.t892 24.9236
R4621 GND.n822 GND.t906 24.9236
R4622 GND.n850 GND.t802 24.9236
R4623 GND.n850 GND.t858 24.9236
R4624 GND.n893 GND.t884 24.9236
R4625 GND.n893 GND.t806 24.9236
R4626 GND.n900 GND.t842 24.9236
R4627 GND.n900 GND.t896 24.9236
R4628 GND.n904 GND.t794 24.9236
R4629 GND.n904 GND.t846 24.9236
R4630 GND.n910 GND.t834 24.9236
R4631 GND.n910 GND.t872 24.9236
R4632 GND.n916 GND.t788 24.9236
R4633 GND.n916 GND.t818 24.9236
R4634 GND.n922 GND.t854 24.9236
R4635 GND.n922 GND.t908 24.9236
R4636 GND.n835 GND.t870 24.9236
R4637 GND.n835 GND.t860 24.9236
R4638 GND.n840 GND.t886 24.9236
R4639 GND.n840 GND.t830 24.9236
R4640 GND.n883 GND.t864 24.9236
R4641 GND.n883 GND.t888 24.9236
R4642 GND.n878 GND.t812 24.9236
R4643 GND.n878 GND.t848 24.9236
R4644 GND.n872 GND.t900 24.9236
R4645 GND.n872 GND.t816 24.9236
R4646 GND.n866 GND.t852 24.9236
R4647 GND.n866 GND.t904 24.9236
R4648 GND.n860 GND.t798 24.9236
R4649 GND.n860 GND.t792 24.9236
R4650 GND.n1500 GND.t740 24.9236
R4651 GND.n1500 GND.t734 24.9236
R4652 GND.n673 GND.t251 24.9236
R4653 GND.n673 GND.t229 24.9236
R4654 GND.n1460 GND.t243 24.9236
R4655 GND.n1460 GND.t227 24.9236
R4656 GND.n1466 GND.t249 24.9236
R4657 GND.n1466 GND.t221 24.9236
R4658 GND.n1470 GND.t233 24.9236
R4659 GND.n1470 GND.t245 24.9236
R4660 GND.n1476 GND.t223 24.9236
R4661 GND.n1476 GND.t235 24.9236
R4662 GND.n1482 GND.t247 24.9236
R4663 GND.n1482 GND.t225 24.9236
R4664 GND.n1488 GND.t231 24.9236
R4665 GND.n1488 GND.t239 24.9236
R4666 GND.n1403 GND.t215 24.9236
R4667 GND.n1403 GND.t113 24.9236
R4668 GND.n1447 GND.t163 24.9236
R4669 GND.n1447 GND.t199 24.9236
R4670 GND.n1440 GND.t141 24.9236
R4671 GND.n1440 GND.t167 24.9236
R4672 GND.n1436 GND.t203 24.9236
R4673 GND.n1436 GND.t131 24.9236
R4674 GND.n1430 GND.t99 24.9236
R4675 GND.n1430 GND.t145 24.9236
R4676 GND.n1424 GND.t197 24.9236
R4677 GND.n1424 GND.t105 24.9236
R4678 GND.n1418 GND.t149 24.9236
R4679 GND.n1418 GND.t179 24.9236
R4680 GND.n742 GND.t159 24.9236
R4681 GND.n742 GND.t195 24.9236
R4682 GND.n677 GND.t187 24.9236
R4683 GND.n677 GND.t93 24.9236
R4684 GND.n794 GND.t119 24.9236
R4685 GND.n794 GND.t169 24.9236
R4686 GND.n798 GND.t97 24.9236
R4687 GND.n798 GND.t143 24.9236
R4688 GND.n804 GND.t173 24.9236
R4689 GND.n804 GND.t209 24.9236
R4690 GND.n810 GND.t135 24.9236
R4691 GND.n810 GND.t155 24.9236
R4692 GND.n816 GND.t123 24.9236
R4693 GND.n816 GND.t129 24.9236
R4694 GND.n730 GND.t161 24.9236
R4695 GND.n730 GND.t217 24.9236
R4696 GND.n781 GND.t115 24.9236
R4697 GND.n781 GND.t165 24.9236
R4698 GND.n774 GND.t201 24.9236
R4699 GND.n774 GND.t127 24.9236
R4700 GND.n770 GND.t153 24.9236
R4701 GND.n770 GND.t205 24.9236
R4702 GND.n764 GND.t193 24.9236
R4703 GND.n764 GND.t103 24.9236
R4704 GND.n758 GND.t147 24.9236
R4705 GND.n758 GND.t177 24.9236
R4706 GND.n752 GND.t213 24.9236
R4707 GND.n752 GND.t139 24.9236
R4708 GND.n681 GND.t101 24.9236
R4709 GND.n681 GND.t219 24.9236
R4710 GND.n686 GND.t117 24.9236
R4711 GND.n686 GND.t189 24.9236
R4712 GND.n695 GND.t95 24.9236
R4713 GND.n695 GND.t121 24.9236
R4714 GND.n700 GND.t171 24.9236
R4715 GND.n700 GND.t207 24.9236
R4716 GND.n706 GND.t133 24.9236
R4717 GND.n706 GND.t175 24.9236
R4718 GND.n712 GND.t211 24.9236
R4719 GND.n712 GND.t137 24.9236
R4720 GND.n718 GND.t157 24.9236
R4721 GND.n718 GND.t151 24.9236
R4722 GND.n353 GND.t601 24.9236
R4723 GND.n353 GND.t599 24.9236
R4724 GND.n416 GND.t508 24.9236
R4725 GND.n416 GND.t506 24.9236
R4726 GND.n406 GND.t514 24.9236
R4727 GND.n406 GND.t520 24.9236
R4728 GND.n399 GND.t516 24.9236
R4729 GND.n399 GND.t522 24.9236
R4730 GND.n395 GND.t510 24.9236
R4731 GND.n395 GND.t518 24.9236
R4732 GND.n389 GND.t528 24.9236
R4733 GND.n389 GND.t524 24.9236
R4734 GND.n383 GND.t534 24.9236
R4735 GND.n383 GND.t530 24.9236
R4736 GND.n376 GND.t526 24.9236
R4737 GND.n376 GND.t536 24.9236
R4738 GND.n272 GND.t714 24.9236
R4739 GND.n272 GND.t696 24.9236
R4740 GND.n266 GND.t672 24.9236
R4741 GND.n266 GND.t706 24.9236
R4742 GND.n452 GND.t690 24.9236
R4743 GND.n452 GND.t720 24.9236
R4744 GND.n447 GND.t616 24.9236
R4745 GND.n447 GND.t604 24.9236
R4746 GND.n440 GND.t724 24.9236
R4747 GND.n440 GND.t712 24.9236
R4748 GND.n434 GND.t608 24.9236
R4749 GND.n434 GND.t632 24.9236
R4750 GND.n427 GND.t622 24.9236
R4751 GND.n427 GND.t640 24.9236
R4752 GND.n247 GND.t624 24.9236
R4753 GND.n247 GND.t658 24.9236
R4754 GND.n253 GND.t644 24.9236
R4755 GND.n253 GND.t628 24.9236
R4756 GND.n260 GND.t662 24.9236
R4757 GND.n260 GND.t648 24.9236
R4758 GND.n301 GND.t676 24.9236
R4759 GND.n301 GND.t650 24.9236
R4760 GND.n294 GND.t680 24.9236
R4761 GND.n294 GND.t666 24.9236
R4762 GND.n288 GND.t654 24.9236
R4763 GND.n288 GND.t684 24.9236
R4764 GND.n282 GND.t668 24.9236
R4765 GND.n282 GND.t700 24.9236
R4766 GND.n199 GND.t688 24.9236
R4767 GND.n199 GND.t708 24.9236
R4768 GND.n205 GND.t730 24.9236
R4769 GND.n205 GND.t718 24.9236
R4770 GND.n211 GND.t614 24.9236
R4771 GND.n211 GND.t692 24.9236
R4772 GND.n215 GND.t722 24.9236
R4773 GND.n215 GND.t618 24.9236
R4774 GND.n221 GND.t606 24.9236
R4775 GND.n221 GND.t630 24.9236
R4776 GND.n229 GND.t620 24.9236
R4777 GND.n229 GND.t610 24.9236
R4778 GND.n235 GND.t634 24.9236
R4779 GND.n235 GND.t612 24.9236
R4780 GND.n167 GND.t638 24.9236
R4781 GND.n167 GND.t626 24.9236
R4782 GND.n175 GND.t660 24.9236
R4783 GND.n175 GND.t646 24.9236
R4784 GND.n181 GND.t674 24.9236
R4785 GND.n181 GND.t704 24.9236
R4786 GND.n185 GND.t678 24.9236
R4787 GND.n185 GND.t664 24.9236
R4788 GND.n328 GND.t652 24.9236
R4789 GND.n328 GND.t682 24.9236
R4790 GND.n322 GND.t710 24.9236
R4791 GND.n322 GND.t698 24.9236
R4792 GND.n316 GND.t726 24.9236
R4793 GND.n316 GND.t670 24.9236
R4794 GND.n84 GND.n75 24.4711
R4795 GND.n57 GND.n53 24.4711
R4796 GND.n17 GND.n16 24.4711
R4797 GND.n640 GND.n631 24.4711
R4798 GND.n590 GND.n586 24.4711
R4799 GND.n139 GND.n138 24.4711
R4800 GND.n1343 GND.n1342 24.4711
R4801 GND.n1056 GND.n1055 24.4711
R4802 GND.n1496 GND.n1495 24.4711
R4803 GND.n357 GND.n336 24.4711
R4804 GND.n23 GND.n7 23.7181
R4805 GND.n145 GND.n129 23.7181
R4806 GND.n80 GND.n79 22.9652
R4807 GND.n474 GND.n473 22.9652
R4808 GND.n52 GND.n48 22.9652
R4809 GND.n30 GND.n28 22.9652
R4810 GND.n35 GND.n34 22.9652
R4811 GND.n636 GND.n635 22.9652
R4812 GND.n555 GND.n554 22.9652
R4813 GND.n585 GND.n581 22.9652
R4814 GND.n152 GND.n150 22.9652
R4815 GND.n157 GND.n156 22.9652
R4816 GND.n86 GND.t589 22.3257
R4817 GND.n1604 GND.t541 22.3257
R4818 GND.n1606 GND.t585 22.3257
R4819 GND.n54 GND.t780 22.3257
R4820 GND.n45 GND.t595 22.3257
R4821 GND.n13 GND.t263 22.3257
R4822 GND.n642 GND.t545 22.3257
R4823 GND.n610 GND.t452 22.3257
R4824 GND.n612 GND.t489 22.3257
R4825 GND.n587 GND.t483 22.3257
R4826 GND.n578 GND.t774 22.3257
R4827 GND.n135 GND.t558 22.3257
R4828 GND.n22 GND.n10 22.2123
R4829 GND.n18 GND.n10 22.2123
R4830 GND.n144 GND.n132 22.2123
R4831 GND.n140 GND.n132 22.2123
R4832 GND.n95 GND.n93 21.4593
R4833 GND.n110 GND.n108 21.4593
R4834 GND.n112 GND.n105 21.4593
R4835 GND.n481 GND.n479 21.4593
R4836 GND.n483 GND.n466 21.4593
R4837 GND.n31 GND.n30 21.4593
R4838 GND.n34 GND.n33 21.4593
R4839 GND.n651 GND.n649 21.4593
R4840 GND.n662 GND.n660 21.4593
R4841 GND.n664 GND.n657 21.4593
R4842 GND.n562 GND.n560 21.4593
R4843 GND.n564 GND.n547 21.4593
R4844 GND.n153 GND.n152 21.4593
R4845 GND.n156 GND.n155 21.4593
R4846 GND.n80 GND.n75 19.9534
R4847 GND.n475 GND.n474 19.9534
R4848 GND.n53 GND.n52 19.9534
R4849 GND.n28 GND.n3 19.9534
R4850 GND.n36 GND.n35 19.9534
R4851 GND.n636 GND.n631 19.9534
R4852 GND.n556 GND.n555 19.9534
R4853 GND.n586 GND.n585 19.9534
R4854 GND.n150 GND.n125 19.9534
R4855 GND.n158 GND.n157 19.9534
R4856 GND.t564 GND.t88 19.2425
R4857 GND.t2 GND.t398 19.2425
R4858 GND.n1260 GND.t380 17.2168
R4859 GND.n31 GND.n27 16.9417
R4860 GND.n33 GND.n7 16.9417
R4861 GND.n153 GND.n149 16.9417
R4862 GND.n155 GND.n129 16.9417
R4863 GND.n1319 GND.n1318 16.9417
R4864 GND.n1271 GND.n1270 16.9417
R4865 GND.n1249 GND.n1248 16.9417
R4866 GND.n1190 GND.n1189 16.9417
R4867 GND.n1164 GND.n1163 16.9417
R4868 GND.n1032 GND.n1031 16.9417
R4869 GND.n983 GND.n982 16.9417
R4870 GND.n961 GND.n960 16.9417
R4871 GND.n906 GND.n905 16.9417
R4872 GND.n880 GND.n879 16.9417
R4873 GND.n1472 GND.n1471 16.9417
R4874 GND.n1438 GND.n1437 16.9417
R4875 GND.n800 GND.n799 16.9417
R4876 GND.n772 GND.n771 16.9417
R4877 GND.n702 GND.n701 16.9417
R4878 GND.n397 GND.n396 16.9417
R4879 GND.n449 GND.n448 16.9417
R4880 GND.n303 GND.n302 16.9417
R4881 GND.n217 GND.n216 16.9417
R4882 GND.n187 GND.n186 16.9417
R4883 GND.n18 GND.n17 16.1887
R4884 GND.n140 GND.n139 16.1887
R4885 GND.t451 GND.t488 14.6672
R4886 GND.t45 GND.t778 14.6672
R4887 GND.t572 GND.t568 14.6672
R4888 GND.t584 GND.t540 14.6672
R4889 GND.t502 GND.t60 14.6672
R4890 GND.t58 GND.t504 14.6672
R4891 GND.n1376 GND.n1352 14.5711
R4892 GND.n1089 GND.n1065 14.5711
R4893 GND.n1529 GND.n1505 14.5711
R4894 GND.n972 GND.t861 14.2308
R4895 GND.n1608 GND.n1605 13.5727
R4896 GND.n614 GND.n611 13.5727
R4897 GND.n1608 GND.n1607 13.5705
R4898 GND.n614 GND.n613 13.5705
R4899 GND.n60 GND.n59 13.5646
R4900 GND.n593 GND.n592 13.5646
R4901 GND.t629 GND.n308 13.4015
R4902 GND.n1315 GND.n1314 11.6711
R4903 GND.n1267 GND.n1266 11.6711
R4904 GND.n1253 GND.n1252 11.6711
R4905 GND.n1186 GND.n1185 11.6711
R4906 GND.n1169 GND.n1168 11.6711
R4907 GND.n1028 GND.n1027 11.6711
R4908 GND.n979 GND.n978 11.6711
R4909 GND.n965 GND.n964 11.6711
R4910 GND.n902 GND.n901 11.6711
R4911 GND.n885 GND.n884 11.6711
R4912 GND.n1468 GND.n1467 11.6711
R4913 GND.n1442 GND.n1441 11.6711
R4914 GND.n796 GND.n795 11.6711
R4915 GND.n776 GND.n775 11.6711
R4916 GND.n697 GND.n696 11.6711
R4917 GND.n401 GND.n400 11.6711
R4918 GND.n454 GND.n453 11.6711
R4919 GND.n262 GND.n261 11.6711
R4920 GND.n213 GND.n212 11.6711
R4921 GND.n183 GND.n182 11.6711
R4922 GND.n1453 GND.t162 11.4291
R4923 GND.n1562 GND.n1561 11.427
R4924 GND.n343 GND.n342 11.427
R4925 GND.n341 GND.n340 11.427
R4926 GND.n500 GND.n499 11.427
R4927 GND.n1325 GND.n1324 10.9181
R4928 GND.n1277 GND.n1276 10.9181
R4929 GND.n1243 GND.n1242 10.9181
R4930 GND.n1196 GND.n1195 10.9181
R4931 GND.n1158 GND.n1157 10.9181
R4932 GND.n1038 GND.n1037 10.9181
R4933 GND.n989 GND.n988 10.9181
R4934 GND.n955 GND.n954 10.9181
R4935 GND.n912 GND.n911 10.9181
R4936 GND.n874 GND.n873 10.9181
R4937 GND.n1478 GND.n1477 10.9181
R4938 GND.n1432 GND.n1431 10.9181
R4939 GND.n806 GND.n805 10.9181
R4940 GND.n766 GND.n765 10.9181
R4941 GND.n708 GND.n707 10.9181
R4942 GND.n391 GND.n390 10.9181
R4943 GND.n442 GND.n441 10.9181
R4944 GND.n296 GND.n295 10.9181
R4945 GND.n223 GND.n222 10.9181
R4946 GND.n330 GND.n329 10.9181
R4947 GND.n344 GND.n343 10.5417
R4948 GND.n87 GND.n85 9.41227
R4949 GND.n56 GND.n55 9.41227
R4950 GND.n643 GND.n641 9.41227
R4951 GND.n589 GND.n588 9.41227
R4952 GND.n1379 GND.t306 7.37892
R4953 GND.n1585 GND.n1557 6.77697
R4954 GND.n1579 GND.n1558 6.77697
R4955 GND.n1573 GND.n1559 6.77697
R4956 GND.n1567 GND.n1560 6.77697
R4957 GND.n1368 GND.n1355 6.77697
R4958 GND.n1081 GND.n1068 6.77697
R4959 GND.n1521 GND.n1508 6.77697
R4960 GND.n523 GND.n495 6.77697
R4961 GND.n517 GND.n496 6.77697
R4962 GND.n511 GND.n497 6.77697
R4963 GND.n505 GND.n498 6.77697
R4964 GND.n309 GND.t701 6.70101
R4965 GND.n88 GND.n87 6.4005
R4966 GND.n1610 GND.n1605 6.4005
R4967 GND.n1607 GND.n1602 6.4005
R4968 GND.n55 GND.n43 6.4005
R4969 GND.n61 GND.n60 6.4005
R4970 GND.n644 GND.n643 6.4005
R4971 GND.n616 GND.n611 6.4005
R4972 GND.n613 GND.n608 6.4005
R4973 GND.n588 GND.n576 6.4005
R4974 GND.n594 GND.n593 6.4005
R4975 GND.n1357 GND.n1356 6.15638
R4976 GND.n1070 GND.n1069 6.15638
R4977 GND.n1510 GND.n1509 6.15638
R4978 GND.n1309 GND.n1308 5.64756
R4979 GND.n1115 GND.n1114 5.64756
R4980 GND.n1227 GND.n1226 5.64756
R4981 GND.n1179 GND.n1178 5.64756
R4982 GND.n1127 GND.n1126 5.64756
R4983 GND.n1022 GND.n1021 5.64756
R4984 GND.n830 GND.n829 5.64756
R4985 GND.n943 GND.n942 5.64756
R4986 GND.n895 GND.n894 5.64756
R4987 GND.n842 GND.n841 5.64756
R4988 GND.n1462 GND.n1461 5.64756
R4989 GND.n1449 GND.n1448 5.64756
R4990 GND.n679 GND.n678 5.64756
R4991 GND.n783 GND.n782 5.64756
R4992 GND.n688 GND.n687 5.64756
R4993 GND.n408 GND.n407 5.64756
R4994 GND.n268 GND.n267 5.64756
R4995 GND.n255 GND.n254 5.64756
R4996 GND.n207 GND.n206 5.64756
R4997 GND.n177 GND.n176 5.64756
R4998 GND.n1331 GND.n1330 4.89462
R4999 GND.n1283 GND.n1282 4.89462
R5000 GND.n1237 GND.n1236 4.89462
R5001 GND.n1202 GND.n1201 4.89462
R5002 GND.n1152 GND.n1151 4.89462
R5003 GND.n1044 GND.n1043 4.89462
R5004 GND.n995 GND.n994 4.89462
R5005 GND.n949 GND.n948 4.89462
R5006 GND.n918 GND.n917 4.89462
R5007 GND.n868 GND.n867 4.89462
R5008 GND.n1484 GND.n1483 4.89462
R5009 GND.n1426 GND.n1425 4.89462
R5010 GND.n812 GND.n811 4.89462
R5011 GND.n760 GND.n759 4.89462
R5012 GND.n714 GND.n713 4.89462
R5013 GND.n385 GND.n384 4.89462
R5014 GND.n436 GND.n435 4.89462
R5015 GND.n290 GND.n289 4.89462
R5016 GND.n231 GND.n230 4.89462
R5017 GND.n324 GND.n323 4.89462
R5018 GND.n1564 GND.n1563 4.6505
R5019 GND.n1566 GND.n1565 4.6505
R5020 GND.n1568 GND.n1567 4.6505
R5021 GND.n1570 GND.n1569 4.6505
R5022 GND.n1572 GND.n1571 4.6505
R5023 GND.n1574 GND.n1573 4.6505
R5024 GND.n1576 GND.n1575 4.6505
R5025 GND.n1578 GND.n1577 4.6505
R5026 GND.n1580 GND.n1579 4.6505
R5027 GND.n1582 GND.n1581 4.6505
R5028 GND.n1584 GND.n1583 4.6505
R5029 GND.n1586 GND.n1585 4.6505
R5030 GND.n82 GND.n75 4.6505
R5031 GND.n93 GND.n72 4.6505
R5032 GND.n92 GND.n91 4.6505
R5033 GND.n90 GND.n73 4.6505
R5034 GND.n89 GND.n88 4.6505
R5035 GND.n85 GND.n74 4.6505
R5036 GND.n84 GND.n83 4.6505
R5037 GND.n81 GND.n80 4.6505
R5038 GND.n115 GND.n114 4.6505
R5039 GND.n113 GND.n103 4.6505
R5040 GND.n112 GND.n111 4.6505
R5041 GND.n111 GND.n110 4.6505
R5042 GND.n109 GND.n103 4.6505
R5043 GND.n115 GND.n102 4.6505
R5044 GND.n117 GND.n116 4.6505
R5045 GND.n474 GND.n469 4.6505
R5046 GND.n476 GND.n475 4.6505
R5047 GND.n483 GND.n482 4.6505
R5048 GND.n484 GND.n464 4.6505
R5049 GND.n486 GND.n485 4.6505
R5050 GND.n479 GND.n467 4.6505
R5051 GND.n482 GND.n481 4.6505
R5052 GND.n480 GND.n464 4.6505
R5053 GND.n486 GND.n463 4.6505
R5054 GND.n488 GND.n487 4.6505
R5055 GND.n1603 GND.n1602 4.6505
R5056 GND.n1614 GND.n1613 4.6505
R5057 GND.n1610 GND.n1609 4.6505
R5058 GND.n1612 GND.n1611 4.6505
R5059 GND.n62 GND.n61 4.6505
R5060 GND.n53 GND.n46 4.6505
R5061 GND.n52 GND.n51 4.6505
R5062 GND.n58 GND.n57 4.6505
R5063 GND.n56 GND.n44 4.6505
R5064 GND.n62 GND.n43 4.6505
R5065 GND.n64 GND.n63 4.6505
R5066 GND.n17 GND.n11 4.6505
R5067 GND.n20 GND.n10 4.6505
R5068 GND.n8 GND.n7 4.6505
R5069 GND.n34 GND.n5 4.6505
R5070 GND.n16 GND.n15 4.6505
R5071 GND.n19 GND.n18 4.6505
R5072 GND.n22 GND.n21 4.6505
R5073 GND.n24 GND.n23 4.6505
R5074 GND.n33 GND.n32 4.6505
R5075 GND.n35 GND.n2 4.6505
R5076 GND.n37 GND.n36 4.6505
R5077 GND.n30 GND.n5 4.6505
R5078 GND.n32 GND.n31 4.6505
R5079 GND.n28 GND.n2 4.6505
R5080 GND.n37 GND.n3 4.6505
R5081 GND.n638 GND.n631 4.6505
R5082 GND.n649 GND.n628 4.6505
R5083 GND.n648 GND.n647 4.6505
R5084 GND.n646 GND.n629 4.6505
R5085 GND.n645 GND.n644 4.6505
R5086 GND.n641 GND.n630 4.6505
R5087 GND.n640 GND.n639 4.6505
R5088 GND.n637 GND.n636 4.6505
R5089 GND.n667 GND.n666 4.6505
R5090 GND.n665 GND.n655 4.6505
R5091 GND.n664 GND.n663 4.6505
R5092 GND.n663 GND.n662 4.6505
R5093 GND.n661 GND.n655 4.6505
R5094 GND.n667 GND.n654 4.6505
R5095 GND.n669 GND.n668 4.6505
R5096 GND.n555 GND.n550 4.6505
R5097 GND.n557 GND.n556 4.6505
R5098 GND.n564 GND.n563 4.6505
R5099 GND.n565 GND.n545 4.6505
R5100 GND.n567 GND.n566 4.6505
R5101 GND.n560 GND.n548 4.6505
R5102 GND.n563 GND.n562 4.6505
R5103 GND.n561 GND.n545 4.6505
R5104 GND.n567 GND.n544 4.6505
R5105 GND.n569 GND.n568 4.6505
R5106 GND.n609 GND.n608 4.6505
R5107 GND.n620 GND.n619 4.6505
R5108 GND.n616 GND.n615 4.6505
R5109 GND.n618 GND.n617 4.6505
R5110 GND.n595 GND.n594 4.6505
R5111 GND.n586 GND.n579 4.6505
R5112 GND.n585 GND.n584 4.6505
R5113 GND.n591 GND.n590 4.6505
R5114 GND.n589 GND.n577 4.6505
R5115 GND.n595 GND.n576 4.6505
R5116 GND.n597 GND.n596 4.6505
R5117 GND.n139 GND.n133 4.6505
R5118 GND.n142 GND.n132 4.6505
R5119 GND.n130 GND.n129 4.6505
R5120 GND.n156 GND.n127 4.6505
R5121 GND.n138 GND.n137 4.6505
R5122 GND.n141 GND.n140 4.6505
R5123 GND.n144 GND.n143 4.6505
R5124 GND.n146 GND.n145 4.6505
R5125 GND.n155 GND.n154 4.6505
R5126 GND.n157 GND.n124 4.6505
R5127 GND.n159 GND.n158 4.6505
R5128 GND.n152 GND.n127 4.6505
R5129 GND.n154 GND.n153 4.6505
R5130 GND.n150 GND.n124 4.6505
R5131 GND.n159 GND.n125 4.6505
R5132 GND.n1141 GND.n1131 4.6505
R5133 GND.n1140 GND.n1132 4.6505
R5134 GND.n1213 GND.n1212 4.6505
R5135 GND.n1215 GND.n1214 4.6505
R5136 GND.n1392 GND.n1111 4.6505
R5137 GND.n1391 GND.n1112 4.6505
R5138 GND.n1294 GND.n1293 4.6505
R5139 GND.n1296 GND.n1295 4.6505
R5140 GND.n1342 GND.n1341 4.6505
R5141 GND.n1344 GND.n1343 4.6505
R5142 GND.n1354 GND.n1353 4.6505
R5143 GND.n1124 GND.n1123 4.6505
R5144 GND.n1128 GND.n1127 4.6505
R5145 GND.n1130 GND.n1129 4.6505
R5146 GND.n1170 GND.n1169 4.6505
R5147 GND.n1165 GND.n1164 4.6505
R5148 GND.n1161 GND.n1160 4.6505
R5149 GND.n1159 GND.n1158 4.6505
R5150 GND.n1155 GND.n1154 4.6505
R5151 GND.n1153 GND.n1152 4.6505
R5152 GND.n1149 GND.n1148 4.6505
R5153 GND.n1147 GND.n1146 4.6505
R5154 GND.n1143 GND.n1142 4.6505
R5155 GND.n1139 GND.n1138 4.6505
R5156 GND.n1137 GND.n1136 4.6505
R5157 GND.n1118 GND.n1117 4.6505
R5158 GND.n1180 GND.n1179 4.6505
R5159 GND.n1183 GND.n1182 4.6505
R5160 GND.n1187 GND.n1186 4.6505
R5161 GND.n1191 GND.n1190 4.6505
R5162 GND.n1193 GND.n1192 4.6505
R5163 GND.n1197 GND.n1196 4.6505
R5164 GND.n1199 GND.n1198 4.6505
R5165 GND.n1203 GND.n1202 4.6505
R5166 GND.n1205 GND.n1204 4.6505
R5167 GND.n1209 GND.n1208 4.6505
R5168 GND.n1211 GND.n1210 4.6505
R5169 GND.n1217 GND.n1216 4.6505
R5170 GND.n1221 GND.n1220 4.6505
R5171 GND.n1223 GND.n1222 4.6505
R5172 GND.n1228 GND.n1227 4.6505
R5173 GND.n1257 GND.n1256 4.6505
R5174 GND.n1254 GND.n1253 4.6505
R5175 GND.n1250 GND.n1249 4.6505
R5176 GND.n1246 GND.n1245 4.6505
R5177 GND.n1244 GND.n1243 4.6505
R5178 GND.n1240 GND.n1239 4.6505
R5179 GND.n1238 GND.n1237 4.6505
R5180 GND.n1234 GND.n1233 4.6505
R5181 GND.n1232 GND.n1231 4.6505
R5182 GND.n1110 GND.n1109 4.6505
R5183 GND.n1390 GND.n1389 4.6505
R5184 GND.n1388 GND.n1387 4.6505
R5185 GND.n1383 GND.n1382 4.6505
R5186 GND.n1116 GND.n1115 4.6505
R5187 GND.n1264 GND.n1263 4.6505
R5188 GND.n1268 GND.n1267 4.6505
R5189 GND.n1272 GND.n1271 4.6505
R5190 GND.n1274 GND.n1273 4.6505
R5191 GND.n1278 GND.n1277 4.6505
R5192 GND.n1280 GND.n1279 4.6505
R5193 GND.n1284 GND.n1283 4.6505
R5194 GND.n1286 GND.n1285 4.6505
R5195 GND.n1290 GND.n1289 4.6505
R5196 GND.n1292 GND.n1291 4.6505
R5197 GND.n1298 GND.n1297 4.6505
R5198 GND.n1302 GND.n1301 4.6505
R5199 GND.n1305 GND.n1304 4.6505
R5200 GND.n1310 GND.n1309 4.6505
R5201 GND.n1312 GND.n1311 4.6505
R5202 GND.n1316 GND.n1315 4.6505
R5203 GND.n1320 GND.n1319 4.6505
R5204 GND.n1322 GND.n1321 4.6505
R5205 GND.n1326 GND.n1325 4.6505
R5206 GND.n1328 GND.n1327 4.6505
R5207 GND.n1332 GND.n1331 4.6505
R5208 GND.n1334 GND.n1333 4.6505
R5209 GND.n1338 GND.n1337 4.6505
R5210 GND.n1340 GND.n1339 4.6505
R5211 GND.n1346 GND.n1345 4.6505
R5212 GND.n1349 GND.n1348 4.6505
R5213 GND.n1351 GND.n1350 4.6505
R5214 GND.n1374 GND.n1373 4.6505
R5215 GND.n1371 GND.n1370 4.6505
R5216 GND.n1369 GND.n1368 4.6505
R5217 GND.n1367 GND.n1366 4.6505
R5218 GND.n1365 GND.n1364 4.6505
R5219 GND.n1363 GND.n1362 4.6505
R5220 GND.n1359 GND.n1358 4.6505
R5221 GND.n857 GND.n847 4.6505
R5222 GND.n856 GND.n848 4.6505
R5223 GND.n929 GND.n928 4.6505
R5224 GND.n931 GND.n930 4.6505
R5225 GND.n1105 GND.n826 4.6505
R5226 GND.n1104 GND.n827 4.6505
R5227 GND.n1006 GND.n1005 4.6505
R5228 GND.n1008 GND.n1007 4.6505
R5229 GND.n1055 GND.n1054 4.6505
R5230 GND.n1057 GND.n1056 4.6505
R5231 GND.n1067 GND.n1066 4.6505
R5232 GND.n839 GND.n838 4.6505
R5233 GND.n843 GND.n842 4.6505
R5234 GND.n846 GND.n845 4.6505
R5235 GND.n886 GND.n885 4.6505
R5236 GND.n881 GND.n880 4.6505
R5237 GND.n877 GND.n876 4.6505
R5238 GND.n875 GND.n874 4.6505
R5239 GND.n871 GND.n870 4.6505
R5240 GND.n869 GND.n868 4.6505
R5241 GND.n865 GND.n864 4.6505
R5242 GND.n863 GND.n862 4.6505
R5243 GND.n859 GND.n858 4.6505
R5244 GND.n855 GND.n854 4.6505
R5245 GND.n853 GND.n852 4.6505
R5246 GND.n833 GND.n832 4.6505
R5247 GND.n896 GND.n895 4.6505
R5248 GND.n899 GND.n898 4.6505
R5249 GND.n903 GND.n902 4.6505
R5250 GND.n907 GND.n906 4.6505
R5251 GND.n909 GND.n908 4.6505
R5252 GND.n913 GND.n912 4.6505
R5253 GND.n915 GND.n914 4.6505
R5254 GND.n919 GND.n918 4.6505
R5255 GND.n921 GND.n920 4.6505
R5256 GND.n925 GND.n924 4.6505
R5257 GND.n927 GND.n926 4.6505
R5258 GND.n933 GND.n932 4.6505
R5259 GND.n937 GND.n936 4.6505
R5260 GND.n939 GND.n938 4.6505
R5261 GND.n944 GND.n943 4.6505
R5262 GND.n969 GND.n968 4.6505
R5263 GND.n966 GND.n965 4.6505
R5264 GND.n962 GND.n961 4.6505
R5265 GND.n958 GND.n957 4.6505
R5266 GND.n956 GND.n955 4.6505
R5267 GND.n952 GND.n951 4.6505
R5268 GND.n950 GND.n949 4.6505
R5269 GND.n946 GND.n945 4.6505
R5270 GND.n825 GND.n824 4.6505
R5271 GND.n1107 GND.n1106 4.6505
R5272 GND.n1103 GND.n1102 4.6505
R5273 GND.n1101 GND.n1100 4.6505
R5274 GND.n1096 GND.n1095 4.6505
R5275 GND.n831 GND.n830 4.6505
R5276 GND.n976 GND.n975 4.6505
R5277 GND.n980 GND.n979 4.6505
R5278 GND.n984 GND.n983 4.6505
R5279 GND.n986 GND.n985 4.6505
R5280 GND.n990 GND.n989 4.6505
R5281 GND.n992 GND.n991 4.6505
R5282 GND.n996 GND.n995 4.6505
R5283 GND.n998 GND.n997 4.6505
R5284 GND.n1002 GND.n1001 4.6505
R5285 GND.n1004 GND.n1003 4.6505
R5286 GND.n1010 GND.n1009 4.6505
R5287 GND.n1015 GND.n1014 4.6505
R5288 GND.n1018 GND.n1017 4.6505
R5289 GND.n1023 GND.n1022 4.6505
R5290 GND.n1025 GND.n1024 4.6505
R5291 GND.n1029 GND.n1028 4.6505
R5292 GND.n1033 GND.n1032 4.6505
R5293 GND.n1035 GND.n1034 4.6505
R5294 GND.n1039 GND.n1038 4.6505
R5295 GND.n1041 GND.n1040 4.6505
R5296 GND.n1045 GND.n1044 4.6505
R5297 GND.n1047 GND.n1046 4.6505
R5298 GND.n1051 GND.n1050 4.6505
R5299 GND.n1053 GND.n1052 4.6505
R5300 GND.n1059 GND.n1058 4.6505
R5301 GND.n1062 GND.n1061 4.6505
R5302 GND.n1064 GND.n1063 4.6505
R5303 GND.n1087 GND.n1086 4.6505
R5304 GND.n1084 GND.n1083 4.6505
R5305 GND.n1082 GND.n1081 4.6505
R5306 GND.n1080 GND.n1079 4.6505
R5307 GND.n1078 GND.n1077 4.6505
R5308 GND.n1076 GND.n1075 4.6505
R5309 GND.n1072 GND.n1071 4.6505
R5310 GND.n725 GND.n724 4.6505
R5311 GND.n727 GND.n726 4.6505
R5312 GND.n749 GND.n737 4.6505
R5313 GND.n748 GND.n738 4.6505
R5314 GND.n1398 GND.n1397 4.6505
R5315 GND.n1400 GND.n1399 4.6505
R5316 GND.n1415 GND.n1410 4.6505
R5317 GND.n1414 GND.n1411 4.6505
R5318 GND.n1495 GND.n1494 4.6505
R5319 GND.n1497 GND.n1496 4.6505
R5320 GND.n1507 GND.n1506 4.6505
R5321 GND.n685 GND.n684 4.6505
R5322 GND.n689 GND.n688 4.6505
R5323 GND.n691 GND.n690 4.6505
R5324 GND.n698 GND.n697 4.6505
R5325 GND.n703 GND.n702 4.6505
R5326 GND.n705 GND.n704 4.6505
R5327 GND.n709 GND.n708 4.6505
R5328 GND.n711 GND.n710 4.6505
R5329 GND.n715 GND.n714 4.6505
R5330 GND.n717 GND.n716 4.6505
R5331 GND.n721 GND.n720 4.6505
R5332 GND.n723 GND.n722 4.6505
R5333 GND.n729 GND.n728 4.6505
R5334 GND.n733 GND.n732 4.6505
R5335 GND.n736 GND.n735 4.6505
R5336 GND.n784 GND.n783 4.6505
R5337 GND.n779 GND.n778 4.6505
R5338 GND.n777 GND.n776 4.6505
R5339 GND.n773 GND.n772 4.6505
R5340 GND.n769 GND.n768 4.6505
R5341 GND.n767 GND.n766 4.6505
R5342 GND.n763 GND.n762 4.6505
R5343 GND.n761 GND.n760 4.6505
R5344 GND.n757 GND.n756 4.6505
R5345 GND.n755 GND.n754 4.6505
R5346 GND.n751 GND.n750 4.6505
R5347 GND.n747 GND.n746 4.6505
R5348 GND.n745 GND.n744 4.6505
R5349 GND.n741 GND.n740 4.6505
R5350 GND.n680 GND.n679 4.6505
R5351 GND.n792 GND.n791 4.6505
R5352 GND.n797 GND.n796 4.6505
R5353 GND.n801 GND.n800 4.6505
R5354 GND.n803 GND.n802 4.6505
R5355 GND.n807 GND.n806 4.6505
R5356 GND.n809 GND.n808 4.6505
R5357 GND.n813 GND.n812 4.6505
R5358 GND.n815 GND.n814 4.6505
R5359 GND.n819 GND.n818 4.6505
R5360 GND.n821 GND.n820 4.6505
R5361 GND.n1402 GND.n1401 4.6505
R5362 GND.n1406 GND.n1405 4.6505
R5363 GND.n1409 GND.n1408 4.6505
R5364 GND.n1450 GND.n1449 4.6505
R5365 GND.n1445 GND.n1444 4.6505
R5366 GND.n1443 GND.n1442 4.6505
R5367 GND.n1439 GND.n1438 4.6505
R5368 GND.n1435 GND.n1434 4.6505
R5369 GND.n1433 GND.n1432 4.6505
R5370 GND.n1429 GND.n1428 4.6505
R5371 GND.n1427 GND.n1426 4.6505
R5372 GND.n1423 GND.n1422 4.6505
R5373 GND.n1421 GND.n1420 4.6505
R5374 GND.n1417 GND.n1416 4.6505
R5375 GND.n1413 GND.n1412 4.6505
R5376 GND.n676 GND.n675 4.6505
R5377 GND.n1458 GND.n1457 4.6505
R5378 GND.n1463 GND.n1462 4.6505
R5379 GND.n1465 GND.n1464 4.6505
R5380 GND.n1469 GND.n1468 4.6505
R5381 GND.n1473 GND.n1472 4.6505
R5382 GND.n1475 GND.n1474 4.6505
R5383 GND.n1479 GND.n1478 4.6505
R5384 GND.n1481 GND.n1480 4.6505
R5385 GND.n1485 GND.n1484 4.6505
R5386 GND.n1487 GND.n1486 4.6505
R5387 GND.n1491 GND.n1490 4.6505
R5388 GND.n1493 GND.n1492 4.6505
R5389 GND.n1499 GND.n1498 4.6505
R5390 GND.n1502 GND.n1501 4.6505
R5391 GND.n1504 GND.n1503 4.6505
R5392 GND.n1527 GND.n1526 4.6505
R5393 GND.n1524 GND.n1523 4.6505
R5394 GND.n1522 GND.n1521 4.6505
R5395 GND.n1520 GND.n1519 4.6505
R5396 GND.n1518 GND.n1517 4.6505
R5397 GND.n1516 GND.n1515 4.6505
R5398 GND.n1512 GND.n1511 4.6505
R5399 GND.n346 GND.n339 4.6505
R5400 GND.n356 GND.n337 4.6505
R5401 GND.n350 GND.n338 4.6505
R5402 GND.n355 GND.n354 4.6505
R5403 GND.n352 GND.n351 4.6505
R5404 GND.n348 GND.n347 4.6505
R5405 GND.n345 GND.n344 4.6505
R5406 GND.n358 GND.n357 4.6505
R5407 GND.n170 GND.n169 4.6505
R5408 GND.n173 GND.n172 4.6505
R5409 GND.n178 GND.n177 4.6505
R5410 GND.n180 GND.n179 4.6505
R5411 GND.n184 GND.n183 4.6505
R5412 GND.n188 GND.n187 4.6505
R5413 GND.n190 GND.n189 4.6505
R5414 GND.n331 GND.n330 4.6505
R5415 GND.n327 GND.n326 4.6505
R5416 GND.n325 GND.n324 4.6505
R5417 GND.n321 GND.n320 4.6505
R5418 GND.n319 GND.n318 4.6505
R5419 GND.n194 GND.n191 4.6505
R5420 GND.n196 GND.n195 4.6505
R5421 GND.n242 GND.n241 4.6505
R5422 GND.n244 GND.n243 4.6505
R5423 GND.n279 GND.n264 4.6505
R5424 GND.n278 GND.n265 4.6505
R5425 GND.n313 GND.n312 4.6505
R5426 GND.n198 GND.n197 4.6505
R5427 GND.n202 GND.n201 4.6505
R5428 GND.n204 GND.n203 4.6505
R5429 GND.n208 GND.n207 4.6505
R5430 GND.n210 GND.n209 4.6505
R5431 GND.n214 GND.n213 4.6505
R5432 GND.n218 GND.n217 4.6505
R5433 GND.n220 GND.n219 4.6505
R5434 GND.n224 GND.n223 4.6505
R5435 GND.n227 GND.n226 4.6505
R5436 GND.n232 GND.n231 4.6505
R5437 GND.n234 GND.n233 4.6505
R5438 GND.n238 GND.n237 4.6505
R5439 GND.n240 GND.n239 4.6505
R5440 GND.n246 GND.n245 4.6505
R5441 GND.n250 GND.n249 4.6505
R5442 GND.n252 GND.n251 4.6505
R5443 GND.n256 GND.n255 4.6505
R5444 GND.n258 GND.n257 4.6505
R5445 GND.n263 GND.n262 4.6505
R5446 GND.n304 GND.n303 4.6505
R5447 GND.n299 GND.n298 4.6505
R5448 GND.n297 GND.n296 4.6505
R5449 GND.n293 GND.n292 4.6505
R5450 GND.n291 GND.n290 4.6505
R5451 GND.n287 GND.n286 4.6505
R5452 GND.n285 GND.n284 4.6505
R5453 GND.n281 GND.n280 4.6505
R5454 GND.n277 GND.n276 4.6505
R5455 GND.n275 GND.n274 4.6505
R5456 GND.n271 GND.n270 4.6505
R5457 GND.n269 GND.n268 4.6505
R5458 GND.n162 GND.n161 4.6505
R5459 GND.n455 GND.n454 4.6505
R5460 GND.n450 GND.n449 4.6505
R5461 GND.n445 GND.n444 4.6505
R5462 GND.n443 GND.n442 4.6505
R5463 GND.n439 GND.n438 4.6505
R5464 GND.n437 GND.n436 4.6505
R5465 GND.n432 GND.n431 4.6505
R5466 GND.n430 GND.n429 4.6505
R5467 GND.n426 GND.n425 4.6505
R5468 GND.n423 GND.n334 4.6505
R5469 GND.n422 GND.n335 4.6505
R5470 GND.n360 GND.n336 4.6505
R5471 GND.n421 GND.n420 4.6505
R5472 GND.n419 GND.n418 4.6505
R5473 GND.n414 GND.n413 4.6505
R5474 GND.n409 GND.n408 4.6505
R5475 GND.n404 GND.n403 4.6505
R5476 GND.n402 GND.n401 4.6505
R5477 GND.n398 GND.n397 4.6505
R5478 GND.n394 GND.n393 4.6505
R5479 GND.n392 GND.n391 4.6505
R5480 GND.n388 GND.n387 4.6505
R5481 GND.n386 GND.n385 4.6505
R5482 GND.n382 GND.n381 4.6505
R5483 GND.n379 GND.n378 4.6505
R5484 GND.n363 GND.n362 4.6505
R5485 GND.n502 GND.n501 4.6505
R5486 GND.n504 GND.n503 4.6505
R5487 GND.n506 GND.n505 4.6505
R5488 GND.n508 GND.n507 4.6505
R5489 GND.n510 GND.n509 4.6505
R5490 GND.n512 GND.n511 4.6505
R5491 GND.n514 GND.n513 4.6505
R5492 GND.n516 GND.n515 4.6505
R5493 GND.n518 GND.n517 4.6505
R5494 GND.n520 GND.n519 4.6505
R5495 GND.n522 GND.n521 4.6505
R5496 GND.n524 GND.n523 4.6505
R5497 GND.n1122 GND.n1121 4.45136
R5498 GND.n837 GND.n836 4.45136
R5499 GND.n683 GND.n682 4.45136
R5500 GND.n372 GND.n371 4.25025
R5501 GND.n96 GND.n95 4.06709
R5502 GND.n652 GND.n651 4.06709
R5503 GND.n106 GND.n105 4.06409
R5504 GND.n658 GND.n657 4.06409
R5505 GND.n108 GND.n106 4.0631
R5506 GND.n660 GND.n658 4.0631
R5507 GND.n477 GND.n466 4.05611
R5508 GND.n558 GND.n547 4.05611
R5509 GND.n27 GND.n25 3.98881
R5510 GND.n149 GND.n147 3.98881
R5511 GND.n473 GND.n472 3.80559
R5512 GND.n50 GND.n48 3.80559
R5513 GND.n554 GND.n553 3.80559
R5514 GND.n583 GND.n581 3.80559
R5515 GND.n79 GND.n77 3.80083
R5516 GND.n635 GND.n633 3.80083
R5517 GND.n1092 GND.t803 2.84655
R5518 GND.n1362 GND.n1361 2.25932
R5519 GND.n1075 GND.n1074 2.25932
R5520 GND.n1515 GND.n1514 2.25932
R5521 GND.n1337 GND.n1336 1.12991
R5522 GND.n1289 GND.n1288 1.12991
R5523 GND.n1231 GND.n1230 1.12991
R5524 GND.n1208 GND.n1207 1.12991
R5525 GND.n1146 GND.n1145 1.12991
R5526 GND.n1050 GND.n1049 1.12991
R5527 GND.n1001 GND.n1000 1.12991
R5528 GND.n824 GND.n823 1.12991
R5529 GND.n924 GND.n923 1.12991
R5530 GND.n862 GND.n861 1.12991
R5531 GND.n1490 GND.n1489 1.12991
R5532 GND.n1420 GND.n1419 1.12991
R5533 GND.n818 GND.n817 1.12991
R5534 GND.n754 GND.n753 1.12991
R5535 GND.n720 GND.n719 1.12991
R5536 GND.n378 GND.n377 1.12991
R5537 GND.n429 GND.n428 1.12991
R5538 GND.n284 GND.n283 1.12991
R5539 GND.n237 GND.n236 1.12991
R5540 GND.n318 GND.n317 1.12991
R5541 GND.n1396 GND.n1395 0.735503
R5542 GND.n166 GND.n165 0.705542
R5543 GND.n333 GND.n332 0.53211
R5544 GND.n1394 GND.n1393 0.48654
R5545 GND.n1395 GND.n1108 0.479239
R5546 GND.n1592 GND.n97 0.411604
R5547 GND.n1537 GND.n1536 0.411604
R5548 GND.n1301 GND.n1300 0.376971
R5549 GND.n1387 GND.n1386 0.376971
R5550 GND.n1220 GND.n1219 0.376971
R5551 GND.n1136 GND.n1135 0.376971
R5552 GND.n1014 GND.n1013 0.376971
R5553 GND.n1100 GND.n1099 0.376971
R5554 GND.n936 GND.n935 0.376971
R5555 GND.n852 GND.n851 0.376971
R5556 GND.n675 GND.n674 0.376971
R5557 GND.n1405 GND.n1404 0.376971
R5558 GND.n744 GND.n743 0.376971
R5559 GND.n732 GND.n731 0.376971
R5560 GND.n418 GND.n417 0.376971
R5561 GND.n274 GND.n273 0.376971
R5562 GND.n249 GND.n248 0.376971
R5563 GND.n201 GND.n200 0.376971
R5564 GND.n169 GND.n168 0.376971
R5565 GND.n1593 GND.n71 0.375505
R5566 GND.n1538 GND.n627 0.375505
R5567 GND.n1594 GND.n69 0.33677
R5568 GND.n1540 GND.n1539 0.33677
R5569 GND.n1394 GND.n0 0.336652
R5570 GND.n1588 GND 0.327423
R5571 GND.n526 GND 0.327423
R5572 GND.n1620 GND.n66 0.326891
R5573 GND.n600 GND.n599 0.326891
R5574 GND.n1621 GND.n40 0.325812
R5575 GND.n539 GND.n98 0.325812
R5576 GND.n333 GND.n0 0.31982
R5577 GND GND.n96 0.295209
R5578 GND GND.n652 0.295209
R5579 GND.n1395 GND.n1394 0.282159
R5580 GND.n1619 GND.n1618 0.279127
R5581 GND.n625 GND.n624 0.279127
R5582 GND.n446 GND 0.228789
R5583 GND.n81 GND.n77 0.226583
R5584 GND.n637 GND.n633 0.226583
R5585 GND.n174 GND 0.209082
R5586 GND.n472 GND.n469 0.189094
R5587 GND.n51 GND.n50 0.189094
R5588 GND.n553 GND.n550 0.189094
R5589 GND.n584 GND.n583 0.189094
R5590 GND.n1622 GND 0.165163
R5591 GND.n1588 GND.n1587 0.15606
R5592 GND.n526 GND.n525 0.15606
R5593 GND.n1589 GND 0.140869
R5594 GND.n527 GND 0.140869
R5595 GND.n97 GND 0.134333
R5596 GND.n1536 GND 0.134333
R5597 GND.n1587 GND.n1586 0.12814
R5598 GND.n525 GND.n524 0.12814
R5599 GND.n1583 GND.n1582 0.1155
R5600 GND.n1582 GND.n1580 0.1155
R5601 GND.n1577 GND.n1576 0.1155
R5602 GND.n1576 GND.n1574 0.1155
R5603 GND.n1571 GND.n1570 0.1155
R5604 GND.n1570 GND.n1568 0.1155
R5605 GND.n1565 GND.n1564 0.1155
R5606 GND.n1564 GND.n1562 0.1155
R5607 GND.n521 GND.n520 0.1155
R5608 GND.n520 GND.n518 0.1155
R5609 GND.n515 GND.n514 0.1155
R5610 GND.n514 GND.n512 0.1155
R5611 GND.n509 GND.n508 0.1155
R5612 GND.n508 GND.n506 0.1155
R5613 GND.n503 GND.n502 0.1155
R5614 GND.n502 GND.n500 0.1155
R5615 GND.n96 GND.n72 0.110055
R5616 GND.n652 GND.n628 0.110055
R5617 GND.n71 GND.n70 0.102077
R5618 GND.n627 GND.n626 0.102077
R5619 GND.n478 GND 0.101889
R5620 GND.n559 GND 0.101889
R5621 GND.n82 GND.n81 0.0963333
R5622 GND.n83 GND.n74 0.0963333
R5623 GND.n89 GND.n74 0.0963333
R5624 GND.n90 GND.n89 0.0963333
R5625 GND.n91 GND.n90 0.0963333
R5626 GND.n638 GND.n637 0.0963333
R5627 GND.n639 GND.n630 0.0963333
R5628 GND.n645 GND.n630 0.0963333
R5629 GND.n646 GND.n645 0.0963333
R5630 GND.n647 GND.n646 0.0963333
R5631 GND.n1124 GND.n1122 0.0894537
R5632 GND.n839 GND.n837 0.0894537
R5633 GND.n685 GND.n683 0.0894537
R5634 GND.n66 GND 0.0824444
R5635 GND.n599 GND 0.0824444
R5636 GND.n1622 GND.n0 0.0795145
R5637 GND.n1619 GND.n1594 0.0740087
R5638 GND.n1539 GND.n625 0.0740087
R5639 GND.n1620 GND.n1619 0.0732412
R5640 GND.n625 GND.n600 0.0732412
R5641 GND.n1621 GND.n1620 0.0727407
R5642 GND.n600 GND.n98 0.0727407
R5643 GND.n1591 GND.n98 0.0696756
R5644 GND.n1590 GND.n1556 0.0696598
R5645 GND.n529 GND.n528 0.0696598
R5646 GND.n1594 GND.n1593 0.0692593
R5647 GND.n1539 GND.n1538 0.0692593
R5648 GND.n111 GND.n106 0.0659695
R5649 GND.n663 GND.n658 0.0659695
R5650 GND.n111 GND.n103 0.0643889
R5651 GND.n115 GND.n103 0.0643889
R5652 GND.n116 GND.n115 0.0643889
R5653 GND.n476 GND.n469 0.0643889
R5654 GND.n482 GND.n467 0.0643889
R5655 GND.n482 GND.n464 0.0643889
R5656 GND.n486 GND.n464 0.0643889
R5657 GND.n487 GND.n486 0.0643889
R5658 GND.n51 GND.n46 0.0643889
R5659 GND.n62 GND.n44 0.0643889
R5660 GND.n63 GND.n62 0.0643889
R5661 GND.n663 GND.n655 0.0643889
R5662 GND.n667 GND.n655 0.0643889
R5663 GND.n668 GND.n667 0.0643889
R5664 GND.n557 GND.n550 0.0643889
R5665 GND.n563 GND.n548 0.0643889
R5666 GND.n563 GND.n545 0.0643889
R5667 GND.n567 GND.n545 0.0643889
R5668 GND.n568 GND.n567 0.0643889
R5669 GND.n584 GND.n579 0.0643889
R5670 GND.n595 GND.n577 0.0643889
R5671 GND.n596 GND.n595 0.0643889
R5672 GND.n358 GND.n356 0.0643889
R5673 GND.n356 GND.n355 0.0643889
R5674 GND.n355 GND.n352 0.0643889
R5675 GND.n352 GND.n350 0.0643889
R5676 GND.n672 GND.n671 0.0636834
R5677 GND.n121 GND.n119 0.0636834
R5678 GND.n1593 GND 0.0628765
R5679 GND.n1538 GND 0.0628765
R5680 GND.n15 GND.n11 0.0610263
R5681 GND.n19 GND.n11 0.0610263
R5682 GND.n20 GND.n19 0.0610263
R5683 GND.n21 GND.n20 0.0610263
R5684 GND.n32 GND.n8 0.0610263
R5685 GND.n32 GND.n5 0.0610263
R5686 GND.n5 GND.n2 0.0610263
R5687 GND.n37 GND.n2 0.0610263
R5688 GND.n137 GND.n133 0.0610263
R5689 GND.n141 GND.n133 0.0610263
R5690 GND.n142 GND.n141 0.0610263
R5691 GND.n143 GND.n142 0.0610263
R5692 GND.n154 GND.n130 0.0610263
R5693 GND.n154 GND.n127 0.0610263
R5694 GND.n127 GND.n124 0.0610263
R5695 GND.n159 GND.n124 0.0610263
R5696 GND.n1622 GND.n1621 0.0593951
R5697 GND.n1609 GND.n1608 0.0580634
R5698 GND.n615 GND.n614 0.0580634
R5699 GND.n118 GND.n101 0.0580441
R5700 GND.n489 GND.n462 0.0580441
R5701 GND.n59 GND.n58 0.0580441
R5702 GND.n65 GND.n42 0.0580441
R5703 GND.n670 GND.n653 0.0580441
R5704 GND.n570 GND.n543 0.0580441
R5705 GND.n592 GND.n591 0.0580441
R5706 GND.n598 GND.n575 0.0580441
R5707 GND.n1583 GND 0.058
R5708 GND.n1577 GND 0.058
R5709 GND.n1565 GND 0.058
R5710 GND.n521 GND 0.058
R5711 GND.n515 GND 0.058
R5712 GND.n503 GND 0.058
R5713 GND.n1612 GND.n1603 0.05675
R5714 GND.n1613 GND.n1601 0.05675
R5715 GND.n618 GND.n609 0.05675
R5716 GND.n619 GND.n607 0.05675
R5717 GND.n478 GND.n477 0.0567153
R5718 GND.n559 GND.n558 0.0567153
R5719 GND.n1590 GND.n1589 0.0558279
R5720 GND.n528 GND.n527 0.0558279
R5721 GND.n1571 GND 0.0555
R5722 GND.n509 GND 0.0555
R5723 GND.n25 GND.n24 0.052907
R5724 GND.n147 GND.n146 0.052907
R5725 GND GND.n1622 0.049821
R5726 GND.n1592 GND.n1591 0.0490741
R5727 GND GND.n14 0.0490201
R5728 GND GND.n136 0.0490201
R5729 GND.n83 GND 0.0484167
R5730 GND GND.n72 0.0484167
R5731 GND.n639 GND 0.0484167
R5732 GND GND.n628 0.0484167
R5733 GND.n490 GND 0.04425
R5734 GND.n571 GND 0.04425
R5735 GND.n119 GND.n71 0.0356562
R5736 GND.n671 GND.n627 0.0356562
R5737 GND.n38 GND 0.0353684
R5738 GND.n160 GND 0.0353684
R5739 GND.n346 GND.n345 0.0352222
R5740 GND.n1616 GND 0.033625
R5741 GND.n622 GND 0.033625
R5742 GND.n58 GND 0.0324444
R5743 GND.n591 GND 0.0324444
R5744 GND GND.n358 0.0324444
R5745 GND GND.n348 0.0324444
R5746 GND.n491 GND.n490 0.03175
R5747 GND.n1541 GND.n571 0.03175
R5748 GND.n15 GND 0.0307632
R5749 GND.n24 GND 0.0307632
R5750 GND.n137 GND 0.0307632
R5751 GND.n146 GND 0.0307632
R5752 GND.n198 GND.n196 0.0307632
R5753 GND.n202 GND.n198 0.0307632
R5754 GND.n204 GND.n202 0.0307632
R5755 GND.n208 GND.n204 0.0307632
R5756 GND.n210 GND.n208 0.0307632
R5757 GND.n214 GND.n210 0.0307632
R5758 GND.n218 GND.n214 0.0307632
R5759 GND.n220 GND.n218 0.0307632
R5760 GND.n224 GND.n220 0.0307632
R5761 GND.n234 GND.n232 0.0307632
R5762 GND.n238 GND.n234 0.0307632
R5763 GND.n240 GND.n238 0.0307632
R5764 GND.n242 GND.n240 0.0307632
R5765 GND.n246 GND.n244 0.0307632
R5766 GND.n250 GND.n246 0.0307632
R5767 GND.n252 GND.n250 0.0307632
R5768 GND.n256 GND.n252 0.0307632
R5769 GND.n258 GND.n256 0.0307632
R5770 GND.n299 GND.n297 0.0307632
R5771 GND.n297 GND.n293 0.0307632
R5772 GND.n293 GND.n291 0.0307632
R5773 GND.n291 GND.n287 0.0307632
R5774 GND.n287 GND.n285 0.0307632
R5775 GND.n285 GND.n281 0.0307632
R5776 GND.n281 GND.n279 0.0307632
R5777 GND.n278 GND.n277 0.0307632
R5778 GND.n277 GND.n275 0.0307632
R5779 GND.n275 GND.n271 0.0307632
R5780 GND.n271 GND.n269 0.0307632
R5781 GND.n269 GND.n162 0.0307632
R5782 GND.n422 GND.n421 0.0307632
R5783 GND.n421 GND.n419 0.0307632
R5784 GND.n404 GND.n402 0.0307632
R5785 GND.n402 GND.n398 0.0307632
R5786 GND.n398 GND.n394 0.0307632
R5787 GND.n394 GND.n392 0.0307632
R5788 GND.n392 GND.n388 0.0307632
R5789 GND.n388 GND.n386 0.0307632
R5790 GND.n386 GND.n382 0.0307632
R5791 GND.n39 GND.n38 0.0301053
R5792 GND.n538 GND.n160 0.0301053
R5793 GND.n348 GND.n346 0.0296667
R5794 GND.n345 GND.n341 0.0296667
R5795 GND.n450 GND.n446 0.0294474
R5796 GND.n1617 GND.n1616 0.028625
R5797 GND.n1618 GND.n1617 0.028625
R5798 GND.n623 GND.n622 0.028625
R5799 GND.n624 GND.n623 0.028625
R5800 GND.n361 GND.n360 0.0284605
R5801 GND.n225 GND.n224 0.0282663
R5802 GND.n119 GND 0.0268889
R5803 GND.n671 GND 0.0268889
R5804 GND.n456 GND.n162 0.0262926
R5805 GND.n419 GND.n415 0.0238553
R5806 GND.n259 GND.n258 0.0231974
R5807 GND.n311 GND.n191 0.0225395
R5808 GND.n300 GND.n299 0.0225395
R5809 GND.n405 GND.n404 0.0218816
R5810 GND.n1586 GND 0.02175
R5811 GND.n1580 GND 0.02175
R5812 GND.n1574 GND 0.02175
R5813 GND.n1568 GND 0.02175
R5814 GND.n1562 GND 0.02175
R5815 GND.n524 GND 0.02175
R5816 GND.n518 GND 0.02175
R5817 GND.n512 GND 0.02175
R5818 GND.n506 GND 0.02175
R5819 GND.n500 GND 0.02175
R5820 GND.n375 GND.n363 0.0212237
R5821 GND.n1556 GND.n1555 0.0209918
R5822 GND.n530 GND.n529 0.0209918
R5823 GND.n228 GND.n227 0.0205658
R5824 GND.n455 GND.n451 0.0185921
R5825 GND.n91 GND 0.0182083
R5826 GND.n647 GND 0.0182083
R5827 GND GND.n349 0.0178611
R5828 GND.n382 GND.n380 0.0172763
R5829 GND GND.n82 0.0171667
R5830 GND GND.n638 0.0171667
R5831 GND.n445 GND.n443 0.0171667
R5832 GND.n443 GND.n439 0.0171667
R5833 GND.n439 GND.n437 0.0171667
R5834 GND.n432 GND.n430 0.0171667
R5835 GND.n430 GND.n426 0.0171667
R5836 GND.n414 GND.n412 0.0166184
R5837 GND.n305 GND.n263 0.0159605
R5838 GND.n314 GND 0.0158101
R5839 GND.n426 GND.n424 0.0157174
R5840 GND.n196 GND 0.0156316
R5841 GND.n244 GND 0.0156316
R5842 GND GND.n278 0.0156316
R5843 GND GND.n422 0.0156316
R5844 GND.n305 GND.n304 0.0153026
R5845 GND.n412 GND.n409 0.0146447
R5846 GND.n173 GND.n171 0.0146077
R5847 GND.n380 GND.n379 0.0139868
R5848 GND.n1128 GND.n1124 0.012734
R5849 GND.n1130 GND.n1128 0.012734
R5850 GND.n1165 GND.n1161 0.012734
R5851 GND.n1161 GND.n1159 0.012734
R5852 GND.n1159 GND.n1155 0.012734
R5853 GND.n1155 GND.n1153 0.012734
R5854 GND.n1153 GND.n1149 0.012734
R5855 GND.n1149 GND.n1147 0.012734
R5856 GND.n1147 GND.n1143 0.012734
R5857 GND.n1143 GND.n1141 0.012734
R5858 GND.n1140 GND.n1139 0.012734
R5859 GND.n1139 GND.n1137 0.012734
R5860 GND.n1187 GND.n1183 0.012734
R5861 GND.n1191 GND.n1187 0.012734
R5862 GND.n1193 GND.n1191 0.012734
R5863 GND.n1197 GND.n1193 0.012734
R5864 GND.n1199 GND.n1197 0.012734
R5865 GND.n1203 GND.n1199 0.012734
R5866 GND.n1205 GND.n1203 0.012734
R5867 GND.n1209 GND.n1205 0.012734
R5868 GND.n1211 GND.n1209 0.012734
R5869 GND.n1212 GND.n1211 0.012734
R5870 GND.n1217 GND.n1215 0.012734
R5871 GND.n1221 GND.n1217 0.012734
R5872 GND.n1223 GND.n1221 0.012734
R5873 GND.n1254 GND.n1250 0.012734
R5874 GND.n1250 GND.n1246 0.012734
R5875 GND.n1246 GND.n1244 0.012734
R5876 GND.n1244 GND.n1240 0.012734
R5877 GND.n1240 GND.n1238 0.012734
R5878 GND.n1238 GND.n1234 0.012734
R5879 GND.n1234 GND.n1232 0.012734
R5880 GND.n1232 GND.n1110 0.012734
R5881 GND.n1391 GND.n1390 0.012734
R5882 GND.n1390 GND.n1388 0.012734
R5883 GND.n1268 GND.n1264 0.012734
R5884 GND.n1272 GND.n1268 0.012734
R5885 GND.n1274 GND.n1272 0.012734
R5886 GND.n1278 GND.n1274 0.012734
R5887 GND.n1280 GND.n1278 0.012734
R5888 GND.n1284 GND.n1280 0.012734
R5889 GND.n1286 GND.n1284 0.012734
R5890 GND.n1290 GND.n1286 0.012734
R5891 GND.n1292 GND.n1290 0.012734
R5892 GND.n1293 GND.n1292 0.012734
R5893 GND.n1298 GND.n1296 0.012734
R5894 GND.n1302 GND.n1298 0.012734
R5895 GND.n1312 GND.n1310 0.012734
R5896 GND.n1316 GND.n1312 0.012734
R5897 GND.n1320 GND.n1316 0.012734
R5898 GND.n1322 GND.n1320 0.012734
R5899 GND.n1326 GND.n1322 0.012734
R5900 GND.n1328 GND.n1326 0.012734
R5901 GND.n1332 GND.n1328 0.012734
R5902 GND.n1334 GND.n1332 0.012734
R5903 GND.n1338 GND.n1334 0.012734
R5904 GND.n1340 GND.n1338 0.012734
R5905 GND.n1341 GND.n1340 0.012734
R5906 GND.n1346 GND.n1344 0.012734
R5907 GND.n1349 GND.n1346 0.012734
R5908 GND.n1351 GND.n1349 0.012734
R5909 GND.n1371 GND.n1369 0.012734
R5910 GND.n1366 GND.n1365 0.012734
R5911 GND.n1365 GND.n1363 0.012734
R5912 GND.n1363 GND.n1359 0.012734
R5913 GND.n1359 GND.n1357 0.012734
R5914 GND.n843 GND.n839 0.012734
R5915 GND.n881 GND.n877 0.012734
R5916 GND.n877 GND.n875 0.012734
R5917 GND.n875 GND.n871 0.012734
R5918 GND.n871 GND.n869 0.012734
R5919 GND.n869 GND.n865 0.012734
R5920 GND.n865 GND.n863 0.012734
R5921 GND.n863 GND.n859 0.012734
R5922 GND.n859 GND.n857 0.012734
R5923 GND.n856 GND.n855 0.012734
R5924 GND.n855 GND.n853 0.012734
R5925 GND.n903 GND.n899 0.012734
R5926 GND.n907 GND.n903 0.012734
R5927 GND.n909 GND.n907 0.012734
R5928 GND.n913 GND.n909 0.012734
R5929 GND.n915 GND.n913 0.012734
R5930 GND.n919 GND.n915 0.012734
R5931 GND.n921 GND.n919 0.012734
R5932 GND.n925 GND.n921 0.012734
R5933 GND.n927 GND.n925 0.012734
R5934 GND.n928 GND.n927 0.012734
R5935 GND.n933 GND.n931 0.012734
R5936 GND.n937 GND.n933 0.012734
R5937 GND.n939 GND.n937 0.012734
R5938 GND.n966 GND.n962 0.012734
R5939 GND.n962 GND.n958 0.012734
R5940 GND.n958 GND.n956 0.012734
R5941 GND.n956 GND.n952 0.012734
R5942 GND.n952 GND.n950 0.012734
R5943 GND.n950 GND.n946 0.012734
R5944 GND.n946 GND.n825 0.012734
R5945 GND.n1107 GND.n1105 0.012734
R5946 GND.n1104 GND.n1103 0.012734
R5947 GND.n1103 GND.n1101 0.012734
R5948 GND.n980 GND.n976 0.012734
R5949 GND.n984 GND.n980 0.012734
R5950 GND.n986 GND.n984 0.012734
R5951 GND.n990 GND.n986 0.012734
R5952 GND.n992 GND.n990 0.012734
R5953 GND.n996 GND.n992 0.012734
R5954 GND.n998 GND.n996 0.012734
R5955 GND.n1002 GND.n998 0.012734
R5956 GND.n1004 GND.n1002 0.012734
R5957 GND.n1005 GND.n1004 0.012734
R5958 GND.n1010 GND.n1008 0.012734
R5959 GND.n1025 GND.n1023 0.012734
R5960 GND.n1029 GND.n1025 0.012734
R5961 GND.n1033 GND.n1029 0.012734
R5962 GND.n1035 GND.n1033 0.012734
R5963 GND.n1039 GND.n1035 0.012734
R5964 GND.n1041 GND.n1039 0.012734
R5965 GND.n1045 GND.n1041 0.012734
R5966 GND.n1047 GND.n1045 0.012734
R5967 GND.n1051 GND.n1047 0.012734
R5968 GND.n1053 GND.n1051 0.012734
R5969 GND.n1054 GND.n1053 0.012734
R5970 GND.n1059 GND.n1057 0.012734
R5971 GND.n1062 GND.n1059 0.012734
R5972 GND.n1064 GND.n1062 0.012734
R5973 GND.n1084 GND.n1082 0.012734
R5974 GND.n1079 GND.n1078 0.012734
R5975 GND.n1078 GND.n1076 0.012734
R5976 GND.n1076 GND.n1072 0.012734
R5977 GND.n1072 GND.n1070 0.012734
R5978 GND.n689 GND.n685 0.012734
R5979 GND.n691 GND.n689 0.012734
R5980 GND.n705 GND.n703 0.012734
R5981 GND.n709 GND.n705 0.012734
R5982 GND.n711 GND.n709 0.012734
R5983 GND.n715 GND.n711 0.012734
R5984 GND.n717 GND.n715 0.012734
R5985 GND.n721 GND.n717 0.012734
R5986 GND.n723 GND.n721 0.012734
R5987 GND.n724 GND.n723 0.012734
R5988 GND.n729 GND.n727 0.012734
R5989 GND.n733 GND.n729 0.012734
R5990 GND.n779 GND.n777 0.012734
R5991 GND.n777 GND.n773 0.012734
R5992 GND.n773 GND.n769 0.012734
R5993 GND.n769 GND.n767 0.012734
R5994 GND.n767 GND.n763 0.012734
R5995 GND.n763 GND.n761 0.012734
R5996 GND.n761 GND.n757 0.012734
R5997 GND.n757 GND.n755 0.012734
R5998 GND.n755 GND.n751 0.012734
R5999 GND.n751 GND.n749 0.012734
R6000 GND.n748 GND.n747 0.012734
R6001 GND.n747 GND.n745 0.012734
R6002 GND.n745 GND.n741 0.012734
R6003 GND.n801 GND.n797 0.012734
R6004 GND.n803 GND.n801 0.012734
R6005 GND.n807 GND.n803 0.012734
R6006 GND.n809 GND.n807 0.012734
R6007 GND.n813 GND.n809 0.012734
R6008 GND.n815 GND.n813 0.012734
R6009 GND.n819 GND.n815 0.012734
R6010 GND.n821 GND.n819 0.012734
R6011 GND.n1402 GND.n1400 0.012734
R6012 GND.n1406 GND.n1402 0.012734
R6013 GND.n1445 GND.n1443 0.012734
R6014 GND.n1443 GND.n1439 0.012734
R6015 GND.n1439 GND.n1435 0.012734
R6016 GND.n1435 GND.n1433 0.012734
R6017 GND.n1433 GND.n1429 0.012734
R6018 GND.n1429 GND.n1427 0.012734
R6019 GND.n1427 GND.n1423 0.012734
R6020 GND.n1423 GND.n1421 0.012734
R6021 GND.n1421 GND.n1417 0.012734
R6022 GND.n1417 GND.n1415 0.012734
R6023 GND.n1414 GND.n1413 0.012734
R6024 GND.n1413 GND.n676 0.012734
R6025 GND.n1465 GND.n1463 0.012734
R6026 GND.n1469 GND.n1465 0.012734
R6027 GND.n1473 GND.n1469 0.012734
R6028 GND.n1475 GND.n1473 0.012734
R6029 GND.n1479 GND.n1475 0.012734
R6030 GND.n1481 GND.n1479 0.012734
R6031 GND.n1485 GND.n1481 0.012734
R6032 GND.n1487 GND.n1485 0.012734
R6033 GND.n1491 GND.n1487 0.012734
R6034 GND.n1493 GND.n1491 0.012734
R6035 GND.n1494 GND.n1493 0.012734
R6036 GND.n1499 GND.n1497 0.012734
R6037 GND.n1502 GND.n1499 0.012734
R6038 GND.n1504 GND.n1502 0.012734
R6039 GND.n1524 GND.n1522 0.012734
R6040 GND.n1519 GND.n1518 0.012734
R6041 GND.n1518 GND.n1516 0.012734
R6042 GND.n1516 GND.n1512 0.012734
R6043 GND.n1512 GND.n1510 0.012734
R6044 GND.n451 GND.n450 0.0126711
R6045 GND.n1393 GND.n1392 0.0126011
R6046 GND.n844 GND.n843 0.0126011
R6047 GND.n1397 GND.n1396 0.0126011
R6048 GND.n21 GND 0.0123421
R6049 GND.n143 GND 0.0123421
R6050 GND.n1108 GND.n825 0.0123351
R6051 GND.n1011 GND.n1010 0.0123351
R6052 GND GND.n118 0.0123056
R6053 GND GND.n489 0.0123056
R6054 GND GND.n65 0.0123056
R6055 GND GND.n670 0.0123056
R6056 GND GND.n570 0.0123056
R6057 GND GND.n598 0.0123056
R6058 GND.n350 GND 0.0123056
R6059 GND GND.n341 0.0123056
R6060 GND.n342 GND 0.0123056
R6061 GND.n1137 GND.n1133 0.0120691
R6062 GND.n734 GND.n733 0.0120691
R6063 GND.n433 GND.n432 0.0117319
R6064 GND GND.n476 0.0116111
R6065 GND.n46 GND 0.0116111
R6066 GND GND.n557 0.0116111
R6067 GND.n579 GND 0.0116111
R6068 GND.n853 GND.n849 0.0115372
R6069 GND GND.n37 0.0110263
R6070 GND GND.n159 0.0110263
R6071 GND.n1352 GND.n1351 0.0107394
R6072 GND.n967 GND.n966 0.0107394
R6073 GND.n976 GND.n974 0.0107394
R6074 GND.n1505 GND.n1504 0.0107394
R6075 GND.n1171 GND.n1130 0.0107015
R6076 GND.n694 GND.n691 0.0107015
R6077 GND.n232 GND.n228 0.0106974
R6078 GND.n1303 GND.n1302 0.0104355
R6079 GND.n1456 GND.n676 0.0104355
R6080 GND.n1255 GND.n1254 0.0102074
R6081 GND.n1264 GND.n1262 0.0102074
R6082 GND.n1065 GND.n1064 0.0102074
R6083 GND.n797 GND.n793 0.0102074
R6084 GND.n1446 GND.n1445 0.0102074
R6085 GND.n379 GND.n375 0.0100395
R6086 GND.n170 GND.n166 0.0100149
R6087 GND GND.n1615 0.009875
R6088 GND GND.n621 0.009875
R6089 GND.n887 GND.n846 0.00967553
R6090 GND.n25 GND.n8 0.00950855
R6091 GND.n147 GND.n130 0.00950855
R6092 GND.n180 GND.n178 0.00941473
R6093 GND.n184 GND.n180 0.00941473
R6094 GND.n188 GND.n184 0.00941473
R6095 GND.n190 GND.n188 0.00941473
R6096 GND.n331 GND.n327 0.00941473
R6097 GND.n327 GND.n325 0.00941473
R6098 GND.n325 GND.n321 0.00941473
R6099 GND.n321 GND.n319 0.00941473
R6100 GND.n1016 GND.n1015 0.00940957
R6101 GND.n409 GND.n405 0.00938158
R6102 GND.n1176 GND.n1118 0.00914362
R6103 GND.n785 GND.n736 0.00914362
R6104 GND.n477 GND.n467 0.00906279
R6105 GND.n558 GND.n548 0.00906279
R6106 GND.n1 GND 0.00898993
R6107 GND.n1224 GND.n1223 0.00887766
R6108 GND.n1388 GND.n1384 0.00887766
R6109 GND.n1085 GND.n1084 0.00887766
R6110 GND.n741 GND.n739 0.00887766
R6111 GND.n1407 GND.n1406 0.00887766
R6112 GND.n313 GND.n311 0.00872368
R6113 GND.n304 GND.n300 0.00872368
R6114 GND.n892 GND.n833 0.0086117
R6115 GND.n1372 GND.n1371 0.00834574
R6116 GND.n940 GND.n939 0.00834574
R6117 GND.n1101 GND.n1097 0.00834574
R6118 GND.n1525 GND.n1524 0.00834574
R6119 GND.n263 GND.n259 0.00806579
R6120 GND GND.n359 0.00806579
R6121 GND.n970 GND.n969 0.00781383
R6122 GND.n1094 GND.n831 0.00781383
R6123 GND.n116 GND.n101 0.00775202
R6124 GND.n487 GND.n462 0.00775202
R6125 GND.n59 GND.n44 0.00775202
R6126 GND.n63 GND.n42 0.00775202
R6127 GND.n668 GND.n653 0.00775202
R6128 GND.n568 GND.n543 0.00775202
R6129 GND.n592 GND.n577 0.00775202
R6130 GND.n596 GND.n575 0.00775202
R6131 GND.n899 GND.n897 0.00754787
R6132 GND.n415 GND.n414 0.00740789
R6133 GND.n1170 GND.n1166 0.00728191
R6134 GND.n1258 GND.n1257 0.00728191
R6135 GND.n1381 GND.n1116 0.00728191
R6136 GND.n699 GND.n698 0.00728191
R6137 GND.n792 GND.n790 0.00728191
R6138 GND.n1451 GND.n1450 0.00728191
R6139 GND.n314 GND.n313 0.00707895
R6140 GND.n1183 GND.n1181 0.00701596
R6141 GND.n1306 GND.n1305 0.00701596
R6142 GND.n780 GND.n779 0.00701596
R6143 GND.n1459 GND.n1458 0.00701596
R6144 GND.n886 GND.n882 0.00675
R6145 GND.n1023 GND.n1019 0.00675
R6146 GND GND.n1140 0.00661702
R6147 GND.n1215 GND 0.00661702
R6148 GND GND.n1391 0.00661702
R6149 GND.n1296 GND 0.00661702
R6150 GND.n1344 GND 0.00661702
R6151 GND.n1366 GND 0.00661702
R6152 GND GND.n856 0.00661702
R6153 GND.n931 GND 0.00661702
R6154 GND GND.n1104 0.00661702
R6155 GND.n1008 GND 0.00661702
R6156 GND.n1057 GND 0.00661702
R6157 GND.n1079 GND 0.00661702
R6158 GND.n727 GND 0.00661702
R6159 GND GND.n748 0.00661702
R6160 GND.n1400 GND 0.00661702
R6161 GND GND.n1414 0.00661702
R6162 GND.n1497 GND 0.00661702
R6163 GND.n1519 GND 0.00661702
R6164 GND.n882 GND.n881 0.00648404
R6165 GND.n1019 GND.n1018 0.00648404
R6166 GND.n174 GND.n173 0.00647015
R6167 GND.n178 GND.n174 0.00631395
R6168 GND.n1181 GND.n1180 0.00621809
R6169 GND.n1310 GND.n1306 0.00621809
R6170 GND.n784 GND.n780 0.00621809
R6171 GND.n1463 GND.n1459 0.00621809
R6172 GND GND.n242 0.00609211
R6173 GND.n279 GND 0.00609211
R6174 GND.n423 GND 0.00609211
R6175 GND.n360 GND 0.00609211
R6176 GND.n1166 GND.n1165 0.00595213
R6177 GND.n1258 GND.n1228 0.00595213
R6178 GND.n1383 GND.n1381 0.00595213
R6179 GND.n1088 GND.n1087 0.00595213
R6180 GND.n703 GND.n699 0.00595213
R6181 GND.n790 GND.n680 0.00595213
R6182 GND.n1451 GND.n1409 0.00595213
R6183 GND.n437 GND.n433 0.00593478
R6184 GND.n456 GND.n455 0.00593421
R6185 GND.n897 GND.n896 0.00568617
R6186 GND.n1375 GND.n1374 0.00542021
R6187 GND.n970 GND.n944 0.00542021
R6188 GND.n1096 GND.n1094 0.00542021
R6189 GND.n1528 GND.n1527 0.00542021
R6190 GND.n332 GND.n331 0.00534496
R6191 GND GND.n193 0.00510526
R6192 GND.n319 GND.n315 0.00505426
R6193 GND.n424 GND 0.00502899
R6194 GND.n1374 GND.n1372 0.0048883
R6195 GND.n944 GND.n940 0.0048883
R6196 GND.n1097 GND.n1096 0.0048883
R6197 GND.n1527 GND.n1525 0.0048883
R6198 GND.n359 GND 0.00466667
R6199 GND.n896 GND.n892 0.00462234
R6200 GND.n332 GND.n190 0.00456977
R6201 GND.n1537 GND 0.00456173
R6202 GND.n171 GND.n170 0.00454478
R6203 GND.n1228 GND.n1224 0.00435638
R6204 GND.n1384 GND.n1383 0.00435638
R6205 GND.n1087 GND.n1085 0.00435638
R6206 GND.n739 GND.n680 0.00435638
R6207 GND.n1409 GND.n1407 0.00435638
R6208 GND.n1180 GND.n1176 0.00409043
R6209 GND.n785 GND.n784 0.00409043
R6210 GND.n227 GND.n225 0.00396053
R6211 GND.n1018 GND.n1016 0.00382447
R6212 GND.n1305 GND.n1303 0.00379255
R6213 GND.n1458 GND.n1456 0.00379255
R6214 GND.n887 GND.n886 0.00355851
R6215 GND.n1171 GND.n1170 0.0035266
R6216 GND.n698 GND.n694 0.0035266
R6217 GND.n528 GND.n1 0.00349775
R6218 GND GND.n1592 0.00340123
R6219 GND GND.n1537 0.00340123
R6220 GND.n349 GND 0.00327778
R6221 GND.n342 GND 0.00327778
R6222 GND.n1622 GND.n1 0.00323583
R6223 GND.n424 GND.n423 0.00313158
R6224 GND.n1554 GND.n1553 0.00307458
R6225 GND.n1257 GND.n1255 0.0030266
R6226 GND.n1262 GND.n1116 0.0030266
R6227 GND.n1067 GND.n1065 0.0030266
R6228 GND.n793 GND.n792 0.0030266
R6229 GND.n1450 GND.n1446 0.0030266
R6230 GND.n315 GND.n314 0.00292248
R6231 GND.n1589 GND.n1588 0.00290385
R6232 GND.n527 GND.n526 0.00290385
R6233 GND.n363 GND.n361 0.00280263
R6234 GND.n1600 GND.n1597 0.00277946
R6235 GND.n606 GND.n603 0.00277946
R6236 GND.n1141 GND 0.00276064
R6237 GND.n1212 GND 0.00276064
R6238 GND.n1392 GND 0.00276064
R6239 GND.n1293 GND 0.00276064
R6240 GND.n1341 GND 0.00276064
R6241 GND GND.n1354 0.00276064
R6242 GND.n1369 GND 0.00276064
R6243 GND.n1357 GND 0.00276064
R6244 GND.n857 GND 0.00276064
R6245 GND.n928 GND 0.00276064
R6246 GND.n1105 GND 0.00276064
R6247 GND.n1005 GND 0.00276064
R6248 GND.n1054 GND 0.00276064
R6249 GND GND.n1067 0.00276064
R6250 GND.n1082 GND 0.00276064
R6251 GND.n1070 GND 0.00276064
R6252 GND.n724 GND 0.00276064
R6253 GND.n749 GND 0.00276064
R6254 GND.n1397 GND 0.00276064
R6255 GND.n1415 GND 0.00276064
R6256 GND.n1494 GND 0.00276064
R6257 GND GND.n1507 0.00276064
R6258 GND.n1522 GND 0.00276064
R6259 GND.n1510 GND 0.00276064
R6260 GND.n1591 GND.n1590 0.00249812
R6261 GND.n1354 GND.n1352 0.00249468
R6262 GND.n969 GND.n967 0.00249468
R6263 GND.n974 GND.n831 0.00249468
R6264 GND.n1507 GND.n1505 0.00249468
R6265 GND.n359 GND 0.00247368
R6266 GND.n532 GND.n531 0.00207681
R6267 GND.n606 GND.n605 0.00193331
R6268 GND.n1600 GND.n1599 0.00193331
R6269 GND.n1609 GND.n1603 0.00175
R6270 GND.n1613 GND.n1612 0.00175
R6271 GND.n1615 GND.n1601 0.00175
R6272 GND.n615 GND.n609 0.00175
R6273 GND.n619 GND.n618 0.00175
R6274 GND.n621 GND.n607 0.00175
R6275 GND.n1375 GND 0.00169681
R6276 GND.n849 GND.n833 0.00169681
R6277 GND.n1528 GND 0.00169681
R6278 GND.n530 GND.n494 0.00150013
R6279 GND.n193 GND.n191 0.00148684
R6280 GND.n446 GND.n445 0.00122464
R6281 GND.n1133 GND.n1118 0.00116489
R6282 GND.n1088 GND 0.00116489
R6283 GND.n736 GND.n734 0.00116489
R6284 GND.n534 GND.n532 0.00115206
R6285 GND.n534 GND.n533 0.00115206
R6286 GND.n1551 GND.n1550 0.00109111
R6287 GND.n1617 GND.n1600 0.00108327
R6288 GND.n623 GND.n606 0.00108327
R6289 GND.n1552 GND.n1551 0.00107707
R6290 GND.n120 GND.n97 0.00106078
R6291 GND.n1536 GND.n1535 0.00106078
R6292 GND.n69 GND.n68 0.00100171
R6293 GND.n365 GND.n40 0.00100171
R6294 GND.n1540 GND.n573 0.00100171
R6295 GND.n540 GND.n539 0.00100171
R6296 GND.n491 GND.n69 0.00100166
R6297 GND.n40 GND.n39 0.00100166
R6298 GND.n1541 GND.n1540 0.00100166
R6299 GND.n539 GND.n538 0.00100166
R6300 GND.n1172 GND.n1171 0.00100097
R6301 GND.n1303 GND.n1261 0.00100097
R6302 GND.n694 GND.n693 0.00100097
R6303 GND.n1456 GND.n1455 0.00100097
R6304 GND.n171 GND.n164 0.00100097
R6305 GND.n225 GND.n192 0.00100097
R6306 GND.n457 GND.n456 0.00100097
R6307 GND.n1555 GND.n1554 0.00100086
R6308 GND.n1555 GND.n1552 0.00100017
R6309 GND.n531 GND.n530 0.001
R6310 GND.n66 GND.n41 0.001
R6311 GND.n599 GND.n574 0.001
R6312 GND.n535 GND.n534 0.001
R6313 GND.n1108 GND.n1107 0.000898936
R6314 GND.n1015 GND.n1011 0.000898936
R6315 GND.n1393 GND.n1110 0.000632979
R6316 GND.n846 GND.n844 0.000632979
R6317 GND.n1396 GND.n821 0.000632979
R6318 GND.n492 GND.n491 0.000560793
R6319 GND.n1542 GND.n1541 0.000560793
R6320 GND.n538 GND.n537 0.000560793
R6321 GND.n541 GND.n540 0.000557763
R6322 GND.n573 GND.n572 0.000557763
R6323 GND.n366 GND.n365 0.000557763
R6324 GND.n68 GND.n67 0.000557763
R6325 GND.n603 GND.n602 0.000528881
R6326 GND.n602 GND.n601 0.000528881
R6327 GND.n605 GND.n604 0.000528881
R6328 GND.n1597 GND.n1596 0.000528881
R6329 GND.n1596 GND.n1595 0.000528881
R6330 GND.n1599 GND.n1598 0.000528881
R6331 GND.n374 GND.n373 0.000506774
R6332 GND.n411 GND.n410 0.000506774
R6333 GND.n308 GND.n192 0.000506774
R6334 GND.n458 GND.n457 0.000506774
R6335 GND.n164 GND.n163 0.000506774
R6336 GND.n310 GND.n309 0.000506774
R6337 GND.n307 GND.n306 0.000506774
R6338 GND.n1173 GND.n1172 0.000506774
R6339 GND.n1175 GND.n1174 0.000506774
R6340 GND.n1378 GND.n1261 0.000506774
R6341 GND.n1377 GND.n1376 0.000506774
R6342 GND.n1380 GND.n1379 0.000506774
R6343 GND.n1260 GND.n1259 0.000506774
R6344 GND.n889 GND.n888 0.000506774
R6345 GND.n891 GND.n890 0.000506774
R6346 GND.n1091 GND.n973 0.000506774
R6347 GND.n1090 GND.n1089 0.000506774
R6348 GND.n1093 GND.n1092 0.000506774
R6349 GND.n972 GND.n971 0.000506774
R6350 GND.n693 GND.n692 0.000506774
R6351 GND.n787 GND.n786 0.000506774
R6352 GND.n1455 GND.n1454 0.000506774
R6353 GND.n1530 GND.n1529 0.000506774
R6354 GND.n1453 GND.n1452 0.000506774
R6355 GND.n789 GND.n788 0.000506774
R6356 GND.n412 GND.n411 0.00050097
R6357 GND.n311 GND.n310 0.00050097
R6358 GND.n306 GND.n305 0.00050097
R6359 GND.n1176 GND.n1175 0.00050097
R6360 GND.n1376 GND.n1375 0.00050097
R6361 GND.n1381 GND.n1380 0.00050097
R6362 GND.n1259 GND.n1258 0.00050097
R6363 GND.n888 GND.n887 0.00050097
R6364 GND.n892 GND.n891 0.00050097
R6365 GND.n1016 GND.n973 0.00050097
R6366 GND.n1089 GND.n1088 0.00050097
R6367 GND.n1094 GND.n1093 0.00050097
R6368 GND.n971 GND.n970 0.00050097
R6369 GND.n786 GND.n785 0.00050097
R6370 GND.n1529 GND.n1528 0.00050097
R6371 GND.n1452 GND.n1451 0.00050097
R6372 GND.n790 GND.n789 0.00050097
R6373 GND.n375 GND.n374 0.00050097
R6374 GND.n433 GND.n333 0.00050016
R6375 A0.n82 A0.n80 145.809
R6376 A0.n25 A0.n23 145.809
R6377 A0.n124 A0.n122 145.809
R6378 A0.n62 A0.n60 145.808
R6379 A0.n25 A0.n24 107.409
R6380 A0.n27 A0.n26 107.409
R6381 A0.n29 A0.n28 107.409
R6382 A0.n31 A0.n30 107.409
R6383 A0.n33 A0.n32 107.409
R6384 A0.n35 A0.n34 107.409
R6385 A0.n124 A0.n123 107.409
R6386 A0.n126 A0.n125 107.409
R6387 A0.n128 A0.n127 107.409
R6388 A0.n130 A0.n129 107.409
R6389 A0.n132 A0.n131 107.409
R6390 A0.n134 A0.n133 107.409
R6391 A0.n82 A0.n81 107.407
R6392 A0.n84 A0.n83 107.407
R6393 A0.n86 A0.n85 107.407
R6394 A0.n88 A0.n87 107.407
R6395 A0.n90 A0.n89 107.407
R6396 A0.n92 A0.n91 107.407
R6397 A0.n62 A0.n61 107.407
R6398 A0.n64 A0.n63 107.407
R6399 A0.n66 A0.n65 107.407
R6400 A0.n68 A0.n67 107.407
R6401 A0.n70 A0.n69 107.407
R6402 A0.n72 A0.n71 107.407
R6403 A0.n98 A0.n96 87.1779
R6404 A0.n43 A0.n41 87.1779
R6405 A0.n4 A0.n2 87.1779
R6406 A0.n142 A0.n140 87.1779
R6407 A0.n14 A0.n13 52.82
R6408 A0.n152 A0.n151 52.82
R6409 A0.n98 A0.n97 52.82
R6410 A0.n100 A0.n99 52.82
R6411 A0.n102 A0.n101 52.82
R6412 A0.n104 A0.n103 52.82
R6413 A0.n106 A0.n105 52.82
R6414 A0.n108 A0.n107 52.82
R6415 A0.n43 A0.n42 52.82
R6416 A0.n45 A0.n44 52.82
R6417 A0.n47 A0.n46 52.82
R6418 A0.n49 A0.n48 52.82
R6419 A0.n51 A0.n50 52.82
R6420 A0.n53 A0.n52 52.82
R6421 A0.n4 A0.n3 52.82
R6422 A0.n6 A0.n5 52.82
R6423 A0.n8 A0.n7 52.82
R6424 A0.n10 A0.n9 52.82
R6425 A0.n12 A0.n11 52.82
R6426 A0.n142 A0.n141 52.82
R6427 A0.n144 A0.n143 52.82
R6428 A0.n146 A0.n145 52.82
R6429 A0.n148 A0.n147 52.82
R6430 A0.n150 A0.n149 52.82
R6431 A0 A0.n109 51.0745
R6432 A0 A0.n54 51.0745
R6433 A0.n84 A0.n82 38.4005
R6434 A0.n86 A0.n84 38.4005
R6435 A0.n88 A0.n86 38.4005
R6436 A0.n90 A0.n88 38.4005
R6437 A0.n92 A0.n90 38.4005
R6438 A0.n93 A0.n92 38.4005
R6439 A0.n64 A0.n62 38.4005
R6440 A0.n66 A0.n64 38.4005
R6441 A0.n68 A0.n66 38.4005
R6442 A0.n70 A0.n68 38.4005
R6443 A0.n72 A0.n70 38.4005
R6444 A0.n73 A0.n72 38.4005
R6445 A0.n27 A0.n25 38.4005
R6446 A0.n29 A0.n27 38.4005
R6447 A0.n31 A0.n29 38.4005
R6448 A0.n33 A0.n31 38.4005
R6449 A0.n35 A0.n33 38.4005
R6450 A0.n36 A0.n35 38.4005
R6451 A0.n126 A0.n124 38.4005
R6452 A0.n128 A0.n126 38.4005
R6453 A0.n130 A0.n128 38.4005
R6454 A0.n132 A0.n130 38.4005
R6455 A0.n134 A0.n132 38.4005
R6456 A0.n135 A0.n134 38.4005
R6457 A0.n100 A0.n98 34.3584
R6458 A0.n102 A0.n100 34.3584
R6459 A0.n104 A0.n102 34.3584
R6460 A0.n106 A0.n104 34.3584
R6461 A0.n108 A0.n106 34.3584
R6462 A0.n110 A0.n108 34.3584
R6463 A0.n45 A0.n43 34.3584
R6464 A0.n47 A0.n45 34.3584
R6465 A0.n49 A0.n47 34.3584
R6466 A0.n51 A0.n49 34.3584
R6467 A0.n53 A0.n51 34.3584
R6468 A0.n55 A0.n53 34.3584
R6469 A0.n6 A0.n4 34.3584
R6470 A0.n8 A0.n6 34.3584
R6471 A0.n10 A0.n8 34.3584
R6472 A0.n12 A0.n10 34.3584
R6473 A0.n14 A0.n12 34.3584
R6474 A0.n18 A0.n14 34.3584
R6475 A0.n144 A0.n142 34.3584
R6476 A0.n146 A0.n144 34.3584
R6477 A0.n148 A0.n146 34.3584
R6478 A0.n150 A0.n148 34.3584
R6479 A0.n152 A0.n150 34.3584
R6480 A0.n153 A0.n152 34.3584
R6481 A0.n78 A0.t108 26.5955
R6482 A0.n78 A0.t123 26.5955
R6483 A0.n80 A0.t105 26.5955
R6484 A0.n80 A0.t78 26.5955
R6485 A0.n81 A0.t68 26.5955
R6486 A0.n81 A0.t90 26.5955
R6487 A0.n83 A0.t88 26.5955
R6488 A0.n83 A0.t114 26.5955
R6489 A0.n85 A0.t80 26.5955
R6490 A0.n85 A0.t65 26.5955
R6491 A0.n87 A0.t99 26.5955
R6492 A0.n87 A0.t117 26.5955
R6493 A0.n89 A0.t115 26.5955
R6494 A0.n89 A0.t86 26.5955
R6495 A0.n91 A0.t72 26.5955
R6496 A0.n91 A0.t97 26.5955
R6497 A0.n59 A0.t70 26.5955
R6498 A0.n59 A0.t95 26.5955
R6499 A0.n60 A0.t84 26.5955
R6500 A0.n60 A0.t69 26.5955
R6501 A0.n61 A0.t93 26.5955
R6502 A0.n61 A0.t77 26.5955
R6503 A0.n63 A0.t120 26.5955
R6504 A0.n63 A0.t82 26.5955
R6505 A0.n65 A0.t87 26.5955
R6506 A0.n65 A0.t102 26.5955
R6507 A0.n67 A0.t100 26.5955
R6508 A0.n67 A0.t64 26.5955
R6509 A0.n69 A0.t126 26.5955
R6510 A0.n69 A0.t75 26.5955
R6511 A0.n71 A0.t113 26.5955
R6512 A0.n71 A0.t109 26.5955
R6513 A0.n22 A0.t71 26.5955
R6514 A0.n22 A0.t96 26.5955
R6515 A0.n23 A0.t85 26.5955
R6516 A0.n23 A0.t106 26.5955
R6517 A0.n24 A0.t104 26.5955
R6518 A0.n24 A0.t122 26.5955
R6519 A0.n26 A0.t67 26.5955
R6520 A0.n26 A0.t89 26.5955
R6521 A0.n28 A0.t118 26.5955
R6522 A0.n28 A0.t112 26.5955
R6523 A0.n30 A0.t79 26.5955
R6524 A0.n30 A0.t92 26.5955
R6525 A0.n32 A0.t98 26.5955
R6526 A0.n32 A0.t116 26.5955
R6527 A0.n34 A0.t124 26.5955
R6528 A0.n34 A0.t73 26.5955
R6529 A0.n121 A0.t111 26.5955
R6530 A0.n121 A0.t66 26.5955
R6531 A0.n122 A0.t91 26.5955
R6532 A0.n122 A0.t107 26.5955
R6533 A0.n123 A0.t83 26.5955
R6534 A0.n123 A0.t94 26.5955
R6535 A0.n125 A0.t103 26.5955
R6536 A0.n125 A0.t121 26.5955
R6537 A0.n127 A0.t119 26.5955
R6538 A0.n127 A0.t81 26.5955
R6539 A0.n129 A0.t76 26.5955
R6540 A0.n129 A0.t101 26.5955
R6541 A0.n131 A0.t110 26.5955
R6542 A0.n131 A0.t127 26.5955
R6543 A0.n133 A0.t125 26.5955
R6544 A0.n133 A0.t74 26.5955
R6545 A0.n109 A0.t46 24.9236
R6546 A0.n109 A0.t61 24.9236
R6547 A0.n96 A0.t43 24.9236
R6548 A0.n96 A0.t16 24.9236
R6549 A0.n97 A0.t6 24.9236
R6550 A0.n97 A0.t28 24.9236
R6551 A0.n99 A0.t26 24.9236
R6552 A0.n99 A0.t52 24.9236
R6553 A0.n101 A0.t18 24.9236
R6554 A0.n101 A0.t3 24.9236
R6555 A0.n103 A0.t37 24.9236
R6556 A0.n103 A0.t55 24.9236
R6557 A0.n105 A0.t53 24.9236
R6558 A0.n105 A0.t24 24.9236
R6559 A0.n107 A0.t10 24.9236
R6560 A0.n107 A0.t35 24.9236
R6561 A0.n54 A0.t8 24.9236
R6562 A0.n54 A0.t33 24.9236
R6563 A0.n41 A0.t22 24.9236
R6564 A0.n41 A0.t7 24.9236
R6565 A0.n42 A0.t31 24.9236
R6566 A0.n42 A0.t15 24.9236
R6567 A0.n44 A0.t58 24.9236
R6568 A0.n44 A0.t20 24.9236
R6569 A0.n46 A0.t25 24.9236
R6570 A0.n46 A0.t40 24.9236
R6571 A0.n48 A0.t38 24.9236
R6572 A0.n48 A0.t2 24.9236
R6573 A0.n50 A0.t0 24.9236
R6574 A0.n50 A0.t13 24.9236
R6575 A0.n52 A0.t51 24.9236
R6576 A0.n52 A0.t47 24.9236
R6577 A0.n15 A0.t9 24.9236
R6578 A0.n15 A0.t34 24.9236
R6579 A0.n2 A0.t23 24.9236
R6580 A0.n2 A0.t44 24.9236
R6581 A0.n3 A0.t42 24.9236
R6582 A0.n3 A0.t60 24.9236
R6583 A0.n5 A0.t5 24.9236
R6584 A0.n5 A0.t27 24.9236
R6585 A0.n7 A0.t56 24.9236
R6586 A0.n7 A0.t50 24.9236
R6587 A0.n9 A0.t17 24.9236
R6588 A0.n9 A0.t30 24.9236
R6589 A0.n11 A0.t36 24.9236
R6590 A0.n11 A0.t54 24.9236
R6591 A0.n13 A0.t62 24.9236
R6592 A0.n13 A0.t11 24.9236
R6593 A0.n154 A0.t49 24.9236
R6594 A0.n154 A0.t4 24.9236
R6595 A0.n140 A0.t29 24.9236
R6596 A0.n140 A0.t45 24.9236
R6597 A0.n141 A0.t21 24.9236
R6598 A0.n141 A0.t32 24.9236
R6599 A0.n143 A0.t41 24.9236
R6600 A0.n143 A0.t59 24.9236
R6601 A0.n145 A0.t57 24.9236
R6602 A0.n145 A0.t19 24.9236
R6603 A0.n147 A0.t14 24.9236
R6604 A0.n147 A0.t39 24.9236
R6605 A0.n149 A0.t48 24.9236
R6606 A0.n149 A0.t1 24.9236
R6607 A0.n151 A0.t63 24.9236
R6608 A0.n151 A0.t12 24.9236
R6609 A0 A0.n110 11.4429
R6610 A0 A0.n55 11.4429
R6611 A0 A0.n18 11.4429
R6612 A0.n37 A0.n22 8.55118
R6613 A0.n136 A0.n121 8.55118
R6614 A0.n74 A0.n59 8.55117
R6615 A0.n79 A0.n78 8.47293
R6616 A0.n16 A0.n15 7.80093
R6617 A0.n155 A0.n154 7.80093
R6618 A0.n38 A0.n37 3.20954
R6619 A0.n137 A0.n136 3.20953
R6620 A0.n75 A0.n74 3.20289
R6621 A0.n111 A0 3.10353
R6622 A0.n56 A0 3.10353
R6623 A0.n19 A0 3.10353
R6624 A0 A0.n159 3.10353
R6625 A0.n95 A0.n94 3.1005
R6626 A0.n17 A0.n1 3.1005
R6627 A0.n157 A0.n156 3.1005
R6628 A0.n94 A0.n93 2.71565
R6629 A0.n74 A0.n73 2.13383
R6630 A0.n37 A0.n36 2.13383
R6631 A0.n136 A0.n135 2.13383
R6632 A0.n110 A0 1.74595
R6633 A0.n55 A0 1.74595
R6634 A0.n18 A0.n17 1.16414
R6635 A0.n156 A0.n153 1.16414
R6636 A0.n117 A0.n116 1.07337
R6637 A0.n118 A0.n117 0.69375
R6638 A0.n119 A0.n118 0.68905
R6639 A0.n16 A0 0.488972
R6640 A0.n155 A0 0.488972
R6641 A0.n118 A0.n39 0.414635
R6642 A0.n117 A0.n76 0.382465
R6643 A0.n119 A0 0.380486
R6644 A0.n120 A0.n119 0.368576
R6645 A0.n94 A0.n79 0.196887
R6646 A0.n39 A0.n38 0.157252
R6647 A0.n137 A0.n120 0.139891
R6648 A0.n116 A0.n115 0.139389
R6649 A0.n76 A0.n75 0.132946
R6650 A0.n20 A0.n1 0.113
R6651 A0.n158 A0.n157 0.113
R6652 A0.n114 A0.n95 0.101889
R6653 A0.n17 A0.n16 0.0893205
R6654 A0.n156 A0.n155 0.0893205
R6655 A0.n114 A0.n112 0.0282778
R6656 A0.n95 A0.n77 0.0268889
R6657 A0.n58 A0.n57 0.0213333
R6658 A0.n21 A0.n20 0.0143889
R6659 A0.n158 A0.n139 0.0143889
R6660 A0.n75 A0.n58 0.00100004
R6661 A0.n139 A0.n137 0.00100004
R6662 A0.n38 A0.n21 0.00100004
R6663 A0.n112 A0.n111 0.000513335
R6664 A0.n57 A0.n56 0.000513335
R6665 A0.n20 A0.n19 0.000513218
R6666 A0.n159 A0.n158 0.000513218
R6667 A0.n58 A0.n40 0.00050517
R6668 A0.n114 A0.n113 0.000504838
R6669 A0.n21 A0.n0 0.000504838
R6670 A0.n139 A0.n138 0.000504838
R6671 A0.n115 A0.n114 0.000501713
R6672 I12.n12 I12.t0 260.435
R6673 I12.n2 I12.t3 230.576
R6674 I12.n5 I12.t5 196.549
R6675 I12.n2 I12.t1 158.275
R6676 I12.n12 I12.t4 156.403
R6677 I12.n5 I12.t2 148.35
R6678 I12.n6 I12.n5 9.49829
R6679 I12.n3 I12.n2 8.76429
R6680 I12.n7 I12.n6 7.9582
R6681 I12.n4 I12.n3 7.74345
R6682 I12.n13 I12.n12 7.60183
R6683 I12.n3 I12 6.66717
R6684 I12.n6 I12 6.44139
R6685 I12 I12.n13 4.8645
R6686 I12.n9 I12.n8 2.33638
R6687 I12.n7 I12.n4 1.0005
R6688 I12.n8 I12 0.590013
R6689 I12.n8 I12.n7 0.446956
R6690 I12.n4 I12 0.380411
R6691 I12.n10 I12.n0 0.0344286
R6692 I12.n9 I12.n1 0.00182856
R6693 I12.n10 I12.n9 0.00149885
R6694 I12.n13 I12.n11 0.00133362
R6695 I12.n11 I12.n10 0.00100077
R6696 A1.n82 A1.n80 145.809
R6697 A1.n25 A1.n23 145.809
R6698 A1.n124 A1.n122 145.809
R6699 A1.n62 A1.n60 145.808
R6700 A1.n25 A1.n24 107.409
R6701 A1.n27 A1.n26 107.409
R6702 A1.n29 A1.n28 107.409
R6703 A1.n31 A1.n30 107.409
R6704 A1.n33 A1.n32 107.409
R6705 A1.n35 A1.n34 107.409
R6706 A1.n124 A1.n123 107.409
R6707 A1.n126 A1.n125 107.409
R6708 A1.n128 A1.n127 107.409
R6709 A1.n130 A1.n129 107.409
R6710 A1.n132 A1.n131 107.409
R6711 A1.n134 A1.n133 107.409
R6712 A1.n82 A1.n81 107.407
R6713 A1.n84 A1.n83 107.407
R6714 A1.n86 A1.n85 107.407
R6715 A1.n88 A1.n87 107.407
R6716 A1.n90 A1.n89 107.407
R6717 A1.n92 A1.n91 107.407
R6718 A1.n62 A1.n61 107.407
R6719 A1.n64 A1.n63 107.407
R6720 A1.n66 A1.n65 107.407
R6721 A1.n68 A1.n67 107.407
R6722 A1.n70 A1.n69 107.407
R6723 A1.n72 A1.n71 107.407
R6724 A1.n98 A1.n96 87.1779
R6725 A1.n43 A1.n41 87.1779
R6726 A1.n4 A1.n2 87.1779
R6727 A1.n142 A1.n140 87.1779
R6728 A1.n14 A1.n13 52.82
R6729 A1.n152 A1.n151 52.82
R6730 A1.n98 A1.n97 52.82
R6731 A1.n100 A1.n99 52.82
R6732 A1.n102 A1.n101 52.82
R6733 A1.n104 A1.n103 52.82
R6734 A1.n106 A1.n105 52.82
R6735 A1.n108 A1.n107 52.82
R6736 A1.n43 A1.n42 52.82
R6737 A1.n45 A1.n44 52.82
R6738 A1.n47 A1.n46 52.82
R6739 A1.n49 A1.n48 52.82
R6740 A1.n51 A1.n50 52.82
R6741 A1.n53 A1.n52 52.82
R6742 A1.n4 A1.n3 52.82
R6743 A1.n6 A1.n5 52.82
R6744 A1.n8 A1.n7 52.82
R6745 A1.n10 A1.n9 52.82
R6746 A1.n12 A1.n11 52.82
R6747 A1.n142 A1.n141 52.82
R6748 A1.n144 A1.n143 52.82
R6749 A1.n146 A1.n145 52.82
R6750 A1.n148 A1.n147 52.82
R6751 A1.n150 A1.n149 52.82
R6752 A1 A1.n109 51.0745
R6753 A1 A1.n54 51.0745
R6754 A1.n84 A1.n82 38.4005
R6755 A1.n86 A1.n84 38.4005
R6756 A1.n88 A1.n86 38.4005
R6757 A1.n90 A1.n88 38.4005
R6758 A1.n92 A1.n90 38.4005
R6759 A1.n93 A1.n92 38.4005
R6760 A1.n64 A1.n62 38.4005
R6761 A1.n66 A1.n64 38.4005
R6762 A1.n68 A1.n66 38.4005
R6763 A1.n70 A1.n68 38.4005
R6764 A1.n72 A1.n70 38.4005
R6765 A1.n73 A1.n72 38.4005
R6766 A1.n27 A1.n25 38.4005
R6767 A1.n29 A1.n27 38.4005
R6768 A1.n31 A1.n29 38.4005
R6769 A1.n33 A1.n31 38.4005
R6770 A1.n35 A1.n33 38.4005
R6771 A1.n36 A1.n35 38.4005
R6772 A1.n126 A1.n124 38.4005
R6773 A1.n128 A1.n126 38.4005
R6774 A1.n130 A1.n128 38.4005
R6775 A1.n132 A1.n130 38.4005
R6776 A1.n134 A1.n132 38.4005
R6777 A1.n135 A1.n134 38.4005
R6778 A1.n100 A1.n98 34.3584
R6779 A1.n102 A1.n100 34.3584
R6780 A1.n104 A1.n102 34.3584
R6781 A1.n106 A1.n104 34.3584
R6782 A1.n108 A1.n106 34.3584
R6783 A1.n110 A1.n108 34.3584
R6784 A1.n45 A1.n43 34.3584
R6785 A1.n47 A1.n45 34.3584
R6786 A1.n49 A1.n47 34.3584
R6787 A1.n51 A1.n49 34.3584
R6788 A1.n53 A1.n51 34.3584
R6789 A1.n55 A1.n53 34.3584
R6790 A1.n6 A1.n4 34.3584
R6791 A1.n8 A1.n6 34.3584
R6792 A1.n10 A1.n8 34.3584
R6793 A1.n12 A1.n10 34.3584
R6794 A1.n14 A1.n12 34.3584
R6795 A1.n18 A1.n14 34.3584
R6796 A1.n144 A1.n142 34.3584
R6797 A1.n146 A1.n144 34.3584
R6798 A1.n148 A1.n146 34.3584
R6799 A1.n150 A1.n148 34.3584
R6800 A1.n152 A1.n150 34.3584
R6801 A1.n153 A1.n152 34.3584
R6802 A1.n78 A1.t103 26.5955
R6803 A1.n78 A1.t117 26.5955
R6804 A1.n80 A1.t91 26.5955
R6805 A1.n80 A1.t85 26.5955
R6806 A1.n81 A1.t83 26.5955
R6807 A1.n81 A1.t76 26.5955
R6808 A1.n83 A1.t74 26.5955
R6809 A1.n83 A1.t67 26.5955
R6810 A1.n85 A1.t73 26.5955
R6811 A1.n85 A1.t81 26.5955
R6812 A1.n87 A1.t127 26.5955
R6813 A1.n87 A1.t79 26.5955
R6814 A1.n89 A1.t77 26.5955
R6815 A1.n89 A1.t112 26.5955
R6816 A1.n91 A1.t69 26.5955
R6817 A1.n91 A1.t125 26.5955
R6818 A1.n59 A1.t89 26.5955
R6819 A1.n59 A1.t84 26.5955
R6820 A1.n60 A1.t116 26.5955
R6821 A1.n60 A1.t123 26.5955
R6822 A1.n61 A1.t64 26.5955
R6823 A1.n61 A1.t102 26.5955
R6824 A1.n63 A1.t121 26.5955
R6825 A1.n63 A1.t114 26.5955
R6826 A1.n65 A1.t93 26.5955
R6827 A1.n65 A1.t106 26.5955
R6828 A1.n67 A1.t104 26.5955
R6829 A1.n67 A1.t100 26.5955
R6830 A1.n69 A1.t98 26.5955
R6831 A1.n69 A1.t110 26.5955
R6832 A1.n71 A1.t95 26.5955
R6833 A1.n71 A1.t87 26.5955
R6834 A1.n22 A1.t68 26.5955
R6835 A1.n22 A1.t124 26.5955
R6836 A1.n23 A1.t96 26.5955
R6837 A1.n23 A1.t92 26.5955
R6838 A1.n24 A1.t90 26.5955
R6839 A1.n24 A1.t101 26.5955
R6840 A1.n26 A1.t82 26.5955
R6841 A1.n26 A1.t75 26.5955
R6842 A1.n28 A1.t80 26.5955
R6843 A1.n28 A1.t65 26.5955
R6844 A1.n30 A1.t72 26.5955
R6845 A1.n30 A1.t86 26.5955
R6846 A1.n32 A1.t126 26.5955
R6847 A1.n32 A1.t78 26.5955
R6848 A1.n34 A1.t118 26.5955
R6849 A1.n34 A1.t70 26.5955
R6850 A1.n121 A1.t94 26.5955
R6851 A1.n121 A1.t108 26.5955
R6852 A1.n122 A1.t119 26.5955
R6853 A1.n122 A1.t71 26.5955
R6854 A1.n123 A1.t115 26.5955
R6855 A1.n123 A1.t66 26.5955
R6856 A1.n125 A1.t107 26.5955
R6857 A1.n125 A1.t122 26.5955
R6858 A1.n127 A1.t120 26.5955
R6859 A1.n127 A1.t113 26.5955
R6860 A1.n129 A1.t111 26.5955
R6861 A1.n129 A1.t105 26.5955
R6862 A1.n131 A1.t88 26.5955
R6863 A1.n131 A1.t99 26.5955
R6864 A1.n133 A1.t97 26.5955
R6865 A1.n133 A1.t109 26.5955
R6866 A1.n109 A1.t22 24.9236
R6867 A1.n109 A1.t37 24.9236
R6868 A1.n96 A1.t19 24.9236
R6869 A1.n96 A1.t56 24.9236
R6870 A1.n97 A1.t46 24.9236
R6871 A1.n97 A1.t4 24.9236
R6872 A1.n99 A1.t2 24.9236
R6873 A1.n99 A1.t28 24.9236
R6874 A1.n101 A1.t58 24.9236
R6875 A1.n101 A1.t43 24.9236
R6876 A1.n103 A1.t13 24.9236
R6877 A1.n103 A1.t31 24.9236
R6878 A1.n105 A1.t29 24.9236
R6879 A1.n105 A1.t0 24.9236
R6880 A1.n107 A1.t50 24.9236
R6881 A1.n107 A1.t11 24.9236
R6882 A1.n54 A1.t48 24.9236
R6883 A1.n54 A1.t9 24.9236
R6884 A1.n41 A1.t62 24.9236
R6885 A1.n41 A1.t47 24.9236
R6886 A1.n42 A1.t7 24.9236
R6887 A1.n42 A1.t55 24.9236
R6888 A1.n44 A1.t34 24.9236
R6889 A1.n44 A1.t60 24.9236
R6890 A1.n46 A1.t1 24.9236
R6891 A1.n46 A1.t16 24.9236
R6892 A1.n48 A1.t14 24.9236
R6893 A1.n48 A1.t42 24.9236
R6894 A1.n50 A1.t40 24.9236
R6895 A1.n50 A1.t53 24.9236
R6896 A1.n52 A1.t27 24.9236
R6897 A1.n52 A1.t23 24.9236
R6898 A1.n15 A1.t49 24.9236
R6899 A1.n15 A1.t10 24.9236
R6900 A1.n2 A1.t63 24.9236
R6901 A1.n2 A1.t20 24.9236
R6902 A1.n3 A1.t18 24.9236
R6903 A1.n3 A1.t36 24.9236
R6904 A1.n5 A1.t45 24.9236
R6905 A1.n5 A1.t3 24.9236
R6906 A1.n7 A1.t32 24.9236
R6907 A1.n7 A1.t26 24.9236
R6908 A1.n9 A1.t57 24.9236
R6909 A1.n9 A1.t6 24.9236
R6910 A1.n11 A1.t12 24.9236
R6911 A1.n11 A1.t30 24.9236
R6912 A1.n13 A1.t38 24.9236
R6913 A1.n13 A1.t51 24.9236
R6914 A1.n154 A1.t25 24.9236
R6915 A1.n154 A1.t44 24.9236
R6916 A1.n140 A1.t5 24.9236
R6917 A1.n140 A1.t21 24.9236
R6918 A1.n141 A1.t61 24.9236
R6919 A1.n141 A1.t8 24.9236
R6920 A1.n143 A1.t17 24.9236
R6921 A1.n143 A1.t35 24.9236
R6922 A1.n145 A1.t33 24.9236
R6923 A1.n145 A1.t59 24.9236
R6924 A1.n147 A1.t54 24.9236
R6925 A1.n147 A1.t15 24.9236
R6926 A1.n149 A1.t24 24.9236
R6927 A1.n149 A1.t41 24.9236
R6928 A1.n151 A1.t39 24.9236
R6929 A1.n151 A1.t52 24.9236
R6930 A1 A1.n110 11.4429
R6931 A1 A1.n55 11.4429
R6932 A1 A1.n18 11.4429
R6933 A1.n37 A1.n22 8.55024
R6934 A1.n136 A1.n121 8.55024
R6935 A1.n74 A1.n59 8.55024
R6936 A1.n79 A1.n78 8.46262
R6937 A1.n16 A1.n15 7.77479
R6938 A1.n155 A1.n154 7.77479
R6939 A1.n95 A1.n94 4.6505
R6940 A1.n111 A1 3.29747
R6941 A1.n56 A1 3.29747
R6942 A1.n38 A1.n37 3.20821
R6943 A1.n137 A1.n136 3.2082
R6944 A1.n75 A1.n74 3.20156
R6945 A1.n19 A1 3.10353
R6946 A1 A1.n159 3.10353
R6947 A1.n17 A1.n1 3.1005
R6948 A1.n157 A1.n156 3.1005
R6949 A1.n94 A1.n93 2.71565
R6950 A1.n74 A1.n73 2.32777
R6951 A1.n37 A1.n36 2.32777
R6952 A1.n136 A1.n135 2.32777
R6953 A1.n110 A1 1.74595
R6954 A1.n55 A1 1.74595
R6955 A1.n117 A1.n116 1.07337
R6956 A1.n18 A1.n17 0.970197
R6957 A1.n156 A1.n153 0.970197
R6958 A1.n118 A1.n117 0.69375
R6959 A1.n119 A1.n118 0.68905
R6960 A1.n16 A1 0.649449
R6961 A1.n155 A1 0.649449
R6962 A1.n118 A1.n39 0.414635
R6963 A1.n117 A1.n76 0.382465
R6964 A1.n119 A1 0.378606
R6965 A1.n120 A1.n119 0.368576
R6966 A1.n94 A1.n79 0.207197
R6967 A1.n39 A1.n38 0.157252
R6968 A1.n137 A1.n120 0.139891
R6969 A1.n116 A1.n115 0.139389
R6970 A1.n76 A1.n75 0.132946
R6971 A1.n17 A1.n16 0.118507
R6972 A1.n156 A1.n155 0.118507
R6973 A1.n20 A1.n1 0.111611
R6974 A1.n158 A1.n157 0.111611
R6975 A1.n114 A1.n95 0.0991111
R6976 A1.n114 A1.n112 0.0296667
R6977 A1.n95 A1.n77 0.0282778
R6978 A1.n58 A1.n57 0.0227222
R6979 A1.n21 A1.n20 0.0171667
R6980 A1.n158 A1.n139 0.0171667
R6981 A1.n75 A1.n58 0.00100004
R6982 A1.n139 A1.n137 0.00100004
R6983 A1.n38 A1.n21 0.00100004
R6984 A1.n112 A1.n111 0.000513563
R6985 A1.n57 A1.n56 0.000513563
R6986 A1.n20 A1.n19 0.000513218
R6987 A1.n159 A1.n158 0.000513218
R6988 A1.n58 A1.n40 0.00050517
R6989 A1.n114 A1.n113 0.000504838
R6990 A1.n21 A1.n0 0.000504838
R6991 A1.n139 A1.n138 0.000504838
R6992 A1.n115 A1.n114 0.000501713
R6993 I15.n3 I15.t2 261.116
R6994 I15.n0 I15.t3 186.03
R6995 I15.n3 I15.t0 155.746
R6996 I15.n0 I15.t1 137.829
R6997 I15 I15.n0 78.5605
R6998 I15.n9 I15 47.2619
R6999 I15.n4 I15.n3 7.65549
R7000 I15.n9 I15.n8 4.04922
R7001 I15.n5 I15 2.46419
R7002 I15.n10 I15 0.893416
R7003 I15.n5 I15.n4 0.754023
R7004 I15 I15.n10 0.70184
R7005 I15.n10 I15.n9 0.585321
R7006 I15.n7 I15.n6 0.0326429
R7007 I15.n7 I15.n2 0.0197253
R7008 I15.n8 I15.n1 0.00182856
R7009 I15.n8 I15.n7 0.00149885
R7010 I15.n7 I15.n5 0.00125261
R7011 EI.n29 EI.t14 330.12
R7012 EI.n30 EI.t8 330.002
R7013 EI.n38 EI.t20 323.342
R7014 EI.n1 EI.t9 260.435
R7015 EI.n27 EI.t2 256.07
R7016 EI.n24 EI.t21 256.07
R7017 EI.n22 EI.t15 256.07
R7018 EI.n19 EI.t16 256.07
R7019 EI.n44 EI.t6 251.637
R7020 EI.n10 EI.t12 229.433
R7021 EI.n29 EI.t5 201.587
R7022 EI.n30 EI.t19 200.782
R7023 EI.n38 EI.t13 194.809
R7024 EI.n40 EI.t0 168.561
R7025 EI.n40 EI.t1 166.328
R7026 EI.n10 EI.t7 158.885
R7027 EI.n1 EI.t3 156.403
R7028 EI.n27 EI.t17 150.03
R7029 EI.n24 EI.t11 150.03
R7030 EI.n22 EI.t4 150.03
R7031 EI.n19 EI.t10 150.03
R7032 EI.n42 EI.t18 145.043
R7033 EI EI.n38 79.5475
R7034 EI EI.n29 78.5148
R7035 EI.n28 EI.n27 77.1383
R7036 EI.n25 EI.n24 76.0005
R7037 EI.n23 EI.n22 76.0005
R7038 EI.n20 EI.n19 76.0005
R7039 EI.n51 EI 26.615
R7040 EI.n55 EI.n21 22.5125
R7041 EI.n49 EI 17.4176
R7042 EI.n54 EI 14.551
R7043 EI.n53 EI.n26 13.4428
R7044 EI.n52 EI 13.4235
R7045 EI.n3 EI 9.58775
R7046 EI EI.n23 9.22489
R7047 EI.n41 EI.n40 9.0245
R7048 EI.n47 EI.n44 8.76429
R7049 EI.n23 EI 7.6805
R7050 EI.n2 EI.n1 7.60183
R7051 EI.n11 EI.n10 7.39171
R7052 EI.n31 EI.n30 7.27155
R7053 EI.n20 EI 6.73734
R7054 EI.n41 EI.n39 6.23487
R7055 EI.n47 EI 5.65631
R7056 EI.n26 EI 5.65631
R7057 EI.n21 EI 5.31371
R7058 EI.n48 EI.n47 4.99699
R7059 EI.n43 EI.n42 4.98671
R7060 EI EI.n2 4.8645
R7061 EI.n48 EI.n41 4.61128
R7062 EI.n44 EI.n43 4.43268
R7063 EI.n28 EI 4.26717
R7064 EI.n21 EI.n20 4.04261
R7065 EI.n33 EI.n32 3.88621
R7066 EI.n13 EI.n12 3.46717
R7067 EI.n14 EI.n13 3.03311
R7068 EI EI.n8 3.02091
R7069 EI EI.n28 2.13383
R7070 EI.n39 EI 2.11184
R7071 EI.n50 EI.n37 1.59861
R7072 EI.n25 EI 1.53093
R7073 EI.n56 EI.n55 1.43354
R7074 EI.n46 EI.n45 1.25267
R7075 EI.n50 EI.n49 1.21925
R7076 EI.n47 EI.n46 1.11354
R7077 EI.n26 EI.n25 1.11354
R7078 EI.n57 EI.n18 1.10387
R7079 EI.n56 EI 1.07862
R7080 EI.n13 EI.n11 1.06717
R7081 EI.n12 EI 1.06717
R7082 EI.n39 EI 0.970197
R7083 EI.n2 EI.n0 0.7685
R7084 EI.n33 EI.n31 0.686214
R7085 EI.n52 EI.n51 0.683536
R7086 EI.n53 EI.n52 0.571929
R7087 EI.n55 EI.n54 0.558536
R7088 EI.n54 EI.n53 0.549607
R7089 EI.n49 EI.n48 0.464786
R7090 EI.n32 EI 0.457643
R7091 EI.n57 EI.n56 0.424377
R7092 EI.n51 EI.n50 0.384429
R7093 EI.n45 EI 0.278761
R7094 EI EI.n57 0.0604792
R7095 EI.n35 EI.n34 0.0308571
R7096 EI.n8 EI.n7 0.0205312
R7097 EI.n18 EI.n16 0.0127256
R7098 EI.n16 EI.n14 0.0125192
R7099 EI.n4 EI.n3 0.0051875
R7100 EI.n16 EI.n15 0.00410577
R7101 EI.n14 EI.n9 0.00339649
R7102 EI.n7 EI.n6 0.00111657
R7103 EI.n18 EI.n17 0.00107203
R7104 EI.n37 EI.n36 0.00107006
R7105 EI.n6 EI.n5 0.00100057
R7106 EI.n36 EI.n35 0.00100008
R7107 EI.n35 EI.n33 0.000834423
R7108 EI.n7 EI.n4 0.000625544
R7109 EI.n4 EI.n0 0.000625542
R7110 I3.n3 I3.t1 334.723
R7111 I3.n2 I3.t2 323.342
R7112 I3.n3 I3.t4 206.19
R7113 I3.n2 I3.t0 194.809
R7114 I3.n0 I3.t5 186.03
R7115 I3.n0 I3.t3 137.829
R7116 I3 I3.n3 84.2291
R7117 I3 I3.n2 82.1338
R7118 I3.n1 I3.n0 76.0005
R7119 I3.n6 I3 66.7187
R7120 I3.n4 I3 26.4877
R7121 I3.n1 I3 7.31479
R7122 I3.n4 I3 4.36044
R7123 I3 I3.n1 4.02336
R7124 I3.n5 I3.n4 2.61211
R7125 I3.n6 I3.n5 1.25943
R7126 I3 I3.n6 0.969697
R7127 I3.n5 I3 0.522827
R7128 I1.t0 I1.t2 618.109
R7129 I1.n0 I1.t1 334.723
R7130 I1 I1.t0 253.56
R7131 I1.n0 I1.t3 206.19
R7132 I1 I1.n0 90.4462
R7133 I1.n3 I1 39.0702
R7134 I1.n1 I1 7.13193
R7135 I1.n1 I1 5.30336
R7136 I1.n2 I1.n1 5.16688
R7137 I1.n3 I1.n2 2.29514
R7138 I1 I1.n3 0.692911
R7139 I1.n2 I1 0.375952
R7140 A3.n134 A3.n132 145.809
R7141 A3.n83 A3.n81 145.809
R7142 A3.n45 A3.n43 145.809
R7143 A3.n23 A3.n21 145.809
R7144 A3.n83 A3.n82 107.409
R7145 A3.n85 A3.n84 107.409
R7146 A3.n87 A3.n86 107.409
R7147 A3.n89 A3.n88 107.409
R7148 A3.n91 A3.n90 107.409
R7149 A3.n93 A3.n92 107.409
R7150 A3.n45 A3.n44 107.409
R7151 A3.n47 A3.n46 107.409
R7152 A3.n49 A3.n48 107.409
R7153 A3.n51 A3.n50 107.409
R7154 A3.n53 A3.n52 107.409
R7155 A3.n55 A3.n54 107.409
R7156 A3.n23 A3.n22 107.409
R7157 A3.n25 A3.n24 107.409
R7158 A3.n27 A3.n26 107.409
R7159 A3.n29 A3.n28 107.409
R7160 A3.n31 A3.n30 107.409
R7161 A3.n33 A3.n32 107.409
R7162 A3.n134 A3.n133 107.407
R7163 A3.n136 A3.n135 107.407
R7164 A3.n138 A3.n137 107.407
R7165 A3.n140 A3.n139 107.407
R7166 A3.n142 A3.n141 107.407
R7167 A3.n144 A3.n143 107.407
R7168 A3.n152 A3.n150 87.1779
R7169 A3.n106 A3.n104 87.1779
R7170 A3.n64 A3.n62 87.1779
R7171 A3.n3 A3.n1 87.1779
R7172 A3.n152 A3.n151 52.82
R7173 A3.n154 A3.n153 52.82
R7174 A3.n156 A3.n155 52.82
R7175 A3.n158 A3.n157 52.82
R7176 A3.n160 A3.n159 52.82
R7177 A3.n162 A3.n161 52.82
R7178 A3.n106 A3.n105 52.82
R7179 A3.n108 A3.n107 52.82
R7180 A3.n110 A3.n109 52.82
R7181 A3.n112 A3.n111 52.82
R7182 A3.n114 A3.n113 52.82
R7183 A3.n116 A3.n115 52.82
R7184 A3.n64 A3.n63 52.82
R7185 A3.n66 A3.n65 52.82
R7186 A3.n68 A3.n67 52.82
R7187 A3.n70 A3.n69 52.82
R7188 A3.n72 A3.n71 52.82
R7189 A3.n74 A3.n73 52.82
R7190 A3.n3 A3.n2 52.82
R7191 A3.n5 A3.n4 52.82
R7192 A3.n7 A3.n6 52.82
R7193 A3.n9 A3.n8 52.82
R7194 A3.n11 A3.n10 52.82
R7195 A3.n13 A3.n12 52.82
R7196 A3.n136 A3.n134 38.4005
R7197 A3.n138 A3.n136 38.4005
R7198 A3.n140 A3.n138 38.4005
R7199 A3.n142 A3.n140 38.4005
R7200 A3.n144 A3.n142 38.4005
R7201 A3.n145 A3.n144 38.4005
R7202 A3.n85 A3.n83 38.4005
R7203 A3.n87 A3.n85 38.4005
R7204 A3.n89 A3.n87 38.4005
R7205 A3.n91 A3.n89 38.4005
R7206 A3.n93 A3.n91 38.4005
R7207 A3.n94 A3.n93 38.4005
R7208 A3.n47 A3.n45 38.4005
R7209 A3.n49 A3.n47 38.4005
R7210 A3.n51 A3.n49 38.4005
R7211 A3.n53 A3.n51 38.4005
R7212 A3.n55 A3.n53 38.4005
R7213 A3.n56 A3.n55 38.4005
R7214 A3.n25 A3.n23 38.4005
R7215 A3.n27 A3.n25 38.4005
R7216 A3.n29 A3.n27 38.4005
R7217 A3.n31 A3.n29 38.4005
R7218 A3.n33 A3.n31 38.4005
R7219 A3.n34 A3.n33 38.4005
R7220 A3.n154 A3.n152 34.3584
R7221 A3.n156 A3.n154 34.3584
R7222 A3.n158 A3.n156 34.3584
R7223 A3.n160 A3.n158 34.3584
R7224 A3.n162 A3.n160 34.3584
R7225 A3.n166 A3.n162 34.3584
R7226 A3.n108 A3.n106 34.3584
R7227 A3.n110 A3.n108 34.3584
R7228 A3.n112 A3.n110 34.3584
R7229 A3.n114 A3.n112 34.3584
R7230 A3.n116 A3.n114 34.3584
R7231 A3.n121 A3.n116 34.3584
R7232 A3.n66 A3.n64 34.3584
R7233 A3.n68 A3.n66 34.3584
R7234 A3.n70 A3.n68 34.3584
R7235 A3.n72 A3.n70 34.3584
R7236 A3.n74 A3.n72 34.3584
R7237 A3.n75 A3.n74 34.3584
R7238 A3.n5 A3.n3 34.3584
R7239 A3.n7 A3.n5 34.3584
R7240 A3.n9 A3.n7 34.3584
R7241 A3.n11 A3.n9 34.3584
R7242 A3.n13 A3.n11 34.3584
R7243 A3.n183 A3.n13 34.3584
R7244 A3.n127 A3.t105 26.5955
R7245 A3.n127 A3.t119 26.5955
R7246 A3.n132 A3.t82 26.5955
R7247 A3.n132 A3.t120 26.5955
R7248 A3.n133 A3.t78 26.5955
R7249 A3.n133 A3.t73 26.5955
R7250 A3.n135 A3.t118 26.5955
R7251 A3.n135 A3.t66 26.5955
R7252 A3.n137 A3.t64 26.5955
R7253 A3.n137 A3.t124 26.5955
R7254 A3.n139 A3.t122 26.5955
R7255 A3.n139 A3.t70 26.5955
R7256 A3.n141 A3.t115 26.5955
R7257 A3.n141 A3.t107 26.5955
R7258 A3.n143 A3.t110 26.5955
R7259 A3.n143 A3.t99 26.5955
R7260 A3.n81 A3.t112 26.5955
R7261 A3.n81 A3.t126 26.5955
R7262 A3.n82 A3.t104 26.5955
R7263 A3.n82 A3.t96 26.5955
R7264 A3.n84 A3.t95 26.5955
R7265 A3.n84 A3.t89 26.5955
R7266 A3.n86 A3.t87 26.5955
R7267 A3.n86 A3.t102 26.5955
R7268 A3.n88 A3.t86 26.5955
R7269 A3.n88 A3.t100 26.5955
R7270 A3.n90 A3.t76 26.5955
R7271 A3.n90 A3.t93 26.5955
R7272 A3.n92 A3.t91 26.5955
R7273 A3.n92 A3.t84 26.5955
R7274 A3.n43 A3.t68 26.5955
R7275 A3.n43 A3.t83 26.5955
R7276 A3.n44 A3.t67 26.5955
R7277 A3.n44 A3.t79 26.5955
R7278 A3.n46 A3.t77 26.5955
R7279 A3.n46 A3.t72 26.5955
R7280 A3.n48 A3.t71 26.5955
R7281 A3.n48 A3.t65 26.5955
R7282 A3.n50 A3.t108 26.5955
R7283 A3.n50 A3.t123 26.5955
R7284 A3.n52 A3.t121 26.5955
R7285 A3.n52 A3.t69 26.5955
R7286 A3.n54 A3.t114 26.5955
R7287 A3.n54 A3.t127 26.5955
R7288 A3.n17 A3.t90 26.5955
R7289 A3.n17 A3.t81 26.5955
R7290 A3.n21 A3.t97 26.5955
R7291 A3.n21 A3.t113 26.5955
R7292 A3.n22 A3.t111 26.5955
R7293 A3.n22 A3.t125 26.5955
R7294 A3.n24 A3.t103 26.5955
R7295 A3.n24 A3.t117 26.5955
R7296 A3.n26 A3.t94 26.5955
R7297 A3.n26 A3.t88 26.5955
R7298 A3.n28 A3.t116 26.5955
R7299 A3.n28 A3.t101 26.5955
R7300 A3.n30 A3.t85 26.5955
R7301 A3.n30 A3.t98 26.5955
R7302 A3.n32 A3.t75 26.5955
R7303 A3.n32 A3.t92 26.5955
R7304 A3.n38 A3.t109 25.6105
R7305 A3.n163 A3.t41 24.9236
R7306 A3.n163 A3.t55 24.9236
R7307 A3.n150 A3.t18 24.9236
R7308 A3.n150 A3.t56 24.9236
R7309 A3.n151 A3.t14 24.9236
R7310 A3.n151 A3.t9 24.9236
R7311 A3.n153 A3.t54 24.9236
R7312 A3.n153 A3.t2 24.9236
R7313 A3.n155 A3.t0 24.9236
R7314 A3.n155 A3.t60 24.9236
R7315 A3.n157 A3.t58 24.9236
R7316 A3.n157 A3.t6 24.9236
R7317 A3.n159 A3.t52 24.9236
R7318 A3.n159 A3.t43 24.9236
R7319 A3.n161 A3.t46 24.9236
R7320 A3.n161 A3.t34 24.9236
R7321 A3.n104 A3.t48 24.9236
R7322 A3.n104 A3.t62 24.9236
R7323 A3.n105 A3.t40 24.9236
R7324 A3.n105 A3.t32 24.9236
R7325 A3.n107 A3.t31 24.9236
R7326 A3.n107 A3.t25 24.9236
R7327 A3.n109 A3.t23 24.9236
R7328 A3.n109 A3.t38 24.9236
R7329 A3.n111 A3.t22 24.9236
R7330 A3.n111 A3.t36 24.9236
R7331 A3.n113 A3.t12 24.9236
R7332 A3.n113 A3.t29 24.9236
R7333 A3.n115 A3.t27 24.9236
R7334 A3.n115 A3.t20 24.9236
R7335 A3.n62 A3.t4 24.9236
R7336 A3.n62 A3.t19 24.9236
R7337 A3.n63 A3.t3 24.9236
R7338 A3.n63 A3.t15 24.9236
R7339 A3.n65 A3.t13 24.9236
R7340 A3.n65 A3.t8 24.9236
R7341 A3.n67 A3.t7 24.9236
R7342 A3.n67 A3.t1 24.9236
R7343 A3.n69 A3.t44 24.9236
R7344 A3.n69 A3.t59 24.9236
R7345 A3.n71 A3.t57 24.9236
R7346 A3.n71 A3.t5 24.9236
R7347 A3.n73 A3.t51 24.9236
R7348 A3.n73 A3.t63 24.9236
R7349 A3.n14 A3.t26 24.9236
R7350 A3.n14 A3.t17 24.9236
R7351 A3.n1 A3.t33 24.9236
R7352 A3.n1 A3.t49 24.9236
R7353 A3.n2 A3.t47 24.9236
R7354 A3.n2 A3.t61 24.9236
R7355 A3.n4 A3.t39 24.9236
R7356 A3.n4 A3.t53 24.9236
R7357 A3.n6 A3.t30 24.9236
R7358 A3.n6 A3.t24 24.9236
R7359 A3.n8 A3.t50 24.9236
R7360 A3.n8 A3.t37 24.9236
R7361 A3.n10 A3.t21 24.9236
R7362 A3.n10 A3.t35 24.9236
R7363 A3.n12 A3.t11 24.9236
R7364 A3.n12 A3.t28 24.9236
R7365 A3.n60 A3.t45 24.7196
R7366 A3.n97 A3.t80 24.6255
R7367 A3.n60 A3.t42 23.9564
R7368 A3.n119 A3.t16 23.1655
R7369 A3.n95 A3.t74 19.1164
R7370 A3.n118 A3.n117 13.8467
R7371 A3 A3.n166 11.4429
R7372 A3 A3.n121 11.4429
R7373 A3 A3.n75 11.4429
R7374 A3 A3.n183 11.4429
R7375 A3.n117 A3.t10 11.0774
R7376 A3.n39 A3.t106 10.8355
R7377 A3.n98 A3.n97 9.3005
R7378 A3.n102 A3.n101 9.3005
R7379 A3.n120 A3.n119 8.77252
R7380 A3.n128 A3.n127 8.76605
R7381 A3.n18 A3.n17 8.76605
R7382 A3.n42 A3.n41 8.70762
R7383 A3.n41 A3.n40 8.69892
R7384 A3.n164 A3.n163 7.87147
R7385 A3.n15 A3.n14 7.87147
R7386 A3.n40 A3.n39 7.77627
R7387 A3.n96 A3.n95 7.29637
R7388 A3.n61 A3.n60 6.88889
R7389 A3.n77 A3.n61 4.758
R7390 A3.n120 A3.n103 4.6505
R7391 A3.n99 A3.n98 4.6505
R7392 A3.n182 A3.n181 4.6505
R7393 A3.n36 A3.n35 4.6505
R7394 A3.n19 A3.n18 4.26717
R7395 A3.n167 A3 3.10353
R7396 A3.n122 A3 3.10353
R7397 A3.n76 A3 3.10353
R7398 A3 A3.n0 3.10353
R7399 A3.n165 A3.n149 3.1005
R7400 A3.n129 A3.n128 3.1005
R7401 A3.n147 A3.n146 3.1005
R7402 A3.n58 A3.n57 2.75
R7403 A3.n146 A3.n145 2.71565
R7404 A3.n98 A3.n94 2.71565
R7405 A3.n57 A3.n56 2.71565
R7406 A3.n35 A3.n34 2.71565
R7407 A3.n58 A3.n42 2.69896
R7408 A3.n97 A3.n96 1.9705
R7409 A3.n166 A3 1.74595
R7410 A3 A3.n165 1.74595
R7411 A3.n121 A3 1.74595
R7412 A3 A3.n120 1.74595
R7413 A3.n75 A3 1.74595
R7414 A3.n183 A3 1.74595
R7415 A3 A3.n182 1.74595
R7416 A3.n119 A3.n118 1.74224
R7417 A3.n173 A3.n172 0.810582
R7418 A3.n175 A3 0.696701
R7419 A3.n175 A3.n174 0.531962
R7420 A3.n174 A3.n173 0.531962
R7421 A3.n174 A3.n78 0.475506
R7422 A3 A3.n61 0.388379
R7423 A3.n165 A3.n164 0.300854
R7424 A3.n182 A3.n15 0.300854
R7425 A3.n176 A3.n175 0.275505
R7426 A3.n173 A3.n126 0.263005
R7427 A3.n172 A3.n171 0.1755
R7428 A3.n126 A3.n125 0.1755
R7429 A3.n177 A3.n176 0.1755
R7430 A3.n168 A3.n149 0.11675
R7431 A3.n123 A3.n103 0.11675
R7432 A3.n181 A3.n179 0.11675
R7433 A3.n124 A3.n99 0.10425
R7434 A3.n170 A3.n147 0.09175
R7435 A3.n178 A3.n36 0.09175
R7436 A3.n78 A3.n58 0.0855244
R7437 A3.n41 A3.n38 0.0578287
R7438 A3.n78 A3.n77 0.0505
R7439 A3.n147 A3.n131 0.04425
R7440 A3.n36 A3.n20 0.04425
R7441 A3.n99 A3.n80 0.043
R7442 A3.n103 A3.n102 0.03175
R7443 A3.n131 A3.n129 0.028
R7444 A3.n20 A3.n16 0.028
R7445 A3.n170 A3.n168 0.0255
R7446 A3.n149 A3.n148 0.0255
R7447 A3.n179 A3.n178 0.0255
R7448 A3.n181 A3.n180 0.0255
R7449 A3.n124 A3.n123 0.013
R7450 A3.n80 A3.n79 0.00450862
R7451 A3.n131 A3.n130 0.0025557
R7452 A3.n20 A3.n19 0.0025557
R7453 A3.n168 A3.n167 0.00053521
R7454 A3.n123 A3.n122 0.00053521
R7455 A3.n77 A3.n76 0.00053521
R7456 A3.n179 A3.n0 0.00053521
R7457 A3.n170 A3.n169 0.00050852
R7458 A3.n124 A3.n100 0.00050852
R7459 A3.n78 A3.n59 0.00050852
R7460 A3.n178 A3.n37 0.00050852
R7461 A3.n171 A3.n170 0.000500999
R7462 A3.n125 A3.n124 0.000500999
R7463 A3.n178 A3.n177 0.000500999
R7464 I14.n16 I14.t1 260.435
R7465 I14.n2 I14.t5 229.433
R7466 I14.n11 I14.t0 196.549
R7467 I14.n2 I14.t3 158.885
R7468 I14.n16 I14.t4 156.403
R7469 I14.n11 I14.t2 148.35
R7470 I14.n12 I14.n11 76.0005
R7471 I14 I14.n15 9.3005
R7472 I14.n17 I14.n16 7.60183
R7473 I14.n3 I14.n2 7.39171
R7474 I14.n21 I14.n13 6.24391
R7475 I14.n12 I14 5.78114
R7476 I14.n17 I14 4.8645
R7477 I14.n6 I14.n5 4.5005
R7478 I14.n21 I14.n20 3.53643
R7479 I14.n13 I14.n12 3.51018
R7480 I14.n5 I14.n4 3.46717
R7481 I14.n23 I14.n10 1.11384
R7482 I14.n5 I14.n3 1.06717
R7483 I14.n4 I14 1.06717
R7484 I14.n23 I14.n22 0.767464
R7485 I14.n22 I14 0.736889
R7486 I14 I14.n23 0.372375
R7487 I14.n22 I14.n21 0.321929
R7488 I14.n13 I14 0.206952
R7489 I14.n19 I14.n15 0.0344286
R7490 I14.n10 I14.n9 0.028
R7491 I14.n8 I14.n7 0.0142363
R7492 I14.n8 I14.n6 0.00599451
R7493 I14.n1 I14.n0 0.00484776
R7494 I14.n6 I14.n1 0.00226981
R7495 I14.n20 I14.n14 0.00182856
R7496 I14.n20 I14.n19 0.00149885
R7497 I14.n18 I14.n17 0.00133362
R7498 I14.n19 I14.n18 0.00100077
R7499 I14.n9 I14.n8 0.000617139
R7500 I4.n12 I4.t5 260.435
R7501 I4.n2 I4.t3 230.576
R7502 I4.n5 I4.t2 196.549
R7503 I4.n2 I4.t1 158.275
R7504 I4.n12 I4.t0 156.403
R7505 I4.n5 I4.t4 148.35
R7506 I4.n6 I4.n5 9.49829
R7507 I4.n3 I4.n2 8.76429
R7508 I4.n7 I4.n6 7.9582
R7509 I4.n4 I4.n3 7.74345
R7510 I4.n13 I4.n12 7.60183
R7511 I4.n3 I4 6.66717
R7512 I4.n6 I4 6.44139
R7513 I4 I4.n13 4.8645
R7514 I4.n9 I4.n8 2.33148
R7515 I4.n7 I4.n4 1.0005
R7516 I4.n8 I4 0.591367
R7517 I4.n8 I4.n7 0.446956
R7518 I4.n4 I4 0.380411
R7519 I4.n10 I4.n0 0.0344286
R7520 I4.n9 I4.n1 0.00182856
R7521 I4.n10 I4.n9 0.00149885
R7522 I4.n13 I4.n11 0.00133362
R7523 I4.n11 I4.n10 0.00100077
R7524 I10.n4 I10.t5 323.342
R7525 I10.n0 I10.t3 228.927
R7526 I10.n2 I10.t4 196.549
R7527 I10.n4 I10.t2 194.809
R7528 I10.n0 I10.t1 159.391
R7529 I10.n2 I10.t0 148.35
R7530 I10.n5 I10.n4 76.0005
R7531 I10.n3 I10.n2 76.0005
R7532 I10.n6 I10.n5 29.3651
R7533 I10.n7 I10 9.11
R7534 I10.n1 I10.n0 8.68501
R7535 I10.n3 I10 5.78114
R7536 I10.n8 I10.n1 4.26764
R7537 I10 I10.n3 3.71663
R7538 I10.n1 I10 1.99697
R7539 I10.n5 I10 1.92927
R7540 I10.n7 I10.n6 1.69246
R7541 I10.n8 I10.n7 0.570143
R7542 I10.n6 I10 0.457435
R7543 I10 I10.n8 0.221483
R7544 I9.t2 I9.t1 618.109
R7545 I9.n0 I9.t3 334.723
R7546 I9 I9.t2 253.56
R7547 I9.n0 I9.t0 206.19
R7548 I9 I9.n0 90.4462
R7549 I9.n3 I9 39.0702
R7550 I9.n1 I9 7.13193
R7551 I9.n1 I9 5.30336
R7552 I9.n2 I9.n1 5.27402
R7553 I9.n3 I9.n2 2.188
R7554 I9 I9.n3 0.692911
R7555 I9.n2 I9 0.369702
R7556 I0.n0 I0.t1 196.549
R7557 I0.n0 I0.t0 148.35
R7558 I0.n1 I0.n0 9.49592
R7559 I0.n2 I0.n1 7.58085
R7560 I0.n1 I0 6.44187
R7561 I0.n2 I0 2.72484
R7562 I0 I0.n2 0.88934
R7563 I7.n3 I7.t3 261.116
R7564 I7.n0 I7.t0 186.03
R7565 I7.n3 I7.t2 155.746
R7566 I7.n0 I7.t1 137.829
R7567 I7 I7.n0 78.5605
R7568 I7.n9 I7 47.2619
R7569 I7.n4 I7.n3 7.65549
R7570 I7.n9 I7.n8 4.04922
R7571 I7.n5 I7 2.46419
R7572 I7.n10 I7 0.899666
R7573 I7 I7.n10 0.808983
R7574 I7.n5 I7.n4 0.754023
R7575 I7.n10 I7.n9 0.478179
R7576 I7.n7 I7.n6 0.0326429
R7577 I7.n7 I7.n2 0.0197253
R7578 I7.n8 I7.n1 0.00182856
R7579 I7.n8 I7.n7 0.00149885
R7580 I7.n7 I7.n5 0.00125261
R7581 I5.t1 I5.t3 618.109
R7582 I5.n12 I5.t2 259.74
R7583 I5 I5.t1 253.56
R7584 I5.n3 I5.t4 228.899
R7585 I5.n18 I5.t5 180.286
R7586 I5.n3 I5.t0 159.411
R7587 I5.n12 I5.t7 157.083
R7588 I5.n20 I5.n19 152
R7589 I5.n20 I5.t6 111.091
R7590 I5.n18 I5.n17 74.4551
R7591 I5 I5.n24 37.6855
R7592 I5.n6 I5.n2 9.3005
R7593 I5.n6 I5.n5 9.3005
R7594 I5.n21 I5.n20 9.3005
R7595 I5.n14 I5 9.3005
R7596 I5.n22 I5.n21 7.80966
R7597 I5.n13 I5.n12 7.57248
R7598 I5.n5 I5.n3 7.36978
R7599 I5.n20 I5.n18 6.53562
R7600 I5 I5.n13 4.8645
R7601 I5.n14 I5.n10 4.50988
R7602 I5.n4 I5.n2 3.46717
R7603 I5.n4 I5.n1 3.03286
R7604 I5.n19 I5.n17 2.32777
R7605 I5.n8 I5.n0 2.26553
R7606 I5.n7 I5.n1 2.26468
R7607 I5.n16 I5.n15 2.251
R7608 I5.n22 I5.n16 2.19001
R7609 I5.n19 I5 1.4966
R7610 I5.n23 I5.n9 1.36032
R7611 I5.n23 I5.n22 1.07639
R7612 I5.n5 I5.n4 1.06717
R7613 I5.n2 I5 1.06717
R7614 I5.n9 I5.n8 0.71595
R7615 I5.n24 I5 0.657683
R7616 I5.n21 I5.n17 0.499201
R7617 I5.n9 I5 0.221483
R7618 I5.n15 I5.n14 0.0301875
R7619 I5.n16 I5.n10 0.0205312
R7620 I5.n6 I5.n0 0.00618182
R7621 I5.n1 I5.n0 0.00555107
R7622 I5.n7 I5.n6 0.00530477
R7623 I5.n11 I5.n10 0.00210765
R7624 I5.n13 I5.n11 0.00133438
R7625 I5.n8 I5.n7 0.00101192
R7626 I5.n15 I5.n11 0.00100001
R7627 I5.n24 I5.n23 0.000507778
R7628 I13.t6 I13.t0 618.109
R7629 I13.n11 I13.t7 259.74
R7630 I13 I13.t6 253.56
R7631 I13.n0 I13.t4 228.899
R7632 I13.n18 I13.t5 180.286
R7633 I13.n0 I13.t2 159.411
R7634 I13.n11 I13.t1 157.083
R7635 I13.n19 I13.t3 111.091
R7636 I13.n22 I13 37.7071
R7637 I13.n20 I13.n19 9.3005
R7638 I13 I13.n10 9.3005
R7639 I13.n21 I13.n20 7.80966
R7640 I13.n12 I13.n11 7.57248
R7641 I13.n1 I13.n0 7.36978
R7642 I13.n19 I13.n18 6.53562
R7643 I13.n12 I13 4.8645
R7644 I13.n3 I13.n2 3.46717
R7645 I13.n4 I13.n3 3.03286
R7646 I13.n17 I13.n16 2.32777
R7647 I13.n21 I13.n15 2.19001
R7648 I13.n16 I13 1.4966
R7649 I13.n24 I13.n23 1.16836
R7650 I13.n22 I13.n21 1.07639
R7651 I13.n3 I13.n1 1.06717
R7652 I13.n2 I13 1.06717
R7653 I13.n24 I13.n8 0.71595
R7654 I13.n23 I13 0.663452
R7655 I13.n20 I13.n17 0.499201
R7656 I13 I13.n24 0.221483
R7657 I13.n23 I13.n22 0.192464
R7658 I13.n10 I13.n9 0.0301875
R7659 I13.n15 I13.n14 0.0205312
R7660 I13.n6 I13.n5 0.00618182
R7661 I13.n5 I13.n4 0.00555107
R7662 I13.n7 I13.n6 0.00530477
R7663 I13.n14 I13.n13 0.00210765
R7664 I13.n13 I13.n12 0.00133438
R7665 I13.n8 I13.n7 0.00101192
R7666 I13.n13 I13.n9 0.00100001
R7667 I8.n0 I8.t0 196.549
R7668 I8.n0 I8.t1 148.35
R7669 I8.n1 I8.n0 9.49592
R7670 I8.n2 I8.n1 7.58085
R7671 I8.n1 I8 6.44187
R7672 I8.n2 I8 2.61769
R7673 I8 I8.n2 0.88934
R7674 I6.n16 I6.t1 260.435
R7675 I6.n2 I6.t5 229.433
R7676 I6.n11 I6.t0 196.549
R7677 I6.n2 I6.t2 158.885
R7678 I6.n16 I6.t4 156.403
R7679 I6.n11 I6.t3 148.35
R7680 I6.n12 I6.n11 76.0005
R7681 I6 I6.n15 9.3005
R7682 I6.n17 I6.n16 7.60183
R7683 I6.n3 I6.n2 7.39171
R7684 I6.n21 I6.n13 6.24391
R7685 I6.n12 I6 5.78114
R7686 I6.n17 I6 4.8645
R7687 I6.n6 I6.n5 4.5005
R7688 I6.n21 I6.n20 3.53643
R7689 I6.n13 I6.n12 3.51018
R7690 I6.n5 I6.n4 3.46717
R7691 I6.n23 I6.n10 1.11384
R7692 I6.n5 I6.n3 1.06717
R7693 I6.n4 I6 1.06717
R7694 I6.n23 I6.n22 0.874607
R7695 I6.n22 I6 0.743139
R7696 I6 I6.n23 0.372375
R7697 I6.n22 I6.n21 0.214786
R7698 I6.n13 I6 0.206952
R7699 I6.n19 I6.n15 0.0344286
R7700 I6.n10 I6.n9 0.028
R7701 I6.n8 I6.n7 0.0142363
R7702 I6.n8 I6.n6 0.00599451
R7703 I6.n1 I6.n0 0.00484776
R7704 I6.n6 I6.n1 0.00226981
R7705 I6.n20 I6.n14 0.00182856
R7706 I6.n20 I6.n19 0.00149885
R7707 I6.n18 I6.n17 0.00133362
R7708 I6.n19 I6.n18 0.00100077
R7709 I6.n9 I6.n8 0.000617139
R7710 I11.n3 I11.t3 334.723
R7711 I11.n2 I11.t0 323.342
R7712 I11.n3 I11.t2 206.19
R7713 I11.n2 I11.t4 194.809
R7714 I11.n0 I11.t1 186.03
R7715 I11.n0 I11.t5 137.829
R7716 I11 I11.n3 84.2291
R7717 I11 I11.n2 82.1338
R7718 I11.n1 I11.n0 76.0005
R7719 I11.n6 I11 66.7187
R7720 I11.n4 I11 26.4877
R7721 I11.n1 I11 7.31479
R7722 I11.n4 I11 4.36044
R7723 I11 I11.n1 4.02336
R7724 I11.n5 I11.n4 2.71925
R7725 I11.n6 I11.n5 1.15229
R7726 I11 I11.n6 0.969697
R7727 I11.n5 I11 0.516577
C0 VDD I3 0.476f
C1 I11 I8 0.659f
C2 x43.A x43.Y 1.52f
C3 VDD x3.x21.B 0.713f
C4 I0 x3.x16.C 0.12f
C5 x3.EI x3.GS 0.123f
C6 a_5475_n13205# x3.x16.X 0.0121f
C7 x3.x18.C I1 0.495f
C8 I5 I13 0.0641f
C9 VDD a_5967_n7607# 0.222f
C10 I1 I3 1.71f
C11 I6 I0 0.342f
C12 x3.x22.A x3.x16.X 0.0732f
C13 x5.x15.X x1.A 0.0206f
C14 VDD I11 0.475f
C15 x3.EO x3.GS 0.9f
C16 I5 x3.x22.A 0.066f
C17 x5.x21.B EI 0.187f
C18 a_5475_n1939# x5.x2.X 0.134f
C19 a_5475_n7635# I13 0.193f
C20 I7 I4 0.767f
C21 x3.A1 x3.x16.X 0.0159f
C22 x3.A2 x3.EO 0.162f
C23 VDD a_6519_n9437# 0.233f
C24 I13 x5.x18.C 0.3f
C25 x5.x22.A x5.x16.X 0.0732f
C26 x3.EI x3.x18.C 1.56f
C27 x3.x19.C x3.x16.C 1.95f
C28 EI I15 4.8f
C29 a_5475_n1175# x5.x2.X 0.0313f
C30 x5.x21.B x5.x19.X 0.262f
C31 x3.EI a_5507_n11927# 0.0878f
C32 x3.EI I3 1.97f
C33 x5.x22.A x5.x19.D 0.0292f
C34 I6 x3.x19.C 0.304f
C35 I6 x3.x17.A 0.0474f
C36 I13 x5.x19.D 0.551f
C37 I10 x5.x16.C 0.925f
C38 x3.EI x3.x21.B 0.187f
C39 x3.x22.A x3.x21.X 0.0749f
C40 x5.x19.X x5.x21.X 0.131f
C41 a_6395_n7385# x5.x20.X 0.0765f
C42 VDD x3.x16.C 0.663f
C43 VDD a_5509_n12251# 0.221f
C44 a_5967_n15647# x3.x21.X 0.109f
C45 x3.x19.X x3.x20.X 0.145f
C46 a_5475_n6649# x5.x19.D 0.148f
C47 I12 I11 1.58f
C48 a_5475_n14689# x3.x19.D 0.148f
C49 VDD I6 0.634f
C50 VDD x35.A 0.537f
C51 I9 I11 1.72f
C52 I8 a_5475_n1175# 0.211f
C53 I2 x3.x19.D 0.196f
C54 I1 x3.x16.C 0.0914f
C55 VDD x5.x20.X 0.251f
C56 a_5475_n5165# I10 0.167f
C57 x5.x22.A x5.x17.A 1.27f
C58 x5.x14.A x5.x17.A 0.105f
C59 VDD a_5475_n1939# 0.153f
C60 I6 I1 0.257f
C61 x5.A2 x1.A 0.38f
C62 x3.EI a_6519_n9437# 0.181f
C63 I13 I8 0.323f
C64 x5.x22.A a_6395_n7385# 0.209f
C65 VDD a_5475_n1175# 0.148f
C66 x5.GS x42.A 0.098f
C67 a_5475_n13205# x3.x19.C 0.173f
C68 x5.x16.X x5.x16.C 0.07f
C69 x5.x21.B x5.x21.X 0.0197f
C70 x5.x4.A x5.EO 0.0491f
C71 x3.x15.X x3.x16.X 0.253f
C72 x3.EI x3.x16.C 2.08f
C73 x3.EI a_5509_n12251# 0.088f
C74 a_6519_n9437# x3.EO 0.135f
C75 I10 EI 1.27f
C76 a_6029_n9459# x3.x1.X 0.192f
C77 x5.x16.X a_5475_n5415# 0.102f
C78 a_5475_n14689# x3.x19.X 0.0873f
C79 VDD x5.x22.A 2.77f
C80 VDD x5.x14.A 0.437f
C81 x3.x22.A x3.x17.A 1.27f
C82 x3.x14.A x3.x17.A 0.105f
C83 x5.x16.C x5.x19.D 1.24f
C84 VDD I13 0.839f
C85 x3.EI I6 2.13f
C86 a_6395_n7385# x2.A 0.148f
C87 a_5475_n1939# I12 0.208f
C88 x1.X x28.A 0.0747f
C89 VDD a_5475_n13205# 0.423f
C90 x3.x20.X x3.x21.X 0.122f
C91 I11 x5.x19.C 0.921f
C92 x5.A2 a_10776_n5725# 0.208f
C93 VDD a_5475_n6649# 0.434f
C94 a_5507_n2647# x5.x14.A 0.135f
C95 A0 x22.Y 8.67f
C96 VDD x3.x22.A 2.78f
C97 VDD x3.x14.A 0.439f
C98 a_5475_n5165# x5.x16.X 0.0121f
C99 VDD x29.A 1.5f
C100 x3.A1 x3.x17.A 0.115f
C101 VDD a_5967_n15647# 0.219f
C102 I9 a_5475_n1175# 0.159f
C103 VDD a_5509_n4211# 0.221f
C104 VDD x2.A 1.26f
C105 A3 x43.Y 7.92f
C106 I5 I2 0.645f
C107 VDD x3.A1 1.58f
C108 x2.A x21.A 0.0121f
C109 x5.x14.A I12 0.0493f
C110 a_5475_n7635# EI 0.343f
C111 I8 x5.x16.C 0.12f
C112 x36.A x36.Y 1.51f
C113 I12 I13 2.92f
C114 VDD a_6519_n1397# 0.233f
C115 EI x5.x18.C 1.56f
C116 I13 I9 0.375f
C117 x3.x4.A a_5475_n9215# 0.0112f
C118 x3.EI x5.x22.A 0.208f
C119 x3.x19.D x3.x2.X 0.014f
C120 x3.EI x5.x14.A 0.0145f
C121 x5.x16.X EI 0.076f
C122 a_5507_n10687# x3.x14.A 0.135f
C123 VDD x3.x1.X 0.389f
C124 I6 a_5475_n9979# 0.214f
C125 x22.A x22.Y 1.51f
C126 VDD x5.GS 0.706f
C127 EI x5.x19.D 1.93f
C128 x3.EI a_5475_n13205# 0.122f
C129 x5.x11.X a_5935_n3179# 0.202f
C130 VDD x5.x16.C 0.663f
C131 x3.EI x3.x22.A 0.0483f
C132 x3.EI x3.x14.A 0.0111f
C133 VDD a_5475_n5415# 0.426f
C134 I3 x3.x4.A 0.0406f
C135 x3.EI a_5967_n15647# 0.106f
C136 I14 I11 0.78f
C137 x3.x22.A x3.A0 0.132f
C138 x3.EI x2.A 0.645f
C139 x5.x19.X x5.x19.D 0.0195f
C140 a_5507_n2957# x5.x11.X 0.109f
C141 x3.x19.X x3.x19.D 0.0195f
C142 x5.x16.X x1.A 0.0159f
C143 x5.x15.X x5.x16.X 0.253f
C144 x3.x18.C I4 0.432f
C145 x2.A x3.A0 0.398f
C146 I10 I15 0.444f
C147 VDD a_10776_n9865# 0.178f
C148 VDD x3.x20.X 0.242f
C149 I0 I2 2.43f
C150 I3 I4 1.6f
C151 VDD A1 6.55f
C152 x5.x17.A EI 0.02f
C153 VDD a_5475_n5165# 0.423f
C154 x3.x17.A x3.x15.X 0.0789f
C155 x29.Y x29.A 1.51f
C156 x3.x11.X a_5935_n11219# 0.202f
C157 x2.A x3.EO 0.02f
C158 EI I8 0.365f
C159 x3.x18.C I7 0.229f
C160 I3 I7 1.25f
C161 x5.x17.A a_5507_n3887# 0.14f
C162 I13 x5.x19.C 0.407f
C163 I12 x5.x16.C 0.202f
C164 x3.x22.A a_6219_n12955# 0.17f
C165 VDD x3.x15.X 0.239f
C166 I9 x5.x16.C 0.0914f
C167 x3.A2 a_5935_n11219# 0.144f
C168 a_5507_n10997# x3.x11.X 0.109f
C169 I5 x3.x19.D 0.551f
C170 a_5475_n6649# x5.x19.C 0.102f
C171 x5.x21.B x5.x18.C 0.014f
C172 x5.x17.A x1.A 0.115f
C173 x5.x17.A x5.x15.X 0.0789f
C174 a_5475_n14689# x3.x19.C 0.102f
C175 x3.x22.A a_6395_n15425# 0.209f
C176 x5.x1.X x5.x2.X 0.129f
C177 x5.x21.B x5.x16.X 0.0218f
C178 x5.x19.X a_6395_n7385# 0.193f
C179 VDD EI 2.3f
C180 I2 x3.x19.C 0.447f
C181 a_5475_n15675# x3.x20.X 0.0895f
C182 x3.A1 a_6219_n12955# 0.151f
C183 a_5475_n1939# I14 0.214f
C184 a_5475_n14437# x3.x19.D 0.14f
C185 x5.x21.B x5.x19.D 0.151f
C186 VDD x36.A 1.51f
C187 I15 x5.x18.C 0.229f
C188 x3.EI x3.x20.X 0.208f
C189 VDD a_5475_n14689# 0.434f
C190 VDD a_5507_n3887# 0.223f
C191 a_5507_n2647# EI 0.0883f
C192 VDD I2 0.448f
C193 x3.x20.X x3.A0 0.0149f
C194 VDD x5.x19.X 0.898f
C195 I15 x5.x19.D 0.244f
C196 I4 x3.x16.C 0.202f
C197 VDD x1.A 1.84f
C198 VDD x5.x15.X 0.239f
C199 I6 I4 2.38f
C200 I1 I2 3.98f
C201 x5.x22.A I14 0.0536f
C202 x3.EI x3.x15.X 0.0245f
C203 I15 x5.x2.X 0.0129f
C204 I13 I14 4.48f
C205 I12 EI 1.81f
C206 A1 x29.Y 8.66f
C207 x5.GS x43.A 0.0166f
C208 I0 x3.x19.D 0.122f
C209 I7 x3.x16.C 0.26f
C210 I7 a_5509_n12251# 0.192f
C211 EI I9 0.403f
C212 x5.x19.C x5.x16.C 1.95f
C213 x5.x22.A a_6219_n4915# 0.17f
C214 a_5475_n5415# x5.x19.C 0.176f
C215 x3.EI EI 0.791f
C216 VDD x5.x1.X 0.389f
C217 a_6029_n9459# x3.x2.X 0.121f
C218 I6 I7 2.18f
C219 I0 x3.x2.X 0.0265f
C220 a_6395_n7385# x5.x21.X 0.202f
C221 I8 I15 0.341f
C222 x3.EI a_5475_n14689# 0.175f
C223 x5.x17.A x5.A2 0.047f
C224 a_6395_n15425# x3.x20.X 0.0765f
C225 x3.x19.X x3.x21.X 0.131f
C226 x3.EI I2 1.27f
C227 a_5475_n5165# x5.x19.C 0.173f
C228 VDD x5.x21.B 0.716f
C229 VDD a_10776_n5725# 0.18f
C230 I10 x5.x18.C 0.341f
C231 a_6219_n12955# x3.x15.X 0.219f
C232 x3.x19.C x3.x19.D 0.996f
C233 x3.EI x1.A 0.534f
C234 VDD x5.x21.X 0.506f
C235 VDD I15 0.204f
C236 I10 x5.x19.D 0.196f
C237 x3.x16.X a_5475_n13455# 0.102f
C238 I11 x5.x4.A 0.0406f
C239 VDD x3.x19.D 1.27f
C240 x3.x14.A I4 0.0493f
C241 VDD x5.A2 2.06f
C242 EI x5.x19.C 1.71f
C243 I14 x5.x16.C 0.491f
C244 VDD x3.x2.X 0.361f
C245 x34.A x35.A 0.0737f
C246 a_6519_n1397# x5.EO 0.135f
C247 I1 x3.x19.D 0.937f
C248 VDD x2.X 0.35f
C249 a_6029_n1419# x5.x1.X 0.192f
C250 I7 x3.x22.A 0.0853f
C251 x5.x14.A a_5935_n3179# 0.197f
C252 x5.x22.A a_5935_n3179# 0.077f
C253 x3.x4.A x3.x1.X 0.118f
C254 I5 I0 0.321f
C255 x5.EO x5.GS 0.927f
C256 x2.X x21.A 0.0749f
C257 I3 a_5475_n9215# 0.0597f
C258 I12 I15 0.784f
C259 a_10776_n9865# x1.X 0.12f
C260 I10 I8 2.42f
C261 I9 I15 0.29f
C262 a_5475_n7635# x5.x19.D 0.0838f
C263 a_5507_n2957# x5.x22.A 0.0288f
C264 a_5475_n15675# x3.x19.D 0.0838f
C265 a_5507_n2957# I13 0.194f
C266 x5.x18.C x5.x19.D 0.491f
C267 x3.x18.C I3 0.251f
C268 VDD x3.x19.X 0.891f
C269 x3.EI x3.x19.D 1.93f
C270 a_6519_n9437# x3.GS 0.136f
C271 x3.x17.A x3.x16.X 0.0198f
C272 x3.EI x5.A2 0.507f
C273 x3.x18.C x3.x21.B 0.014f
C274 x3.x22.A a_5935_n11219# 0.077f
C275 x3.x14.A a_5935_n11219# 0.197f
C276 VDD I10 0.448f
C277 I3 x3.x21.B 0.0112f
C278 x2.A a_10776_n13515# 0.207f
C279 I5 x3.x19.C 0.407f
C280 I14 EI 2.22f
C281 VDD x3.x16.X 0.465f
C282 x5.x19.D x5.x2.X 0.014f
C283 x5.x4.A a_5475_n1175# 0.0112f
C284 a_5507_n10997# x3.x22.A 0.0288f
C285 a_5475_n14437# x3.x19.C 0.157f
C286 x5.x21.B x5.x19.C 0.0127f
C287 x5.x17.A x5.x16.X 0.0198f
C288 a_5507_n3887# I14 0.186f
C289 VDD I5 0.828f
C290 I8 x5.x18.C 0.119f
C291 x3.x2.X x3.EO 0.0749f
C292 I13 x5.x4.A 0.0107f
C293 VDD x36.Y 16.6f
C294 VDD a_5475_n14437# 0.428f
C295 EI x5.EO 0.18f
C296 I8 x5.x19.D 0.122f
C297 x3.EI x3.x19.X 0.0149f
C298 I15 x5.x19.C 0.239f
C299 a_5475_n13455# x3.x19.C 0.176f
C300 I10 I12 0.838f
C301 I5 I1 0.375f
C302 x1.A x1.X 0.0412f
C303 VDD a_5475_n7635# 0.205f
C304 x3.x19.X x3.A0 0.0123f
C305 I10 I9 3.97f
C306 x5.x11.X x5.x22.A 0.0936f
C307 x5.x14.A x5.x11.X 0.0721f
C308 a_6219_n4915# x1.A 0.151f
C309 a_6219_n4915# x5.x15.X 0.219f
C310 I8 x5.x2.X 0.0265f
C311 x5.x11.X I13 0.0201f
C312 I2 x3.x4.A 0.0109f
C313 VDD x5.x18.C 0.547f
C314 VDD x3.x21.X 0.501f
C315 I1 a_5475_n14437# 0.147f
C316 VDD x5.x16.X 0.463f
C317 VDD a_5475_n13455# 0.426f
C318 I0 x3.x19.C 0.12f
C319 I3 x3.x16.C 0.132f
C320 VDD x42.A 0.536f
C321 x3.x2.X a_5475_n9979# 0.134f
C322 x3.x18.C I6 0.3f
C323 x3.EI x3.x16.X 0.076f
C324 I5 a_5475_n15675# 0.193f
C325 I6 a_5507_n11927# 0.186f
C326 VDD x5.x19.D 1.28f
C327 I6 I3 0.6f
C328 I2 I4 0.839f
C329 VDD a_6029_n9459# 0.15f
C330 x3.EI I5 3.69f
C331 VDD I0 0.0984f
C332 VDD x5.x2.X 0.361f
C333 x3.x11.X x3.x22.A 0.0936f
C334 x3.x14.A x3.x11.X 0.0721f
C335 I7 I2 0.468f
C336 x28.A x29.A 0.392f
C337 a_5967_n7607# x5.x20.X 0.137f
C338 I1 I0 2.1f
C339 I12 x5.x18.C 0.432f
C340 x3.x19.X a_6395_n15425# 0.193f
C341 VDD x5.x17.A 1.17f
C342 x2.A x3.GS 0.0652f
C343 I14 I15 2.16f
C344 I9 x5.x18.C 0.495f
C345 x3.A2 x3.x14.A 0.074f
C346 x3.A2 x3.x22.A 0.0408f
C347 VDD I8 0.0984f
C348 I12 x5.x19.D 0.206f
C349 I10 x5.x19.C 0.447f
C350 a_6219_n12955# x3.x16.X 0.0673f
C351 x3.EI a_5475_n13455# 0.14f
C352 a_5507_n2957# EI 0.0829f
C353 VDD a_6395_n7385# 0.158f
C354 x3.A2 x2.A 0.401f
C355 I9 x5.x19.D 0.937f
C356 VDD x3.x17.A 1.17f
C357 VDD x3.x19.C 1f
C358 I12 x5.x2.X 0.0262f
C359 x3.A2 x3.A1 0.787f
C360 I11 a_5475_n1175# 0.0597f
C361 x3.EI I0 0.365f
C362 I5 a_5475_n9979# 0.16f
C363 I6 x3.x16.C 0.491f
C364 I1 x3.x19.C 0.347f
C365 a_5475_n6397# x5.x21.B 0.116f
C366 x3.x19.D x3.x4.A 0.0516f
C367 x3.x22.A x3.x21.B 0.064f
C368 x5.A2 x5.EO 0.136f
C369 a_6029_n1419# x5.x2.X 0.121f
C370 a_5967_n15647# x3.x21.B 0.186f
C371 VDD x21.A 0.537f
C372 I12 I8 0.553f
C373 I13 I11 1.27f
C374 a_6029_n9459# x3.EO 0.128f
C375 x3.EI x5.x17.A 0.0296f
C376 x3.x4.A x3.x2.X 0.125f
C377 a_5475_n9215# x3.x1.X 0.0991f
C378 VDD I1 1.21f
C379 VDD a_5507_n2647# 0.227f
C380 I9 I8 2.06f
C381 I4 x3.x19.D 0.206f
C382 EI x5.x4.A 0.547f
C383 a_5475_n6649# I11 0.15f
C384 x5.x18.C x5.x19.C 2.6f
C385 a_6395_n15425# x3.x21.X 0.202f
C386 I4 x3.x2.X 0.0262f
C387 x3.EI x3.x19.C 1.71f
C388 x3.EI x3.x17.A 0.02f
C389 I10 I14 0.441f
C390 VDD a_5507_n10687# 0.227f
C391 x42.A x43.A 0.392f
C392 I7 x3.x19.D 0.244f
C393 x5.x19.C x5.x19.D 0.996f
C394 VDD a_5475_n15675# 0.201f
C395 VDD I12 0.691f
C396 VDD I9 1.21f
C397 I7 x3.x2.X 0.0129f
C398 VDD x3.EI 4.87f
C399 a_5475_n13205# x3.x16.C 0.0949f
C400 a_5507_n2647# I12 0.188f
C401 VDD x3.A0 0.816f
C402 a_5935_n3179# x5.A2 0.144f
C403 x3.x22.A a_5509_n12251# 0.155f
C404 VDD a_6029_n1419# 0.15f
C405 x3.EI I1 0.437f
C406 a_5475_n1939# I13 0.16f
C407 I6 x3.x22.A 0.0536f
C408 VDD x3.EO 0.73f
C409 a_10776_n5725# x34.A 0.12f
C410 x3.x17.A a_6219_n12955# 0.213f
C411 VDD x29.Y 16.5f
C412 x3.x20.X x3.x21.B 0.0561f
C413 x5.x4.A x5.x1.X 0.118f
C414 I11 x5.x16.C 0.132f
C415 I8 x5.x19.C 0.12f
C416 a_5475_n5415# I11 0.162f
C417 I5 x3.x4.A 0.0107f
C418 I12 I9 0.427f
C419 I14 x5.x18.C 0.301f
C420 x3.EI a_5507_n10687# 0.0883f
C421 x36.Y A2 8.67f
C422 x5.x20.X x2.A 0.0148f
C423 a_10776_n13515# x2.X 0.12f
C424 x3.EI a_5475_n15675# 0.343f
C425 VDD a_6219_n12955# 0.155f
C426 x1.A x28.A 0.0126f
C427 I14 x5.x19.D 0.464f
C428 x5.A2 x34.A 0.0422f
C429 x5.x14.A x5.x22.A 0.0179f
C430 I5 I4 2.94f
C431 x5.x22.A I13 0.066f
C432 a_6219_n4915# x5.x16.X 0.0673f
C433 VDD x5.x19.C 1f
C434 I2 a_5475_n9215# 0.216f
C435 VDD a_5475_n9979# 0.153f
C436 VDD a_6395_n15425# 0.151f
C437 x5.A2 x43.Y 0.0114f
C438 I14 x5.x2.X 0.0177f
C439 VDD x43.A 1.46f
C440 x3.A2 x1.A 1.46f
C441 I5 I7 1.11f
C442 x3.x18.C I2 0.341f
C443 I3 a_5475_n14689# 0.15f
C444 x3.EI x3.EO 0.187f
C445 a_5967_n7607# EI 0.106f
C446 x5.x22.A a_5509_n4211# 0.155f
C447 x5.x22.A x2.A 0.132f
C448 I3 I2 2.81f
C449 x3.x22.A a_5475_n13205# 0.0116f
C450 x5.x17.A I14 0.0474f
C451 a_5475_n14689# x3.x21.B 0.0141f
C452 x3.x4.A a_6029_n9459# 0.299f
C453 x3.x14.A x3.x22.A 0.0179f
C454 I14 I8 0.353f
C455 EI I11 1.96f
C456 a_5475_n6397# x5.x18.C 0.117f
C457 x5.x17.A a_6219_n4915# 0.213f
C458 x5.x2.X x5.EO 0.0749f
C459 I12 x5.x19.C 0.405f
C460 I9 x5.x19.C 0.347f
C461 a_5475_n6397# x5.x19.D 0.14f
C462 I0 I4 0.553f
C463 VDD A0 6.58f
C464 x3.A2 a_10776_n5725# 0.119f
C465 x3.A1 x3.x22.A 0.519f
C466 x3.x15.X x3.x16.C 0.0319f
C467 a_6395_n15425# x3.A0 0.149f
C468 VDD I14 0.633f
C469 x2.A x3.A1 1.21f
C470 VDD x1.X 0.345f
C471 I0 I7 0.375f
C472 I13 x5.x16.C 0.415f
C473 VDD a_6219_n4915# 0.155f
C474 I5 a_5507_n10997# 0.194f
C475 x5.A2 x3.A2 0.358f
C476 VDD A2 6.58f
C477 I10 x5.x4.A 0.0109f
C478 x5.x20.X EI 0.208f
C479 I2 x3.x16.C 0.925f
C480 I4 x3.x19.C 0.405f
C481 x35.A x36.A 0.392f
C482 VDD x3.x4.A 1.38f
C483 x5.x22.A a_5475_n5165# 0.0116f
C484 VDD x22.A 1.51f
C485 VDD x5.EO 0.868f
C486 x5.x21.B a_5967_n7607# 0.186f
C487 a_5475_n9215# x3.x2.X 0.0313f
C488 I6 I2 0.439f
C489 x3.x18.C x3.x19.D 0.491f
C490 I12 I14 2.35f
C491 a_6519_n1397# x5.GS 0.136f
C492 I7 x3.x19.C 0.239f
C493 I1 x3.x4.A 0.0154f
C494 I3 x3.x19.D 1.27f
C495 x21.A x22.A 0.392f
C496 a_5967_n7607# x5.x21.X 0.109f
C497 VDD I4 0.692f
C498 x5.x19.X x5.x20.X 0.145f
C499 x5.x21.B I11 0.0112f
C500 I14 I9 0.258f
C501 x5.x17.A a_5935_n3179# 0.2f
C502 a_5967_n15647# x3.x20.X 0.137f
C503 x3.x21.B x3.x19.D 0.151f
C504 VDD a_5475_n6397# 0.428f
C505 a_5475_n13205# x3.x15.X 0.0951f
C506 I1 I4 0.428f
C507 x3.A1 a_10776_n9865# 0.121f
C508 VDD I7 0.205f
C509 x5.x14.A EI 0.0111f
C510 x5.x22.A EI 0.0483f
C511 I11 I15 1.03f
C512 I13 EI 3.7f
C513 x3.x22.A x3.x15.X 0.209f
C514 a_5475_n5415# x5.x16.C 0.0677f
C515 I5 x3.x11.X 0.0201f
C516 x3.EI x3.x4.A 0.547f
C517 a_5475_n6649# EI 0.175f
C518 I1 I7 0.24f
C519 a_5507_n10687# I4 0.188f
C520 VDD a_5935_n3179# 0.152f
C521 x5.x22.A x5.x19.X 0.418f
C522 x3.EI x5.EO 0.644f
C523 x3.x17.A a_5935_n11219# 0.2f
C524 x5.x19.D x5.x4.A 0.0516f
C525 x3.A1 x3.x15.X 0.0206f
C526 a_5509_n4211# EI 0.088f
C527 VDD A3 6.95f
C528 a_5475_n13205# I2 0.167f
C529 x5.x22.A x1.A 0.492f
C530 x5.x22.A x5.x15.X 0.209f
C531 x3.EI I4 1.8f
C532 a_6029_n1419# x5.EO 0.128f
C533 a_5475_n5165# x5.x16.C 0.0949f
C534 x5.x4.A x5.x2.X 0.125f
C535 a_5475_n1175# x5.x1.X 0.0991f
C536 VDD a_10776_n13515# 0.18f
C537 x3.x19.X x3.x21.B 0.262f
C538 x5.x21.B x5.x20.X 0.0561f
C539 a_5475_n6397# I9 0.147f
C540 a_5475_n6649# x5.x19.X 0.0873f
C541 x3.x4.A x3.EO 0.0491f
C542 VDD a_5935_n11219# 0.152f
C543 VDD a_5507_n2957# 0.215f
C544 I14 x5.x19.C 0.305f
C545 x3.x16.C x3.x19.D 1.24f
C546 x5.x19.X x2.A 0.0122f
C547 x5.x20.X x5.x21.X 0.122f
C548 EI a_6519_n1397# 0.18f
C549 x3.EI I7 4.77f
C550 I3 x3.x16.X 0.0148f
C551 I6 x3.x19.D 0.464f
C552 x5.A2 x35.A 0.0138f
C553 x3.x18.C I5 0.299f
C554 x2.A x1.A 0.304f
C555 VDD a_5507_n10997# 0.215f
C556 x3.x16.X x3.x21.B 0.0218f
C557 a_5475_n1939# I15 0.0614f
C558 VDD x34.A 0.346f
C559 EI x5.GS 0.0608f
C560 I5 I3 1.27f
C561 I6 x3.x2.X 0.0177f
C562 VDD x43.Y 11.3f
C563 I10 I11 2.81f
C564 EI x5.x16.C 2.08f
C565 x5.x11.X x5.x17.A 0.125f
C566 x3.A1 x1.A 0.426f
C567 x3.x18.C a_5475_n14437# 0.117f
C568 a_5475_n5415# EI 0.14f
C569 x5.x22.A x5.x21.B 0.064f
C570 a_5475_n14437# x3.x21.B 0.116f
C571 x5.x22.A x5.x21.X 0.0749f
C572 I4 a_5475_n9979# 0.208f
C573 x5.x21.B a_5475_n6649# 0.0141f
C574 VDD x5.x4.A 1.37f
C575 x5.x22.A I15 0.0853f
C576 a_10776_n13515# x3.A0 0.119f
C577 I0 a_5475_n9215# 0.211f
C578 a_5475_n5165# EI 0.122f
C579 I13 I15 1.13f
C580 a_5475_n6397# x5.x19.C 0.157f
C581 I3 a_5475_n13455# 0.162f
C582 x3.x21.X x3.x21.B 0.0197f
C583 x5.x15.X x5.x16.C 0.0319f
C584 x5.x14.A x5.A2 0.074f
C585 x5.x22.A x5.A2 0.0408f
C586 I7 a_5475_n9979# 0.0614f
C587 VDD x5.x11.X 0.501f
C588 x3.x11.X x3.x17.A 0.125f
C589 x3.EI a_5507_n10997# 0.0829f
C590 x3.x18.C I0 0.119f
C591 I3 I0 0.654f
C592 x3.x16.X x3.x16.C 0.07f
C593 x3.x22.A x3.x19.D 0.0292f
C594 a_5509_n4211# I15 0.192f
C595 x1.A a_10776_n9865# 0.206f
C596 I11 x5.x18.C 0.251f
C597 x3.A2 x3.x17.A 0.047f
C598 VDD x3.x11.X 0.501f
C599 a_5475_n5165# x5.x15.X 0.0951f
C600 x5.x16.X I11 0.0148f
C601 I5 x3.x16.C 0.415f
C602 VDD x3.GS 0.565f
C603 VDD x28.A 0.534f
C604 I9 x5.x4.A 0.0154f
C605 I11 x5.x19.D 1.27f
C606 I5 I6 4.51f
C607 I10 a_5475_n1175# 0.216f
C608 VDD x3.A2 1.41f
C609 a_5507_n3887# EI 0.0878f
C610 x2.A x2.X 0.0402f
C611 x5.x19.X EI 0.0149f
C612 x3.x18.C x3.x19.C 2.6f
C613 VDD a_5475_n9215# 0.148f
C614 x3.x17.A a_5507_n11927# 0.14f
C615 I3 x3.x19.C 0.921f
C616 VDD x22.Y 16.6f
C617 x5.x4.A a_6029_n1419# 0.299f
C618 x5.x15.X EI 0.0245f
C619 x3.x21.B x3.x19.C 0.0127f
C620 I15 x5.x16.C 0.26f
C621 a_5475_n13455# x3.x16.C 0.0677f
C622 I10 I13 0.641f
C623 x3.x22.A x3.x19.X 0.418f
C624 I1 a_5475_n9215# 0.159f
C625 a_5475_n7635# x5.x20.X 0.0895f
C626 VDD x3.x18.C 0.547f
C627 x3.x1.X x3.x2.X 0.129f
C628 VDD a_5507_n11927# 0.223f
C629 A0 GND 13.2f
C630 A1 GND 13.3f
C631 I7 GND 5.05f
C632 I0 GND 4.86f
C633 I3 GND 5.85f
C634 I1 GND 4.62f
C635 I6 GND 5.22f
C636 I5 GND 6.69f
C637 I4 GND 4.06f
C638 I2 GND 5f
C639 A2 GND 13.2f
C640 I15 GND 5f
C641 A3 GND 17.2f
C642 I8 GND 4.83f
C643 I11 GND 5.85f
C644 I9 GND 4.64f
C645 EI GND 19.1f
C646 I14 GND 5.24f
C647 I13 GND 6.7f
C648 I12 GND 4.06f
C649 I10 GND 4.84f
C650 VDD GND 0.223p
C651 x3.x21.X GND 0.241f
C652 x3.x20.X GND 0.683f
C653 a_6395_n15425# GND 0.362f
C654 a_5967_n15647# GND 0.217f
C655 a_5475_n15675# GND 0.292f
C656 x3.x19.X GND 0.432f
C657 a_5475_n14689# GND 0.293f
C658 x3.x21.B GND 0.656f
C659 a_5475_n14437# GND 0.295f
C660 x3.A0 GND 5.13f
C661 a_5475_n13455# GND 0.297f
C662 x22.Y GND 9.83f
C663 x22.A GND 2.12f
C664 x21.A GND 0.661f
C665 x2.X GND 0.381f
C666 a_10776_n13515# GND 0.263f
C667 x3.x16.X GND 0.871f
C668 x3.x15.X GND 0.334f
C669 a_6219_n12955# GND 0.369f
C670 a_5475_n13205# GND 0.296f
C671 a_5509_n12251# GND 0.286f
C672 a_5507_n11927# GND 0.288f
C673 a_5935_n11219# GND 0.367f
C674 x3.x17.A GND 0.917f
C675 x3.x22.A GND 2.01f
C676 x3.x11.X GND 0.263f
C677 a_5507_n10997# GND 0.28f
C678 x3.x14.A GND 0.978f
C679 a_5507_n10687# GND 0.289f
C680 x3.A1 GND 5.12f
C681 x29.Y GND 9.87f
C682 x29.A GND 2.13f
C683 x28.A GND 0.665f
C684 x1.X GND 0.383f
C685 a_10776_n9865# GND 0.265f
C686 a_5475_n9979# GND 0.388f
C687 x3.GS GND 2.06f
C688 x3.EO GND 2.32f
C689 x3.x2.X GND 0.676f
C690 x3.x1.X GND 0.162f
C691 a_6519_n9437# GND 0.258f
C692 a_6029_n9459# GND 0.343f
C693 a_5475_n9215# GND 0.379f
C694 x3.x4.A GND 1.07f
C695 x3.x19.D GND 4.1f
C696 x3.x16.C GND 1.84f
C697 x3.x19.C GND 4.41f
C698 x3.x18.C GND 1.88f
C699 x2.A GND 6.64f
C700 x5.x21.X GND 0.242f
C701 x5.x20.X GND 0.684f
C702 a_6395_n7385# GND 0.364f
C703 a_5967_n7607# GND 0.217f
C704 a_5475_n7635# GND 0.291f
C705 x5.x19.X GND 0.434f
C706 a_5475_n6649# GND 0.293f
C707 x5.x21.B GND 0.652f
C708 a_5475_n6397# GND 0.295f
C709 x3.A2 GND 7.64f
C710 x36.Y GND 9.83f
C711 x36.A GND 2.12f
C712 x35.A GND 0.662f
C713 x34.A GND 0.379f
C714 a_10776_n5725# GND 0.263f
C715 a_5475_n5415# GND 0.297f
C716 x1.A GND 5.67f
C717 x5.x16.X GND 0.871f
C718 x5.x15.X GND 0.334f
C719 a_6219_n4915# GND 0.369f
C720 a_5475_n5165# GND 0.296f
C721 a_5509_n4211# GND 0.286f
C722 a_5507_n3887# GND 0.288f
C723 x5.A2 GND 5.29f
C724 a_5935_n3179# GND 0.367f
C725 x5.x17.A GND 0.876f
C726 x5.x22.A GND 1.77f
C727 x5.x11.X GND 0.263f
C728 a_5507_n2957# GND 0.28f
C729 x5.x14.A GND 0.958f
C730 a_5507_n2647# GND 0.289f
C731 x3.EI GND 18.4f
C732 a_5475_n1939# GND 0.391f
C733 x43.Y GND 9.88f
C734 x43.A GND 2.02f
C735 x42.A GND 0.633f
C736 x5.GS GND 2.5f
C737 x5.EO GND 2.62f
C738 x5.x2.X GND 0.684f
C739 x5.x1.X GND 0.166f
C740 a_6519_n1397# GND 0.262f
C741 a_6029_n1419# GND 0.347f
C742 a_5475_n1175# GND 0.384f
C743 x5.x4.A GND 1.5f
C744 x5.x19.D GND 4.1f
C745 x5.x16.C GND 1.84f
C746 x5.x19.C GND 4.41f
C747 x5.x18.C GND 1.88f
C748 I11.n2 GND 0.0117f
C749 I11.n4 GND 0.99f
C750 I11.n5 GND 0.565f
C751 I11.n6 GND 0.552f
C752 I6.n0 GND 0.0245f
C753 I6.t2 GND 0.0182f
C754 I6.t5 GND 0.0289f
C755 I6.n2 GND 0.0547f
C756 I6.n3 GND 0.0117f
C757 I6.n7 GND 0.0198f
C758 I6.n9 GND 0.0394f
C759 I6.n10 GND 0.484f
C760 I6.t0 GND 0.0156f
C761 I6.t3 GND 0.0129f
C762 I6.n11 GND 0.0354f
C763 I6.n12 GND 0.0362f
C764 I6.n13 GND 0.633f
C765 I6.n14 GND 0.0212f
C766 I6.n15 GND 0.0138f
C767 I6.t1 GND 0.0193f
C768 I6.t4 GND 0.0135f
C769 I6.n16 GND 0.0463f
C770 I6.n17 GND 0.0116f
C771 I6.n18 GND 0.0167f
C772 I6.n20 GND 1.52f
C773 I6.n21 GND 2.47f
C774 I6.n22 GND 2.08f
C775 I6.n23 GND 1.23f
C776 I8.n0 GND 0.0213f
C777 I8.n1 GND 0.647f
C778 I8.n2 GND 1.81f
C779 I13.t2 GND 0.0113f
C780 I13.t4 GND 0.0178f
C781 I13.n0 GND 0.0337f
C782 I13.n7 GND 0.015f
C783 I13.n8 GND 0.376f
C784 I13.t0 GND 0.0162f
C785 I13.t6 GND 0.0307f
C786 I13.t7 GND 0.0119f
C787 I13.n11 GND 0.0286f
C788 I13.n14 GND 0.0243f
C789 I13.n15 GND 0.535f
C790 I13.n18 GND 0.024f
C791 I13.n19 GND 0.0156f
C792 I13.n20 GND 1.42f
C793 I13.n21 GND 3.36f
C794 I13.n22 GND 1.57f
C795 I13.n23 GND 1.29f
C796 I13.n24 GND 0.878f
C797 I5.t3 GND 0.0162f
C798 I5.t1 GND 0.0307f
C799 I5.t0 GND 0.0113f
C800 I5.t4 GND 0.0177f
C801 I5.n3 GND 0.0337f
C802 I5.n7 GND 0.015f
C803 I5.n8 GND 0.376f
C804 I5.n9 GND 0.937f
C805 I5.n10 GND 0.0242f
C806 I5.t2 GND 0.0119f
C807 I5.n12 GND 0.0286f
C808 I5.n16 GND 0.534f
C809 I5.n18 GND 0.024f
C810 I5.n20 GND 0.0156f
C811 I5.n21 GND 1.42f
C812 I5.n22 GND 3.36f
C813 I5.n23 GND 0.763f
C814 I5.n24 GND 2.06f
C815 I7.n0 GND 0.0323f
C816 I7.n1 GND 0.0136f
C817 I7.t3 GND 0.0125f
C818 I7.n3 GND 0.0299f
C819 I7.n8 GND 1.17f
C820 I7.n9 GND 2.51f
C821 I7.n10 GND 1.35f
C822 I0.n0 GND 0.021f
C823 I0.n1 GND 0.638f
C824 I0.n2 GND 1.81f
C825 I9.t1 GND 0.0133f
C826 I9.t2 GND 0.0251f
C827 I9.t3 GND 0.012f
C828 I9.n0 GND 0.0268f
C829 I9.n1 GND 1.15f
C830 I9.n2 GND 2.34f
C831 I9.n3 GND 1.49f
C832 I10.t1 GND 0.0128f
C833 I10.t3 GND 0.0201f
C834 I10.n0 GND 0.0386f
C835 I10.n1 GND 0.28f
C836 I10.t4 GND 0.0109f
C837 I10.n2 GND 0.0247f
C838 I10.n3 GND 0.0257f
C839 I10.t5 GND 0.0161f
C840 I10.t2 GND 0.0109f
C841 I10.n4 GND 0.0441f
C842 I10.n5 GND 0.206f
C843 I10.n6 GND 3.85f
C844 I10.n7 GND 1.41f
C845 I10.n8 GND 0.569f
C846 I4.n1 GND 0.0115f
C847 I4.t3 GND 0.0157f
C848 I4.n2 GND 0.0293f
C849 I4.n3 GND 0.0804f
C850 I4.n4 GND 0.873f
C851 I4.n5 GND 0.0203f
C852 I4.n6 GND 0.38f
C853 I4.n7 GND 0.81f
C854 I4.n8 GND 1.42f
C855 I4.n9 GND 0.496f
C856 I4.t5 GND 0.0104f
C857 I4.n12 GND 0.025f
C858 I14.n0 GND 0.0248f
C859 I14.t3 GND 0.0184f
C860 I14.t5 GND 0.0291f
C861 I14.n2 GND 0.0552f
C862 I14.n3 GND 0.0118f
C863 I14.n7 GND 0.02f
C864 I14.n9 GND 0.0398f
C865 I14.n10 GND 0.489f
C866 I14.t0 GND 0.0158f
C867 I14.t2 GND 0.013f
C868 I14.n11 GND 0.0358f
C869 I14.n12 GND 0.0365f
C870 I14.n13 GND 0.64f
C871 I14.n14 GND 0.0214f
C872 I14.n15 GND 0.014f
C873 I14.t1 GND 0.0195f
C874 I14.t4 GND 0.0136f
C875 I14.n16 GND 0.0468f
C876 I14.n17 GND 0.0117f
C877 I14.n18 GND 0.0169f
C878 I14.n20 GND 1.53f
C879 I14.n21 GND 2.55f
C880 I14.n22 GND 2.09f
C881 I14.n23 GND 1.18f
C882 A3.n1 GND 0.03f
C883 A3.n2 GND 0.0161f
C884 A3.n3 GND 0.0635f
C885 A3.n4 GND 0.0161f
C886 A3.n5 GND 0.0422f
C887 A3.n6 GND 0.0161f
C888 A3.n7 GND 0.0422f
C889 A3.n8 GND 0.0161f
C890 A3.n9 GND 0.0422f
C891 A3.n10 GND 0.0161f
C892 A3.n11 GND 0.0422f
C893 A3.n12 GND 0.0161f
C894 A3.n13 GND 0.0422f
C895 A3.n14 GND 0.0139f
C896 A3.n15 GND 0.0138f
C897 A3.n16 GND 0.0143f
C898 A3.n17 GND 0.0208f
C899 A3.n18 GND 0.0272f
C900 A3.n20 GND 0.0104f
C901 A3.n21 GND 0.0367f
C902 A3.n22 GND 0.0238f
C903 A3.n23 GND 0.0915f
C904 A3.n24 GND 0.0238f
C905 A3.n25 GND 0.0553f
C906 A3.n26 GND 0.0238f
C907 A3.n27 GND 0.0553f
C908 A3.n28 GND 0.0238f
C909 A3.n29 GND 0.0553f
C910 A3.n30 GND 0.0238f
C911 A3.n31 GND 0.0553f
C912 A3.n32 GND 0.0238f
C913 A3.n33 GND 0.0553f
C914 A3.n34 GND 0.0151f
C915 A3.n36 GND 0.0197f
C916 A3.n42 GND 0.0267f
C917 A3.n43 GND 0.0367f
C918 A3.n44 GND 0.0238f
C919 A3.n45 GND 0.0915f
C920 A3.n46 GND 0.0238f
C921 A3.n47 GND 0.0553f
C922 A3.n48 GND 0.0238f
C923 A3.n49 GND 0.0553f
C924 A3.n50 GND 0.0238f
C925 A3.n51 GND 0.0553f
C926 A3.n52 GND 0.0238f
C927 A3.n53 GND 0.0553f
C928 A3.n54 GND 0.0238f
C929 A3.n55 GND 0.0553f
C930 A3.n56 GND 0.0127f
C931 A3.n58 GND 0.0472f
C932 A3.n60 GND 0.0152f
C933 A3.n61 GND 0.0223f
C934 A3.n62 GND 0.03f
C935 A3.n63 GND 0.0161f
C936 A3.n64 GND 0.0635f
C937 A3.n65 GND 0.0161f
C938 A3.n66 GND 0.0422f
C939 A3.n67 GND 0.0161f
C940 A3.n68 GND 0.0422f
C941 A3.n69 GND 0.0161f
C942 A3.n70 GND 0.0422f
C943 A3.n71 GND 0.0161f
C944 A3.n72 GND 0.0422f
C945 A3.n73 GND 0.0161f
C946 A3.n74 GND 0.0422f
C947 A3.n75 GND 0.0153f
C948 A3.n77 GND 0.0451f
C949 A3.n78 GND 0.143f
C950 A3.n79 GND 0.0334f
C951 A3.n80 GND 0.025f
C952 A3.n81 GND 0.0367f
C953 A3.n82 GND 0.0238f
C954 A3.n83 GND 0.0915f
C955 A3.n84 GND 0.0238f
C956 A3.n85 GND 0.0553f
C957 A3.n86 GND 0.0238f
C958 A3.n87 GND 0.0553f
C959 A3.n88 GND 0.0238f
C960 A3.n89 GND 0.0553f
C961 A3.n90 GND 0.0238f
C962 A3.n91 GND 0.0553f
C963 A3.n92 GND 0.0238f
C964 A3.n93 GND 0.0553f
C965 A3.n94 GND 0.0163f
C966 A3.n99 GND 0.0214f
C967 A3.n101 GND 0.0185f
C968 A3.n102 GND 0.0144f
C969 A3.n103 GND 0.0216f
C970 A3.n104 GND 0.03f
C971 A3.n105 GND 0.0161f
C972 A3.n106 GND 0.0635f
C973 A3.n107 GND 0.0161f
C974 A3.n108 GND 0.0422f
C975 A3.n109 GND 0.0161f
C976 A3.n110 GND 0.0422f
C977 A3.n111 GND 0.0161f
C978 A3.n112 GND 0.0422f
C979 A3.n113 GND 0.0161f
C980 A3.n114 GND 0.0422f
C981 A3.n115 GND 0.0161f
C982 A3.n116 GND 0.0422f
C983 A3.n121 GND 0.0153f
C984 A3.n123 GND 0.0188f
C985 A3.n124 GND 0.017f
C986 A3.n125 GND 0.0846f
C987 A3.n126 GND 0.064f
C988 A3.n127 GND 0.0208f
C989 A3.n128 GND 0.0272f
C990 A3.n129 GND 0.0143f
C991 A3.n131 GND 0.0104f
C992 A3.n132 GND 0.0367f
C993 A3.n133 GND 0.0238f
C994 A3.n134 GND 0.0915f
C995 A3.n135 GND 0.0238f
C996 A3.n136 GND 0.0553f
C997 A3.n137 GND 0.0238f
C998 A3.n138 GND 0.0553f
C999 A3.n139 GND 0.0238f
C1000 A3.n140 GND 0.0553f
C1001 A3.n141 GND 0.0238f
C1002 A3.n142 GND 0.0553f
C1003 A3.n143 GND 0.0238f
C1004 A3.n144 GND 0.0553f
C1005 A3.n145 GND 0.0151f
C1006 A3.n147 GND 0.0197f
C1007 A3.n148 GND 0.0168f
C1008 A3.n149 GND 0.0206f
C1009 A3.n150 GND 0.03f
C1010 A3.n151 GND 0.0161f
C1011 A3.n152 GND 0.0635f
C1012 A3.n153 GND 0.0161f
C1013 A3.n154 GND 0.0422f
C1014 A3.n155 GND 0.0161f
C1015 A3.n156 GND 0.0422f
C1016 A3.n157 GND 0.0161f
C1017 A3.n158 GND 0.0422f
C1018 A3.n159 GND 0.0161f
C1019 A3.n160 GND 0.0422f
C1020 A3.n161 GND 0.0161f
C1021 A3.n162 GND 0.0422f
C1022 A3.n163 GND 0.0139f
C1023 A3.n164 GND 0.0138f
C1024 A3.n166 GND 0.0153f
C1025 A3.n168 GND 0.0206f
C1026 A3.n170 GND 0.017f
C1027 A3.n171 GND 0.081f
C1028 A3.n172 GND 0.356f
C1029 A3.n173 GND 0.912f
C1030 A3.n174 GND 0.791f
C1031 A3.n175 GND 2.38f
C1032 A3.n176 GND 0.0658f
C1033 A3.n177 GND 0.081f
C1034 A3.n178 GND 0.017f
C1035 A3.n179 GND 0.0206f
C1036 A3.n180 GND 0.0132f
C1037 A3.n181 GND 0.0206f
C1038 A3.n183 GND 0.0153f
C1039 I1.t2 GND 0.0133f
C1040 I1.t0 GND 0.0251f
C1041 I1.t1 GND 0.012f
C1042 I1.n0 GND 0.0268f
C1043 I1.n1 GND 1.13f
C1044 I1.n2 GND 2.34f
C1045 I1.n3 GND 1.52f
C1046 I3.n2 GND 0.0117f
C1047 I3.n4 GND 0.98f
C1048 I3.n5 GND 0.567f
C1049 I3.n6 GND 0.561f
C1050 EI.n1 GND 0.0216f
C1051 EI.n7 GND 0.0126f
C1052 EI.n8 GND 0.578f
C1053 EI.t12 GND 0.0134f
C1054 EI.n10 GND 0.0255f
C1055 EI.n15 GND 0.0158f
C1056 EI.n16 GND 0.0188f
C1057 EI.n18 GND 0.19f
C1058 EI.n19 GND 0.026f
C1059 EI.n21 GND 0.0465f
C1060 EI.n22 GND 0.026f
C1061 EI.n24 GND 0.026f
C1062 EI.n26 GND 0.065f
C1063 EI.n27 GND 0.0261f
C1064 EI.n28 GND 0.0132f
C1065 EI.t14 GND 0.0109f
C1066 EI.n29 GND 0.0247f
C1067 EI.t8 GND 0.0109f
C1068 EI.n30 GND 0.0251f
C1069 EI.n31 GND 0.027f
C1070 EI.n37 GND 0.357f
C1071 EI.t20 GND 0.0108f
C1072 EI.n38 GND 0.0305f
C1073 EI.n39 GND 0.0125f
C1074 EI.n40 GND 0.021f
C1075 EI.n41 GND 0.308f
C1076 EI.n42 GND 0.0106f
C1077 EI.n44 GND 0.0138f
C1078 EI.n47 GND 0.273f
C1079 EI.n48 GND 1.21f
C1080 EI.n49 GND 1.01f
C1081 EI.n50 GND 0.725f
C1082 EI.n51 GND 0.931f
C1083 EI.n52 GND 1.15f
C1084 EI.n53 GND 1.14f
C1085 EI.n54 GND 1.03f
C1086 EI.n55 GND 1.19f
C1087 EI.n56 GND 1.06f
C1088 EI.n57 GND 0.462f
C1089 I15.n0 GND 0.0323f
C1090 I15.n1 GND 0.0136f
C1091 I15.t2 GND 0.0125f
C1092 I15.n3 GND 0.03f
C1093 I15.n8 GND 1.17f
C1094 I15.n9 GND 2.55f
C1095 I15.n10 GND 1.35f
C1096 A1.n0 GND 0.0141f
C1097 A1.n1 GND 0.0306f
C1098 A1.n2 GND 0.0442f
C1099 A1.n3 GND 0.0238f
C1100 A1.n4 GND 0.0938f
C1101 A1.n5 GND 0.0238f
C1102 A1.n6 GND 0.0623f
C1103 A1.n7 GND 0.0238f
C1104 A1.n8 GND 0.0623f
C1105 A1.n9 GND 0.0238f
C1106 A1.n10 GND 0.0623f
C1107 A1.n11 GND 0.0238f
C1108 A1.n12 GND 0.0623f
C1109 A1.n13 GND 0.0238f
C1110 A1.n14 GND 0.0623f
C1111 A1.n15 GND 0.0228f
C1112 A1.n18 GND 0.0218f
C1113 A1.n20 GND 0.0223f
C1114 A1.n21 GND 0.0221f
C1115 A1.t68 GND 0.0146f
C1116 A1.t124 GND 0.0146f
C1117 A1.n22 GND 0.0342f
C1118 A1.t96 GND 0.0146f
C1119 A1.t92 GND 0.0146f
C1120 A1.n23 GND 0.0542f
C1121 A1.t90 GND 0.0146f
C1122 A1.t101 GND 0.0146f
C1123 A1.n24 GND 0.0352f
C1124 A1.n25 GND 0.135f
C1125 A1.t82 GND 0.0146f
C1126 A1.t75 GND 0.0146f
C1127 A1.n26 GND 0.0352f
C1128 A1.n27 GND 0.0817f
C1129 A1.t80 GND 0.0146f
C1130 A1.t65 GND 0.0146f
C1131 A1.n28 GND 0.0352f
C1132 A1.n29 GND 0.0817f
C1133 A1.t72 GND 0.0146f
C1134 A1.t86 GND 0.0146f
C1135 A1.n30 GND 0.0352f
C1136 A1.n31 GND 0.0817f
C1137 A1.t126 GND 0.0146f
C1138 A1.t78 GND 0.0146f
C1139 A1.n32 GND 0.0352f
C1140 A1.n33 GND 0.0817f
C1141 A1.t118 GND 0.0146f
C1142 A1.t70 GND 0.0146f
C1143 A1.n34 GND 0.0352f
C1144 A1.n35 GND 0.0817f
C1145 A1.n36 GND 0.0234f
C1146 A1.n37 GND 0.0571f
C1147 A1.n38 GND 0.106f
C1148 A1.n39 GND 0.079f
C1149 A1.n40 GND 0.0139f
C1150 A1.n41 GND 0.0442f
C1151 A1.n42 GND 0.0238f
C1152 A1.n43 GND 0.0938f
C1153 A1.n44 GND 0.0238f
C1154 A1.n45 GND 0.0623f
C1155 A1.n46 GND 0.0238f
C1156 A1.n47 GND 0.0623f
C1157 A1.n48 GND 0.0238f
C1158 A1.n49 GND 0.0623f
C1159 A1.n50 GND 0.0238f
C1160 A1.n51 GND 0.0623f
C1161 A1.n52 GND 0.0238f
C1162 A1.n53 GND 0.0623f
C1163 A1.n54 GND 0.0227f
C1164 A1.n55 GND 0.0226f
C1165 A1.n57 GND 0.0489f
C1166 A1.n58 GND 0.0218f
C1167 A1.t89 GND 0.0146f
C1168 A1.t84 GND 0.0146f
C1169 A1.n59 GND 0.0342f
C1170 A1.t116 GND 0.0146f
C1171 A1.t123 GND 0.0146f
C1172 A1.n60 GND 0.0542f
C1173 A1.t64 GND 0.0146f
C1174 A1.t102 GND 0.0146f
C1175 A1.n61 GND 0.0352f
C1176 A1.n62 GND 0.135f
C1177 A1.t121 GND 0.0146f
C1178 A1.t114 GND 0.0146f
C1179 A1.n63 GND 0.0352f
C1180 A1.n64 GND 0.0817f
C1181 A1.t93 GND 0.0146f
C1182 A1.t106 GND 0.0146f
C1183 A1.n65 GND 0.0352f
C1184 A1.n66 GND 0.0817f
C1185 A1.t104 GND 0.0146f
C1186 A1.t100 GND 0.0146f
C1187 A1.n67 GND 0.0352f
C1188 A1.n68 GND 0.0817f
C1189 A1.t98 GND 0.0146f
C1190 A1.t110 GND 0.0146f
C1191 A1.n69 GND 0.0352f
C1192 A1.n70 GND 0.0817f
C1193 A1.t95 GND 0.0146f
C1194 A1.t87 GND 0.0146f
C1195 A1.n71 GND 0.0352f
C1196 A1.n72 GND 0.0817f
C1197 A1.n73 GND 0.0225f
C1198 A1.n74 GND 0.057f
C1199 A1.n75 GND 0.11f
C1200 A1.n76 GND 0.0907f
C1201 A1.n77 GND 0.0316f
C1202 A1.t103 GND 0.0146f
C1203 A1.t117 GND 0.0146f
C1204 A1.n78 GND 0.0325f
C1205 A1.n79 GND 0.0369f
C1206 A1.t91 GND 0.0146f
C1207 A1.t85 GND 0.0146f
C1208 A1.n80 GND 0.0542f
C1209 A1.t83 GND 0.0146f
C1210 A1.t76 GND 0.0146f
C1211 A1.n81 GND 0.0352f
C1212 A1.n82 GND 0.135f
C1213 A1.t74 GND 0.0146f
C1214 A1.t67 GND 0.0146f
C1215 A1.n83 GND 0.0352f
C1216 A1.n84 GND 0.0817f
C1217 A1.t73 GND 0.0146f
C1218 A1.t81 GND 0.0146f
C1219 A1.n85 GND 0.0352f
C1220 A1.n86 GND 0.0817f
C1221 A1.t127 GND 0.0146f
C1222 A1.t79 GND 0.0146f
C1223 A1.n87 GND 0.0352f
C1224 A1.n88 GND 0.0817f
C1225 A1.t77 GND 0.0146f
C1226 A1.t112 GND 0.0146f
C1227 A1.n89 GND 0.0352f
C1228 A1.n90 GND 0.0817f
C1229 A1.t69 GND 0.0146f
C1230 A1.t125 GND 0.0146f
C1231 A1.n91 GND 0.0352f
C1232 A1.n92 GND 0.0817f
C1233 A1.n93 GND 0.022f
C1234 A1.n95 GND 0.0221f
C1235 A1.n96 GND 0.0442f
C1236 A1.n97 GND 0.0238f
C1237 A1.n98 GND 0.0938f
C1238 A1.n99 GND 0.0238f
C1239 A1.n100 GND 0.0623f
C1240 A1.n101 GND 0.0238f
C1241 A1.n102 GND 0.0623f
C1242 A1.n103 GND 0.0238f
C1243 A1.n104 GND 0.0623f
C1244 A1.n105 GND 0.0238f
C1245 A1.n106 GND 0.0623f
C1246 A1.n107 GND 0.0238f
C1247 A1.n108 GND 0.0623f
C1248 A1.n109 GND 0.0227f
C1249 A1.n110 GND 0.0226f
C1250 A1.n112 GND 0.0501f
C1251 A1.n113 GND 0.0139f
C1252 A1.n114 GND 0.0223f
C1253 A1.n115 GND 0.0792f
C1254 A1.n116 GND 0.421f
C1255 A1.n117 GND 1.07f
C1256 A1.n118 GND 0.872f
C1257 A1.n119 GND 1.61f
C1258 A1.n120 GND 0.0889f
C1259 A1.t94 GND 0.0146f
C1260 A1.t108 GND 0.0146f
C1261 A1.n121 GND 0.0342f
C1262 A1.t119 GND 0.0146f
C1263 A1.t71 GND 0.0146f
C1264 A1.n122 GND 0.0542f
C1265 A1.t115 GND 0.0146f
C1266 A1.t66 GND 0.0146f
C1267 A1.n123 GND 0.0352f
C1268 A1.n124 GND 0.135f
C1269 A1.t107 GND 0.0146f
C1270 A1.t122 GND 0.0146f
C1271 A1.n125 GND 0.0352f
C1272 A1.n126 GND 0.0817f
C1273 A1.t120 GND 0.0146f
C1274 A1.t113 GND 0.0146f
C1275 A1.n127 GND 0.0352f
C1276 A1.n128 GND 0.0817f
C1277 A1.t111 GND 0.0146f
C1278 A1.t105 GND 0.0146f
C1279 A1.n129 GND 0.0352f
C1280 A1.n130 GND 0.0817f
C1281 A1.t88 GND 0.0146f
C1282 A1.t99 GND 0.0146f
C1283 A1.n131 GND 0.0352f
C1284 A1.n132 GND 0.0817f
C1285 A1.t97 GND 0.0146f
C1286 A1.t109 GND 0.0146f
C1287 A1.n133 GND 0.0352f
C1288 A1.n134 GND 0.0817f
C1289 A1.n135 GND 0.0234f
C1290 A1.n136 GND 0.0571f
C1291 A1.n137 GND 0.115f
C1292 A1.n138 GND 0.0141f
C1293 A1.n139 GND 0.0221f
C1294 A1.n140 GND 0.0442f
C1295 A1.n141 GND 0.0238f
C1296 A1.n142 GND 0.0938f
C1297 A1.n143 GND 0.0238f
C1298 A1.n144 GND 0.0623f
C1299 A1.n145 GND 0.0238f
C1300 A1.n146 GND 0.0623f
C1301 A1.n147 GND 0.0238f
C1302 A1.n148 GND 0.0623f
C1303 A1.n149 GND 0.0238f
C1304 A1.n150 GND 0.0623f
C1305 A1.n151 GND 0.0238f
C1306 A1.n152 GND 0.0623f
C1307 A1.n153 GND 0.0218f
C1308 A1.n154 GND 0.0228f
C1309 A1.n157 GND 0.0306f
C1310 A1.n158 GND 0.0223f
C1311 I12.n1 GND 0.0115f
C1312 I12.t3 GND 0.0158f
C1313 I12.n2 GND 0.0295f
C1314 I12.n3 GND 0.0809f
C1315 I12.n4 GND 0.878f
C1316 I12.n5 GND 0.0204f
C1317 I12.n6 GND 0.382f
C1318 I12.n7 GND 0.815f
C1319 I12.n8 GND 1.4f
C1320 I12.n9 GND 0.5f
C1321 I12.t0 GND 0.0105f
C1322 I12.n12 GND 0.0252f
C1323 A0.n0 GND 0.0141f
C1324 A0.n1 GND 0.0313f
C1325 A0.n2 GND 0.0442f
C1326 A0.n3 GND 0.0238f
C1327 A0.n4 GND 0.0938f
C1328 A0.n5 GND 0.0238f
C1329 A0.n6 GND 0.0623f
C1330 A0.n7 GND 0.0238f
C1331 A0.n8 GND 0.0623f
C1332 A0.n9 GND 0.0238f
C1333 A0.n10 GND 0.0623f
C1334 A0.n11 GND 0.0238f
C1335 A0.n12 GND 0.0623f
C1336 A0.n13 GND 0.0238f
C1337 A0.n14 GND 0.0623f
C1338 A0.n15 GND 0.0228f
C1339 A0.n18 GND 0.022f
C1340 A0.n20 GND 0.0221f
C1341 A0.n21 GND 0.0218f
C1342 A0.t71 GND 0.0146f
C1343 A0.t96 GND 0.0146f
C1344 A0.n22 GND 0.0343f
C1345 A0.t85 GND 0.0146f
C1346 A0.t106 GND 0.0146f
C1347 A0.n23 GND 0.0542f
C1348 A0.t104 GND 0.0146f
C1349 A0.t122 GND 0.0146f
C1350 A0.n24 GND 0.0352f
C1351 A0.n25 GND 0.135f
C1352 A0.t67 GND 0.0146f
C1353 A0.t89 GND 0.0146f
C1354 A0.n26 GND 0.0352f
C1355 A0.n27 GND 0.0817f
C1356 A0.t118 GND 0.0146f
C1357 A0.t112 GND 0.0146f
C1358 A0.n28 GND 0.0352f
C1359 A0.n29 GND 0.0817f
C1360 A0.t79 GND 0.0146f
C1361 A0.t92 GND 0.0146f
C1362 A0.n30 GND 0.0352f
C1363 A0.n31 GND 0.0817f
C1364 A0.t98 GND 0.0146f
C1365 A0.t116 GND 0.0146f
C1366 A0.n32 GND 0.0352f
C1367 A0.n33 GND 0.0817f
C1368 A0.t124 GND 0.0146f
C1369 A0.t73 GND 0.0146f
C1370 A0.n34 GND 0.0352f
C1371 A0.n35 GND 0.0817f
C1372 A0.n36 GND 0.0236f
C1373 A0.n37 GND 0.0572f
C1374 A0.n38 GND 0.106f
C1375 A0.n39 GND 0.079f
C1376 A0.n40 GND 0.0141f
C1377 A0.n41 GND 0.0442f
C1378 A0.n42 GND 0.0238f
C1379 A0.n43 GND 0.0938f
C1380 A0.n44 GND 0.0238f
C1381 A0.n45 GND 0.0623f
C1382 A0.n46 GND 0.0238f
C1383 A0.n47 GND 0.0623f
C1384 A0.n48 GND 0.0238f
C1385 A0.n49 GND 0.0623f
C1386 A0.n50 GND 0.0238f
C1387 A0.n51 GND 0.0623f
C1388 A0.n52 GND 0.0238f
C1389 A0.n53 GND 0.0623f
C1390 A0.n54 GND 0.0226f
C1391 A0.n55 GND 0.0226f
C1392 A0.n57 GND 0.0491f
C1393 A0.n58 GND 0.0218f
C1394 A0.t70 GND 0.0146f
C1395 A0.t95 GND 0.0146f
C1396 A0.n59 GND 0.0343f
C1397 A0.t84 GND 0.0146f
C1398 A0.t69 GND 0.0146f
C1399 A0.n60 GND 0.0542f
C1400 A0.t93 GND 0.0146f
C1401 A0.t77 GND 0.0146f
C1402 A0.n61 GND 0.0352f
C1403 A0.n62 GND 0.135f
C1404 A0.t120 GND 0.0146f
C1405 A0.t82 GND 0.0146f
C1406 A0.n63 GND 0.0352f
C1407 A0.n64 GND 0.0817f
C1408 A0.t87 GND 0.0146f
C1409 A0.t102 GND 0.0146f
C1410 A0.n65 GND 0.0352f
C1411 A0.n66 GND 0.0817f
C1412 A0.t100 GND 0.0146f
C1413 A0.t64 GND 0.0146f
C1414 A0.n67 GND 0.0352f
C1415 A0.n68 GND 0.0817f
C1416 A0.t126 GND 0.0146f
C1417 A0.t75 GND 0.0146f
C1418 A0.n69 GND 0.0352f
C1419 A0.n70 GND 0.0817f
C1420 A0.t113 GND 0.0146f
C1421 A0.t109 GND 0.0146f
C1422 A0.n71 GND 0.0352f
C1423 A0.n72 GND 0.0817f
C1424 A0.n73 GND 0.0227f
C1425 A0.n74 GND 0.057f
C1426 A0.n75 GND 0.11f
C1427 A0.n76 GND 0.0907f
C1428 A0.n77 GND 0.0304f
C1429 A0.t108 GND 0.0146f
C1430 A0.t123 GND 0.0146f
C1431 A0.n78 GND 0.0326f
C1432 A0.n79 GND 0.0374f
C1433 A0.t105 GND 0.0146f
C1434 A0.t78 GND 0.0146f
C1435 A0.n80 GND 0.0542f
C1436 A0.t68 GND 0.0146f
C1437 A0.t90 GND 0.0146f
C1438 A0.n81 GND 0.0352f
C1439 A0.n82 GND 0.135f
C1440 A0.t88 GND 0.0146f
C1441 A0.t114 GND 0.0146f
C1442 A0.n83 GND 0.0352f
C1443 A0.n84 GND 0.0817f
C1444 A0.t80 GND 0.0146f
C1445 A0.t65 GND 0.0146f
C1446 A0.n85 GND 0.0352f
C1447 A0.n86 GND 0.0817f
C1448 A0.t99 GND 0.0146f
C1449 A0.t117 GND 0.0146f
C1450 A0.n87 GND 0.0352f
C1451 A0.n88 GND 0.0817f
C1452 A0.t115 GND 0.0146f
C1453 A0.t86 GND 0.0146f
C1454 A0.n89 GND 0.0352f
C1455 A0.n90 GND 0.0817f
C1456 A0.t72 GND 0.0146f
C1457 A0.t97 GND 0.0146f
C1458 A0.n91 GND 0.0352f
C1459 A0.n92 GND 0.0817f
C1460 A0.n93 GND 0.0223f
C1461 A0.n95 GND 0.0223f
C1462 A0.n96 GND 0.0442f
C1463 A0.n97 GND 0.0238f
C1464 A0.n98 GND 0.0938f
C1465 A0.n99 GND 0.0238f
C1466 A0.n100 GND 0.0623f
C1467 A0.n101 GND 0.0238f
C1468 A0.n102 GND 0.0623f
C1469 A0.n103 GND 0.0238f
C1470 A0.n104 GND 0.0623f
C1471 A0.n105 GND 0.0238f
C1472 A0.n106 GND 0.0623f
C1473 A0.n107 GND 0.0238f
C1474 A0.n108 GND 0.0623f
C1475 A0.n109 GND 0.0226f
C1476 A0.n110 GND 0.0226f
C1477 A0.n112 GND 0.0503f
C1478 A0.n113 GND 0.0141f
C1479 A0.n114 GND 0.0226f
C1480 A0.n115 GND 0.0792f
C1481 A0.n116 GND 0.421f
C1482 A0.n117 GND 1.07f
C1483 A0.n118 GND 0.872f
C1484 A0.n119 GND 1.6f
C1485 A0.n120 GND 0.0889f
C1486 A0.t111 GND 0.0146f
C1487 A0.t66 GND 0.0146f
C1488 A0.n121 GND 0.0343f
C1489 A0.t91 GND 0.0146f
C1490 A0.t107 GND 0.0146f
C1491 A0.n122 GND 0.0542f
C1492 A0.t83 GND 0.0146f
C1493 A0.t94 GND 0.0146f
C1494 A0.n123 GND 0.0352f
C1495 A0.n124 GND 0.135f
C1496 A0.t103 GND 0.0146f
C1497 A0.t121 GND 0.0146f
C1498 A0.n125 GND 0.0352f
C1499 A0.n126 GND 0.0817f
C1500 A0.t119 GND 0.0146f
C1501 A0.t81 GND 0.0146f
C1502 A0.n127 GND 0.0352f
C1503 A0.n128 GND 0.0817f
C1504 A0.t76 GND 0.0146f
C1505 A0.t101 GND 0.0146f
C1506 A0.n129 GND 0.0352f
C1507 A0.n130 GND 0.0817f
C1508 A0.t110 GND 0.0146f
C1509 A0.t127 GND 0.0146f
C1510 A0.n131 GND 0.0352f
C1511 A0.n132 GND 0.0817f
C1512 A0.t125 GND 0.0146f
C1513 A0.t74 GND 0.0146f
C1514 A0.n133 GND 0.0352f
C1515 A0.n134 GND 0.0817f
C1516 A0.n135 GND 0.0236f
C1517 A0.n136 GND 0.0572f
C1518 A0.n137 GND 0.115f
C1519 A0.n138 GND 0.0141f
C1520 A0.n139 GND 0.0218f
C1521 A0.n140 GND 0.0442f
C1522 A0.n141 GND 0.0238f
C1523 A0.n142 GND 0.0938f
C1524 A0.n143 GND 0.0238f
C1525 A0.n144 GND 0.0623f
C1526 A0.n145 GND 0.0238f
C1527 A0.n146 GND 0.0623f
C1528 A0.n147 GND 0.0238f
C1529 A0.n148 GND 0.0623f
C1530 A0.n149 GND 0.0238f
C1531 A0.n150 GND 0.0623f
C1532 A0.n151 GND 0.0238f
C1533 A0.n152 GND 0.0623f
C1534 A0.n153 GND 0.022f
C1535 A0.n154 GND 0.0228f
C1536 A0.n157 GND 0.0313f
C1537 A0.n158 GND 0.0221f
C1538 I2.t4 GND 0.0142f
C1539 I2.t0 GND 0.0224f
C1540 I2.n0 GND 0.0431f
C1541 I2.n1 GND 0.312f
C1542 I2.t2 GND 0.01f
C1543 I2.t5 GND 0.0121f
C1544 I2.n2 GND 0.0275f
C1545 I2.n3 GND 0.0287f
C1546 I2.t3 GND 0.018f
C1547 I2.t1 GND 0.0122f
C1548 I2.n4 GND 0.0493f
C1549 I2.n5 GND 0.22f
C1550 I2.n6 GND 4.32f
C1551 I2.n7 GND 1.62f
C1552 I2.n8 GND 0.635f
C1553 A2.n0 GND 0.0141f
C1554 A2.n1 GND 0.0313f
C1555 A2.n2 GND 0.0442f
C1556 A2.n3 GND 0.0238f
C1557 A2.n4 GND 0.0938f
C1558 A2.n5 GND 0.0238f
C1559 A2.n6 GND 0.0623f
C1560 A2.n7 GND 0.0238f
C1561 A2.n8 GND 0.0623f
C1562 A2.n9 GND 0.0238f
C1563 A2.n10 GND 0.0623f
C1564 A2.n11 GND 0.0238f
C1565 A2.n12 GND 0.0623f
C1566 A2.n13 GND 0.0238f
C1567 A2.n14 GND 0.0623f
C1568 A2.n15 GND 0.0228f
C1569 A2.n18 GND 0.022f
C1570 A2.n20 GND 0.0221f
C1571 A2.n21 GND 0.0218f
C1572 A2.t82 GND 0.0146f
C1573 A2.t74 GND 0.0146f
C1574 A2.n22 GND 0.0343f
C1575 A2.t110 GND 0.0146f
C1576 A2.t106 GND 0.0146f
C1577 A2.n23 GND 0.0542f
C1578 A2.t104 GND 0.0146f
C1579 A2.t115 GND 0.0146f
C1580 A2.n24 GND 0.0352f
C1581 A2.n25 GND 0.135f
C1582 A2.t96 GND 0.0146f
C1583 A2.t89 GND 0.0146f
C1584 A2.n26 GND 0.0352f
C1585 A2.n27 GND 0.0817f
C1586 A2.t94 GND 0.0146f
C1587 A2.t79 GND 0.0146f
C1588 A2.n28 GND 0.0352f
C1589 A2.n29 GND 0.0817f
C1590 A2.t86 GND 0.0146f
C1591 A2.t101 GND 0.0146f
C1592 A2.n30 GND 0.0352f
C1593 A2.n31 GND 0.0817f
C1594 A2.t76 GND 0.0146f
C1595 A2.t92 GND 0.0146f
C1596 A2.n32 GND 0.0352f
C1597 A2.n33 GND 0.0817f
C1598 A2.t68 GND 0.0146f
C1599 A2.t84 GND 0.0146f
C1600 A2.n34 GND 0.0352f
C1601 A2.n35 GND 0.0817f
C1602 A2.n36 GND 0.0236f
C1603 A2.n37 GND 0.0572f
C1604 A2.n38 GND 0.106f
C1605 A2.n39 GND 0.079f
C1606 A2.n40 GND 0.0141f
C1607 A2.n41 GND 0.0442f
C1608 A2.n42 GND 0.0238f
C1609 A2.n43 GND 0.0938f
C1610 A2.n44 GND 0.0238f
C1611 A2.n45 GND 0.0623f
C1612 A2.n46 GND 0.0238f
C1613 A2.n47 GND 0.0623f
C1614 A2.n48 GND 0.0238f
C1615 A2.n49 GND 0.0623f
C1616 A2.n50 GND 0.0238f
C1617 A2.n51 GND 0.0623f
C1618 A2.n52 GND 0.0238f
C1619 A2.n53 GND 0.0623f
C1620 A2.n54 GND 0.0226f
C1621 A2.n55 GND 0.0226f
C1622 A2.n57 GND 0.0491f
C1623 A2.n58 GND 0.0218f
C1624 A2.t103 GND 0.0146f
C1625 A2.t98 GND 0.0146f
C1626 A2.n59 GND 0.0343f
C1627 A2.t66 GND 0.0146f
C1628 A2.t73 GND 0.0146f
C1629 A2.n60 GND 0.0542f
C1630 A2.t78 GND 0.0146f
C1631 A2.t116 GND 0.0146f
C1632 A2.n61 GND 0.0352f
C1633 A2.n62 GND 0.135f
C1634 A2.t71 GND 0.0146f
C1635 A2.t64 GND 0.0146f
C1636 A2.n63 GND 0.0352f
C1637 A2.n64 GND 0.0817f
C1638 A2.t107 GND 0.0146f
C1639 A2.t120 GND 0.0146f
C1640 A2.n65 GND 0.0352f
C1641 A2.n66 GND 0.0817f
C1642 A2.t118 GND 0.0146f
C1643 A2.t114 GND 0.0146f
C1644 A2.n67 GND 0.0352f
C1645 A2.n68 GND 0.0817f
C1646 A2.t112 GND 0.0146f
C1647 A2.t60 GND 0.0146f
C1648 A2.n69 GND 0.0352f
C1649 A2.n70 GND 0.0817f
C1650 A2.t109 GND 0.0146f
C1651 A2.t100 GND 0.0146f
C1652 A2.n71 GND 0.0352f
C1653 A2.n72 GND 0.0817f
C1654 A2.n73 GND 0.0227f
C1655 A2.n74 GND 0.057f
C1656 A2.n75 GND 0.11f
C1657 A2.n76 GND 0.0907f
C1658 A2.n77 GND 0.0304f
C1659 A2.t117 GND 0.0146f
C1660 A2.t67 GND 0.0146f
C1661 A2.n78 GND 0.0326f
C1662 A2.n79 GND 0.0374f
C1663 A2.t105 GND 0.0146f
C1664 A2.t99 GND 0.0146f
C1665 A2.n80 GND 0.0542f
C1666 A2.t97 GND 0.0146f
C1667 A2.t90 GND 0.0146f
C1668 A2.n81 GND 0.0352f
C1669 A2.n82 GND 0.135f
C1670 A2.t88 GND 0.0146f
C1671 A2.t80 GND 0.0146f
C1672 A2.n83 GND 0.0352f
C1673 A2.n84 GND 0.0817f
C1674 A2.t87 GND 0.0146f
C1675 A2.t95 GND 0.0146f
C1676 A2.n85 GND 0.0352f
C1677 A2.n86 GND 0.0817f
C1678 A2.t77 GND 0.0146f
C1679 A2.t93 GND 0.0146f
C1680 A2.n87 GND 0.0352f
C1681 A2.n88 GND 0.0817f
C1682 A2.t91 GND 0.0146f
C1683 A2.t62 GND 0.0146f
C1684 A2.n89 GND 0.0352f
C1685 A2.n90 GND 0.0817f
C1686 A2.t83 GND 0.0146f
C1687 A2.t75 GND 0.0146f
C1688 A2.n91 GND 0.0352f
C1689 A2.n92 GND 0.0817f
C1690 A2.n93 GND 0.0223f
C1691 A2.n95 GND 0.0223f
C1692 A2.n96 GND 0.0442f
C1693 A2.n97 GND 0.0238f
C1694 A2.n98 GND 0.0938f
C1695 A2.n99 GND 0.0238f
C1696 A2.n100 GND 0.0623f
C1697 A2.n101 GND 0.0238f
C1698 A2.n102 GND 0.0623f
C1699 A2.n103 GND 0.0238f
C1700 A2.n104 GND 0.0623f
C1701 A2.n105 GND 0.0238f
C1702 A2.n106 GND 0.0623f
C1703 A2.n107 GND 0.0238f
C1704 A2.n108 GND 0.0623f
C1705 A2.n109 GND 0.0226f
C1706 A2.n110 GND 0.0226f
C1707 A2.n112 GND 0.0503f
C1708 A2.n113 GND 0.0141f
C1709 A2.n114 GND 0.0226f
C1710 A2.n115 GND 0.0792f
C1711 A2.n116 GND 0.421f
C1712 A2.n117 GND 1.07f
C1713 A2.n118 GND 0.872f
C1714 A2.n119 GND 1.6f
C1715 A2.n120 GND 0.0889f
C1716 A2.t108 GND 0.0146f
C1717 A2.t58 GND 0.0146f
C1718 A2.n121 GND 0.0343f
C1719 A2.t69 GND 0.0146f
C1720 A2.t85 GND 0.0146f
C1721 A2.n122 GND 0.0542f
C1722 A2.t65 GND 0.0146f
C1723 A2.t81 GND 0.0146f
C1724 A2.n123 GND 0.0352f
C1725 A2.n124 GND 0.135f
C1726 A2.t57 GND 0.0146f
C1727 A2.t72 GND 0.0146f
C1728 A2.n125 GND 0.0352f
C1729 A2.n126 GND 0.0817f
C1730 A2.t70 GND 0.0146f
C1731 A2.t63 GND 0.0146f
C1732 A2.n127 GND 0.0352f
C1733 A2.n128 GND 0.0817f
C1734 A2.t61 GND 0.0146f
C1735 A2.t119 GND 0.0146f
C1736 A2.n129 GND 0.0352f
C1737 A2.n130 GND 0.0817f
C1738 A2.t102 GND 0.0146f
C1739 A2.t113 GND 0.0146f
C1740 A2.n131 GND 0.0352f
C1741 A2.n132 GND 0.0817f
C1742 A2.t111 GND 0.0146f
C1743 A2.t59 GND 0.0146f
C1744 A2.n133 GND 0.0352f
C1745 A2.n134 GND 0.0817f
C1746 A2.n135 GND 0.0236f
C1747 A2.n136 GND 0.0572f
C1748 A2.n137 GND 0.115f
C1749 A2.n138 GND 0.0141f
C1750 A2.n139 GND 0.0218f
C1751 A2.n140 GND 0.0442f
C1752 A2.n141 GND 0.0238f
C1753 A2.n142 GND 0.0938f
C1754 A2.n143 GND 0.0238f
C1755 A2.n144 GND 0.0623f
C1756 A2.n145 GND 0.0238f
C1757 A2.n146 GND 0.0623f
C1758 A2.n147 GND 0.0238f
C1759 A2.n148 GND 0.0623f
C1760 A2.n149 GND 0.0238f
C1761 A2.n150 GND 0.0623f
C1762 A2.n151 GND 0.0238f
C1763 A2.n152 GND 0.0623f
C1764 A2.n153 GND 0.022f
C1765 A2.n154 GND 0.0228f
C1766 A2.n157 GND 0.0313f
C1767 A2.n158 GND 0.0221f
C1768 VDD.n0 GND 0.0156f
C1769 VDD.n3 GND 0.0168f
C1770 VDD.n8 GND 0.0189f
C1771 VDD.n9 GND 0.0763f
C1772 VDD.n11 GND 0.0126f
C1773 VDD.n15 GND 0.0168f
C1774 VDD.n16 GND 0.0168f
C1775 VDD.n17 GND 0.0101f
C1776 VDD.n21 GND 0.044f
C1777 VDD.n54 GND 0.0325f
C1778 VDD.n55 GND 0.0114f
C1779 VDD.n57 GND 0.0112f
C1780 VDD.t257 GND 0.014f
C1781 VDD.t463 GND 0.0351f
C1782 VDD.t786 GND 0.0338f
C1783 VDD.t768 GND 0.0411f
C1784 VDD.t480 GND 0.0354f
C1785 VDD.t767 GND 0.0307f
C1786 VDD.t38 GND 0.0256f
C1787 VDD.t42 GND 0.0405f
C1788 VDD.t83 GND 0.0354f
C1789 VDD.t799 GND 0.0307f
C1790 VDD.t39 GND 0.0307f
C1791 VDD.t764 GND 0.0292f
C1792 VDD.t485 GND 0.0314f
C1793 VDD.t253 GND 0.0312f
C1794 VDD.t592 GND 0.0314f
C1795 VDD.t506 GND 0.0314f
C1796 VDD.t752 GND 0.0397f
C1797 VDD.n58 GND 0.096f
C1798 VDD.n60 GND 0.0106f
C1799 VDD.n62 GND 0.0266f
C1800 VDD.n63 GND 0.64f
C1801 VDD.n66 GND 0.0265f
C1802 VDD.n68 GND 0.181f
C1803 VDD.n72 GND 0.0383f
C1804 VDD.n73 GND 2.87f
C1805 VDD.n77 GND 0.0409f
C1806 VDD.n81 GND 0.0143f
C1807 VDD.n84 GND 0.0169f
C1808 VDD.t541 GND 0.0324f
C1809 VDD.t537 GND 0.0324f
C1810 VDD.t547 GND 0.0297f
C1811 VDD.n87 GND 0.0171f
C1812 VDD.n89 GND 0.0229f
C1813 VDD.n92 GND 0.0229f
C1814 VDD.n94 GND 0.0229f
C1815 VDD.n96 GND 0.0127f
C1816 VDD.n101 GND 0.0142f
C1817 VDD.n103 GND 0.015f
C1818 VDD.n104 GND 0.0131f
C1819 VDD.n108 GND 0.0143f
C1820 VDD.t446 GND 0.0401f
C1821 VDD.n109 GND 0.0409f
C1822 VDD.t620 GND 0.0307f
C1823 VDD.t616 GND 0.0324f
C1824 VDD.t618 GND 0.0324f
C1825 VDD.t614 GND 0.0419f
C1826 VDD.t543 GND 0.0178f
C1827 VDD.n110 GND 0.0243f
C1828 VDD.n111 GND 0.0143f
C1829 VDD.n112 GND 0.0138f
C1830 VDD.n115 GND 0.0131f
C1831 VDD.n119 GND 0.0163f
C1832 VDD.n121 GND 0.0229f
C1833 VDD.n125 GND 0.0229f
C1834 VDD.n127 GND 0.0229f
C1835 VDD.n131 GND 0.018f
C1836 VDD.n132 GND 0.0131f
C1837 VDD.t531 GND 0.0324f
C1838 VDD.t527 GND 0.0324f
C1839 VDD.t533 GND 0.0324f
C1840 VDD.t521 GND 0.0274f
C1841 VDD.t545 GND 0.0324f
C1842 VDD.t535 GND 0.0324f
C1843 VDD.t539 GND 0.0324f
C1844 VDD.t529 GND 0.0212f
C1845 VDD.n135 GND 0.0243f
C1846 VDD.n136 GND 0.0143f
C1847 VDD.n144 GND 0.0164f
C1848 VDD.n148 GND 0.0211f
C1849 VDD.n150 GND 0.0229f
C1850 VDD.n154 GND 0.0229f
C1851 VDD.n156 GND 0.0229f
C1852 VDD.n160 GND 0.0188f
C1853 VDD.n161 GND 0.0131f
C1854 VDD.t708 GND 0.0324f
C1855 VDD.t738 GND 0.0324f
C1856 VDD.t630 GND 0.0324f
C1857 VDD.t622 GND 0.0309f
C1858 VDD.n164 GND 0.0243f
C1859 VDD.t742 GND 0.0178f
C1860 VDD.t730 GND 0.0324f
C1861 VDD.t626 GND 0.0324f
C1862 VDD.t650 GND 0.0324f
C1863 VDD.t642 GND 0.0324f
C1864 VDD.t658 GND 0.0324f
C1865 VDD.t734 GND 0.0313f
C1866 VDD.t525 GND 0.0324f
C1867 VDD.t517 GND 0.0324f
C1868 VDD.t519 GND 0.0324f
C1869 VDD.t523 GND 0.017f
C1870 VDD.n165 GND 0.0339f
C1871 VDD.n166 GND 0.0143f
C1872 VDD.n171 GND 0.0107f
C1873 VDD.n172 GND 0.0135f
C1874 VDD.n174 GND 0.0229f
C1875 VDD.n178 GND 0.0229f
C1876 VDD.n180 GND 0.0229f
C1877 VDD.n184 GND 0.0229f
C1878 VDD.n186 GND 0.0162f
C1879 VDD.n187 GND 0.0164f
C1880 VDD.n196 GND 0.0219f
C1881 VDD.n200 GND 0.0229f
C1882 VDD.n204 GND 0.0229f
C1883 VDD.n206 GND 0.0229f
C1884 VDD.n210 GND 0.0229f
C1885 VDD.n212 GND 0.0229f
C1886 VDD.n216 GND 0.0236f
C1887 VDD.t636 GND 0.0324f
C1888 VDD.t624 GND 0.0324f
C1889 VDD.t648 GND 0.0324f
C1890 VDD.t638 GND 0.0324f
C1891 VDD.t628 GND 0.0324f
C1892 VDD.t652 GND 0.0324f
C1893 VDD.t632 GND 0.0324f
C1894 VDD.t660 GND 0.0282f
C1895 VDD.n220 GND 0.0361f
C1896 VDD.n224 GND 0.0496f
C1897 VDD.n228 GND 0.0496f
C1898 VDD.n230 GND 0.0496f
C1899 VDD.n234 GND 0.0464f
C1900 VDD.n235 GND 0.163f
C1901 VDD.n237 GND 0.0129f
C1902 VDD.n241 GND 0.0229f
C1903 VDD.n243 GND 0.0229f
C1904 VDD.n247 GND 0.0229f
C1905 VDD.n249 GND 0.0183f
C1906 VDD.n250 GND 0.0131f
C1907 VDD.t674 GND 0.0745f
C1908 VDD.t656 GND 0.0324f
C1909 VDD.t646 GND 0.0324f
C1910 VDD.t678 GND 0.0324f
C1911 VDD.t664 GND 0.0324f
C1912 VDD.t690 GND 0.0324f
C1913 VDD.t724 GND 0.0324f
C1914 VDD.t696 GND 0.0324f
C1915 VDD.t682 GND 0.0324f
C1916 VDD.t670 GND 0.0324f
C1917 VDD.t700 GND 0.0324f
C1918 VDD.t728 GND 0.0324f
C1919 VDD.t716 GND 0.0324f
C1920 VDD.t744 GND 0.0324f
C1921 VDD.t688 GND 0.0324f
C1922 VDD.t720 GND 0.0313f
C1923 VDD.t740 GND 0.0324f
C1924 VDD.t710 GND 0.0324f
C1925 VDD.t634 GND 0.0324f
C1926 VDD.t736 GND 0.0324f
C1927 VDD.t748 GND 0.0324f
C1928 VDD.t722 GND 0.0324f
C1929 VDD.t706 GND 0.0324f
C1930 VDD.t712 GND 0.039f
C1931 VDD.n253 GND 0.0339f
C1932 VDD.n254 GND 0.0143f
C1933 VDD.n258 GND 0.0164f
C1934 VDD.n260 GND 0.0209f
C1935 VDD.n264 GND 0.0229f
C1936 VDD.n266 GND 0.0229f
C1937 VDD.n270 GND 0.0229f
C1938 VDD.n272 GND 0.0229f
C1939 VDD.n276 GND 0.0229f
C1940 VDD.n280 GND 0.0229f
C1941 VDD.n282 GND 0.0229f
C1942 VDD.n286 GND 0.0229f
C1943 VDD.n288 GND 0.0229f
C1944 VDD.n292 GND 0.0229f
C1945 VDD.n294 GND 0.0229f
C1946 VDD.n298 GND 0.0229f
C1947 VDD.n300 GND 0.0143f
C1948 VDD.n301 GND 0.0131f
C1949 VDD.n308 GND 0.0671f
C1950 VDD.n310 GND 0.0671f
C1951 VDD.n314 GND 0.0671f
C1952 VDD.n316 GND 0.0671f
C1953 VDD.n320 GND 0.199f
C1954 VDD.n322 GND 0.0229f
C1955 VDD.n323 GND 0.0134f
C1956 VDD.n324 GND 0.0107f
C1957 VDD.n328 GND 0.0143f
C1958 VDD.n329 GND 0.0231f
C1959 VDD.t654 GND 0.0421f
C1960 VDD.t644 GND 0.0326f
C1961 VDD.t676 GND 0.0723f
C1962 VDD.t662 GND 0.0719f
C1963 VDD.t640 GND 0.0719f
C1964 VDD.t680 GND 0.0719f
C1965 VDD.t666 GND 0.0719f
C1966 VDD.t694 GND 0.0719f
C1967 VDD.t668 GND 0.0719f
C1968 VDD.t698 GND 0.0719f
C1969 VDD.t684 GND 0.0719f
C1970 VDD.t672 GND 0.0719f
C1971 VDD.t702 GND 0.0711f
C1972 VDD.t686 GND 0.0497f
C1973 VDD.t718 GND 0.0324f
C1974 VDD.t746 GND 0.0313f
C1975 VDD.t704 GND 0.0332f
C1976 VDD.t726 GND 0.0324f
C1977 VDD.t692 GND 0.0324f
C1978 VDD.t714 GND 0.0324f
C1979 VDD.t732 GND 0.0251f
C1980 VDD.n330 GND 0.0243f
C1981 VDD.n331 GND 0.0143f
C1982 VDD.n334 GND 0.0119f
C1983 VDD.n336 GND 0.021f
C1984 VDD.n337 GND 0.0135f
C1985 VDD.n339 GND 0.0229f
C1986 VDD.n343 GND 0.0179f
C1987 VDD.n344 GND 0.124f
C1988 VDD.n345 GND 0.0482f
C1989 VDD.n349 GND 0.0671f
C1990 VDD.n351 GND 0.0671f
C1991 VDD.n355 GND 0.0671f
C1992 VDD.n357 GND 0.0598f
C1993 VDD.n358 GND 0.563f
C1994 VDD.n359 GND 2.39f
C1995 VDD.n360 GND 1.92f
C1996 VDD.n361 GND 1.13f
C1997 VDD.t784 GND 0.0444f
C1998 VDD.n365 GND 0.0641f
C1999 VDD.n369 GND 0.157f
C2000 VDD.t53 GND 0.0172f
C2001 VDD.t511 GND 0.0165f
C2002 VDD.t85 GND 0.0144f
C2003 VDD.t87 GND 0.0124f
C2004 VDD.t445 GND 0.0183f
C2005 VDD.t612 GND 0.0164f
C2006 VDD.t795 GND 0.023f
C2007 VDD.t388 GND 0.0634f
C2008 VDD.n385 GND 0.0209f
C2009 VDD.n386 GND 0.351f
C2010 VDD.t395 GND 0.0615f
C2011 VDD.t54 GND 0.0213f
C2012 VDD.t56 GND 0.0472f
C2013 VDD.t598 GND 0.088f
C2014 VDD.t439 GND 0.0374f
C2015 VDD.n387 GND 0.0282f
C2016 VDD.n416 GND 0.0158f
C2017 VDD.n417 GND 0.218f
C2018 VDD.t58 GND 0.0171f
C2019 VDD.t490 GND 0.0169f
C2020 VDD.t78 GND 0.0142f
C2021 VDD.t62 GND 0.0176f
C2022 VDD.t4 GND 0.0183f
C2023 VDD.t554 GND 0.0146f
C2024 VDD.t936 GND 0.0383f
C2025 VDD.t40 GND 0.0661f
C2026 VDD.t564 GND 0.0271f
C2027 VDD.t549 GND 0.0285f
C2028 VDD.t394 GND 0.0285f
C2029 VDD.t502 GND 0.0329f
C2030 VDD.t51 GND 0.0534f
C2031 VDD.n420 GND 0.0262f
C2032 VDD.n446 GND 0.0421f
C2033 VDD.n447 GND 0.0177f
C2034 VDD.n448 GND 0.0117f
C2035 VDD.n451 GND 0.0162f
C2036 VDD.n452 GND 0.162f
C2037 VDD.n453 GND 0.0234f
C2038 VDD.n456 GND 0.0389f
C2039 VDD.n460 GND 0.0247f
C2040 VDD.n461 GND 0.0197f
C2041 VDD.n462 GND 0.0247f
C2042 VDD.n465 GND 0.0462f
C2043 VDD.n468 GND 0.0462f
C2044 VDD.n474 GND 0.0462f
C2045 VDD.n475 GND 0.0274f
C2046 VDD.n476 GND 0.0347f
C2047 VDD.n478 GND 0.0176f
C2048 VDD.n479 GND 0.0231f
C2049 VDD.n480 GND 0.0247f
C2050 VDD.t266 GND 0.0154f
C2051 VDD.n481 GND 0.0247f
C2052 VDD.n482 GND 0.0231f
C2053 VDD.n483 GND 0.0176f
C2054 VDD.n484 GND 0.0462f
C2055 VDD.n488 GND 0.0462f
C2056 VDD.n491 GND 0.0462f
C2057 VDD.n494 GND 0.0462f
C2058 VDD.n498 GND 0.0462f
C2059 VDD.n501 GND 0.0235f
C2060 VDD.n502 GND 0.0173f
C2061 VDD.t362 GND 0.0571f
C2062 VDD.t262 GND 0.0249f
C2063 VDD.t368 GND 0.0249f
C2064 VDD.t264 GND 0.0249f
C2065 VDD.t350 GND 0.0249f
C2066 VDD.t372 GND 0.0175f
C2067 VDD.n503 GND 0.0247f
C2068 VDD.n504 GND 0.0231f
C2069 VDD.n505 GND 0.0176f
C2070 VDD.n506 GND 0.0462f
C2071 VDD.n510 GND 0.0294f
C2072 VDD.n514 GND 0.184f
C2073 VDD.n515 GND 0.0419f
C2074 VDD.n517 GND 0.0176f
C2075 VDD.n524 GND 0.0462f
C2076 VDD.n528 GND 0.0462f
C2077 VDD.n529 GND 0.0274f
C2078 VDD.n530 GND 0.0347f
C2079 VDD.n532 GND 0.0455f
C2080 VDD.n542 GND 0.0462f
C2081 VDD.n543 GND 0.0462f
C2082 VDD.n544 GND 0.0462f
C2083 VDD.n550 GND 0.0462f
C2084 VDD.n551 GND 0.0462f
C2085 VDD.n556 GND 0.0462f
C2086 VDD.n557 GND 0.0462f
C2087 VDD.n562 GND 0.0384f
C2088 VDD.n563 GND 0.0247f
C2089 VDD.n564 GND 0.0197f
C2090 VDD.n565 GND 0.0201f
C2091 VDD.t268 GND 0.0198f
C2092 VDD.t384 GND 0.0249f
C2093 VDD.t286 GND 0.0249f
C2094 VDD.t272 GND 0.0249f
C2095 VDD.t260 GND 0.0249f
C2096 VDD.t290 GND 0.0249f
C2097 VDD.t276 GND 0.0249f
C2098 VDD.t308 GND 0.0249f
C2099 VDD.t284 GND 0.0249f
C2100 VDD.t316 GND 0.024f
C2101 VDD.t310 GND 0.0323f
C2102 VDD.t294 GND 0.0249f
C2103 VDD.t282 GND 0.0249f
C2104 VDD.t314 GND 0.0249f
C2105 VDD.t298 GND 0.0207f
C2106 VDD.t370 GND 0.0249f
C2107 VDD.t346 GND 0.0249f
C2108 VDD.t364 GND 0.0249f
C2109 VDD.t342 GND 0.0249f
C2110 VDD.t352 GND 0.0323f
C2111 VDD.t358 GND 0.024f
C2112 VDD.t366 GND 0.0249f
C2113 VDD.t376 GND 0.0249f
C2114 VDD.t354 GND 0.0249f
C2115 VDD.t326 GND 0.0249f
C2116 VDD.t338 GND 0.0249f
C2117 VDD.t304 GND 0.0249f
C2118 VDD.t334 GND 0.0249f
C2119 VDD.t348 GND 0.0249f
C2120 VDD.t318 GND 0.0249f
C2121 VDD.t332 GND 0.0166f
C2122 VDD.n566 GND 0.0201f
C2123 VDD.n567 GND 0.0197f
C2124 VDD.n568 GND 0.0247f
C2125 VDD.n569 GND 0.0309f
C2126 VDD.n570 GND 0.0462f
C2127 VDD.n575 GND 0.0462f
C2128 VDD.n576 GND 0.0462f
C2129 VDD.n581 GND 0.0462f
C2130 VDD.n582 GND 0.0462f
C2131 VDD.n586 GND 0.0274f
C2132 VDD.n587 GND 0.0347f
C2133 VDD.n588 GND 0.0462f
C2134 VDD.n593 GND 0.0462f
C2135 VDD.n594 GND 0.0384f
C2136 VDD.n596 GND 0.0176f
C2137 VDD.n603 GND 0.0462f
C2138 VDD.n609 GND 0.0462f
C2139 VDD.n610 GND 0.0462f
C2140 VDD.n615 GND 0.0462f
C2141 VDD.n616 GND 0.0462f
C2142 VDD.n621 GND 0.0419f
C2143 VDD.n622 GND 0.0247f
C2144 VDD.n623 GND 0.0197f
C2145 VDD.n624 GND 0.0201f
C2146 VDD.t382 GND 0.0219f
C2147 VDD.t374 GND 0.0249f
C2148 VDD.t360 GND 0.0249f
C2149 VDD.t386 GND 0.0249f
C2150 VDD.t288 GND 0.0249f
C2151 VDD.t274 GND 0.0249f
C2152 VDD.t302 GND 0.0249f
C2153 VDD.t378 GND 0.0249f
C2154 VDD.t278 GND 0.0249f
C2155 VDD.t292 GND 0.024f
C2156 VDD.t380 GND 0.0323f
C2157 VDD.t280 GND 0.0249f
C2158 VDD.t312 GND 0.0249f
C2159 VDD.t296 GND 0.0133f
C2160 VDD.n625 GND 0.0201f
C2161 VDD.t330 GND 0.024f
C2162 VDD.t270 GND 0.0249f
C2163 VDD.t300 GND 0.0249f
C2164 VDD.t320 GND 0.0249f
C2165 VDD.t324 GND 0.0249f
C2166 VDD.t336 GND 0.0249f
C2167 VDD.t322 GND 0.0249f
C2168 VDD.t306 GND 0.0249f
C2169 VDD.t340 GND 0.0249f
C2170 VDD.t328 GND 0.0249f
C2171 VDD.t356 GND 0.0249f
C2172 VDD.t344 GND 0.024f
C2173 VDD.t402 GND 0.0323f
C2174 VDD.t416 GND 0.0246f
C2175 VDD.t60 GND 0.0263f
C2176 VDD.t450 GND 0.025f
C2177 VDD.t500 GND 0.0417f
C2178 VDD.t452 GND 0.0308f
C2179 VDD.n627 GND 0.0247f
C2180 VDD.n629 GND 0.0462f
C2181 VDD.n632 GND 0.0462f
C2182 VDD.n636 GND 0.0462f
C2183 VDD.n639 GND 0.0462f
C2184 VDD.n644 GND 0.0176f
C2185 VDD.n648 GND 0.0414f
C2186 VDD.n649 GND 0.0462f
C2187 VDD.n656 GND 0.0462f
C2188 VDD.n657 GND 0.0462f
C2189 VDD.n658 GND 0.0462f
C2190 VDD.n663 GND 0.0462f
C2191 VDD.n664 GND 0.0462f
C2192 VDD.n669 GND 0.0462f
C2193 VDD.n670 GND 0.0274f
C2194 VDD.n671 GND 0.0347f
C2195 VDD.n675 GND 0.0462f
C2196 VDD.n676 GND 0.0462f
C2197 VDD.n677 GND 0.0269f
C2198 VDD.n683 GND 0.0691f
C2199 VDD.n684 GND 0.0538f
C2200 VDD.n685 GND 0.0347f
C2201 VDD.n688 GND 0.0274f
C2202 VDD.n689 GND 0.0304f
C2203 VDD.n692 GND 0.0176f
C2204 VDD.n693 GND 0.0116f
C2205 VDD.n694 GND 0.0197f
C2206 VDD.n695 GND 0.0328f
C2207 VDD.t437 GND 0.0235f
C2208 VDD.t431 GND 0.0249f
C2209 VDD.t433 GND 0.0249f
C2210 VDD.t435 GND 0.0321f
C2211 VDD.t398 GND 0.024f
C2212 VDD.t400 GND 0.0249f
C2213 VDD.t396 GND 0.0249f
C2214 VDD.t422 GND 0.0249f
C2215 VDD.t426 GND 0.0249f
C2216 VDD.t414 GND 0.0249f
C2217 VDD.t420 GND 0.0249f
C2218 VDD.t424 GND 0.0249f
C2219 VDD.t412 GND 0.0249f
C2220 VDD.t418 GND 0.0249f
C2221 VDD.t406 GND 0.0249f
C2222 VDD.t408 GND 0.0249f
C2223 VDD.t404 GND 0.0249f
C2224 VDD.t410 GND 0.0127f
C2225 VDD.n696 GND 0.0201f
C2226 VDD.n697 GND 0.0197f
C2227 VDD.n698 GND 0.0247f
C2228 VDD.n699 GND 0.0389f
C2229 VDD.n705 GND 0.0462f
C2230 VDD.n706 GND 0.0462f
C2231 VDD.n711 GND 0.0462f
C2232 VDD.n712 GND 0.0462f
C2233 VDD.n713 GND 0.0462f
C2234 VDD.n718 GND 0.0462f
C2235 VDD.n719 GND 0.0414f
C2236 VDD.n722 GND 0.0176f
C2237 VDD.n723 GND 0.0231f
C2238 VDD.n724 GND 0.0176f
C2239 VDD.n729 GND 0.0462f
C2240 VDD.n730 GND 0.0347f
C2241 VDD.n731 GND 0.0271f
C2242 VDD.n732 GND 11.2f
C2243 VDD.n756 GND 0.0148f
C2244 VDD.t608 GND 0.157f
C2245 VDD.t2 GND 0.0759f
C2246 VDD.t44 GND 0.159f
C2247 VDD.t76 GND 0.0601f
C2248 VDD.n757 GND 0.0645f
C2249 VDD.n758 GND 0.0928f
C2250 VDD.t494 GND 0.026f
C2251 VDD.t791 GND 0.0174f
C2252 VDD.t930 GND 0.0162f
C2253 VDD.t473 GND 0.0181f
C2254 VDD.t80 GND 0.0166f
C2255 VDD.t475 GND 0.015f
C2256 VDD.t789 GND 0.0215f
C2257 VDD.t47 GND 0.0176f
C2258 VDD.t390 GND 0.0216f
C2259 VDD.t782 GND 0.0335f
C2260 VDD.t606 GND 0.0482f
C2261 VDD.t461 GND 0.0279f
C2262 VDD.t444 GND 0.0293f
C2263 VDD.t505 GND 0.0293f
C2264 VDD.t392 GND 0.0338f
C2265 VDD.t454 GND 0.0557f
C2266 VDD.n763 GND 0.01f
C2267 VDD.n772 GND 0.0187f
C2268 VDD.n780 GND 0.0125f
C2269 VDD.n804 GND 0.0172f
C2270 VDD.n805 GND 0.117f
C2271 VDD.n806 GND 0.0156f
C2272 VDD.n809 GND 0.0168f
C2273 VDD.n814 GND 0.0189f
C2274 VDD.n815 GND 0.0763f
C2275 VDD.n817 GND 0.0126f
C2276 VDD.n821 GND 0.0168f
C2277 VDD.n822 GND 0.0168f
C2278 VDD.n823 GND 0.0101f
C2279 VDD.n827 GND 0.044f
C2280 VDD.n828 GND 0.0112f
C2281 VDD.t570 GND 0.014f
C2282 VDD.t572 GND 0.0351f
C2283 VDD.t478 GND 0.0338f
C2284 VDD.t251 GND 0.0411f
C2285 VDD.t556 GND 0.0354f
C2286 VDD.t611 GND 0.0307f
C2287 VDD.t477 GND 0.0256f
C2288 VDD.t797 GND 0.0405f
C2289 VDD.t552 GND 0.0354f
C2290 VDD.t562 GND 0.0307f
C2291 VDD.t259 GND 0.0307f
C2292 VDD.t510 GND 0.0292f
C2293 VDD.t456 GND 0.0314f
C2294 VDD.t568 GND 0.0312f
C2295 VDD.t64 GND 0.0314f
C2296 VDD.t428 GND 0.0314f
C2297 VDD.t582 GND 0.0397f
C2298 VDD.n831 GND 0.096f
C2299 VDD.n864 GND 0.0325f
C2300 VDD.n865 GND 0.0114f
C2301 VDD.n866 GND 0.0106f
C2302 VDD.n868 GND 0.0266f
C2303 VDD.n869 GND 0.64f
C2304 VDD.n870 GND 0.0455f
C2305 VDD.n871 GND 0.0274f
C2306 VDD.n873 GND 0.0347f
C2307 VDD.n875 GND 0.0176f
C2308 VDD.n876 GND 0.0231f
C2309 VDD.n877 GND 0.0247f
C2310 VDD.t894 GND 0.0148f
C2311 VDD.n878 GND 0.0247f
C2312 VDD.n879 GND 0.0231f
C2313 VDD.n880 GND 0.0176f
C2314 VDD.n881 GND 0.0462f
C2315 VDD.n885 GND 0.0462f
C2316 VDD.n888 GND 0.0462f
C2317 VDD.n891 GND 0.0462f
C2318 VDD.n895 GND 0.0462f
C2319 VDD.n898 GND 0.0223f
C2320 VDD.n899 GND 0.0185f
C2321 VDD.t862 GND 0.0583f
C2322 VDD.t890 GND 0.0249f
C2323 VDD.t868 GND 0.0249f
C2324 VDD.t892 GND 0.0249f
C2325 VDD.t850 GND 0.0249f
C2326 VDD.t872 GND 0.0169f
C2327 VDD.n900 GND 0.0247f
C2328 VDD.n901 GND 0.0231f
C2329 VDD.n902 GND 0.0176f
C2330 VDD.n903 GND 0.0462f
C2331 VDD.n907 GND 0.0297f
C2332 VDD.n911 GND 0.186f
C2333 VDD.n912 GND 0.0409f
C2334 VDD.n914 GND 0.0176f
C2335 VDD.n921 GND 0.0462f
C2336 VDD.n925 GND 0.0462f
C2337 VDD.n926 GND 0.0274f
C2338 VDD.n927 GND 0.0347f
C2339 VDD.n929 GND 0.0445f
C2340 VDD.n939 GND 0.0462f
C2341 VDD.n940 GND 0.0462f
C2342 VDD.n941 GND 0.0462f
C2343 VDD.n947 GND 0.0462f
C2344 VDD.n948 GND 0.0462f
C2345 VDD.n953 GND 0.0462f
C2346 VDD.n954 GND 0.0462f
C2347 VDD.n959 GND 0.0394f
C2348 VDD.n960 GND 0.0247f
C2349 VDD.n961 GND 0.0197f
C2350 VDD.n962 GND 0.0201f
C2351 VDD.t896 GND 0.0204f
C2352 VDD.t886 GND 0.0249f
C2353 VDD.t914 GND 0.0249f
C2354 VDD.t900 GND 0.0249f
C2355 VDD.t888 GND 0.0249f
C2356 VDD.t918 GND 0.0249f
C2357 VDD.t906 GND 0.0249f
C2358 VDD.t806 GND 0.0249f
C2359 VDD.t912 GND 0.0249f
C2360 VDD.t816 GND 0.024f
C2361 VDD.t810 GND 0.0323f
C2362 VDD.t922 GND 0.0249f
C2363 VDD.t910 GND 0.0249f
C2364 VDD.t814 GND 0.0249f
C2365 VDD.t926 GND 0.0201f
C2366 VDD.t870 GND 0.0249f
C2367 VDD.t848 GND 0.0249f
C2368 VDD.t864 GND 0.0249f
C2369 VDD.t842 GND 0.0249f
C2370 VDD.t852 GND 0.0323f
C2371 VDD.t858 GND 0.024f
C2372 VDD.t866 GND 0.0249f
C2373 VDD.t876 GND 0.0249f
C2374 VDD.t854 GND 0.0249f
C2375 VDD.t824 GND 0.0249f
C2376 VDD.t838 GND 0.0249f
C2377 VDD.t804 GND 0.0249f
C2378 VDD.t834 GND 0.0249f
C2379 VDD.t846 GND 0.0249f
C2380 VDD.t818 GND 0.0249f
C2381 VDD.t830 GND 0.0172f
C2382 VDD.n963 GND 0.0201f
C2383 VDD.n964 GND 0.0197f
C2384 VDD.n965 GND 0.0247f
C2385 VDD.n966 GND 0.0319f
C2386 VDD.n967 GND 0.0462f
C2387 VDD.n972 GND 0.0462f
C2388 VDD.n973 GND 0.0462f
C2389 VDD.n978 GND 0.0462f
C2390 VDD.n979 GND 0.0462f
C2391 VDD.n983 GND 0.0274f
C2392 VDD.n984 GND 0.0347f
C2393 VDD.n985 GND 0.0462f
C2394 VDD.n990 GND 0.0462f
C2395 VDD.n991 GND 0.0374f
C2396 VDD.n993 GND 0.0176f
C2397 VDD.n1000 GND 0.0462f
C2398 VDD.n1004 GND 0.0462f
C2399 VDD.n1009 GND 0.0462f
C2400 VDD.n1010 GND 0.0462f
C2401 VDD.n1015 GND 0.0429f
C2402 VDD.n1016 GND 0.0247f
C2403 VDD.n1017 GND 0.0197f
C2404 VDD.n1018 GND 0.0201f
C2405 VDD.t882 GND 0.0225f
C2406 VDD.t874 GND 0.0249f
C2407 VDD.t860 GND 0.0249f
C2408 VDD.t884 GND 0.0249f
C2409 VDD.t916 GND 0.0249f
C2410 VDD.t902 GND 0.0249f
C2411 VDD.t802 GND 0.0249f
C2412 VDD.t878 GND 0.0249f
C2413 VDD.t904 GND 0.0249f
C2414 VDD.t920 GND 0.024f
C2415 VDD.t880 GND 0.0323f
C2416 VDD.t908 GND 0.0249f
C2417 VDD.t812 GND 0.0249f
C2418 VDD.t924 GND 0.0127f
C2419 VDD.n1019 GND 0.0197f
C2420 VDD.t46 GND 0.0263f
C2421 VDD.t49 GND 0.025f
C2422 VDD.t496 GND 0.0417f
C2423 VDD.t565 GND 0.0314f
C2424 VDD.n1021 GND 0.0247f
C2425 VDD.n1023 GND 0.0462f
C2426 VDD.n1026 GND 0.0462f
C2427 VDD.n1030 GND 0.0462f
C2428 VDD.n1033 GND 0.0462f
C2429 VDD.n1036 GND 0.0231f
C2430 VDD.n1040 GND 0.0462f
C2431 VDD.n1044 GND 0.0462f
C2432 VDD.n1052 GND 0.0176f
C2433 VDD.n1057 GND 0.0424f
C2434 VDD.n1058 GND 0.0462f
C2435 VDD.n1059 GND 0.0462f
C2436 VDD.n1066 GND 0.0462f
C2437 VDD.n1067 GND 0.0462f
C2438 VDD.n1068 GND 0.0462f
C2439 VDD.n1074 GND 0.0462f
C2440 VDD.n1075 GND 0.0462f
C2441 VDD.n1076 GND 0.0274f
C2442 VDD.n1079 GND 0.0347f
C2443 VDD.n1080 GND 0.0379f
C2444 VDD.n1081 GND 0.0247f
C2445 VDD.n1082 GND 0.0176f
C2446 VDD.n1088 GND 0.0176f
C2447 VDD.n1089 GND 0.0247f
C2448 VDD.n1090 GND 0.0424f
C2449 VDD.n1091 GND 0.0462f
C2450 VDD.n1098 GND 0.0462f
C2451 VDD.n1099 GND 0.0462f
C2452 VDD.n1100 GND 0.0462f
C2453 VDD.n1105 GND 0.0462f
C2454 VDD.n1106 GND 0.0462f
C2455 VDD.n1111 GND 0.0462f
C2456 VDD.n1112 GND 0.0274f
C2457 VDD.n1113 GND 0.0347f
C2458 VDD.n1117 GND 0.0462f
C2459 VDD.n1118 GND 0.0462f
C2460 VDD.n1119 GND 0.0259f
C2461 VDD.n1125 GND 0.0691f
C2462 VDD.n1126 GND 0.0538f
C2463 VDD.n1127 GND 0.0347f
C2464 VDD.n1130 GND 0.0274f
C2465 VDD.n1131 GND 0.0314f
C2466 VDD.n1134 GND 0.0176f
C2467 VDD.n1135 GND 0.0116f
C2468 VDD.n1136 GND 0.0197f
C2469 VDD.n1137 GND 0.0328f
C2470 VDD.t776 GND 0.0235f
C2471 VDD.t778 GND 0.0249f
C2472 VDD.t780 GND 0.0249f
C2473 VDD.t774 GND 0.0321f
C2474 VDD.t36 GND 0.024f
C2475 VDD.t6 GND 0.0249f
C2476 VDD.t34 GND 0.0249f
C2477 VDD.t28 GND 0.0249f
C2478 VDD.t32 GND 0.0249f
C2479 VDD.t20 GND 0.0249f
C2480 VDD.t26 GND 0.0249f
C2481 VDD.t30 GND 0.0249f
C2482 VDD.t18 GND 0.0249f
C2483 VDD.t24 GND 0.0249f
C2484 VDD.t12 GND 0.0249f
C2485 VDD.t14 GND 0.0249f
C2486 VDD.t10 GND 0.0249f
C2487 VDD.t16 GND 0.0133f
C2488 VDD.n1138 GND 0.0201f
C2489 VDD.t22 GND 0.024f
C2490 VDD.t8 GND 0.0323f
C2491 VDD.t844 GND 0.024f
C2492 VDD.t856 GND 0.0249f
C2493 VDD.t826 GND 0.0249f
C2494 VDD.t840 GND 0.0249f
C2495 VDD.t808 GND 0.0249f
C2496 VDD.t822 GND 0.0249f
C2497 VDD.t836 GND 0.0249f
C2498 VDD.t820 GND 0.0249f
C2499 VDD.t832 GND 0.0249f
C2500 VDD.t928 GND 0.0249f
C2501 VDD.t898 GND 0.0249f
C2502 VDD.t828 GND 0.0246f
C2503 VDD.n1139 GND 0.0201f
C2504 VDD.n1140 GND 0.0197f
C2505 VDD.n1141 GND 0.0247f
C2506 VDD.n1142 GND 0.0379f
C2507 VDD.n1143 GND 0.0462f
C2508 VDD.n1148 GND 0.0239f
C2509 VDD.n1149 GND 11.2f
C2510 VDD.t61 GND 0.0172f
C2511 VDD.t580 GND 0.0165f
C2512 VDD.t498 GND 0.0144f
C2513 VDD.t469 GND 0.0124f
C2514 VDD.t430 GND 0.0183f
C2515 VDD.t793 GND 0.0164f
C2516 VDD.t467 GND 0.023f
C2517 VDD.t594 GND 0.0634f
C2518 VDD.n1165 GND 0.0209f
C2519 VDD.n1166 GND 0.351f
C2520 VDD.t484 GND 0.0615f
C2521 VDD.t471 GND 0.0213f
C2522 VDD.t255 GND 0.0472f
C2523 VDD.t492 GND 0.088f
C2524 VDD.t459 GND 0.0374f
C2525 VDD.n1167 GND 0.0282f
C2526 VDD.n1196 GND 0.0158f
C2527 VDD.n1197 GND 0.218f
C2528 VDD.t442 GND 0.0171f
C2529 VDD.t574 GND 0.0169f
C2530 VDD.t600 GND 0.0142f
C2531 VDD.t513 GND 0.0176f
C2532 VDD.t933 GND 0.0183f
C2533 VDD.t448 GND 0.0146f
C2534 VDD.t576 GND 0.0383f
C2535 VDD.t68 GND 0.0661f
C2536 VDD.t770 GND 0.0271f
C2537 VDD.t86 GND 0.0285f
C2538 VDD.t773 GND 0.0285f
C2539 VDD.t482 GND 0.0329f
C2540 VDD.t765 GND 0.0534f
C2541 VDD.n1200 GND 0.0262f
C2542 VDD.n1226 GND 0.0421f
C2543 VDD.n1227 GND 0.0177f
C2544 VDD.n1228 GND 0.0117f
C2545 VDD.n1231 GND 0.0162f
C2546 VDD.n1232 GND 0.162f
C2547 VDD.n1233 GND 0.0234f
C2548 VDD.n1236 GND 0.0389f
C2549 VDD.n1240 GND 0.0247f
C2550 VDD.n1241 GND 0.0197f
C2551 VDD.n1242 GND 0.0247f
C2552 VDD.n1245 GND 0.0462f
C2553 VDD.n1248 GND 0.0462f
C2554 VDD.n1254 GND 0.0462f
C2555 VDD.n1255 GND 0.0274f
C2556 VDD.n1256 GND 0.0347f
C2557 VDD.n1258 GND 0.0176f
C2558 VDD.n1259 GND 0.0231f
C2559 VDD.n1260 GND 0.0247f
C2560 VDD.t113 GND 0.0154f
C2561 VDD.n1261 GND 0.0247f
C2562 VDD.n1262 GND 0.0231f
C2563 VDD.n1263 GND 0.0176f
C2564 VDD.n1264 GND 0.0462f
C2565 VDD.n1268 GND 0.0462f
C2566 VDD.n1271 GND 0.0462f
C2567 VDD.n1274 GND 0.0462f
C2568 VDD.n1278 GND 0.0462f
C2569 VDD.n1281 GND 0.0235f
C2570 VDD.n1282 GND 0.0173f
C2571 VDD.t187 GND 0.0571f
C2572 VDD.t95 GND 0.0249f
C2573 VDD.t213 GND 0.0249f
C2574 VDD.t111 GND 0.0249f
C2575 VDD.t185 GND 0.0249f
C2576 VDD.t217 GND 0.0175f
C2577 VDD.n1283 GND 0.0247f
C2578 VDD.n1284 GND 0.0231f
C2579 VDD.n1285 GND 0.0176f
C2580 VDD.n1286 GND 0.0462f
C2581 VDD.n1290 GND 0.0294f
C2582 VDD.n1294 GND 0.184f
C2583 VDD.n1295 GND 0.0419f
C2584 VDD.n1297 GND 0.0176f
C2585 VDD.n1304 GND 0.0462f
C2586 VDD.n1308 GND 0.0462f
C2587 VDD.n1309 GND 0.0274f
C2588 VDD.n1310 GND 0.0347f
C2589 VDD.n1312 GND 0.0455f
C2590 VDD.n1322 GND 0.0462f
C2591 VDD.n1323 GND 0.0462f
C2592 VDD.n1324 GND 0.0462f
C2593 VDD.n1330 GND 0.0462f
C2594 VDD.n1331 GND 0.0462f
C2595 VDD.n1336 GND 0.0462f
C2596 VDD.n1337 GND 0.0462f
C2597 VDD.n1342 GND 0.0384f
C2598 VDD.n1343 GND 0.0247f
C2599 VDD.n1344 GND 0.0197f
C2600 VDD.n1345 GND 0.0201f
C2601 VDD.t115 GND 0.0198f
C2602 VDD.t165 GND 0.0249f
C2603 VDD.t201 GND 0.0249f
C2604 VDD.t125 GND 0.0249f
C2605 VDD.t169 GND 0.0249f
C2606 VDD.t205 GND 0.0249f
C2607 VDD.t129 GND 0.0249f
C2608 VDD.t151 GND 0.0249f
C2609 VDD.t145 GND 0.0249f
C2610 VDD.t177 GND 0.024f
C2611 VDD.t105 GND 0.0323f
C2612 VDD.t155 GND 0.0249f
C2613 VDD.t211 GND 0.0249f
C2614 VDD.t109 GND 0.0249f
C2615 VDD.t159 GND 0.0207f
C2616 VDD.t215 GND 0.0249f
C2617 VDD.t183 GND 0.0249f
C2618 VDD.t191 GND 0.0249f
C2619 VDD.t153 GND 0.0249f
C2620 VDD.t103 GND 0.0323f
C2621 VDD.t175 GND 0.024f
C2622 VDD.t133 GND 0.0249f
C2623 VDD.t207 GND 0.0249f
C2624 VDD.t171 GND 0.0249f
C2625 VDD.t141 GND 0.0249f
C2626 VDD.t97 GND 0.0249f
C2627 VDD.t189 GND 0.0249f
C2628 VDD.t199 GND 0.0249f
C2629 VDD.t147 GND 0.0249f
C2630 VDD.t121 GND 0.0249f
C2631 VDD.t181 GND 0.0166f
C2632 VDD.n1346 GND 0.0201f
C2633 VDD.n1347 GND 0.0197f
C2634 VDD.n1348 GND 0.0247f
C2635 VDD.n1349 GND 0.0309f
C2636 VDD.n1350 GND 0.0462f
C2637 VDD.n1355 GND 0.0462f
C2638 VDD.n1356 GND 0.0462f
C2639 VDD.n1361 GND 0.0462f
C2640 VDD.n1362 GND 0.0462f
C2641 VDD.n1366 GND 0.0274f
C2642 VDD.n1367 GND 0.0347f
C2643 VDD.n1368 GND 0.0462f
C2644 VDD.n1373 GND 0.0462f
C2645 VDD.n1374 GND 0.0384f
C2646 VDD.n1376 GND 0.0176f
C2647 VDD.n1383 GND 0.0462f
C2648 VDD.n1389 GND 0.0462f
C2649 VDD.n1390 GND 0.0462f
C2650 VDD.n1395 GND 0.0462f
C2651 VDD.n1396 GND 0.0462f
C2652 VDD.n1401 GND 0.0419f
C2653 VDD.n1402 GND 0.0247f
C2654 VDD.n1403 GND 0.0197f
C2655 VDD.n1404 GND 0.0201f
C2656 VDD.t163 GND 0.0219f
C2657 VDD.t91 GND 0.0249f
C2658 VDD.t137 GND 0.0249f
C2659 VDD.t167 GND 0.0249f
C2660 VDD.t203 GND 0.0249f
C2661 VDD.t127 GND 0.0249f
C2662 VDD.t149 GND 0.0249f
C2663 VDD.t117 GND 0.0249f
C2664 VDD.t131 GND 0.0249f
C2665 VDD.t101 GND 0.024f
C2666 VDD.t179 GND 0.0323f
C2667 VDD.t209 GND 0.0249f
C2668 VDD.t107 GND 0.0249f
C2669 VDD.t157 GND 0.0133f
C2670 VDD.n1405 GND 0.0201f
C2671 VDD.t195 GND 0.024f
C2672 VDD.t135 GND 0.0249f
C2673 VDD.t161 GND 0.0249f
C2674 VDD.t197 GND 0.0249f
C2675 VDD.t123 GND 0.0249f
C2676 VDD.t93 GND 0.0249f
C2677 VDD.t139 GND 0.0249f
C2678 VDD.t193 GND 0.0249f
C2679 VDD.t99 GND 0.0249f
C2680 VDD.t143 GND 0.0249f
C2681 VDD.t173 GND 0.0249f
C2682 VDD.t119 GND 0.024f
C2683 VDD.t237 GND 0.0323f
C2684 VDD.t247 GND 0.0246f
C2685 VDD.t563 GND 0.0263f
C2686 VDD.t465 GND 0.025f
C2687 VDD.t750 GND 0.0417f
C2688 VDD.t560 GND 0.0308f
C2689 VDD.n1407 GND 0.0247f
C2690 VDD.n1409 GND 0.0462f
C2691 VDD.n1412 GND 0.0462f
C2692 VDD.n1416 GND 0.0462f
C2693 VDD.n1419 GND 0.0462f
C2694 VDD.n1424 GND 0.0176f
C2695 VDD.n1428 GND 0.0414f
C2696 VDD.n1429 GND 0.0462f
C2697 VDD.n1436 GND 0.0462f
C2698 VDD.n1437 GND 0.0462f
C2699 VDD.n1438 GND 0.0462f
C2700 VDD.n1443 GND 0.0462f
C2701 VDD.n1444 GND 0.0462f
C2702 VDD.n1449 GND 0.0462f
C2703 VDD.n1450 GND 0.0274f
C2704 VDD.n1451 GND 0.0347f
C2705 VDD.n1455 GND 0.0462f
C2706 VDD.n1456 GND 0.0462f
C2707 VDD.n1457 GND 0.0269f
C2708 VDD.n1463 GND 0.0691f
C2709 VDD.n1464 GND 0.0538f
C2710 VDD.n1465 GND 0.0347f
C2711 VDD.n1468 GND 0.0274f
C2712 VDD.n1469 GND 0.0304f
C2713 VDD.n1472 GND 0.0176f
C2714 VDD.n1473 GND 0.0116f
C2715 VDD.n1474 GND 0.0197f
C2716 VDD.n1475 GND 0.0328f
C2717 VDD.t758 GND 0.0235f
C2718 VDD.t754 GND 0.0249f
C2719 VDD.t760 GND 0.0249f
C2720 VDD.t756 GND 0.0321f
C2721 VDD.t233 GND 0.024f
C2722 VDD.t235 GND 0.0249f
C2723 VDD.t227 GND 0.0249f
C2724 VDD.t221 GND 0.0249f
C2725 VDD.t243 GND 0.0249f
C2726 VDD.t231 GND 0.0249f
C2727 VDD.t219 GND 0.0249f
C2728 VDD.t241 GND 0.0249f
C2729 VDD.t229 GND 0.0249f
C2730 VDD.t249 GND 0.0249f
C2731 VDD.t245 GND 0.0249f
C2732 VDD.t223 GND 0.0249f
C2733 VDD.t239 GND 0.0249f
C2734 VDD.t225 GND 0.0127f
C2735 VDD.n1476 GND 0.0201f
C2736 VDD.n1477 GND 0.0197f
C2737 VDD.n1478 GND 0.0247f
C2738 VDD.n1479 GND 0.0389f
C2739 VDD.n1485 GND 0.0462f
C2740 VDD.n1486 GND 0.0462f
C2741 VDD.n1491 GND 0.0462f
C2742 VDD.n1492 GND 0.0462f
C2743 VDD.n1493 GND 0.0462f
C2744 VDD.n1498 GND 0.0462f
C2745 VDD.n1499 GND 0.0414f
C2746 VDD.n1502 GND 0.0176f
C2747 VDD.n1503 GND 0.0231f
C2748 VDD.n1504 GND 0.0176f
C2749 VDD.n1509 GND 0.0462f
C2750 VDD.n1510 GND 0.0347f
C2751 VDD.n1511 GND 0.0271f
C2752 VDD.n1512 GND 11.2f
C2753 VDD.n1536 GND 0.0148f
C2754 VDD.t939 GND 0.157f
C2755 VDD.t508 GND 0.0759f
C2756 VDD.t89 GND 0.159f
C2757 VDD.t72 GND 0.0601f
C2758 VDD.n1537 GND 0.0645f
C2759 VDD.n1538 GND 0.0928f
C2760 VDD.t66 GND 0.026f
C2761 VDD.t70 GND 0.0174f
C2762 VDD.t596 GND 0.0162f
C2763 VDD.t578 GND 0.0181f
C2764 VDD.t602 GND 0.0166f
C2765 VDD.t550 GND 0.015f
C2766 VDD.t74 GND 0.0215f
C2767 VDD.t590 GND 0.0176f
C2768 VDD.t587 GND 0.0216f
C2769 VDD.t0 GND 0.0335f
C2770 VDD.t558 GND 0.0482f
C2771 VDD.t499 GND 0.0279f
C2772 VDD.t441 GND 0.0293f
C2773 VDD.t489 GND 0.0293f
C2774 VDD.t771 GND 0.0338f
C2775 VDD.t762 GND 0.0557f
C2776 VDD.n1543 GND 0.01f
C2777 VDD.n1552 GND 0.0187f
C2778 VDD.n1560 GND 0.0125f
C2779 VDD.n1584 GND 0.0172f
C2780 VDD.n1585 GND 0.117f
C2781 VDD.n1586 GND 0.637f
C2782 VDD.n1587 GND 0.994f
C2783 VDD.n1588 GND 1.5f
C2784 VDD.n1589 GND 0.632f
C2785 VDD.n1590 GND 1.1f
C2786 VDD.n1591 GND 0.812f
C2787 VDD.n1592 GND 1.52f
C2788 VDD.n1593 GND 0.798f
C2789 VDD.n1594 GND 1.15f
C2790 VDD.n1595 GND 0.912f
C2791 VDD.n1596 GND 1.5f
C2792 VDD.n1597 GND 0.714f
C2793 VDD.n1598 GND 1.1f
C2794 VDD.n1599 GND 0.79f
C2795 VDD.n1600 GND 0.607f
C2796 VDD.n1601 GND 2.85f
.ends

