magic
tech sky130A
magscale 1 2
timestamp 1717121788
<< nwell >>
rect 747 -340 4700 68
rect 1250 -1394 5200 -952
<< pwell >>
rect 884 -578 5032 -510
rect 884 -680 5050 -578
rect 884 -850 5032 -680
<< psubdiff >>
rect 1476 -646 1500 -612
rect 1600 -646 1624 -612
rect 2326 -646 2350 -612
rect 2450 -646 2474 -612
rect 3176 -646 3200 -612
rect 3300 -646 3324 -612
rect 4026 -646 4050 -612
rect 4150 -646 4174 -612
rect 4876 -646 4900 -612
rect 5000 -646 5024 -612
rect 920 -680 960 -656
rect 920 -744 960 -720
<< nsubdiff >>
rect 1500 -34 1550 0
rect 1600 -34 1650 0
rect 1950 -34 2000 0
rect 2050 -34 2100 0
rect 2400 -34 2450 0
rect 2500 -34 2550 0
rect 2850 -34 2900 0
rect 2950 -34 3000 0
rect 3300 -34 3350 0
rect 3400 -34 3450 0
rect 3750 -34 3800 0
rect 3850 -34 3900 0
rect 4200 -34 4250 0
rect 4300 -34 4350 0
rect 1400 -1292 1450 -1258
rect 1500 -1292 1550 -1258
rect 1850 -1292 1900 -1258
rect 1950 -1292 2000 -1258
rect 2300 -1292 2350 -1258
rect 2400 -1292 2450 -1258
rect 2750 -1292 2800 -1258
rect 2850 -1292 2900 -1258
rect 3200 -1292 3250 -1258
rect 3300 -1292 3350 -1258
rect 3650 -1292 3700 -1258
rect 3750 -1292 3800 -1258
rect 4100 -1292 4150 -1258
rect 4200 -1292 4250 -1258
rect 4678 -1284 4728 -1250
rect 4778 -1284 4828 -1250
<< psubdiffcont >>
rect 1500 -646 1600 -612
rect 2350 -646 2450 -612
rect 3200 -646 3300 -612
rect 4050 -646 4150 -612
rect 4900 -646 5000 -612
rect 920 -720 960 -680
<< nsubdiffcont >>
rect 1550 -34 1600 0
rect 2000 -34 2050 0
rect 2450 -34 2500 0
rect 2900 -34 2950 0
rect 3350 -34 3400 0
rect 3800 -34 3850 0
rect 4250 -34 4300 0
rect 1450 -1292 1500 -1258
rect 1900 -1292 1950 -1258
rect 2350 -1292 2400 -1258
rect 2800 -1292 2850 -1258
rect 3250 -1292 3300 -1258
rect 3700 -1292 3750 -1258
rect 4150 -1292 4200 -1258
rect 4728 -1284 4778 -1250
<< locali >>
rect 1500 0 1650 34
rect 1500 -34 1550 0
rect 1600 -34 1650 0
rect 1950 0 2100 34
rect 1950 -34 2000 0
rect 2050 -34 2100 0
rect 2400 0 2550 34
rect 2400 -34 2450 0
rect 2500 -34 2550 0
rect 2850 0 3000 34
rect 2850 -34 2900 0
rect 2950 -34 3000 0
rect 3300 0 3450 34
rect 3300 -34 3350 0
rect 3400 -34 3450 0
rect 3750 0 3900 34
rect 3750 -34 3800 0
rect 3850 -34 3900 0
rect 4200 0 4350 34
rect 4200 -34 4250 0
rect 4300 -34 4350 0
rect 1250 -331 1450 -325
rect 1250 -369 1256 -331
rect 1294 -369 1406 -331
rect 1444 -369 1450 -331
rect 1250 -375 1450 -369
rect 920 -680 960 -600
rect 1450 -612 1650 -578
rect 1450 -646 1500 -612
rect 1600 -646 1650 -612
rect 1450 -680 1650 -646
rect 2300 -612 2500 -578
rect 2300 -646 2350 -612
rect 2450 -646 2500 -612
rect 2300 -680 2500 -646
rect 3150 -612 3350 -578
rect 3150 -646 3200 -612
rect 3300 -646 3350 -612
rect 3150 -680 3350 -646
rect 4000 -612 4200 -578
rect 4000 -646 4050 -612
rect 4150 -646 4200 -612
rect 4000 -680 4200 -646
rect 4850 -612 5050 -578
rect 4850 -646 4900 -612
rect 5000 -646 5050 -612
rect 4850 -680 5050 -646
rect 920 -736 960 -720
rect 1400 -1258 1550 -1224
rect 1400 -1292 1450 -1258
rect 1500 -1292 1550 -1258
rect 1850 -1258 2000 -1224
rect 1850 -1292 1900 -1258
rect 1950 -1292 2000 -1258
rect 2300 -1258 2450 -1224
rect 2300 -1292 2350 -1258
rect 2400 -1292 2450 -1258
rect 2750 -1258 2900 -1224
rect 2750 -1292 2800 -1258
rect 2850 -1292 2900 -1258
rect 3200 -1258 3350 -1224
rect 3200 -1292 3250 -1258
rect 3300 -1292 3350 -1258
rect 3650 -1258 3800 -1224
rect 3650 -1292 3700 -1258
rect 3750 -1292 3800 -1258
rect 4100 -1258 4250 -1224
rect 4100 -1292 4150 -1258
rect 4200 -1292 4250 -1258
rect 4678 -1250 4828 -1216
rect 4678 -1284 4728 -1250
rect 4778 -1284 4828 -1250
<< viali >>
rect 1707 -318 1744 -281
rect 1081 -369 1119 -331
rect 1256 -369 1294 -331
rect 1406 -369 1444 -331
rect 1855 -370 1895 -330
rect 2206 -368 2243 -331
rect 2531 -369 2569 -331
rect 2831 -369 2869 -331
rect 3151 -374 3199 -327
rect 3406 -369 3444 -331
rect 3556 -369 3594 -331
rect 3976 -374 4024 -327
rect 4231 -369 4269 -331
rect 4406 -369 4444 -331
rect 1051 -849 1099 -801
rect 1201 -924 1249 -876
rect 1355 -945 1395 -905
rect 1855 -945 1895 -905
rect 2306 -943 2344 -905
rect 2555 -945 2595 -905
rect 2705 -945 2745 -905
rect 3006 -944 3044 -906
rect 3355 -945 3395 -905
rect 3556 -944 3594 -906
rect 1700 -1000 1750 -950
rect 3856 -969 3894 -931
rect 4026 -948 4074 -901
rect 4406 -944 4444 -906
rect 4655 -945 4695 -905
rect 4805 -945 4845 -905
<< metal1 >>
rect 1594 -150 1600 -50
rect 1700 -150 1706 -50
rect 1700 -250 2250 -200
rect 1700 -281 1750 -250
rect 1700 -318 1707 -281
rect 1744 -318 1750 -281
rect 1075 -331 1125 -319
rect 1700 -325 1750 -318
rect 1075 -369 1081 -331
rect 1119 -369 1125 -331
rect 1075 -425 1125 -369
rect 1244 -331 1456 -325
rect 1701 -330 1750 -325
rect 1244 -369 1256 -331
rect 1294 -369 1406 -331
rect 1444 -369 1456 -331
rect 1244 -375 1456 -369
rect 1843 -376 1849 -324
rect 1901 -376 1907 -324
rect 2200 -325 2250 -250
rect 3400 -275 4450 -225
rect 2693 -325 2699 -324
rect 2200 -331 2249 -325
rect 2200 -368 2206 -331
rect 2243 -368 2249 -331
rect 2200 -380 2249 -368
rect 2519 -331 2699 -325
rect 2519 -369 2531 -331
rect 2569 -369 2699 -331
rect 2519 -375 2699 -369
rect 2693 -376 2699 -375
rect 2751 -376 2757 -324
rect 2825 -331 2875 -319
rect 2825 -369 2831 -331
rect 2869 -369 2875 -331
rect 1343 -425 1349 -424
rect 1075 -475 1349 -425
rect 1343 -476 1349 -475
rect 1401 -476 1407 -424
rect 2543 -476 2549 -424
rect 2601 -425 2607 -424
rect 2825 -425 2875 -369
rect 3139 -380 3145 -320
rect 3205 -380 3211 -320
rect 3400 -331 3450 -275
rect 3400 -369 3406 -331
rect 3444 -369 3450 -331
rect 3400 -381 3450 -369
rect 3550 -331 3600 -319
rect 3550 -369 3556 -331
rect 3594 -369 3600 -331
rect 2601 -475 2875 -425
rect 2601 -476 2607 -475
rect 3343 -476 3349 -424
rect 3401 -425 3407 -424
rect 3550 -425 3600 -369
rect 3964 -380 3970 -320
rect 4030 -380 4036 -320
rect 4225 -331 4275 -319
rect 4225 -369 4231 -331
rect 4269 -369 4275 -331
rect 3401 -475 3600 -425
rect 4225 -425 4275 -369
rect 4400 -331 4450 -275
rect 4400 -369 4406 -331
rect 4444 -369 4450 -331
rect 4400 -381 4450 -369
rect 4799 -424 4851 -418
rect 4225 -475 4799 -425
rect 3401 -476 3407 -475
rect 4799 -482 4851 -476
rect 990 -700 1000 -600
rect 1100 -700 1110 -600
rect 1025 -795 1125 -775
rect 1025 -855 1045 -795
rect 1105 -855 1125 -795
rect 1025 -875 1125 -855
rect 3850 -850 4450 -800
rect 1189 -930 1195 -870
rect 1255 -930 1261 -870
rect 1343 -951 1349 -899
rect 1401 -951 1407 -899
rect 1688 -950 1762 -944
rect 1688 -1000 1700 -950
rect 1750 -1000 1762 -950
rect 1843 -951 1849 -899
rect 1901 -951 1907 -899
rect 2300 -905 2350 -893
rect 2300 -943 2306 -905
rect 2344 -943 2350 -905
rect 2300 -1000 2350 -943
rect 2543 -951 2549 -899
rect 2601 -951 2607 -899
rect 2693 -951 2699 -899
rect 2751 -951 2757 -899
rect 3000 -906 3050 -894
rect 3000 -944 3006 -906
rect 3044 -944 3050 -906
rect 1688 -1006 2350 -1000
rect 1700 -1050 2350 -1006
rect 2550 -1000 2600 -951
rect 3000 -1000 3050 -944
rect 3343 -951 3349 -899
rect 3401 -951 3407 -899
rect 3550 -906 3600 -894
rect 3550 -944 3556 -906
rect 3594 -944 3600 -906
rect 3550 -1000 3600 -944
rect 3850 -931 3900 -850
rect 3850 -969 3856 -931
rect 3894 -969 3900 -931
rect 4014 -955 4020 -895
rect 4080 -955 4086 -895
rect 4400 -906 4450 -850
rect 4400 -944 4406 -906
rect 4444 -944 4450 -906
rect 4400 -956 4450 -944
rect 4643 -951 4649 -899
rect 4701 -951 4707 -899
rect 4793 -951 4799 -899
rect 4851 -951 4857 -899
rect 3850 -981 3900 -969
rect 2550 -1050 3600 -1000
rect 1590 -1300 1600 -1200
rect 1700 -1300 1710 -1200
<< via1 >>
rect 1600 -150 1700 -50
rect 1849 -330 1901 -324
rect 1849 -370 1855 -330
rect 1855 -370 1895 -330
rect 1895 -370 1901 -330
rect 1849 -376 1901 -370
rect 2699 -376 2751 -324
rect 1349 -476 1401 -424
rect 2549 -476 2601 -424
rect 3145 -327 3205 -320
rect 3145 -374 3151 -327
rect 3151 -374 3199 -327
rect 3199 -374 3205 -327
rect 3145 -380 3205 -374
rect 3349 -476 3401 -424
rect 3970 -327 4030 -320
rect 3970 -374 3976 -327
rect 3976 -374 4024 -327
rect 4024 -374 4030 -327
rect 3970 -380 4030 -374
rect 4799 -476 4851 -424
rect 1000 -700 1100 -600
rect 1045 -801 1105 -795
rect 1045 -849 1051 -801
rect 1051 -849 1099 -801
rect 1099 -849 1105 -801
rect 1045 -855 1105 -849
rect 1195 -876 1255 -870
rect 1195 -924 1201 -876
rect 1201 -924 1249 -876
rect 1249 -924 1255 -876
rect 1195 -930 1255 -924
rect 1349 -905 1401 -899
rect 1349 -945 1355 -905
rect 1355 -945 1395 -905
rect 1395 -945 1401 -905
rect 1349 -951 1401 -945
rect 1849 -905 1901 -899
rect 1849 -945 1855 -905
rect 1855 -945 1895 -905
rect 1895 -945 1901 -905
rect 1849 -951 1901 -945
rect 2549 -905 2601 -899
rect 2549 -945 2555 -905
rect 2555 -945 2595 -905
rect 2595 -945 2601 -905
rect 2549 -951 2601 -945
rect 2699 -905 2751 -899
rect 2699 -945 2705 -905
rect 2705 -945 2745 -905
rect 2745 -945 2751 -905
rect 2699 -951 2751 -945
rect 3349 -905 3401 -899
rect 3349 -945 3355 -905
rect 3355 -945 3395 -905
rect 3395 -945 3401 -905
rect 3349 -951 3401 -945
rect 4020 -901 4080 -895
rect 4020 -948 4026 -901
rect 4026 -948 4074 -901
rect 4074 -948 4080 -901
rect 4020 -955 4080 -948
rect 4649 -905 4701 -899
rect 4649 -945 4655 -905
rect 4655 -945 4695 -905
rect 4695 -945 4701 -905
rect 4649 -951 4701 -945
rect 4799 -905 4851 -899
rect 4799 -945 4805 -905
rect 4805 -945 4845 -905
rect 4845 -945 4851 -905
rect 4799 -951 4851 -945
rect 1600 -1300 1700 -1200
<< metal2 >>
rect 1600 2250 1700 2259
rect 1600 -50 1700 2150
rect 1300 -400 1400 -390
rect 1400 -424 1425 -400
rect 1401 -475 1425 -424
rect 1400 -482 1401 -476
rect 1300 -510 1400 -500
rect 1000 -600 1100 -590
rect 1000 -710 1100 -700
rect 1025 -795 1125 -775
rect 1025 -855 1045 -795
rect 1105 -855 1125 -795
rect 1025 -875 1125 -855
rect 1195 -870 1255 -864
rect 1350 -893 1400 -510
rect 1195 -967 1255 -930
rect 1349 -899 1401 -893
rect 1349 -957 1401 -951
rect 1195 -1023 1197 -967
rect 1253 -1023 1255 -967
rect 1195 -1025 1255 -1023
rect 1197 -1032 1253 -1025
rect 1600 -1200 1700 -150
rect 1849 -324 1901 -318
rect 1849 -382 1901 -376
rect 2699 -324 2751 -318
rect 2699 -382 2751 -376
rect 3145 -320 3205 -314
rect 1850 -786 1900 -382
rect 2549 -424 2601 -418
rect 2549 -482 2601 -476
rect 1845 -795 1905 -786
rect 1845 -864 1905 -855
rect 1850 -893 1900 -864
rect 2550 -893 2600 -482
rect 2700 -893 2750 -382
rect 1849 -899 1901 -893
rect 1849 -957 1901 -951
rect 2549 -899 2601 -893
rect 2549 -957 2601 -951
rect 2699 -899 2751 -893
rect 2699 -957 2751 -951
rect 3145 -967 3205 -380
rect 3970 -320 4030 -314
rect 3349 -424 3401 -418
rect 3349 -482 3401 -476
rect 3350 -893 3400 -482
rect 3970 -522 4030 -380
rect 4800 -400 4900 -390
rect 4793 -476 4799 -424
rect 4800 -510 4900 -500
rect 4645 -520 4705 -511
rect 3963 -578 3972 -522
rect 4028 -578 4037 -522
rect 3970 -580 4030 -578
rect 4645 -589 4705 -580
rect 3349 -899 3401 -893
rect 3349 -957 3401 -951
rect 4020 -895 4080 -889
rect 4650 -893 4700 -589
rect 4800 -893 4850 -510
rect 4020 -967 4080 -955
rect 4649 -899 4701 -893
rect 4649 -957 4701 -951
rect 4799 -899 4851 -893
rect 4799 -957 4851 -951
rect 3138 -1023 3147 -967
rect 3203 -1023 3212 -967
rect 4020 -1023 4022 -967
rect 4078 -1023 4080 -967
rect 3145 -1025 3205 -1023
rect 4020 -1025 4080 -1023
rect 4022 -1032 4078 -1025
rect 1600 -1310 1700 -1300
<< via2 >>
rect 1600 2150 1700 2250
rect 1300 -424 1400 -400
rect 1300 -476 1349 -424
rect 1349 -476 1400 -424
rect 1300 -500 1400 -476
rect 1000 -700 1100 -600
rect 1047 -853 1103 -797
rect 1197 -1023 1253 -967
rect 1845 -855 1905 -795
rect 4800 -424 4900 -400
rect 4800 -476 4851 -424
rect 4851 -476 4900 -424
rect 4800 -500 4900 -476
rect 3972 -578 4028 -522
rect 4645 -580 4705 -520
rect 3147 -1023 3203 -967
rect 4022 -1023 4078 -967
<< metal3 >>
rect 4500 11400 5300 12200
rect -22500 9800 -21700 10600
rect -4549 9349 -4251 9355
rect -5100 9051 -4549 9300
rect -4251 9051 -4200 9300
rect -5100 8900 -4200 9051
rect 1583 2255 1713 2263
rect 1583 2145 1595 2255
rect 1705 2145 1713 2255
rect 1583 2140 1713 2145
rect -4550 -200 -4250 -194
rect -4250 -400 300 -200
rect 4800 -395 5000 -300
rect 1290 -400 1410 -395
rect -4250 -500 1300 -400
rect 1400 -500 1410 -400
rect -4550 -506 -4250 -500
rect 1290 -505 1410 -500
rect 4790 -400 5000 -395
rect 4790 -500 4800 -400
rect 4900 -500 5000 -400
rect 4790 -505 4910 -500
rect 3967 -520 4033 -517
rect 4640 -520 4710 -515
rect 3967 -522 4645 -520
rect 3967 -578 3972 -522
rect 4028 -578 4645 -522
rect 3967 -580 4645 -578
rect 4705 -580 4710 -520
rect 3967 -583 4033 -580
rect 4640 -585 4710 -580
rect 990 -600 1110 -595
rect -2000 -700 -1950 -600
rect -1850 -700 1000 -600
rect 1100 -700 1110 -600
rect 990 -705 1110 -700
rect 1025 -795 1125 -775
rect 1840 -795 1910 -790
rect 1025 -797 1845 -795
rect 1025 -800 1047 -797
rect 300 -853 1047 -800
rect 1103 -853 1845 -797
rect 300 -855 1845 -853
rect 1905 -855 1910 -795
rect 300 -875 1125 -855
rect 1840 -860 1910 -855
rect 300 -900 1100 -875
rect 300 -1000 500 -900
rect 1192 -965 1258 -962
rect 3142 -965 3208 -962
rect 4017 -965 4083 -962
rect 1192 -967 4083 -965
rect 1192 -1023 1197 -967
rect 1253 -1023 3147 -967
rect 3203 -1023 4022 -967
rect 4078 -1023 4083 -967
rect 1192 -1025 4083 -1023
rect 1192 -1028 1258 -1025
rect 3142 -1028 3208 -1025
rect 4017 -1028 4083 -1025
<< via3 >>
rect -4549 9051 -4251 9349
rect 1595 2250 1705 2255
rect 1595 2150 1600 2250
rect 1600 2150 1700 2250
rect 1700 2150 1705 2250
rect 1595 2145 1705 2150
rect -4550 -500 -4250 -200
rect -1950 -700 -1850 -600
<< metal4 >>
rect -4550 9349 -4250 9350
rect -4550 9051 -4549 9349
rect -4251 9051 -4250 9349
rect -4550 -199 -4250 9051
rect 200 2255 3900 3500
rect 200 2145 1595 2255
rect 1705 2145 3900 2255
rect 200 2000 3900 2145
rect -4551 -200 -4249 -199
rect -4551 -500 -4550 -200
rect -4250 -500 -4249 -200
rect -4551 -501 -4249 -500
rect -1951 -600 -1849 -599
rect -1951 -700 -1950 -600
rect -1850 -700 -1849 -600
rect -1951 -701 -1849 -700
rect -17100 -15200 -12400 -13200
use C2S2_Fingers_Amplifier  C2S2_Fingers_Amplifier_0
timestamp 1716868724
transform 1 0 -52296 0 1 -678100
box 29796 662800 57684 701260
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3430 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x3
timestamp 1701704242
transform -1 0 2974 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x4
timestamp 1701704242
transform 1 0 2142 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x5
timestamp 1701704242
transform -1 0 2146 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x6
timestamp 1701704242
transform 1 0 1314 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 858 0 1 -592
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  x9
timestamp 1701704242
transform 1 0 3802 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x10
timestamp 1701704242
transform 1 0 4258 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x11
timestamp 1701704242
transform 1 0 2974 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  x13
timestamp 1701704242
transform 1 0 2970 0 -1 -683
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  x14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1038 0 -1 -683
box -38 -48 314 592
<< labels >>
rlabel metal3 4800 -500 5000 -300 1 OUT
port 2 n
rlabel metal3 -22500 9800 -21700 10600 1 SIG
port 3 n
rlabel metal3 4500 11400 5300 12200 1 VMID
port 4 n
rlabel metal4 -17100 -15200 -12400 -13200 1 VSS
port 5 n
rlabel metal4 200 2000 3900 3500 1 VDD
port 6 n
rlabel metal3 300 -1000 500 -800 1 CLK
port 7 n
<< end >>
