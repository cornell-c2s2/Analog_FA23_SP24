* NGSPICE file created from RSfetsym-lvs.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_8X7CJE a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_ENQT6S a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_CBNSG2 a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_GNLSML a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_K7FRP5 w_n226_n419# a_30_n200# a_n33_n297# a_n88_n200#
X0 a_30_n200# a_n33_n297# a_n88_n200# w_n226_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
.ends

.subckt sky130_fd_pr__pfet_01v8_GHY9W9 w_n226_n419# a_30_n200# a_n33_n297# a_n88_n200#
X0 a_30_n200# a_n33_n297# a_n88_n200# w_n226_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
.ends

.subckt sky130_fd_pr__pfet_01v8_E3L9V7 a_21_231# a_79_n200# w_n275_n419# a_n87_n297#
+ a_n137_n200# a_n29_n200#
X0 a_n29_n200# a_n87_n297# a_n137_n200# w_n275_n419# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1 a_79_n200# a_21_231# a_n29_n200# w_n275_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
.ends

.subckt sky130_fd_pr__pfet_01v8_EDASV7 a_21_231# a_79_n200# w_n275_n419# a_n87_n297#
+ a_n137_n200# a_n29_n200#
X0 a_n29_n200# a_n87_n297# a_n137_n200# w_n275_n419# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1 a_79_n200# a_21_231# a_n29_n200# w_n275_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
.ends

.subckt sky130_fd_pr__nfet_01v8_4WSMTB a_n185_n374# a_n83_n200# a_25_n200# a_n33_n288#
X0 a_25_n200# a_n33_n288# a_n83_n200# a_n185_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
.ends

.subckt sky130_fd_pr__nfet_01v8_XJSMYS a_n185_n374# a_n83_n200# a_25_n200# a_n33_n288#
X0 a_25_n200# a_n33_n288# a_n83_n200# a_n185_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
.ends

.subckt RSfetsym-lvs VDD S R Q QN GND
Xx1 R GND GND VDD VDD x1/Y sky130_fd_sc_hd__inv_4
Xx2 S GND GND VDD VDD x2/Y sky130_fd_sc_hd__inv_4
XXM1 QN S m1_1070_n1180# GND sky130_fd_pr__nfet_01v8_8X7CJE
XXM2 m1_1070_n1180# Q GND GND sky130_fd_pr__nfet_01v8_ENQT6S
XXM3 Q R m1_1580_n1170# GND sky130_fd_pr__nfet_01v8_CBNSG2
XXM4 m1_1580_n1170# QN GND GND sky130_fd_pr__nfet_01v8_GNLSML
XXM5 VDD QN Q VDD sky130_fd_pr__pfet_01v8_K7FRP5
XXM6 VDD Q QN VDD sky130_fd_pr__pfet_01v8_GHY9W9
XXM7 S VDD VDD S VDD QN sky130_fd_pr__pfet_01v8_E3L9V7
XXM8 R VDD VDD R VDD Q sky130_fd_pr__pfet_01v8_EDASV7
XXM9 GND QN GND x1/Y sky130_fd_pr__nfet_01v8_4WSMTB
XXM10 GND Q GND x2/Y sky130_fd_pr__nfet_01v8_XJSMYS
.ends

