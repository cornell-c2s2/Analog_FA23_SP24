magic
tech sky130A
timestamp 1713142167
<< end >>
