magic
tech sky130A
magscale 1 2
timestamp 1713142632
<< pwell >>
rect -3223 -5974 3223 5974
<< psubdiff >>
rect -3187 5904 -3091 5938
rect 3091 5904 3187 5938
rect -3187 5842 -3153 5904
rect 3153 5842 3187 5904
rect -3187 -5904 -3153 -5842
rect 3153 -5904 3187 -5842
rect -3187 -5938 -3091 -5904
rect 3091 -5938 3187 -5904
<< psubdiffcont >>
rect -3091 5904 3091 5938
rect -3187 -5842 -3153 5842
rect 3153 -5842 3187 5842
rect -3091 -5938 3091 -5904
<< xpolycontact >>
rect 1911 5376 3057 5808
rect -3057 -5808 -1911 -5376
<< xpolyres >>
rect -3057 5271 -1911 5272
rect -1815 5271 -669 5272
rect -3057 4125 -669 5271
rect -3057 -5376 -1911 4125
rect -1815 -4126 -669 4125
rect -573 5271 573 5272
rect 669 5271 1815 5272
rect -573 4125 1815 5271
rect -573 -4126 573 4125
rect -1815 -5272 573 -4126
rect 669 -4126 1815 4125
rect 1911 -4126 3057 5376
rect 669 -5272 3057 -4126
<< locali >>
rect -3187 5904 -3091 5938
rect 3091 5904 3187 5938
rect -3187 5842 -3153 5904
rect 3153 5842 3187 5904
rect -3187 -5904 -3153 -5842
rect 3153 -5904 3187 -5842
rect -3187 -5938 -3091 -5904
rect 3091 -5938 3187 -5904
<< properties >>
string FIXED_BBOX -3170 -5921 3170 5921
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 52.716 m 1 nx 5 wmin 5.730 lmin 0.50 rho 2000 val 100.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
