magic
tech sky130A
magscale 1 2
timestamp 1710000196
<< pwell >>
rect -673 -325 673 325
<< nmos >>
rect -487 -125 -287 125
rect -229 -125 -29 125
rect 29 -125 229 125
rect 287 -125 487 125
<< ndiff >>
rect -545 85 -487 125
rect -545 51 -533 85
rect -499 51 -487 85
rect -545 17 -487 51
rect -545 -17 -533 17
rect -499 -17 -487 17
rect -545 -51 -487 -17
rect -545 -85 -533 -51
rect -499 -85 -487 -51
rect -545 -125 -487 -85
rect -287 85 -229 125
rect -287 51 -275 85
rect -241 51 -229 85
rect -287 17 -229 51
rect -287 -17 -275 17
rect -241 -17 -229 17
rect -287 -51 -229 -17
rect -287 -85 -275 -51
rect -241 -85 -229 -51
rect -287 -125 -229 -85
rect -29 85 29 125
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -125 29 -85
rect 229 85 287 125
rect 229 51 241 85
rect 275 51 287 85
rect 229 17 287 51
rect 229 -17 241 17
rect 275 -17 287 17
rect 229 -51 287 -17
rect 229 -85 241 -51
rect 275 -85 287 -51
rect 229 -125 287 -85
rect 487 85 545 125
rect 487 51 499 85
rect 533 51 545 85
rect 487 17 545 51
rect 487 -17 499 17
rect 533 -17 545 17
rect 487 -51 545 -17
rect 487 -85 499 -51
rect 533 -85 545 -51
rect 487 -125 545 -85
<< ndiffc >>
rect -533 51 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -51
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 499 51 533 85
rect 499 -17 533 17
rect 499 -85 533 -51
<< psubdiff >>
rect -647 265 -527 299
rect -493 265 -459 299
rect -425 265 -391 299
rect -357 265 -323 299
rect -289 265 -255 299
rect -221 265 -187 299
rect -153 265 -119 299
rect -85 265 -51 299
rect -17 265 17 299
rect 51 265 85 299
rect 119 265 153 299
rect 187 265 221 299
rect 255 265 289 299
rect 323 265 357 299
rect 391 265 425 299
rect 459 265 493 299
rect 527 265 647 299
rect -647 187 -613 265
rect -647 119 -613 153
rect 613 187 647 265
rect -647 51 -613 85
rect -647 -17 -613 17
rect -647 -85 -613 -51
rect -647 -153 -613 -119
rect 613 119 647 153
rect 613 51 647 85
rect 613 -17 647 17
rect 613 -85 647 -51
rect -647 -265 -613 -187
rect 613 -153 647 -119
rect 613 -265 647 -187
rect -647 -299 -527 -265
rect -493 -299 -459 -265
rect -425 -299 -391 -265
rect -357 -299 -323 -265
rect -289 -299 -255 -265
rect -221 -299 -187 -265
rect -153 -299 -119 -265
rect -85 -299 -51 -265
rect -17 -299 17 -265
rect 51 -299 85 -265
rect 119 -299 153 -265
rect 187 -299 221 -265
rect 255 -299 289 -265
rect 323 -299 357 -265
rect 391 -299 425 -265
rect 459 -299 493 -265
rect 527 -299 647 -265
<< psubdiffcont >>
rect -527 265 -493 299
rect -459 265 -425 299
rect -391 265 -357 299
rect -323 265 -289 299
rect -255 265 -221 299
rect -187 265 -153 299
rect -119 265 -85 299
rect -51 265 -17 299
rect 17 265 51 299
rect 85 265 119 299
rect 153 265 187 299
rect 221 265 255 299
rect 289 265 323 299
rect 357 265 391 299
rect 425 265 459 299
rect 493 265 527 299
rect -647 153 -613 187
rect 613 153 647 187
rect -647 85 -613 119
rect -647 17 -613 51
rect -647 -51 -613 -17
rect -647 -119 -613 -85
rect 613 85 647 119
rect 613 17 647 51
rect 613 -51 647 -17
rect 613 -119 647 -85
rect -647 -187 -613 -153
rect 613 -187 647 -153
rect -527 -299 -493 -265
rect -459 -299 -425 -265
rect -391 -299 -357 -265
rect -323 -299 -289 -265
rect -255 -299 -221 -265
rect -187 -299 -153 -265
rect -119 -299 -85 -265
rect -51 -299 -17 -265
rect 17 -299 51 -265
rect 85 -299 119 -265
rect 153 -299 187 -265
rect 221 -299 255 -265
rect 289 -299 323 -265
rect 357 -299 391 -265
rect 425 -299 459 -265
rect 493 -299 527 -265
<< poly >>
rect -487 197 -287 213
rect -487 163 -438 197
rect -404 163 -370 197
rect -336 163 -287 197
rect -487 125 -287 163
rect -229 197 -29 213
rect -229 163 -180 197
rect -146 163 -112 197
rect -78 163 -29 197
rect -229 125 -29 163
rect 29 197 229 213
rect 29 163 78 197
rect 112 163 146 197
rect 180 163 229 197
rect 29 125 229 163
rect 287 197 487 213
rect 287 163 336 197
rect 370 163 404 197
rect 438 163 487 197
rect 287 125 487 163
rect -487 -163 -287 -125
rect -487 -197 -438 -163
rect -404 -197 -370 -163
rect -336 -197 -287 -163
rect -487 -213 -287 -197
rect -229 -163 -29 -125
rect -229 -197 -180 -163
rect -146 -197 -112 -163
rect -78 -197 -29 -163
rect -229 -213 -29 -197
rect 29 -163 229 -125
rect 29 -197 78 -163
rect 112 -197 146 -163
rect 180 -197 229 -163
rect 29 -213 229 -197
rect 287 -163 487 -125
rect 287 -197 336 -163
rect 370 -197 404 -163
rect 438 -197 487 -163
rect 287 -213 487 -197
<< polycont >>
rect -438 163 -404 197
rect -370 163 -336 197
rect -180 163 -146 197
rect -112 163 -78 197
rect 78 163 112 197
rect 146 163 180 197
rect 336 163 370 197
rect 404 163 438 197
rect -438 -197 -404 -163
rect -370 -197 -336 -163
rect -180 -197 -146 -163
rect -112 -197 -78 -163
rect 78 -197 112 -163
rect 146 -197 180 -163
rect 336 -197 370 -163
rect 404 -197 438 -163
<< locali >>
rect -647 265 -527 299
rect -493 265 -459 299
rect -425 265 -391 299
rect -357 265 -323 299
rect -289 265 -255 299
rect -221 265 -187 299
rect -153 265 -119 299
rect -85 265 -51 299
rect -17 265 17 299
rect 51 265 85 299
rect 119 265 153 299
rect 187 265 221 299
rect 255 265 289 299
rect 323 265 357 299
rect 391 265 425 299
rect 459 265 493 299
rect 527 265 647 299
rect -647 187 -613 265
rect -487 163 -440 197
rect -404 163 -370 197
rect -334 163 -287 197
rect -229 163 -182 197
rect -146 163 -112 197
rect -76 163 -29 197
rect 29 163 76 197
rect 112 163 146 197
rect 182 163 229 197
rect 287 163 334 197
rect 370 163 404 197
rect 440 163 487 197
rect 613 187 647 265
rect -647 119 -613 153
rect -647 51 -613 85
rect -647 -17 -613 17
rect -647 -85 -613 -51
rect -647 -153 -613 -119
rect -533 89 -499 129
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -129 -499 -89
rect -275 89 -241 129
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -129 -241 -89
rect -17 89 17 129
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -129 17 -89
rect 241 89 275 129
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -129 275 -89
rect 499 89 533 129
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -129 533 -89
rect 613 119 647 153
rect 613 51 647 85
rect 613 -17 647 17
rect 613 -85 647 -51
rect 613 -153 647 -119
rect -647 -265 -613 -187
rect -487 -197 -440 -163
rect -404 -197 -370 -163
rect -334 -197 -287 -163
rect -229 -197 -182 -163
rect -146 -197 -112 -163
rect -76 -197 -29 -163
rect 29 -197 76 -163
rect 112 -197 146 -163
rect 182 -197 229 -163
rect 287 -197 334 -163
rect 370 -197 404 -163
rect 440 -197 487 -163
rect 613 -265 647 -187
rect -647 -299 -527 -265
rect -493 -299 -459 -265
rect -425 -299 -391 -265
rect -357 -299 -323 -265
rect -289 -299 -255 -265
rect -221 -299 -187 -265
rect -153 -299 -119 -265
rect -85 -299 -51 -265
rect -17 -299 17 -265
rect 51 -299 85 -265
rect 119 -299 153 -265
rect 187 -299 221 -265
rect 255 -299 289 -265
rect 323 -299 357 -265
rect 391 -299 425 -265
rect 459 -299 493 -265
rect 527 -299 647 -265
<< viali >>
rect -440 163 -438 197
rect -438 163 -406 197
rect -368 163 -336 197
rect -336 163 -334 197
rect -182 163 -180 197
rect -180 163 -148 197
rect -110 163 -78 197
rect -78 163 -76 197
rect 76 163 78 197
rect 78 163 110 197
rect 148 163 180 197
rect 180 163 182 197
rect 334 163 336 197
rect 336 163 368 197
rect 406 163 438 197
rect 438 163 440 197
rect -533 85 -499 89
rect -533 55 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -55
rect -533 -89 -499 -85
rect -275 85 -241 89
rect -275 55 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -55
rect -275 -89 -241 -85
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect 241 85 275 89
rect 241 55 275 85
rect 241 -17 275 17
rect 241 -85 275 -55
rect 241 -89 275 -85
rect 499 85 533 89
rect 499 55 533 85
rect 499 -17 533 17
rect 499 -85 533 -55
rect 499 -89 533 -85
rect -440 -197 -438 -163
rect -438 -197 -406 -163
rect -368 -197 -336 -163
rect -336 -197 -334 -163
rect -182 -197 -180 -163
rect -180 -197 -148 -163
rect -110 -197 -78 -163
rect -78 -197 -76 -163
rect 76 -197 78 -163
rect 78 -197 110 -163
rect 148 -197 180 -163
rect 180 -197 182 -163
rect 334 -197 336 -163
rect 336 -197 368 -163
rect 406 -197 438 -163
rect 438 -197 440 -163
<< metal1 >>
rect -483 197 -291 203
rect -483 163 -440 197
rect -406 163 -368 197
rect -334 163 -291 197
rect -483 157 -291 163
rect -225 197 -33 203
rect -225 163 -182 197
rect -148 163 -110 197
rect -76 163 -33 197
rect -225 157 -33 163
rect 33 197 225 203
rect 33 163 76 197
rect 110 163 148 197
rect 182 163 225 197
rect 33 157 225 163
rect 291 197 483 203
rect 291 163 334 197
rect 368 163 406 197
rect 440 163 483 197
rect 291 157 483 163
rect -539 89 -493 125
rect -539 55 -533 89
rect -499 55 -493 89
rect -539 17 -493 55
rect -539 -17 -533 17
rect -499 -17 -493 17
rect -539 -55 -493 -17
rect -539 -89 -533 -55
rect -499 -89 -493 -55
rect -539 -125 -493 -89
rect -281 89 -235 125
rect -281 55 -275 89
rect -241 55 -235 89
rect -281 17 -235 55
rect -281 -17 -275 17
rect -241 -17 -235 17
rect -281 -55 -235 -17
rect -281 -89 -275 -55
rect -241 -89 -235 -55
rect -281 -125 -235 -89
rect -23 89 23 125
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -125 23 -89
rect 235 89 281 125
rect 235 55 241 89
rect 275 55 281 89
rect 235 17 281 55
rect 235 -17 241 17
rect 275 -17 281 17
rect 235 -55 281 -17
rect 235 -89 241 -55
rect 275 -89 281 -55
rect 235 -125 281 -89
rect 493 89 539 125
rect 493 55 499 89
rect 533 55 539 89
rect 493 17 539 55
rect 493 -17 499 17
rect 533 -17 539 17
rect 493 -55 539 -17
rect 493 -89 499 -55
rect 533 -89 539 -55
rect 493 -125 539 -89
rect -483 -163 -291 -157
rect -483 -197 -440 -163
rect -406 -197 -368 -163
rect -334 -197 -291 -163
rect -483 -203 -291 -197
rect -225 -163 -33 -157
rect -225 -197 -182 -163
rect -148 -197 -110 -163
rect -76 -197 -33 -163
rect -225 -203 -33 -197
rect 33 -163 225 -157
rect 33 -197 76 -163
rect 110 -197 148 -163
rect 182 -197 225 -163
rect 33 -203 225 -197
rect 291 -163 483 -157
rect 291 -197 334 -163
rect 368 -197 406 -163
rect 440 -197 483 -163
rect 291 -203 483 -197
<< properties >>
string FIXED_BBOX -630 -282 630 282
<< end >>
