magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< pwell >>
rect -739 -850 739 850
<< psubdiff >>
rect -703 780 -607 814
rect 607 780 703 814
rect -703 718 -669 780
rect 669 718 703 780
rect -703 -780 -669 -718
rect 669 -780 703 -718
rect -703 -814 -607 -780
rect 607 -814 703 -780
<< psubdiffcont >>
rect -607 780 607 814
rect -703 -718 -669 718
rect 669 -718 703 718
rect -607 -814 607 -780
<< xpolycontact >>
rect -573 252 573 684
rect -573 -684 573 -252
<< xpolyres >>
rect -573 -252 573 252
<< locali >>
rect -703 780 -607 814
rect 607 780 703 814
rect -703 718 -669 780
rect 669 718 703 780
rect -703 -780 -669 -718
rect 669 -780 703 -718
rect -703 -814 -607 -780
rect 607 -814 703 -780
<< viali >>
rect -557 269 557 666
rect -557 -666 557 -269
<< metal1 >>
rect -569 666 569 672
rect -569 269 -557 666
rect 557 269 569 666
rect -569 263 569 269
rect -569 -269 569 -263
rect -569 -666 -557 -269
rect 557 -666 569 -269
rect -569 -672 569 -666
<< properties >>
string FIXED_BBOX -686 -797 686 797
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 2.677 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 1.0k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
