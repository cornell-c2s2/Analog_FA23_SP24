magic
tech sky130A
magscale 1 2
timestamp 1714231380
<< nwell >>
rect 1766 227 3330 4465
<< pwell >>
rect 1190 -5 1632 322
rect -2527 -1225 6511 -5
rect -2530 -4098 15822 -1248
<< pmoslvt >>
rect 1962 446 2162 4246
rect 2448 446 2648 4246
rect 2934 446 3134 4246
<< nmoslvt >>
rect 1338 96 1422 126
rect -2331 -1015 -2211 -215
rect -1925 -1015 -1805 -215
rect -1519 -1015 -1399 -215
rect -1113 -1015 -993 -215
rect -707 -1015 -587 -215
rect -301 -1015 -181 -215
rect 105 -1015 225 -215
rect 511 -1015 631 -215
rect 917 -1015 1037 -215
rect 1323 -1015 1443 -215
rect 1729 -1015 1849 -215
rect 2135 -1015 2255 -215
rect 2541 -1015 2661 -215
rect 2947 -1015 3067 -215
rect 3353 -1015 3473 -215
rect 3759 -1015 3879 -215
rect 4165 -1015 4285 -215
rect 4571 -1015 4691 -215
rect 4977 -1015 5097 -215
rect 5383 -1015 5503 -215
rect 5789 -1015 5909 -215
rect 6195 -1015 6315 -215
<< ndiff >>
rect 1338 172 1422 184
rect 1338 138 1350 172
rect 1410 138 1422 172
rect 1338 126 1422 138
rect 1338 84 1422 96
rect 1338 50 1350 84
rect 1410 50 1422 84
rect 1338 38 1422 50
rect -2389 -227 -2331 -215
rect -2389 -1003 -2377 -227
rect -2343 -1003 -2331 -227
rect -2389 -1015 -2331 -1003
rect -2211 -227 -2153 -215
rect -2211 -1003 -2199 -227
rect -2165 -1003 -2153 -227
rect -2211 -1015 -2153 -1003
rect -1983 -227 -1925 -215
rect -1983 -1003 -1971 -227
rect -1937 -1003 -1925 -227
rect -1983 -1015 -1925 -1003
rect -1805 -227 -1747 -215
rect -1805 -1003 -1793 -227
rect -1759 -1003 -1747 -227
rect -1805 -1015 -1747 -1003
rect -1577 -227 -1519 -215
rect -1577 -1003 -1565 -227
rect -1531 -1003 -1519 -227
rect -1577 -1015 -1519 -1003
rect -1399 -227 -1341 -215
rect -1399 -1003 -1387 -227
rect -1353 -1003 -1341 -227
rect -1399 -1015 -1341 -1003
rect -1171 -227 -1113 -215
rect -1171 -1003 -1159 -227
rect -1125 -1003 -1113 -227
rect -1171 -1015 -1113 -1003
rect -993 -227 -935 -215
rect -993 -1003 -981 -227
rect -947 -1003 -935 -227
rect -993 -1015 -935 -1003
rect -765 -227 -707 -215
rect -765 -1003 -753 -227
rect -719 -1003 -707 -227
rect -765 -1015 -707 -1003
rect -587 -227 -529 -215
rect -587 -1003 -575 -227
rect -541 -1003 -529 -227
rect -587 -1015 -529 -1003
rect -359 -227 -301 -215
rect -359 -1003 -347 -227
rect -313 -1003 -301 -227
rect -359 -1015 -301 -1003
rect -181 -227 -123 -215
rect -181 -1003 -169 -227
rect -135 -1003 -123 -227
rect -181 -1015 -123 -1003
rect 47 -227 105 -215
rect 47 -1003 59 -227
rect 93 -1003 105 -227
rect 47 -1015 105 -1003
rect 225 -227 283 -215
rect 225 -1003 237 -227
rect 271 -1003 283 -227
rect 225 -1015 283 -1003
rect 453 -227 511 -215
rect 453 -1003 465 -227
rect 499 -1003 511 -227
rect 453 -1015 511 -1003
rect 631 -227 689 -215
rect 631 -1003 643 -227
rect 677 -1003 689 -227
rect 631 -1015 689 -1003
rect 859 -227 917 -215
rect 859 -1003 871 -227
rect 905 -1003 917 -227
rect 859 -1015 917 -1003
rect 1037 -227 1095 -215
rect 1037 -1003 1049 -227
rect 1083 -1003 1095 -227
rect 1037 -1015 1095 -1003
rect 1265 -227 1323 -215
rect 1265 -1003 1277 -227
rect 1311 -1003 1323 -227
rect 1265 -1015 1323 -1003
rect 1443 -227 1501 -215
rect 1443 -1003 1455 -227
rect 1489 -1003 1501 -227
rect 1443 -1015 1501 -1003
rect 1671 -227 1729 -215
rect 1671 -1003 1683 -227
rect 1717 -1003 1729 -227
rect 1671 -1015 1729 -1003
rect 1849 -227 1907 -215
rect 1849 -1003 1861 -227
rect 1895 -1003 1907 -227
rect 1849 -1015 1907 -1003
rect 2077 -227 2135 -215
rect 2077 -1003 2089 -227
rect 2123 -1003 2135 -227
rect 2077 -1015 2135 -1003
rect 2255 -227 2313 -215
rect 2255 -1003 2267 -227
rect 2301 -1003 2313 -227
rect 2255 -1015 2313 -1003
rect 2483 -227 2541 -215
rect 2483 -1003 2495 -227
rect 2529 -1003 2541 -227
rect 2483 -1015 2541 -1003
rect 2661 -227 2719 -215
rect 2661 -1003 2673 -227
rect 2707 -1003 2719 -227
rect 2661 -1015 2719 -1003
rect 2889 -227 2947 -215
rect 2889 -1003 2901 -227
rect 2935 -1003 2947 -227
rect 2889 -1015 2947 -1003
rect 3067 -227 3125 -215
rect 3067 -1003 3079 -227
rect 3113 -1003 3125 -227
rect 3067 -1015 3125 -1003
rect 3295 -227 3353 -215
rect 3295 -1003 3307 -227
rect 3341 -1003 3353 -227
rect 3295 -1015 3353 -1003
rect 3473 -227 3531 -215
rect 3473 -1003 3485 -227
rect 3519 -1003 3531 -227
rect 3473 -1015 3531 -1003
rect 3701 -227 3759 -215
rect 3701 -1003 3713 -227
rect 3747 -1003 3759 -227
rect 3701 -1015 3759 -1003
rect 3879 -227 3937 -215
rect 3879 -1003 3891 -227
rect 3925 -1003 3937 -227
rect 3879 -1015 3937 -1003
rect 4107 -227 4165 -215
rect 4107 -1003 4119 -227
rect 4153 -1003 4165 -227
rect 4107 -1015 4165 -1003
rect 4285 -227 4343 -215
rect 4285 -1003 4297 -227
rect 4331 -1003 4343 -227
rect 4285 -1015 4343 -1003
rect 4513 -227 4571 -215
rect 4513 -1003 4525 -227
rect 4559 -1003 4571 -227
rect 4513 -1015 4571 -1003
rect 4691 -227 4749 -215
rect 4691 -1003 4703 -227
rect 4737 -1003 4749 -227
rect 4691 -1015 4749 -1003
rect 4919 -227 4977 -215
rect 4919 -1003 4931 -227
rect 4965 -1003 4977 -227
rect 4919 -1015 4977 -1003
rect 5097 -227 5155 -215
rect 5097 -1003 5109 -227
rect 5143 -1003 5155 -227
rect 5097 -1015 5155 -1003
rect 5325 -227 5383 -215
rect 5325 -1003 5337 -227
rect 5371 -1003 5383 -227
rect 5325 -1015 5383 -1003
rect 5503 -227 5561 -215
rect 5503 -1003 5515 -227
rect 5549 -1003 5561 -227
rect 5503 -1015 5561 -1003
rect 5731 -227 5789 -215
rect 5731 -1003 5743 -227
rect 5777 -1003 5789 -227
rect 5731 -1015 5789 -1003
rect 5909 -227 5967 -215
rect 5909 -1003 5921 -227
rect 5955 -1003 5967 -227
rect 5909 -1015 5967 -1003
rect 6137 -227 6195 -215
rect 6137 -1003 6149 -227
rect 6183 -1003 6195 -227
rect 6137 -1015 6195 -1003
rect 6315 -227 6373 -215
rect 6315 -1003 6327 -227
rect 6361 -1003 6373 -227
rect 6315 -1015 6373 -1003
<< pdiff >>
rect 1904 4234 1962 4246
rect 1904 458 1916 4234
rect 1950 458 1962 4234
rect 1904 446 1962 458
rect 2162 4234 2220 4246
rect 2162 458 2174 4234
rect 2208 458 2220 4234
rect 2162 446 2220 458
rect 2390 4234 2448 4246
rect 2390 458 2402 4234
rect 2436 458 2448 4234
rect 2390 446 2448 458
rect 2648 4234 2706 4246
rect 2648 458 2660 4234
rect 2694 458 2706 4234
rect 2648 446 2706 458
rect 2876 4234 2934 4246
rect 2876 458 2888 4234
rect 2922 458 2934 4234
rect 2876 446 2934 458
rect 3134 4234 3192 4246
rect 3134 458 3146 4234
rect 3180 458 3192 4234
rect 3134 446 3192 458
<< ndiffc >>
rect 1350 138 1410 172
rect 1350 50 1410 84
rect -2377 -1003 -2343 -227
rect -2199 -1003 -2165 -227
rect -1971 -1003 -1937 -227
rect -1793 -1003 -1759 -227
rect -1565 -1003 -1531 -227
rect -1387 -1003 -1353 -227
rect -1159 -1003 -1125 -227
rect -981 -1003 -947 -227
rect -753 -1003 -719 -227
rect -575 -1003 -541 -227
rect -347 -1003 -313 -227
rect -169 -1003 -135 -227
rect 59 -1003 93 -227
rect 237 -1003 271 -227
rect 465 -1003 499 -227
rect 643 -1003 677 -227
rect 871 -1003 905 -227
rect 1049 -1003 1083 -227
rect 1277 -1003 1311 -227
rect 1455 -1003 1489 -227
rect 1683 -1003 1717 -227
rect 1861 -1003 1895 -227
rect 2089 -1003 2123 -227
rect 2267 -1003 2301 -227
rect 2495 -1003 2529 -227
rect 2673 -1003 2707 -227
rect 2901 -1003 2935 -227
rect 3079 -1003 3113 -227
rect 3307 -1003 3341 -227
rect 3485 -1003 3519 -227
rect 3713 -1003 3747 -227
rect 3891 -1003 3925 -227
rect 4119 -1003 4153 -227
rect 4297 -1003 4331 -227
rect 4525 -1003 4559 -227
rect 4703 -1003 4737 -227
rect 4931 -1003 4965 -227
rect 5109 -1003 5143 -227
rect 5337 -1003 5371 -227
rect 5515 -1003 5549 -227
rect 5743 -1003 5777 -227
rect 5921 -1003 5955 -227
rect 6149 -1003 6183 -227
rect 6327 -1003 6361 -227
<< pdiffc >>
rect 1916 458 1950 4234
rect 2174 458 2208 4234
rect 2402 458 2436 4234
rect 2660 458 2694 4234
rect 2888 458 2922 4234
rect 3146 458 3180 4234
<< psubdiff >>
rect 1226 252 1322 286
rect 1500 252 1596 286
rect 1226 190 1260 252
rect 1562 190 1596 252
rect 1226 -30 1260 32
rect 1562 -30 1596 32
rect 1226 -41 1596 -30
rect -2491 -75 -2395 -41
rect -2147 -75 -1989 -41
rect -1741 -75 -1583 -41
rect -1335 -75 -1177 -41
rect -929 -75 -771 -41
rect -523 -75 -365 -41
rect -117 -75 41 -41
rect 289 -75 447 -41
rect 695 -75 853 -41
rect 1101 -75 1259 -41
rect 1507 -75 1665 -41
rect 1913 -75 2071 -41
rect 2319 -75 2477 -41
rect 2725 -75 2883 -41
rect 3131 -75 3289 -41
rect 3537 -75 3695 -41
rect 3943 -75 4101 -41
rect 4349 -75 4507 -41
rect 4755 -75 4913 -41
rect 5161 -75 5319 -41
rect 5567 -75 5725 -41
rect 5973 -75 6131 -41
rect 6379 -75 6475 -41
rect -2491 -137 -2457 -75
rect -2085 -137 -2051 -75
rect -2491 -1155 -2457 -1093
rect -1679 -137 -1645 -75
rect -2085 -1155 -2051 -1093
rect -1273 -137 -1239 -75
rect -1679 -1155 -1645 -1093
rect -867 -137 -833 -75
rect -1273 -1155 -1239 -1093
rect -461 -137 -427 -75
rect -867 -1155 -833 -1093
rect -55 -137 -21 -75
rect -461 -1155 -427 -1093
rect 351 -137 385 -75
rect -55 -1155 -21 -1093
rect 757 -137 791 -75
rect 351 -1155 385 -1093
rect 1163 -137 1197 -75
rect 757 -1155 791 -1093
rect 1569 -137 1603 -75
rect 1163 -1155 1197 -1093
rect 1975 -137 2009 -75
rect 1569 -1155 1603 -1093
rect 2381 -137 2415 -75
rect 1975 -1155 2009 -1093
rect 2787 -137 2821 -75
rect 2381 -1155 2415 -1093
rect 3193 -137 3227 -75
rect 2787 -1155 2821 -1093
rect 3599 -137 3633 -75
rect 3193 -1155 3227 -1093
rect 4005 -137 4039 -75
rect 3599 -1155 3633 -1093
rect 4411 -137 4445 -75
rect 4005 -1155 4039 -1093
rect 4817 -137 4851 -75
rect 4411 -1155 4445 -1093
rect 5223 -137 5257 -75
rect 4817 -1155 4851 -1093
rect 5629 -137 5663 -75
rect 5223 -1155 5257 -1093
rect 6035 -137 6069 -75
rect 5629 -1155 5663 -1093
rect 6441 -137 6475 -75
rect 6035 -1155 6069 -1093
rect 6441 -1155 6475 -1093
rect -2491 -1189 -2395 -1155
rect -2147 -1189 -1989 -1155
rect -1741 -1189 -1583 -1155
rect -1335 -1189 -1177 -1155
rect -929 -1189 -771 -1155
rect -523 -1189 -365 -1155
rect -117 -1189 41 -1155
rect 289 -1189 447 -1155
rect 695 -1189 853 -1155
rect 1101 -1189 1259 -1155
rect 1507 -1189 1665 -1155
rect 1913 -1189 2071 -1155
rect 2319 -1189 2477 -1155
rect 2725 -1189 2883 -1155
rect 3131 -1189 3289 -1155
rect 3537 -1189 3695 -1155
rect 3943 -1189 4101 -1155
rect 4349 -1189 4507 -1155
rect 4755 -1189 4913 -1155
rect 5161 -1189 5319 -1155
rect 5567 -1189 5725 -1155
rect 5973 -1189 6131 -1155
rect 6379 -1189 6475 -1155
rect -2494 -1318 -2398 -1284
rect 15690 -1318 15786 -1284
rect -2494 -1380 -2460 -1318
rect 15752 -1380 15786 -1318
rect -2494 -2656 -2460 -2594
rect 15752 -2656 15786 -2594
rect -2494 -2690 -2398 -2656
rect 15690 -2690 15786 -2656
rect -2494 -2752 -2460 -2690
rect 15752 -2752 15786 -2690
rect -2494 -4028 -2460 -3966
rect 15752 -4028 15786 -3966
rect -2494 -4062 -2398 -4028
rect 15690 -4062 15786 -4028
<< nsubdiff >>
rect 1802 4395 1898 4429
rect 2226 4395 2384 4429
rect 2712 4395 2870 4429
rect 3198 4395 3294 4429
rect 1802 4333 1836 4395
rect 2288 4333 2322 4395
rect 1802 297 1836 359
rect 2774 4333 2808 4395
rect 2288 297 2322 359
rect 3260 4333 3294 4395
rect 2774 297 2808 359
rect 3260 297 3294 359
rect 1802 263 1898 297
rect 2226 263 2384 297
rect 2712 263 2870 297
rect 3198 263 3294 297
<< psubdiffcont >>
rect 1322 252 1500 286
rect 1226 32 1260 190
rect 1562 32 1596 190
rect -2395 -75 -2147 -41
rect -1989 -75 -1741 -41
rect -1583 -75 -1335 -41
rect -1177 -75 -929 -41
rect -771 -75 -523 -41
rect -365 -75 -117 -41
rect 41 -75 289 -41
rect 447 -75 695 -41
rect 853 -75 1101 -41
rect 1259 -75 1507 -41
rect 1665 -75 1913 -41
rect 2071 -75 2319 -41
rect 2477 -75 2725 -41
rect 2883 -75 3131 -41
rect 3289 -75 3537 -41
rect 3695 -75 3943 -41
rect 4101 -75 4349 -41
rect 4507 -75 4755 -41
rect 4913 -75 5161 -41
rect 5319 -75 5567 -41
rect 5725 -75 5973 -41
rect 6131 -75 6379 -41
rect -2491 -1093 -2457 -137
rect -2085 -1093 -2051 -137
rect -1679 -1093 -1645 -137
rect -1273 -1093 -1239 -137
rect -867 -1093 -833 -137
rect -461 -1093 -427 -137
rect -55 -1093 -21 -137
rect 351 -1093 385 -137
rect 757 -1093 791 -137
rect 1163 -1093 1197 -137
rect 1569 -1093 1603 -137
rect 1975 -1093 2009 -137
rect 2381 -1093 2415 -137
rect 2787 -1093 2821 -137
rect 3193 -1093 3227 -137
rect 3599 -1093 3633 -137
rect 4005 -1093 4039 -137
rect 4411 -1093 4445 -137
rect 4817 -1093 4851 -137
rect 5223 -1093 5257 -137
rect 5629 -1093 5663 -137
rect 6035 -1093 6069 -137
rect 6441 -1093 6475 -137
rect -2395 -1189 -2147 -1155
rect -1989 -1189 -1741 -1155
rect -1583 -1189 -1335 -1155
rect -1177 -1189 -929 -1155
rect -771 -1189 -523 -1155
rect -365 -1189 -117 -1155
rect 41 -1189 289 -1155
rect 447 -1189 695 -1155
rect 853 -1189 1101 -1155
rect 1259 -1189 1507 -1155
rect 1665 -1189 1913 -1155
rect 2071 -1189 2319 -1155
rect 2477 -1189 2725 -1155
rect 2883 -1189 3131 -1155
rect 3289 -1189 3537 -1155
rect 3695 -1189 3943 -1155
rect 4101 -1189 4349 -1155
rect 4507 -1189 4755 -1155
rect 4913 -1189 5161 -1155
rect 5319 -1189 5567 -1155
rect 5725 -1189 5973 -1155
rect 6131 -1189 6379 -1155
rect -2398 -1318 15690 -1284
rect -2494 -2594 -2460 -1380
rect 15752 -2594 15786 -1380
rect -2398 -2690 15690 -2656
rect -2494 -3966 -2460 -2752
rect 15752 -3966 15786 -2752
rect -2398 -4062 15690 -4028
<< nsubdiffcont >>
rect 1898 4395 2226 4429
rect 2384 4395 2712 4429
rect 2870 4395 3198 4429
rect 1802 359 1836 4333
rect 2288 359 2322 4333
rect 2774 359 2808 4333
rect 3260 359 3294 4333
rect 1898 263 2226 297
rect 2384 263 2712 297
rect 2870 263 3198 297
<< poly >>
rect 1962 4327 2162 4343
rect 1962 4293 1978 4327
rect 2146 4293 2162 4327
rect 1962 4246 2162 4293
rect 1962 399 2162 446
rect 1962 365 1978 399
rect 2146 365 2162 399
rect 1962 349 2162 365
rect 2448 4327 2648 4343
rect 2448 4293 2464 4327
rect 2632 4293 2648 4327
rect 2448 4246 2648 4293
rect 2448 399 2648 446
rect 2448 365 2464 399
rect 2632 365 2648 399
rect 2448 349 2648 365
rect 2934 4327 3134 4343
rect 2934 4293 2950 4327
rect 3118 4293 3134 4327
rect 2934 4246 3134 4293
rect 2934 399 3134 446
rect 2934 365 2950 399
rect 3118 365 3134 399
rect 2934 349 3134 365
rect 1444 128 1510 144
rect 1444 126 1460 128
rect 1312 96 1338 126
rect 1422 96 1460 126
rect 1444 94 1460 96
rect 1494 94 1510 128
rect 1444 78 1510 94
rect -2331 -143 -2211 -127
rect -2331 -177 -2315 -143
rect -2227 -177 -2211 -143
rect -2331 -215 -2211 -177
rect -2331 -1053 -2211 -1015
rect -2331 -1087 -2315 -1053
rect -2227 -1087 -2211 -1053
rect -2331 -1103 -2211 -1087
rect -1925 -143 -1805 -127
rect -1925 -177 -1909 -143
rect -1821 -177 -1805 -143
rect -1925 -215 -1805 -177
rect -1925 -1053 -1805 -1015
rect -1925 -1087 -1909 -1053
rect -1821 -1087 -1805 -1053
rect -1925 -1103 -1805 -1087
rect -1519 -143 -1399 -127
rect -1519 -177 -1503 -143
rect -1415 -177 -1399 -143
rect -1519 -215 -1399 -177
rect -1519 -1053 -1399 -1015
rect -1519 -1087 -1503 -1053
rect -1415 -1087 -1399 -1053
rect -1519 -1103 -1399 -1087
rect -1113 -143 -993 -127
rect -1113 -177 -1097 -143
rect -1009 -177 -993 -143
rect -1113 -215 -993 -177
rect -1113 -1053 -993 -1015
rect -1113 -1087 -1097 -1053
rect -1009 -1087 -993 -1053
rect -1113 -1103 -993 -1087
rect -707 -143 -587 -127
rect -707 -177 -691 -143
rect -603 -177 -587 -143
rect -707 -215 -587 -177
rect -707 -1053 -587 -1015
rect -707 -1087 -691 -1053
rect -603 -1087 -587 -1053
rect -707 -1103 -587 -1087
rect -301 -143 -181 -127
rect -301 -177 -285 -143
rect -197 -177 -181 -143
rect -301 -215 -181 -177
rect -301 -1053 -181 -1015
rect -301 -1087 -285 -1053
rect -197 -1087 -181 -1053
rect -301 -1103 -181 -1087
rect 105 -143 225 -127
rect 105 -177 121 -143
rect 209 -177 225 -143
rect 105 -215 225 -177
rect 105 -1053 225 -1015
rect 105 -1087 121 -1053
rect 209 -1087 225 -1053
rect 105 -1103 225 -1087
rect 511 -143 631 -127
rect 511 -177 527 -143
rect 615 -177 631 -143
rect 511 -215 631 -177
rect 511 -1053 631 -1015
rect 511 -1087 527 -1053
rect 615 -1087 631 -1053
rect 511 -1103 631 -1087
rect 917 -143 1037 -127
rect 917 -177 933 -143
rect 1021 -177 1037 -143
rect 917 -215 1037 -177
rect 917 -1053 1037 -1015
rect 917 -1087 933 -1053
rect 1021 -1087 1037 -1053
rect 917 -1103 1037 -1087
rect 1323 -143 1443 -127
rect 1323 -177 1339 -143
rect 1427 -177 1443 -143
rect 1323 -215 1443 -177
rect 1323 -1053 1443 -1015
rect 1323 -1087 1339 -1053
rect 1427 -1087 1443 -1053
rect 1323 -1103 1443 -1087
rect 1729 -143 1849 -127
rect 1729 -177 1745 -143
rect 1833 -177 1849 -143
rect 1729 -215 1849 -177
rect 1729 -1053 1849 -1015
rect 1729 -1087 1745 -1053
rect 1833 -1087 1849 -1053
rect 1729 -1103 1849 -1087
rect 2135 -143 2255 -127
rect 2135 -177 2151 -143
rect 2239 -177 2255 -143
rect 2135 -215 2255 -177
rect 2135 -1053 2255 -1015
rect 2135 -1087 2151 -1053
rect 2239 -1087 2255 -1053
rect 2135 -1103 2255 -1087
rect 2541 -143 2661 -127
rect 2541 -177 2557 -143
rect 2645 -177 2661 -143
rect 2541 -215 2661 -177
rect 2541 -1053 2661 -1015
rect 2541 -1087 2557 -1053
rect 2645 -1087 2661 -1053
rect 2541 -1103 2661 -1087
rect 2947 -143 3067 -127
rect 2947 -177 2963 -143
rect 3051 -177 3067 -143
rect 2947 -215 3067 -177
rect 2947 -1053 3067 -1015
rect 2947 -1087 2963 -1053
rect 3051 -1087 3067 -1053
rect 2947 -1103 3067 -1087
rect 3353 -143 3473 -127
rect 3353 -177 3369 -143
rect 3457 -177 3473 -143
rect 3353 -215 3473 -177
rect 3353 -1053 3473 -1015
rect 3353 -1087 3369 -1053
rect 3457 -1087 3473 -1053
rect 3353 -1103 3473 -1087
rect 3759 -143 3879 -127
rect 3759 -177 3775 -143
rect 3863 -177 3879 -143
rect 3759 -215 3879 -177
rect 3759 -1053 3879 -1015
rect 3759 -1087 3775 -1053
rect 3863 -1087 3879 -1053
rect 3759 -1103 3879 -1087
rect 4165 -143 4285 -127
rect 4165 -177 4181 -143
rect 4269 -177 4285 -143
rect 4165 -215 4285 -177
rect 4165 -1053 4285 -1015
rect 4165 -1087 4181 -1053
rect 4269 -1087 4285 -1053
rect 4165 -1103 4285 -1087
rect 4571 -143 4691 -127
rect 4571 -177 4587 -143
rect 4675 -177 4691 -143
rect 4571 -215 4691 -177
rect 4571 -1053 4691 -1015
rect 4571 -1087 4587 -1053
rect 4675 -1087 4691 -1053
rect 4571 -1103 4691 -1087
rect 4977 -143 5097 -127
rect 4977 -177 4993 -143
rect 5081 -177 5097 -143
rect 4977 -215 5097 -177
rect 4977 -1053 5097 -1015
rect 4977 -1087 4993 -1053
rect 5081 -1087 5097 -1053
rect 4977 -1103 5097 -1087
rect 5383 -143 5503 -127
rect 5383 -177 5399 -143
rect 5487 -177 5503 -143
rect 5383 -215 5503 -177
rect 5383 -1053 5503 -1015
rect 5383 -1087 5399 -1053
rect 5487 -1087 5503 -1053
rect 5383 -1103 5503 -1087
rect 5789 -143 5909 -127
rect 5789 -177 5805 -143
rect 5893 -177 5909 -143
rect 5789 -215 5909 -177
rect 5789 -1053 5909 -1015
rect 5789 -1087 5805 -1053
rect 5893 -1087 5909 -1053
rect 5789 -1103 5909 -1087
rect 6195 -143 6315 -127
rect 6195 -177 6211 -143
rect 6299 -177 6315 -143
rect 6195 -215 6315 -177
rect 6195 -1053 6315 -1015
rect 6195 -1087 6211 -1053
rect 6299 -1087 6315 -1053
rect 6195 -1103 6315 -1087
<< polycont >>
rect 1978 4293 2146 4327
rect 1978 365 2146 399
rect 2464 4293 2632 4327
rect 2464 365 2632 399
rect 2950 4293 3118 4327
rect 2950 365 3118 399
rect 1460 94 1494 128
rect -2315 -177 -2227 -143
rect -2315 -1087 -2227 -1053
rect -1909 -177 -1821 -143
rect -1909 -1087 -1821 -1053
rect -1503 -177 -1415 -143
rect -1503 -1087 -1415 -1053
rect -1097 -177 -1009 -143
rect -1097 -1087 -1009 -1053
rect -691 -177 -603 -143
rect -691 -1087 -603 -1053
rect -285 -177 -197 -143
rect -285 -1087 -197 -1053
rect 121 -177 209 -143
rect 121 -1087 209 -1053
rect 527 -177 615 -143
rect 527 -1087 615 -1053
rect 933 -177 1021 -143
rect 933 -1087 1021 -1053
rect 1339 -177 1427 -143
rect 1339 -1087 1427 -1053
rect 1745 -177 1833 -143
rect 1745 -1087 1833 -1053
rect 2151 -177 2239 -143
rect 2151 -1087 2239 -1053
rect 2557 -177 2645 -143
rect 2557 -1087 2645 -1053
rect 2963 -177 3051 -143
rect 2963 -1087 3051 -1053
rect 3369 -177 3457 -143
rect 3369 -1087 3457 -1053
rect 3775 -177 3863 -143
rect 3775 -1087 3863 -1053
rect 4181 -177 4269 -143
rect 4181 -1087 4269 -1053
rect 4587 -177 4675 -143
rect 4587 -1087 4675 -1053
rect 4993 -177 5081 -143
rect 4993 -1087 5081 -1053
rect 5399 -177 5487 -143
rect 5399 -1087 5487 -1053
rect 5805 -177 5893 -143
rect 5805 -1087 5893 -1053
rect 6211 -177 6299 -143
rect 6211 -1087 6299 -1053
<< xpolycontact >>
rect -2364 -2560 -1932 -1414
rect 15224 -2560 15656 -1414
rect -2364 -3932 -1932 -2786
rect 15224 -3932 15656 -2786
<< xpolyres >>
rect -1932 -2560 15224 -1414
rect -1932 -3932 15224 -2786
<< locali >>
rect 1802 4395 1898 4429
rect 2226 4395 2384 4429
rect 2712 4395 2870 4429
rect 3198 4395 3294 4429
rect 1802 4333 1836 4395
rect 2288 4333 2322 4395
rect 1962 4293 1978 4327
rect 2146 4293 2162 4327
rect 1916 4234 1950 4250
rect 1916 442 1950 458
rect 2174 4234 2208 4250
rect 2774 4333 2808 4395
rect 2448 4293 2464 4327
rect 2632 4293 2648 4327
rect 2402 4234 2436 4250
rect 2174 442 2208 458
rect 1962 365 1978 399
rect 2146 365 2162 399
rect 1802 297 1836 359
rect 2402 442 2436 458
rect 2660 4234 2694 4250
rect 2660 442 2694 458
rect 3260 4333 3294 4395
rect 2934 4293 2950 4327
rect 3118 4293 3134 4327
rect 2888 4234 2922 4250
rect 2448 365 2464 399
rect 2632 365 2648 399
rect 2288 297 2322 359
rect 2888 442 2922 458
rect 3146 4234 3180 4250
rect 3146 442 3180 458
rect 2934 365 2950 399
rect 3118 365 3134 399
rect 2774 297 2808 359
rect 3260 297 3294 359
rect 1226 252 1322 286
rect 1500 252 1596 286
rect 1802 263 1898 297
rect 2226 263 2384 297
rect 2712 263 2870 297
rect 3198 263 3294 297
rect 1226 190 1260 252
rect 1562 190 1596 252
rect 1334 138 1350 172
rect 1410 138 1426 172
rect 1460 128 1494 144
rect 1334 50 1350 84
rect 1410 50 1426 84
rect 1460 78 1494 94
rect 1226 -20 1260 32
rect 1562 -20 1596 32
rect -2491 -80 -2490 -41
rect -2491 -137 -2457 -80
rect -2085 -137 -2051 -80
rect -2331 -177 -2315 -143
rect -2227 -177 -2211 -143
rect -2377 -227 -2343 -211
rect -2377 -1019 -2343 -1003
rect -2199 -227 -2165 -211
rect -2199 -1019 -2165 -1003
rect -2331 -1087 -2315 -1053
rect -2227 -1087 -2211 -1053
rect -2491 -1152 -2457 -1093
rect -1679 -137 -1645 -80
rect -1925 -177 -1909 -143
rect -1821 -177 -1805 -143
rect -1971 -227 -1937 -211
rect -1971 -1019 -1937 -1003
rect -1793 -227 -1759 -211
rect -1793 -1019 -1759 -1003
rect -1925 -1087 -1909 -1053
rect -1821 -1087 -1805 -1053
rect -2085 -1152 -2051 -1093
rect -1273 -137 -1239 -80
rect -1519 -177 -1503 -143
rect -1415 -177 -1399 -143
rect -1565 -227 -1531 -211
rect -1565 -1019 -1531 -1003
rect -1387 -227 -1353 -211
rect -1387 -1019 -1353 -1003
rect -1519 -1087 -1503 -1053
rect -1415 -1087 -1399 -1053
rect -1679 -1152 -1645 -1093
rect -867 -137 -833 -80
rect -1113 -177 -1097 -143
rect -1009 -177 -993 -143
rect -1159 -227 -1125 -211
rect -1159 -1019 -1125 -1003
rect -981 -227 -947 -211
rect -981 -1019 -947 -1003
rect -1113 -1087 -1097 -1053
rect -1009 -1087 -993 -1053
rect -1273 -1152 -1239 -1093
rect -461 -137 -427 -80
rect -707 -177 -691 -143
rect -603 -177 -587 -143
rect -753 -227 -719 -211
rect -753 -1019 -719 -1003
rect -575 -227 -541 -211
rect -575 -1019 -541 -1003
rect -707 -1087 -691 -1053
rect -603 -1087 -587 -1053
rect -867 -1152 -833 -1093
rect -55 -137 -21 -80
rect -301 -177 -285 -143
rect -197 -177 -181 -143
rect -347 -227 -313 -211
rect -347 -1019 -313 -1003
rect -169 -227 -135 -211
rect -169 -1019 -135 -1003
rect -301 -1087 -285 -1053
rect -197 -1087 -181 -1053
rect -461 -1152 -427 -1093
rect 351 -137 385 -80
rect 105 -177 121 -143
rect 209 -177 225 -143
rect 59 -227 93 -211
rect 59 -1019 93 -1003
rect 237 -227 271 -211
rect 237 -1019 271 -1003
rect 105 -1087 121 -1053
rect 209 -1087 225 -1053
rect -55 -1152 -21 -1093
rect 757 -137 791 -80
rect 511 -177 527 -143
rect 615 -177 631 -143
rect 465 -227 499 -211
rect 465 -1019 499 -1003
rect 643 -227 677 -211
rect 643 -1019 677 -1003
rect 511 -1087 527 -1053
rect 615 -1087 631 -1053
rect 351 -1152 385 -1093
rect 1163 -137 1197 -80
rect 917 -177 933 -143
rect 1021 -177 1037 -143
rect 871 -227 905 -211
rect 871 -1019 905 -1003
rect 1049 -227 1083 -211
rect 1049 -1019 1083 -1003
rect 917 -1087 933 -1053
rect 1021 -1087 1037 -1053
rect 757 -1152 791 -1093
rect 1569 -137 1603 -80
rect 1323 -177 1339 -143
rect 1427 -177 1443 -143
rect 1277 -227 1311 -211
rect 1277 -1019 1311 -1003
rect 1455 -227 1489 -211
rect 1455 -1019 1489 -1003
rect 1323 -1087 1339 -1053
rect 1427 -1087 1443 -1053
rect 1163 -1152 1197 -1093
rect 1975 -137 2009 -80
rect 1729 -177 1745 -143
rect 1833 -177 1849 -143
rect 1683 -227 1717 -211
rect 1683 -1019 1717 -1003
rect 1861 -227 1895 -211
rect 1861 -1019 1895 -1003
rect 1729 -1087 1745 -1053
rect 1833 -1087 1849 -1053
rect 1569 -1152 1603 -1093
rect 2381 -137 2415 -80
rect 2135 -177 2151 -143
rect 2239 -177 2255 -143
rect 2089 -227 2123 -211
rect 2089 -1019 2123 -1003
rect 2267 -227 2301 -211
rect 2267 -1019 2301 -1003
rect 2135 -1087 2151 -1053
rect 2239 -1087 2255 -1053
rect 1975 -1152 2009 -1093
rect 2787 -137 2821 -80
rect 2541 -177 2557 -143
rect 2645 -177 2661 -143
rect 2495 -227 2529 -211
rect 2495 -1019 2529 -1003
rect 2673 -227 2707 -211
rect 2673 -1019 2707 -1003
rect 2541 -1087 2557 -1053
rect 2645 -1087 2661 -1053
rect 2381 -1152 2415 -1093
rect 3193 -137 3227 -80
rect 2947 -177 2963 -143
rect 3051 -177 3067 -143
rect 2901 -227 2935 -211
rect 2901 -1019 2935 -1003
rect 3079 -227 3113 -211
rect 3079 -1019 3113 -1003
rect 2947 -1087 2963 -1053
rect 3051 -1087 3067 -1053
rect 2787 -1152 2821 -1093
rect 3599 -137 3633 -80
rect 3353 -177 3369 -143
rect 3457 -177 3473 -143
rect 3307 -227 3341 -211
rect 3307 -1019 3341 -1003
rect 3485 -227 3519 -211
rect 3485 -1019 3519 -1003
rect 3353 -1087 3369 -1053
rect 3457 -1087 3473 -1053
rect 3193 -1152 3227 -1093
rect 4005 -137 4039 -80
rect 3759 -177 3775 -143
rect 3863 -177 3879 -143
rect 3713 -227 3747 -211
rect 3713 -1019 3747 -1003
rect 3891 -227 3925 -211
rect 3891 -1019 3925 -1003
rect 3759 -1087 3775 -1053
rect 3863 -1087 3879 -1053
rect 3599 -1152 3633 -1093
rect 4411 -137 4445 -80
rect 4165 -177 4181 -143
rect 4269 -177 4285 -143
rect 4119 -227 4153 -211
rect 4119 -1019 4153 -1003
rect 4297 -227 4331 -211
rect 4297 -1019 4331 -1003
rect 4165 -1087 4181 -1053
rect 4269 -1087 4285 -1053
rect 4005 -1152 4039 -1093
rect 4817 -137 4851 -80
rect 4571 -177 4587 -143
rect 4675 -177 4691 -143
rect 4525 -227 4559 -211
rect 4525 -1019 4559 -1003
rect 4703 -227 4737 -211
rect 4703 -1019 4737 -1003
rect 4571 -1087 4587 -1053
rect 4675 -1087 4691 -1053
rect 4411 -1152 4445 -1093
rect 5223 -137 5257 -80
rect 4977 -177 4993 -143
rect 5081 -177 5097 -143
rect 4931 -227 4965 -211
rect 4931 -1019 4965 -1003
rect 5109 -227 5143 -211
rect 5109 -1019 5143 -1003
rect 4977 -1087 4993 -1053
rect 5081 -1087 5097 -1053
rect 4817 -1152 4851 -1093
rect 5629 -137 5663 -80
rect 5383 -177 5399 -143
rect 5487 -177 5503 -143
rect 5337 -227 5371 -211
rect 5337 -1019 5371 -1003
rect 5515 -227 5549 -211
rect 5515 -1019 5549 -1003
rect 5383 -1087 5399 -1053
rect 5487 -1087 5503 -1053
rect 5223 -1152 5257 -1093
rect 6035 -137 6069 -80
rect 5789 -177 5805 -143
rect 5893 -177 5909 -143
rect 5743 -227 5777 -211
rect 5743 -1019 5777 -1003
rect 5921 -227 5955 -211
rect 5921 -1019 5955 -1003
rect 5789 -1087 5805 -1053
rect 5893 -1087 5909 -1053
rect 5629 -1152 5663 -1093
rect 6195 -177 6211 -143
rect 6299 -177 6315 -143
rect 6149 -227 6183 -211
rect 6149 -1019 6183 -1003
rect 6327 -227 6361 -211
rect 6327 -1019 6361 -1003
rect 6430 -1047 6432 -174
rect 6195 -1087 6211 -1053
rect 6299 -1087 6315 -1053
rect 6035 -1152 6069 -1093
rect 6430 -1117 6431 -1047
rect -2491 -1189 -2482 -1152
<< viali >>
rect 1978 4293 2146 4327
rect 1916 458 1950 4234
rect 2174 458 2208 4234
rect 2464 4293 2632 4327
rect 2276 483 2288 4213
rect 2288 483 2322 4213
rect 2322 483 2326 4213
rect 1978 365 2146 399
rect 2402 458 2436 4234
rect 2660 458 2694 4234
rect 2950 4293 3118 4327
rect 2776 473 2808 4213
rect 2808 473 2826 4213
rect 2464 365 2632 399
rect 2888 458 2922 4234
rect 3146 458 3180 4234
rect 2950 365 3118 399
rect 1350 138 1410 172
rect 1460 94 1494 128
rect 1350 50 1410 84
rect -2490 -41 6480 -20
rect -2490 -75 -2395 -41
rect -2395 -75 -2147 -41
rect -2147 -75 -1989 -41
rect -1989 -75 -1741 -41
rect -1741 -75 -1583 -41
rect -1583 -75 -1335 -41
rect -1335 -75 -1177 -41
rect -1177 -75 -929 -41
rect -929 -75 -771 -41
rect -771 -75 -523 -41
rect -523 -75 -365 -41
rect -365 -75 -117 -41
rect -117 -75 41 -41
rect 41 -75 289 -41
rect 289 -75 447 -41
rect 447 -75 695 -41
rect 695 -75 853 -41
rect 853 -75 1101 -41
rect 1101 -75 1259 -41
rect 1259 -75 1507 -41
rect 1507 -75 1665 -41
rect 1665 -75 1913 -41
rect 1913 -75 2071 -41
rect 2071 -75 2319 -41
rect 2319 -75 2477 -41
rect 2477 -75 2725 -41
rect 2725 -75 2883 -41
rect 2883 -75 3131 -41
rect 3131 -75 3289 -41
rect 3289 -75 3537 -41
rect 3537 -75 3695 -41
rect 3695 -75 3943 -41
rect 3943 -75 4101 -41
rect 4101 -75 4349 -41
rect 4349 -75 4507 -41
rect 4507 -75 4755 -41
rect 4755 -75 4913 -41
rect 4913 -75 5161 -41
rect 5161 -75 5319 -41
rect 5319 -75 5567 -41
rect 5567 -75 5725 -41
rect 5725 -75 5973 -41
rect 5973 -75 6131 -41
rect 6131 -75 6379 -41
rect 6379 -75 6480 -41
rect -2490 -80 6480 -75
rect -2315 -177 -2227 -143
rect -2377 -1003 -2343 -227
rect -2199 -1003 -2165 -227
rect -2315 -1087 -2227 -1053
rect -1909 -177 -1821 -143
rect -1971 -1003 -1937 -227
rect -1793 -1003 -1759 -227
rect -1909 -1087 -1821 -1053
rect -1503 -177 -1415 -143
rect -1565 -1003 -1531 -227
rect -1387 -1003 -1353 -227
rect -1503 -1087 -1415 -1053
rect -1097 -177 -1009 -143
rect -1159 -1003 -1125 -227
rect -981 -1003 -947 -227
rect -1097 -1087 -1009 -1053
rect -691 -177 -603 -143
rect -753 -1003 -719 -227
rect -575 -1003 -541 -227
rect -691 -1087 -603 -1053
rect -285 -177 -197 -143
rect -347 -1003 -313 -227
rect -169 -1003 -135 -227
rect -285 -1087 -197 -1053
rect 121 -177 209 -143
rect 59 -1003 93 -227
rect 237 -1003 271 -227
rect 121 -1087 209 -1053
rect 527 -177 615 -143
rect 465 -1003 499 -227
rect 643 -1003 677 -227
rect 527 -1087 615 -1053
rect 933 -177 1021 -143
rect 871 -1003 905 -227
rect 1049 -1003 1083 -227
rect 933 -1087 1021 -1053
rect 1339 -177 1427 -143
rect 1277 -1003 1311 -227
rect 1455 -1003 1489 -227
rect 1339 -1087 1427 -1053
rect 1745 -177 1833 -143
rect 1683 -1003 1717 -227
rect 1861 -1003 1895 -227
rect 1745 -1087 1833 -1053
rect 2151 -177 2239 -143
rect 2089 -1003 2123 -227
rect 2267 -1003 2301 -227
rect 2151 -1087 2239 -1053
rect 2557 -177 2645 -143
rect 2495 -1003 2529 -227
rect 2673 -1003 2707 -227
rect 2557 -1087 2645 -1053
rect 2963 -177 3051 -143
rect 2901 -1003 2935 -227
rect 3079 -1003 3113 -227
rect 2963 -1087 3051 -1053
rect 3369 -177 3457 -143
rect 3307 -1003 3341 -227
rect 3485 -1003 3519 -227
rect 3369 -1087 3457 -1053
rect 3775 -177 3863 -143
rect 3713 -1003 3747 -227
rect 3891 -1003 3925 -227
rect 3775 -1087 3863 -1053
rect 4181 -177 4269 -143
rect 4119 -1003 4153 -227
rect 4297 -1003 4331 -227
rect 4181 -1087 4269 -1053
rect 4587 -177 4675 -143
rect 4525 -1003 4559 -227
rect 4703 -1003 4737 -227
rect 4587 -1087 4675 -1053
rect 4993 -177 5081 -143
rect 4931 -1003 4965 -227
rect 5109 -1003 5143 -227
rect 4993 -1087 5081 -1053
rect 5399 -177 5487 -143
rect 5337 -1003 5371 -227
rect 5515 -1003 5549 -227
rect 5399 -1087 5487 -1053
rect 5805 -177 5893 -143
rect 5743 -1003 5777 -227
rect 5921 -1003 5955 -227
rect 5805 -1087 5893 -1053
rect 6430 -137 6480 -80
rect 6211 -177 6299 -143
rect 6430 -174 6441 -137
rect 6149 -1003 6183 -227
rect 6327 -1003 6361 -227
rect 6432 -1047 6441 -174
rect 6211 -1087 6299 -1053
rect 6431 -1093 6441 -1047
rect 6441 -1093 6475 -137
rect 6475 -1093 6480 -137
rect 6431 -1117 6480 -1093
rect 6430 -1152 6480 -1117
rect -2482 -1155 6480 -1152
rect -2482 -1189 -2395 -1155
rect -2395 -1189 -2147 -1155
rect -2147 -1189 -1989 -1155
rect -1989 -1189 -1741 -1155
rect -1741 -1189 -1583 -1155
rect -1583 -1189 -1335 -1155
rect -1335 -1189 -1177 -1155
rect -1177 -1189 -929 -1155
rect -929 -1189 -771 -1155
rect -771 -1189 -523 -1155
rect -523 -1189 -365 -1155
rect -365 -1189 -117 -1155
rect -117 -1189 41 -1155
rect 41 -1189 289 -1155
rect 289 -1189 447 -1155
rect 447 -1189 695 -1155
rect 695 -1189 853 -1155
rect 853 -1189 1101 -1155
rect 1101 -1189 1259 -1155
rect 1259 -1189 1507 -1155
rect 1507 -1189 1665 -1155
rect 1665 -1189 1913 -1155
rect 1913 -1189 2071 -1155
rect 2071 -1189 2319 -1155
rect 2319 -1189 2477 -1155
rect 2477 -1189 2725 -1155
rect 2725 -1189 2883 -1155
rect 2883 -1189 3131 -1155
rect 3131 -1189 3289 -1155
rect 3289 -1189 3537 -1155
rect 3537 -1189 3695 -1155
rect 3695 -1189 3943 -1155
rect 3943 -1189 4101 -1155
rect 4101 -1189 4349 -1155
rect 4349 -1189 4507 -1155
rect 4507 -1189 4755 -1155
rect 4755 -1189 4913 -1155
rect 4913 -1189 5161 -1155
rect 5161 -1189 5319 -1155
rect 5319 -1189 5567 -1155
rect 5567 -1189 5725 -1155
rect 5725 -1189 5973 -1155
rect 5973 -1189 6131 -1155
rect 6131 -1189 6379 -1155
rect 6379 -1189 6480 -1155
rect -2482 -1200 6480 -1189
rect -2482 -1212 6470 -1200
rect -2510 -1284 15790 -1260
rect -2510 -1318 -2398 -1284
rect -2398 -1318 15690 -1284
rect 15690 -1318 15790 -1284
rect -2510 -1320 15790 -1318
rect -2510 -1380 -2440 -1320
rect -2510 -2594 -2494 -1380
rect -2494 -2594 -2460 -1380
rect -2460 -2594 -2440 -1380
rect 15700 -1380 15790 -1320
rect -2346 -2544 -1949 -1430
rect 15241 -2544 15638 -1430
rect -2510 -2640 -2440 -2594
rect 15700 -2594 15752 -1380
rect 15752 -2594 15786 -1380
rect 15786 -2594 15790 -1380
rect 15700 -2640 15790 -2594
rect -2510 -2656 15794 -2640
rect -2510 -2690 -2398 -2656
rect -2398 -2690 15690 -2656
rect 15690 -2690 15794 -2656
rect -2510 -2700 15794 -2690
rect -2510 -2752 -2440 -2700
rect -2510 -3966 -2494 -2752
rect -2494 -3966 -2460 -2752
rect -2460 -3966 -2440 -2752
rect 15700 -2752 15790 -2700
rect -2346 -3916 -1949 -2802
rect 15241 -3916 15638 -2802
rect -2510 -3990 -2440 -3966
rect 15700 -3966 15752 -2752
rect 15752 -3966 15786 -2752
rect 15786 -3966 15790 -2752
rect 15700 -3990 15790 -3966
rect -2510 -4028 15800 -3990
rect -2510 -4062 -2398 -4028
rect -2398 -4062 15690 -4028
rect 15690 -4062 15800 -4028
rect -2510 -4080 15800 -4062
<< metal1 >>
rect 2416 4620 2736 4693
rect 2416 4493 2460 4620
rect 2450 4490 2460 4493
rect 2690 4493 2736 4620
rect 2690 4490 2700 4493
rect 1956 4327 3146 4373
rect 1956 4293 1978 4327
rect 2146 4293 2464 4327
rect 2632 4293 2950 4327
rect 3118 4293 3146 4327
rect 1966 4287 2158 4293
rect 2452 4287 2716 4293
rect 2938 4287 3130 4293
rect 1910 4243 1956 4246
rect 2168 4243 2214 4246
rect 2396 4243 2442 4246
rect 1866 4234 1956 4243
rect 1866 4227 1916 4234
rect 1950 4227 1956 4234
rect 2166 4234 2446 4243
rect 1864 473 1874 4227
rect 1950 473 1958 4227
rect 1866 458 1916 473
rect 1950 458 1956 473
rect 1866 443 1956 458
rect 2166 458 2174 4234
rect 2208 4213 2402 4234
rect 2208 4133 2276 4213
rect 2326 4133 2402 4213
rect 2208 623 2256 4133
rect 2346 623 2402 4133
rect 2208 483 2276 623
rect 2326 483 2402 623
rect 2208 458 2402 483
rect 2436 458 2446 4234
rect 2166 453 2446 458
rect 2626 4234 2716 4287
rect 2882 4243 2928 4246
rect 2626 458 2660 4234
rect 2694 458 2716 4234
rect 2776 4234 2928 4243
rect 2776 4225 2888 4234
rect 2770 4213 2888 4225
rect 2770 473 2776 4213
rect 2826 4133 2888 4213
rect 2886 623 2888 4133
rect 2826 473 2888 623
rect 2770 461 2888 473
rect 2168 446 2214 453
rect 2396 446 2442 453
rect 2626 405 2716 458
rect 2776 458 2888 461
rect 2922 458 2928 4234
rect 3140 4234 3186 4246
rect 3140 4230 3146 4234
rect 3180 4230 3186 4234
rect 3130 470 3140 4230
rect 3210 470 3220 4230
rect 5800 670 6610 720
rect 5790 470 5800 670
rect 6260 470 6610 670
rect 2776 446 2928 458
rect 3140 458 3146 470
rect 3180 458 3186 470
rect 5800 460 6610 470
rect 3140 446 3186 458
rect 2776 443 2926 446
rect 1966 403 2158 405
rect 2452 403 2716 405
rect 2938 403 3130 405
rect 1956 400 3146 403
rect 1450 399 2140 400
rect 2980 399 3146 400
rect 1450 365 1978 399
rect 3118 365 3146 399
rect 1450 330 2140 365
rect 2980 330 3146 365
rect 1450 323 3146 330
rect 1450 320 2050 323
rect 1450 180 1510 320
rect 1350 178 1510 180
rect 1338 172 1510 178
rect 1338 138 1350 172
rect 1410 140 1510 172
rect 1410 138 1422 140
rect 1338 132 1422 138
rect 1450 128 1510 140
rect 1450 94 1460 128
rect 1494 94 1510 128
rect 1338 84 1422 90
rect 1338 80 1350 84
rect 1320 20 1330 80
rect 1410 44 1422 84
rect 1450 80 1510 94
rect 1410 20 1420 44
rect 6424 -14 6486 -8
rect -2502 -20 6492 -14
rect -2502 -80 -2490 -20
rect -2502 -86 6430 -80
rect -2450 -130 6100 -120
rect -2520 -143 6100 -130
rect -2520 -177 -2315 -143
rect -2227 -177 -1909 -143
rect -1821 -177 -1503 -143
rect -1415 -177 -1097 -143
rect -1009 -177 -691 -143
rect -603 -177 -285 -143
rect -197 -177 121 -143
rect 209 -177 527 -143
rect 615 -177 933 -143
rect 1021 -177 1339 -143
rect 1427 -177 1745 -143
rect 1833 -177 2151 -143
rect 2239 -177 2557 -143
rect 2645 -177 2963 -143
rect 3051 -177 3369 -143
rect 3457 -177 3775 -143
rect 3863 -177 4181 -143
rect 4269 -177 4587 -143
rect 4675 -177 4993 -143
rect 5081 -177 5399 -143
rect 5487 -177 5805 -143
rect 5893 -177 6100 -143
rect -2520 -180 6100 -177
rect -2520 -1050 -2450 -180
rect -2327 -183 -2215 -180
rect -1921 -183 -1809 -180
rect -1515 -183 -1403 -180
rect -1109 -183 -997 -180
rect -703 -183 -591 -180
rect -297 -183 -185 -180
rect 109 -183 221 -180
rect 515 -183 627 -180
rect 921 -183 1033 -180
rect 1327 -183 1439 -180
rect 1733 -183 1845 -180
rect 1880 -210 1950 -180
rect 2139 -183 2251 -180
rect 2545 -183 2657 -180
rect 2951 -183 3063 -180
rect 3357 -183 3469 -180
rect 3763 -183 3875 -180
rect 4169 -183 4281 -180
rect 4575 -183 4687 -180
rect 4981 -183 5093 -180
rect 5387 -183 5499 -180
rect 5793 -183 5905 -180
rect 1860 -215 1950 -210
rect -2383 -227 -2337 -215
rect -2205 -227 -2159 -215
rect -1977 -227 -1931 -215
rect -1799 -227 -1753 -215
rect -1571 -227 -1525 -215
rect -1393 -227 -1347 -215
rect -1165 -227 -1119 -215
rect -987 -227 -941 -215
rect -759 -227 -713 -215
rect -581 -227 -535 -215
rect -353 -227 -307 -215
rect -175 -227 -129 -215
rect 53 -227 99 -215
rect 231 -227 277 -215
rect 459 -227 505 -215
rect 637 -227 683 -215
rect 865 -227 911 -215
rect 1043 -227 1089 -215
rect 1271 -227 1317 -215
rect 1449 -227 1495 -215
rect 1677 -227 1723 -215
rect 1855 -227 1950 -215
rect 2083 -227 2129 -215
rect 2261 -227 2307 -215
rect 2489 -227 2535 -215
rect 2667 -227 2713 -215
rect 2895 -227 2941 -215
rect 3073 -227 3119 -215
rect 3301 -227 3347 -215
rect 3479 -227 3525 -215
rect 3707 -227 3753 -215
rect 3885 -227 3931 -215
rect 4113 -227 4159 -215
rect 4291 -227 4337 -215
rect 4519 -227 4565 -215
rect 4697 -227 4743 -215
rect 4925 -227 4971 -215
rect 5103 -227 5149 -215
rect 5331 -227 5377 -215
rect 5509 -227 5555 -215
rect 5737 -227 5783 -215
rect 5915 -227 5961 -215
rect -2413 -1004 -2403 -227
rect -2343 -1003 -2334 -227
rect -2205 -228 -2199 -227
rect -2165 -228 -2159 -227
rect -2344 -1004 -2334 -1003
rect -2383 -1015 -2337 -1004
rect -2210 -1005 -2200 -228
rect -2141 -1005 -2131 -228
rect -2007 -1004 -1997 -227
rect -1937 -1003 -1928 -227
rect -1799 -228 -1793 -227
rect -1759 -228 -1753 -227
rect -1938 -1004 -1928 -1003
rect -2205 -1015 -2159 -1005
rect -1977 -1015 -1931 -1004
rect -1804 -1005 -1794 -228
rect -1735 -1005 -1725 -228
rect -1601 -1004 -1591 -227
rect -1531 -1003 -1522 -227
rect -1393 -228 -1387 -227
rect -1353 -228 -1347 -227
rect -1532 -1004 -1522 -1003
rect -1799 -1015 -1753 -1005
rect -1571 -1015 -1525 -1004
rect -1398 -1005 -1388 -228
rect -1329 -1005 -1319 -228
rect -1195 -1004 -1185 -227
rect -1125 -1003 -1116 -227
rect -987 -228 -981 -227
rect -947 -228 -941 -227
rect -1126 -1004 -1116 -1003
rect -1393 -1015 -1347 -1005
rect -1165 -1015 -1119 -1004
rect -992 -1005 -982 -228
rect -923 -1005 -913 -228
rect -789 -1004 -779 -227
rect -719 -1003 -710 -227
rect -581 -228 -575 -227
rect -541 -228 -535 -227
rect -720 -1004 -710 -1003
rect -987 -1015 -941 -1005
rect -759 -1015 -713 -1004
rect -586 -1005 -576 -228
rect -517 -1005 -507 -228
rect -383 -1004 -373 -227
rect -313 -1003 -304 -227
rect -175 -228 -169 -227
rect -135 -228 -129 -227
rect -314 -1004 -304 -1003
rect -581 -1015 -535 -1005
rect -353 -1015 -307 -1004
rect -180 -1005 -170 -228
rect -111 -1005 -101 -228
rect 23 -1004 33 -227
rect 93 -1003 102 -227
rect 231 -228 237 -227
rect 271 -228 277 -227
rect 92 -1004 102 -1003
rect -175 -1015 -129 -1005
rect 53 -1015 99 -1004
rect 226 -1005 236 -228
rect 295 -1005 305 -228
rect 429 -1004 439 -227
rect 499 -1003 508 -227
rect 637 -228 643 -227
rect 677 -228 683 -227
rect 498 -1004 508 -1003
rect 231 -1015 277 -1005
rect 459 -1015 505 -1004
rect 632 -1005 642 -228
rect 701 -1005 711 -228
rect 835 -1004 845 -227
rect 905 -1003 914 -227
rect 1043 -228 1049 -227
rect 1083 -228 1089 -227
rect 904 -1004 914 -1003
rect 637 -1015 683 -1005
rect 865 -1015 911 -1004
rect 1038 -1005 1048 -228
rect 1107 -1005 1117 -228
rect 1241 -1004 1251 -227
rect 1311 -1003 1320 -227
rect 1449 -228 1455 -227
rect 1489 -228 1495 -227
rect 1310 -1004 1320 -1003
rect 1043 -1015 1089 -1005
rect 1271 -1015 1317 -1004
rect 1444 -1005 1454 -228
rect 1513 -1005 1523 -228
rect 1647 -250 1683 -227
rect 1640 -940 1650 -250
rect 1647 -1003 1683 -940
rect 1717 -1003 1726 -227
rect 1855 -228 1861 -227
rect 1647 -1004 1726 -1003
rect 1850 -1003 1861 -228
rect 1895 -249 1950 -227
rect 1931 -939 1950 -249
rect 1895 -1003 1950 -939
rect 1449 -1015 1495 -1005
rect 1677 -1015 1723 -1004
rect 1850 -1005 1950 -1003
rect 2053 -1004 2063 -227
rect 2123 -1003 2132 -227
rect 2261 -228 2267 -227
rect 2301 -228 2307 -227
rect 2122 -1004 2132 -1003
rect 1855 -1015 1950 -1005
rect 2083 -1015 2129 -1004
rect 2256 -1005 2266 -228
rect 2325 -1005 2335 -228
rect 2459 -1004 2469 -227
rect 2529 -1003 2538 -227
rect 2667 -228 2673 -227
rect 2707 -228 2713 -227
rect 2528 -1004 2538 -1003
rect 2261 -1015 2307 -1005
rect 2489 -1015 2535 -1004
rect 2662 -1005 2672 -228
rect 2731 -1005 2741 -228
rect 2865 -1004 2875 -227
rect 2935 -1003 2944 -227
rect 3073 -228 3079 -227
rect 3113 -228 3119 -227
rect 2934 -1004 2944 -1003
rect 2667 -1015 2713 -1005
rect 2895 -1015 2941 -1004
rect 3068 -1005 3078 -228
rect 3137 -1005 3147 -228
rect 3271 -1004 3281 -227
rect 3341 -1003 3350 -227
rect 3479 -228 3485 -227
rect 3519 -228 3525 -227
rect 3340 -1004 3350 -1003
rect 3073 -1015 3119 -1005
rect 3301 -1015 3347 -1004
rect 3474 -1005 3484 -228
rect 3543 -1005 3553 -228
rect 3677 -1004 3687 -227
rect 3747 -1003 3756 -227
rect 3885 -228 3891 -227
rect 3925 -228 3931 -227
rect 3746 -1004 3756 -1003
rect 3479 -1015 3525 -1005
rect 3707 -1015 3753 -1004
rect 3880 -1005 3890 -228
rect 3949 -1005 3959 -228
rect 4083 -1004 4093 -227
rect 4153 -1003 4162 -227
rect 4291 -228 4297 -227
rect 4331 -228 4337 -227
rect 4152 -1004 4162 -1003
rect 3885 -1015 3931 -1005
rect 4113 -1015 4159 -1004
rect 4286 -1005 4296 -228
rect 4355 -1005 4365 -228
rect 4489 -1004 4499 -227
rect 4559 -1003 4568 -227
rect 4697 -228 4703 -227
rect 4737 -228 4743 -227
rect 4558 -1004 4568 -1003
rect 4291 -1015 4337 -1005
rect 4519 -1015 4565 -1004
rect 4692 -1005 4702 -228
rect 4761 -1005 4771 -228
rect 4895 -1004 4905 -227
rect 4965 -1003 4974 -227
rect 5103 -228 5109 -227
rect 5143 -228 5149 -227
rect 4964 -1004 4974 -1003
rect 4697 -1015 4743 -1005
rect 4925 -1015 4971 -1004
rect 5098 -1005 5108 -228
rect 5167 -1005 5177 -228
rect 5301 -1004 5311 -227
rect 5371 -1003 5380 -227
rect 5509 -228 5515 -227
rect 5549 -228 5555 -227
rect 5370 -1004 5380 -1003
rect 5103 -1015 5149 -1005
rect 5331 -1015 5377 -1004
rect 5504 -1005 5514 -228
rect 5573 -1005 5583 -228
rect 5707 -1004 5717 -227
rect 5777 -1003 5786 -227
rect 5915 -228 5921 -227
rect 5955 -228 5961 -227
rect 5776 -1004 5786 -1003
rect 5509 -1015 5555 -1005
rect 5737 -1015 5783 -1004
rect 5910 -1005 5920 -228
rect 5979 -1005 5989 -228
rect 5915 -1015 5961 -1005
rect 1860 -1020 1950 -1015
rect -2327 -1050 -2215 -1047
rect -1921 -1050 -1809 -1047
rect -1515 -1050 -1403 -1047
rect -1109 -1050 -997 -1047
rect -703 -1050 -591 -1047
rect -297 -1050 -185 -1047
rect 109 -1050 221 -1047
rect 515 -1050 627 -1047
rect 921 -1050 1033 -1047
rect 1327 -1050 1439 -1047
rect 1733 -1050 1845 -1047
rect 1880 -1050 1950 -1020
rect 2139 -1050 2251 -1047
rect 2545 -1050 2657 -1047
rect 2951 -1050 3063 -1047
rect 3357 -1050 3469 -1047
rect 3763 -1050 3875 -1047
rect 4169 -1050 4281 -1047
rect 4575 -1050 4687 -1047
rect 4981 -1050 5093 -1047
rect 5387 -1050 5499 -1047
rect 5793 -1050 5905 -1047
rect -2520 -1051 5910 -1050
rect 6030 -1051 6100 -180
rect 6150 -190 6160 -120
rect 6280 -143 6320 -120
rect 6299 -174 6320 -143
rect 6424 -174 6430 -86
rect 6480 -86 6492 -20
rect 6480 -160 6486 -86
rect 6299 -177 6316 -174
rect 6280 -180 6316 -177
rect 6280 -183 6311 -180
rect 6280 -190 6290 -183
rect 6150 -215 6210 -190
rect 6143 -227 6210 -215
rect 6143 -1003 6149 -227
rect 6183 -1003 6210 -227
rect 6143 -1015 6210 -1003
rect 6321 -227 6367 -215
rect 6321 -1003 6327 -227
rect 6361 -266 6367 -227
rect 6424 -234 6432 -174
rect 6423 -266 6432 -234
rect 6361 -934 6432 -266
rect 6361 -1003 6367 -934
rect 6321 -1015 6367 -1003
rect -2520 -1053 6100 -1051
rect -2520 -1087 -2315 -1053
rect -2227 -1087 -1909 -1053
rect -1821 -1087 -1503 -1053
rect -1415 -1087 -1097 -1053
rect -1009 -1087 -691 -1053
rect -603 -1087 -285 -1053
rect -197 -1087 121 -1053
rect 209 -1087 527 -1053
rect 615 -1087 933 -1053
rect 1021 -1087 1339 -1053
rect 1427 -1087 1745 -1053
rect 1833 -1087 2151 -1053
rect 2239 -1087 2557 -1053
rect 2645 -1087 2963 -1053
rect 3051 -1087 3369 -1053
rect 3457 -1087 3775 -1053
rect 3863 -1087 4181 -1053
rect 4269 -1087 4587 -1053
rect 4675 -1087 4993 -1053
rect 5081 -1087 5399 -1053
rect 5487 -1087 5805 -1053
rect 5893 -1087 6100 -1053
rect 6150 -1047 6210 -1015
rect 6423 -1047 6432 -934
rect 6150 -1053 6311 -1047
rect 6150 -1080 6211 -1053
rect -2520 -1110 6100 -1087
rect 6199 -1087 6211 -1080
rect 6299 -1087 6311 -1053
rect 6199 -1093 6311 -1087
rect 6423 -1117 6431 -1047
rect 6423 -1146 6430 -1117
rect -2494 -1152 6430 -1146
rect -2494 -1212 -2482 -1152
rect 6480 -1200 15800 -160
rect 6470 -1212 15800 -1200
rect -2494 -1218 1640 -1212
rect -2490 -1248 1640 -1218
rect -2516 -1260 1640 -1248
rect 1740 -1260 15800 -1212
rect -2516 -3984 -2510 -1260
rect -2440 -1326 15700 -1320
rect -2440 -2634 -2434 -1326
rect -2352 -1430 -1943 -1418
rect 15230 -1430 15700 -1326
rect -2360 -2540 -2350 -1430
rect -1940 -2540 -1930 -1430
rect -2352 -2544 -2346 -2540
rect -1949 -2544 -1943 -2540
rect -2352 -2556 -1943 -2544
rect 15230 -2544 15241 -1430
rect 15638 -2544 15700 -1430
rect 15230 -2634 15700 -2544
rect -2440 -2640 15700 -2634
rect 15790 -1326 15800 -1260
rect 15790 -2634 15796 -1326
rect 15790 -2640 15806 -2634
rect 15794 -2700 15806 -2640
rect -2522 -4080 -2510 -3984
rect -2440 -2706 15700 -2700
rect -2440 -3984 -2434 -2706
rect -2352 -2802 -1943 -2790
rect -2352 -2810 -2346 -2802
rect -1949 -2810 -1943 -2802
rect 15230 -2802 15700 -2706
rect -2360 -3920 -2350 -2810
rect -1940 -3920 -1930 -2810
rect 15230 -3916 15241 -2802
rect 15638 -3916 15700 -2802
rect -2352 -3928 -1943 -3920
rect 15230 -3984 15700 -3916
rect -2440 -3990 15700 -3984
rect 15790 -2706 15806 -2700
rect 15790 -3984 15796 -2706
rect 15790 -3990 15812 -3984
rect 15800 -4080 15812 -3990
rect -2522 -4086 15812 -4080
<< via1 >>
rect 2460 4490 2690 4620
rect 1874 473 1916 4227
rect 1916 473 1948 4227
rect 2256 623 2276 4133
rect 2276 623 2326 4133
rect 2326 623 2346 4133
rect 2796 623 2826 4133
rect 2826 623 2886 4133
rect 3140 470 3146 4230
rect 3146 470 3180 4230
rect 3180 470 3210 4230
rect 5800 470 6260 670
rect 2140 399 2980 400
rect 2140 365 2146 399
rect 2146 365 2464 399
rect 2464 365 2632 399
rect 2632 365 2950 399
rect 2950 365 2980 399
rect 2140 330 2980 365
rect 1330 50 1350 80
rect 1350 50 1410 80
rect 1330 20 1410 50
rect -2403 -1003 -2377 -227
rect -2377 -1003 -2344 -227
rect -2403 -1004 -2344 -1003
rect -2200 -1003 -2199 -228
rect -2199 -1003 -2165 -228
rect -2165 -1003 -2141 -228
rect -2200 -1005 -2141 -1003
rect -1997 -1003 -1971 -227
rect -1971 -1003 -1938 -227
rect -1997 -1004 -1938 -1003
rect -1794 -1003 -1793 -228
rect -1793 -1003 -1759 -228
rect -1759 -1003 -1735 -228
rect -1794 -1005 -1735 -1003
rect -1591 -1003 -1565 -227
rect -1565 -1003 -1532 -227
rect -1591 -1004 -1532 -1003
rect -1388 -1003 -1387 -228
rect -1387 -1003 -1353 -228
rect -1353 -1003 -1329 -228
rect -1388 -1005 -1329 -1003
rect -1185 -1003 -1159 -227
rect -1159 -1003 -1126 -227
rect -1185 -1004 -1126 -1003
rect -982 -1003 -981 -228
rect -981 -1003 -947 -228
rect -947 -1003 -923 -228
rect -982 -1005 -923 -1003
rect -779 -1003 -753 -227
rect -753 -1003 -720 -227
rect -779 -1004 -720 -1003
rect -576 -1003 -575 -228
rect -575 -1003 -541 -228
rect -541 -1003 -517 -228
rect -576 -1005 -517 -1003
rect -373 -1003 -347 -227
rect -347 -1003 -314 -227
rect -373 -1004 -314 -1003
rect -170 -1003 -169 -228
rect -169 -1003 -135 -228
rect -135 -1003 -111 -228
rect -170 -1005 -111 -1003
rect 33 -1003 59 -227
rect 59 -1003 92 -227
rect 33 -1004 92 -1003
rect 236 -1003 237 -228
rect 237 -1003 271 -228
rect 271 -1003 295 -228
rect 236 -1005 295 -1003
rect 439 -1003 465 -227
rect 465 -1003 498 -227
rect 439 -1004 498 -1003
rect 642 -1003 643 -228
rect 643 -1003 677 -228
rect 677 -1003 701 -228
rect 642 -1005 701 -1003
rect 845 -1003 871 -227
rect 871 -1003 904 -227
rect 845 -1004 904 -1003
rect 1048 -1003 1049 -228
rect 1049 -1003 1083 -228
rect 1083 -1003 1107 -228
rect 1048 -1005 1107 -1003
rect 1251 -1003 1277 -227
rect 1277 -1003 1310 -227
rect 1251 -1004 1310 -1003
rect 1454 -1003 1455 -228
rect 1455 -1003 1489 -228
rect 1489 -1003 1513 -228
rect 1454 -1005 1513 -1003
rect 1650 -940 1683 -250
rect 1683 -940 1710 -250
rect 1871 -939 1895 -249
rect 1895 -939 1931 -249
rect 2063 -1003 2089 -227
rect 2089 -1003 2122 -227
rect 2063 -1004 2122 -1003
rect 2266 -1003 2267 -228
rect 2267 -1003 2301 -228
rect 2301 -1003 2325 -228
rect 2266 -1005 2325 -1003
rect 2469 -1003 2495 -227
rect 2495 -1003 2528 -227
rect 2469 -1004 2528 -1003
rect 2672 -1003 2673 -228
rect 2673 -1003 2707 -228
rect 2707 -1003 2731 -228
rect 2672 -1005 2731 -1003
rect 2875 -1003 2901 -227
rect 2901 -1003 2934 -227
rect 2875 -1004 2934 -1003
rect 3078 -1003 3079 -228
rect 3079 -1003 3113 -228
rect 3113 -1003 3137 -228
rect 3078 -1005 3137 -1003
rect 3281 -1003 3307 -227
rect 3307 -1003 3340 -227
rect 3281 -1004 3340 -1003
rect 3484 -1003 3485 -228
rect 3485 -1003 3519 -228
rect 3519 -1003 3543 -228
rect 3484 -1005 3543 -1003
rect 3687 -1003 3713 -227
rect 3713 -1003 3746 -227
rect 3687 -1004 3746 -1003
rect 3890 -1003 3891 -228
rect 3891 -1003 3925 -228
rect 3925 -1003 3949 -228
rect 3890 -1005 3949 -1003
rect 4093 -1003 4119 -227
rect 4119 -1003 4152 -227
rect 4093 -1004 4152 -1003
rect 4296 -1003 4297 -228
rect 4297 -1003 4331 -228
rect 4331 -1003 4355 -228
rect 4296 -1005 4355 -1003
rect 4499 -1003 4525 -227
rect 4525 -1003 4558 -227
rect 4499 -1004 4558 -1003
rect 4702 -1003 4703 -228
rect 4703 -1003 4737 -228
rect 4737 -1003 4761 -228
rect 4702 -1005 4761 -1003
rect 4905 -1003 4931 -227
rect 4931 -1003 4964 -227
rect 4905 -1004 4964 -1003
rect 5108 -1003 5109 -228
rect 5109 -1003 5143 -228
rect 5143 -1003 5167 -228
rect 5108 -1005 5167 -1003
rect 5311 -1003 5337 -227
rect 5337 -1003 5370 -227
rect 5311 -1004 5370 -1003
rect 5514 -1003 5515 -228
rect 5515 -1003 5549 -228
rect 5549 -1003 5573 -228
rect 5514 -1005 5573 -1003
rect 5717 -1003 5743 -227
rect 5743 -1003 5776 -227
rect 5717 -1004 5776 -1003
rect 5920 -1003 5921 -228
rect 5921 -1003 5955 -228
rect 5955 -1003 5979 -228
rect 5920 -1005 5979 -1003
rect 6160 -143 6280 -120
rect 6160 -177 6211 -143
rect 6211 -177 6280 -143
rect 6160 -190 6280 -177
rect 1640 -1212 1740 -1210
rect 1640 -1260 1740 -1212
rect 1640 -1290 1740 -1260
rect -2350 -2540 -2346 -1430
rect -2346 -2540 -1949 -1430
rect -1949 -2540 -1940 -1430
rect -2350 -3916 -2346 -2810
rect -2346 -3916 -1949 -2810
rect -1949 -3916 -1940 -2810
rect -2350 -3920 -1940 -3916
<< metal2 >>
rect 2226 4620 2926 4633
rect 2226 4490 2460 4620
rect 2690 4490 2926 4620
rect 2226 4423 2926 4490
rect 1874 4227 1948 4237
rect 2226 4133 2376 4423
rect 2226 4073 2256 4133
rect 2346 4073 2376 4133
rect 2786 4133 2926 4423
rect 2786 4073 2796 4133
rect 2256 613 2346 623
rect 2886 4073 2926 4133
rect 3140 4230 3210 4240
rect 2796 613 2886 623
rect 1874 463 1948 473
rect 3210 670 6280 680
rect 3210 470 5800 670
rect 6260 470 6280 670
rect 3140 460 6280 470
rect 2140 400 2980 410
rect 1870 100 1950 110
rect 1320 20 1330 80
rect 1410 20 1870 80
rect 1330 10 1870 20
rect 1870 0 1950 10
rect 2140 -80 2980 330
rect -2200 -120 5980 -80
rect 6160 -120 6280 460
rect -2200 -160 5979 -120
rect -2403 -227 -2344 -217
rect -2403 -1005 -2344 -1004
rect -2404 -1014 -2344 -1005
rect -2200 -228 -2141 -160
rect -1997 -227 -1938 -217
rect -1997 -1005 -1938 -1004
rect -2404 -1060 -2345 -1014
rect -2200 -1015 -2141 -1005
rect -1998 -1014 -1938 -1005
rect -1794 -228 -1735 -160
rect -1591 -227 -1532 -217
rect -1591 -1005 -1532 -1004
rect -1998 -1060 -1939 -1014
rect -1794 -1015 -1735 -1005
rect -1592 -1014 -1532 -1005
rect -1388 -228 -1329 -160
rect -1185 -227 -1126 -217
rect -1185 -1005 -1126 -1004
rect -1592 -1060 -1533 -1014
rect -1388 -1015 -1329 -1005
rect -1186 -1014 -1126 -1005
rect -982 -228 -923 -160
rect -779 -227 -720 -217
rect -779 -1005 -720 -1004
rect -1186 -1060 -1127 -1014
rect -982 -1015 -923 -1005
rect -780 -1014 -720 -1005
rect -576 -228 -517 -160
rect -373 -227 -314 -217
rect -373 -1005 -314 -1004
rect -780 -1060 -721 -1014
rect -576 -1015 -517 -1005
rect -374 -1014 -314 -1005
rect -170 -228 -111 -160
rect 33 -227 92 -217
rect 33 -1005 92 -1004
rect -374 -1060 -315 -1014
rect -170 -1015 -111 -1005
rect 32 -1014 92 -1005
rect 236 -228 295 -160
rect 439 -227 498 -217
rect 439 -1005 498 -1004
rect 32 -1060 91 -1014
rect 236 -1015 295 -1005
rect 438 -1014 498 -1005
rect 642 -228 701 -160
rect 845 -227 904 -217
rect 845 -1005 904 -1004
rect 438 -1060 497 -1014
rect 642 -1015 701 -1005
rect 844 -1014 904 -1005
rect 1048 -228 1107 -160
rect 1251 -227 1310 -217
rect 1251 -1005 1310 -1004
rect 844 -1060 903 -1014
rect 1048 -1015 1107 -1005
rect 1250 -1014 1310 -1005
rect 1454 -228 1513 -160
rect 2063 -227 2122 -217
rect 1650 -250 1710 -240
rect 1650 -950 1710 -940
rect 1871 -249 1931 -239
rect 1871 -949 1931 -939
rect 2063 -1005 2122 -1004
rect 1250 -1060 1309 -1014
rect 1454 -1015 1513 -1005
rect 2062 -1014 2122 -1005
rect 2266 -228 2325 -160
rect 2469 -227 2528 -217
rect 2469 -1005 2528 -1004
rect 2062 -1060 2121 -1014
rect 2266 -1015 2325 -1005
rect 2468 -1014 2528 -1005
rect 2672 -228 2731 -160
rect 2875 -227 2934 -217
rect 2875 -1005 2934 -1004
rect 2468 -1060 2527 -1014
rect 2672 -1015 2731 -1005
rect 2874 -1014 2934 -1005
rect 3078 -228 3137 -160
rect 3281 -227 3340 -217
rect 3281 -1005 3340 -1004
rect 2874 -1060 2933 -1014
rect 3078 -1015 3137 -1005
rect 3280 -1014 3340 -1005
rect 3484 -228 3543 -160
rect 3687 -227 3746 -217
rect 3687 -1005 3746 -1004
rect 3280 -1060 3339 -1014
rect 3484 -1015 3543 -1005
rect 3686 -1014 3746 -1005
rect 3890 -228 3949 -160
rect 4093 -227 4152 -217
rect 4093 -1005 4152 -1004
rect 3686 -1060 3745 -1014
rect 3890 -1015 3949 -1005
rect 4092 -1014 4152 -1005
rect 4296 -228 4355 -160
rect 4499 -227 4558 -217
rect 4499 -1005 4558 -1004
rect 4092 -1060 4151 -1014
rect 4296 -1015 4355 -1005
rect 4498 -1014 4558 -1005
rect 4702 -228 4761 -160
rect 4905 -227 4964 -217
rect 4905 -1005 4964 -1004
rect 4498 -1060 4557 -1014
rect 4702 -1015 4761 -1005
rect 4904 -1014 4964 -1005
rect 5108 -228 5167 -160
rect 5311 -227 5370 -217
rect 5311 -1005 5370 -1004
rect 4904 -1060 4963 -1014
rect 5108 -1015 5167 -1005
rect 5310 -1014 5370 -1005
rect 5514 -228 5573 -160
rect 5717 -227 5776 -217
rect 5717 -1005 5776 -1004
rect 5310 -1060 5369 -1014
rect 5514 -1015 5573 -1005
rect 5716 -1014 5776 -1005
rect 5920 -228 5979 -160
rect 6160 -200 6280 -190
rect 5716 -1060 5775 -1014
rect 5920 -1015 5979 -1005
rect -2404 -1112 5775 -1060
rect -2404 -1152 5776 -1112
rect -2404 -1153 -1930 -1152
rect -1592 -1153 -1533 -1152
rect -1186 -1153 -1127 -1152
rect -780 -1153 -721 -1152
rect -374 -1153 -315 -1152
rect 32 -1153 91 -1152
rect 438 -1153 497 -1152
rect 844 -1153 903 -1152
rect 1250 -1153 1309 -1152
rect 1656 -1153 1715 -1152
rect 2062 -1153 2121 -1152
rect 2468 -1153 2527 -1152
rect 2874 -1153 2933 -1152
rect 3280 -1153 3339 -1152
rect 3686 -1153 3745 -1152
rect 4092 -1153 4151 -1152
rect 4498 -1153 4557 -1152
rect 4904 -1153 4963 -1152
rect 5310 -1153 5369 -1152
rect 5716 -1153 5775 -1152
rect -2400 -1210 -1930 -1153
rect -2340 -1420 -1930 -1210
rect 1640 -1210 1740 -1200
rect 1640 -1300 1740 -1290
rect -2350 -1430 -1930 -1420
rect -1940 -2540 -1930 -1430
rect -2350 -2550 -1930 -2540
rect -2340 -2800 -1930 -2550
rect -2350 -2810 -1930 -2800
rect -1940 -3920 -1930 -2810
rect -2350 -3930 -1940 -3920
<< via2 >>
rect 1874 473 1948 4227
rect 1870 10 1950 100
rect 1650 -940 1710 -250
rect 1871 -939 1931 -249
rect 1640 -1290 1740 -1210
<< metal3 >>
rect 1864 4227 1958 4232
rect 1864 473 1874 4227
rect 1948 473 1958 4227
rect 1864 468 1958 473
rect 1871 105 1947 468
rect 1860 100 1960 105
rect 1860 10 1870 100
rect 1950 10 1960 100
rect 1860 5 1960 10
rect 1871 -130 1947 5
rect 1870 -244 1950 -130
rect 1640 -250 1720 -245
rect 1640 -940 1650 -250
rect 1710 -940 1720 -250
rect 1640 -945 1720 -940
rect 1861 -249 1950 -244
rect 1861 -939 1871 -249
rect 1931 -300 1950 -249
rect 1931 -939 1947 -300
rect 1861 -944 1941 -939
rect 1640 -1205 1710 -945
rect 1630 -1210 1750 -1205
rect 1630 -1290 1640 -1210
rect 1740 -1290 1750 -1210
rect 1630 -1295 1750 -1290
<< labels >>
flabel metal1 2466 4493 2666 4693 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 6380 510 6580 710 0 FreeSans 256 0 0 0 VOUT
port 1 nsew
flabel metal1 9480 -990 9680 -790 0 FreeSans 256 0 0 0 VSS
port 2 nsew
<< end >>
