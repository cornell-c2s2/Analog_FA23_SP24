magic
tech sky130A
magscale 1 2
timestamp 1712613491
<< nwell >>
rect -1630 -250 2190 180
rect 450 -510 2190 -250
rect 450 -1770 2190 -1120
rect 440 -3010 2190 -2360
rect 450 -4250 2190 -3610
rect 440 -5490 2190 -4840
rect 440 -6730 2190 -6070
<< pwell >>
rect -1600 230 170 500
rect 250 -1020 1940 -570
rect 250 -2280 1500 -1830
rect 250 -3550 940 -3070
rect 250 -4790 1690 -4300
rect 250 -6030 1140 -5530
rect 250 -6970 1970 -6760
<< psubdiff >>
rect 20 460 130 480
rect 20 410 50 460
rect 100 410 130 460
rect 20 340 130 410
rect 20 290 50 340
rect 100 290 130 340
rect 20 260 130 290
rect 330 -660 450 -630
rect 330 -720 360 -660
rect 420 -720 450 -660
rect 330 -750 450 -720
rect 330 -860 450 -830
rect 330 -920 360 -860
rect 420 -920 450 -860
rect 330 -950 450 -920
rect 310 -1900 430 -1870
rect 310 -1960 340 -1900
rect 400 -1960 430 -1900
rect 310 -1990 430 -1960
rect 310 -2150 430 -2120
rect 310 -2210 340 -2150
rect 400 -2210 430 -2150
rect 310 -2240 430 -2210
rect 330 -3160 450 -3130
rect 330 -3220 360 -3160
rect 420 -3220 450 -3160
rect 330 -3330 450 -3220
rect 330 -3390 360 -3330
rect 420 -3390 450 -3330
rect 330 -3420 450 -3390
rect 320 -4410 440 -4380
rect 320 -4470 350 -4410
rect 410 -4470 440 -4410
rect 320 -4500 440 -4470
rect 320 -4590 440 -4560
rect 320 -4650 350 -4590
rect 410 -4650 440 -4590
rect 320 -4680 440 -4650
rect 310 -5580 430 -5550
rect 310 -5640 340 -5580
rect 400 -5640 430 -5580
rect 310 -5670 430 -5640
rect 310 -5830 430 -5800
rect 310 -5890 340 -5830
rect 400 -5890 430 -5830
rect 310 -5920 430 -5890
rect 300 -6830 420 -6800
rect 300 -6890 330 -6830
rect 390 -6890 420 -6830
rect 300 -6920 420 -6890
<< nsubdiff >>
rect -160 0 -50 30
rect -160 -50 -130 0
rect -80 -50 -50 0
rect -160 -130 -50 -50
rect -160 -180 -130 -130
rect -80 -180 -50 -130
rect -160 -210 -50 -180
rect 1160 -1420 1270 -1390
rect 1160 -1470 1190 -1420
rect 1240 -1470 1270 -1420
rect 1160 -1500 1270 -1470
rect 1470 -1420 1580 -1390
rect 1470 -1470 1500 -1420
rect 1550 -1470 1580 -1420
rect 1470 -1500 1580 -1470
rect 1710 -1420 1820 -1390
rect 1710 -1470 1740 -1420
rect 1790 -1470 1820 -1420
rect 1710 -1500 1820 -1470
rect 1970 -1420 2080 -1390
rect 1970 -1470 2000 -1420
rect 2050 -1470 2080 -1420
rect 1970 -1500 2080 -1470
rect 1540 -2660 1650 -2630
rect 1540 -2710 1570 -2660
rect 1620 -2710 1650 -2660
rect 1540 -2740 1650 -2710
rect 1760 -2660 1870 -2630
rect 1760 -2710 1790 -2660
rect 1840 -2710 1870 -2660
rect 1760 -2740 1870 -2710
rect 2000 -2660 2110 -2630
rect 2000 -2710 2030 -2660
rect 2080 -2710 2110 -2660
rect 2000 -2740 2110 -2710
rect 1730 -3910 1840 -3880
rect 1730 -3960 1760 -3910
rect 1810 -3960 1840 -3910
rect 1730 -3990 1840 -3960
rect 1960 -3910 2070 -3880
rect 1960 -3960 1990 -3910
rect 2040 -3960 2070 -3910
rect 1960 -3990 2070 -3960
rect 1190 -5140 1300 -5110
rect 1190 -5190 1220 -5140
rect 1270 -5190 1300 -5140
rect 1190 -5220 1300 -5190
rect 1490 -5140 1600 -5110
rect 1490 -5190 1520 -5140
rect 1570 -5190 1600 -5140
rect 1490 -5220 1600 -5190
rect 1790 -5140 1900 -5110
rect 1790 -5190 1820 -5140
rect 1870 -5190 1900 -5140
rect 1790 -5220 1900 -5190
rect 2030 -6380 2140 -6350
rect 2030 -6430 2060 -6380
rect 2110 -6430 2140 -6380
rect 2030 -6460 2140 -6430
<< psubdiffcont >>
rect 50 410 100 460
rect 50 290 100 340
rect 360 -720 420 -660
rect 360 -920 420 -860
rect 340 -1960 400 -1900
rect 340 -2210 400 -2150
rect 360 -3220 420 -3160
rect 360 -3390 420 -3330
rect 350 -4470 410 -4410
rect 350 -4650 410 -4590
rect 340 -5640 400 -5580
rect 340 -5890 400 -5830
rect 330 -6890 390 -6830
<< nsubdiffcont >>
rect -130 -50 -80 0
rect -130 -180 -80 -130
rect 1190 -1470 1240 -1420
rect 1500 -1470 1550 -1420
rect 1740 -1470 1790 -1420
rect 2000 -1470 2050 -1420
rect 1570 -2710 1620 -2660
rect 1790 -2710 1840 -2660
rect 2030 -2710 2080 -2660
rect 1760 -3960 1810 -3910
rect 1990 -3960 2040 -3910
rect 1220 -5190 1270 -5140
rect 1520 -5190 1570 -5140
rect 1820 -5190 1870 -5140
rect 2060 -6430 2110 -6380
<< viali >>
rect 20 460 130 480
rect 20 410 50 460
rect 50 410 100 460
rect 100 410 130 460
rect 20 340 130 410
rect -1420 279 -1386 313
rect -1148 276 -1114 310
rect -873 277 -839 311
rect -598 277 -564 311
rect -322 275 -288 309
rect 20 290 50 340
rect 50 290 100 340
rect 100 290 130 340
rect 20 260 130 290
rect -1510 180 -1470 220
rect -1420 187 -1386 221
rect -1228 193 -1194 227
rect -1143 187 -1109 221
rect -962 186 -928 220
rect -866 186 -832 220
rect -686 187 -652 221
rect -593 187 -559 221
rect -410 187 -376 221
rect -318 186 -284 220
rect -1420 98 -1386 132
rect -1147 93 -1113 127
rect -875 92 -841 126
rect -598 93 -564 127
rect -322 93 -288 127
rect -872 20 -838 54
rect -160 0 -50 30
rect -160 -50 -130 0
rect -130 -50 -80 0
rect -80 -50 -50 0
rect -160 -130 -50 -50
rect -160 -180 -130 -130
rect -130 -180 -80 -130
rect -80 -180 -50 -130
rect -160 -210 -50 -180
rect 330 -660 450 -630
rect 330 -720 360 -660
rect 360 -720 420 -660
rect 420 -720 450 -660
rect 330 -750 450 -720
rect 330 -860 450 -830
rect 330 -920 360 -860
rect 360 -920 420 -860
rect 420 -920 450 -860
rect 330 -950 450 -920
rect 1160 -1420 1270 -1390
rect 1160 -1470 1190 -1420
rect 1190 -1470 1240 -1420
rect 1240 -1470 1270 -1420
rect 1160 -1500 1270 -1470
rect 1470 -1420 1580 -1390
rect 1470 -1470 1500 -1420
rect 1500 -1470 1550 -1420
rect 1550 -1470 1580 -1420
rect 1470 -1500 1580 -1470
rect 1710 -1420 1820 -1390
rect 1710 -1470 1740 -1420
rect 1740 -1470 1790 -1420
rect 1790 -1470 1820 -1420
rect 1710 -1500 1820 -1470
rect 1970 -1420 2080 -1390
rect 1970 -1470 2000 -1420
rect 2000 -1470 2050 -1420
rect 2050 -1470 2080 -1420
rect 1970 -1500 2080 -1470
rect 310 -1900 430 -1870
rect 310 -1960 340 -1900
rect 340 -1960 400 -1900
rect 400 -1960 430 -1900
rect 310 -1990 430 -1960
rect 310 -2150 430 -2120
rect 310 -2210 340 -2150
rect 340 -2210 400 -2150
rect 400 -2210 430 -2150
rect 310 -2240 430 -2210
rect 1540 -2660 1650 -2630
rect 1540 -2710 1570 -2660
rect 1570 -2710 1620 -2660
rect 1620 -2710 1650 -2660
rect 1540 -2740 1650 -2710
rect 1760 -2660 1870 -2630
rect 1760 -2710 1790 -2660
rect 1790 -2710 1840 -2660
rect 1840 -2710 1870 -2660
rect 1760 -2740 1870 -2710
rect 2000 -2660 2110 -2630
rect 2000 -2710 2030 -2660
rect 2030 -2710 2080 -2660
rect 2080 -2710 2110 -2660
rect 2000 -2740 2110 -2710
rect 330 -3160 450 -3130
rect 330 -3220 360 -3160
rect 360 -3220 420 -3160
rect 420 -3220 450 -3160
rect 330 -3330 450 -3220
rect 330 -3390 360 -3330
rect 360 -3390 420 -3330
rect 420 -3390 450 -3330
rect 330 -3420 450 -3390
rect 1730 -3910 1840 -3880
rect 1730 -3960 1760 -3910
rect 1760 -3960 1810 -3910
rect 1810 -3960 1840 -3910
rect 1730 -3990 1840 -3960
rect 1960 -3910 2070 -3880
rect 1960 -3960 1990 -3910
rect 1990 -3960 2040 -3910
rect 2040 -3960 2070 -3910
rect 1960 -3990 2070 -3960
rect 320 -4410 440 -4380
rect 320 -4470 350 -4410
rect 350 -4470 410 -4410
rect 410 -4470 440 -4410
rect 320 -4500 440 -4470
rect 320 -4590 440 -4560
rect 320 -4650 350 -4590
rect 350 -4650 410 -4590
rect 410 -4650 440 -4590
rect 320 -4680 440 -4650
rect 1190 -5140 1300 -5110
rect 1190 -5190 1220 -5140
rect 1220 -5190 1270 -5140
rect 1270 -5190 1300 -5140
rect 1190 -5220 1300 -5190
rect 1490 -5140 1600 -5110
rect 1490 -5190 1520 -5140
rect 1520 -5190 1570 -5140
rect 1570 -5190 1600 -5140
rect 1490 -5220 1600 -5190
rect 1790 -5140 1900 -5110
rect 1790 -5190 1820 -5140
rect 1820 -5190 1870 -5140
rect 1870 -5190 1900 -5140
rect 1790 -5220 1900 -5190
rect 310 -5580 430 -5550
rect 310 -5640 340 -5580
rect 340 -5640 400 -5580
rect 400 -5640 430 -5580
rect 310 -5670 430 -5640
rect 310 -5830 430 -5800
rect 310 -5890 340 -5830
rect 340 -5890 400 -5830
rect 400 -5890 430 -5830
rect 310 -5920 430 -5890
rect 2030 -6380 2140 -6350
rect 2030 -6430 2060 -6380
rect 2060 -6430 2110 -6380
rect 2110 -6430 2140 -6380
rect 2030 -6460 2140 -6430
rect 300 -6830 420 -6800
rect 300 -6890 330 -6830
rect 330 -6890 390 -6830
rect 390 -6890 420 -6830
rect 300 -6920 420 -6890
<< metal1 >>
rect -3910 470 -3710 690
rect -3910 280 -3870 470
rect -3750 280 -3710 470
rect -3910 270 -3710 280
rect -3660 470 -3460 690
rect -3660 280 -3620 470
rect -3500 280 -3460 470
rect -3660 270 -3460 280
rect -3410 470 -3210 690
rect -3410 280 -3370 470
rect -3250 280 -3210 470
rect -3410 270 -3210 280
rect -3160 470 -2960 690
rect -3160 280 -3120 470
rect -3000 280 -2960 470
rect -3160 270 -2960 280
rect -2910 470 -2710 690
rect -2910 280 -2870 470
rect -2750 280 -2710 470
rect -2910 270 -2710 280
rect -2660 470 -2460 690
rect -2660 280 -2620 470
rect -2500 280 -2460 470
rect -2660 270 -2460 280
rect -2410 470 -2210 690
rect -2410 280 -2370 470
rect -2250 280 -2210 470
rect -2410 270 -2210 280
rect -2160 470 -1960 690
rect -2160 280 -2120 470
rect -2000 280 -1960 470
rect -2160 270 -1960 280
rect -1910 470 -1710 690
rect -210 490 170 494
rect -1910 280 -1870 470
rect -1750 280 -1710 470
rect -1590 480 170 490
rect -1590 420 20 480
rect -1590 390 -170 420
rect -1429 330 -1362 336
rect -1910 270 -1710 280
rect -1430 313 -1362 330
rect -1430 279 -1420 313
rect -1386 279 -1362 313
rect -1430 260 -1362 279
rect -1157 310 -1079 338
rect -325 332 -273 338
rect -1157 276 -1148 310
rect -1114 276 -1079 310
rect -1157 260 -1079 276
rect -886 311 -822 327
rect -886 277 -873 311
rect -839 277 -822 311
rect -886 260 -822 277
rect -607 311 -541 324
rect -607 277 -598 311
rect -564 277 -541 311
rect -1690 240 -1610 250
rect -1430 247 -1326 260
rect -1700 234 -1680 240
rect -3380 182 -3367 234
rect -3250 182 -1680 234
rect -1690 180 -1680 182
rect -1620 234 -1600 240
rect -1530 234 -1460 240
rect -1620 220 -1460 234
rect -1620 182 -1510 220
rect -1620 180 -1610 182
rect -1690 170 -1610 180
rect -1530 180 -1510 182
rect -1470 180 -1460 220
rect -1530 160 -1460 180
rect -1430 221 -1417 247
rect -1430 187 -1420 221
rect -1430 169 -1417 187
rect -1339 169 -1326 247
rect -1430 156 -1326 169
rect -1250 248 -1190 249
rect -1250 227 -1188 248
rect -1250 193 -1228 227
rect -1194 193 -1188 227
rect -1250 167 -1188 193
rect -1157 247 -1053 260
rect -1157 169 -1144 247
rect -1066 169 -1053 247
rect -1157 156 -1053 169
rect -988 247 -923 260
rect -886 247 -767 260
rect -607 247 -541 277
rect -331 309 -273 332
rect -331 275 -322 309
rect -288 275 -273 309
rect -331 247 -273 275
rect -208 300 -170 390
rect -30 300 20 420
rect -208 260 20 300
rect 130 260 170 480
rect -208 250 170 260
rect -923 169 -922 234
rect -886 220 -858 247
rect -886 186 -866 220
rect -886 169 -858 186
rect -780 169 -767 247
rect -988 156 -923 169
rect -886 156 -767 169
rect -728 236 -637 247
rect -728 221 -635 236
rect -728 187 -686 221
rect -652 187 -635 221
rect -728 167 -635 187
rect -607 234 -494 247
rect -607 221 -585 234
rect -607 187 -593 221
rect -607 169 -585 187
rect -507 169 -494 234
rect -728 156 -637 167
rect -607 156 -494 169
rect -455 234 -364 247
rect -455 156 -442 234
rect -1430 132 -1362 156
rect -1430 98 -1420 132
rect -1386 98 -1362 132
rect -1430 80 -1362 98
rect -1157 127 -1079 156
rect -1157 93 -1147 127
rect -1113 93 -1079 127
rect -1157 52 -1079 93
rect -886 126 -822 156
rect -886 92 -875 126
rect -841 92 -822 126
rect -886 54 -822 92
rect -607 127 -541 156
rect -455 143 -364 156
rect -331 234 -247 247
rect -331 220 -299 234
rect -331 186 -318 220
rect -331 156 -299 186
rect -331 143 -247 156
rect -607 93 -598 127
rect -564 93 -541 127
rect -607 76 -541 93
rect -331 127 -273 143
rect -331 93 -322 127
rect -288 93 -273 127
rect -331 74 -273 93
rect -886 20 -872 54
rect -838 20 -822 54
rect -886 7 -822 20
rect -325 0 -273 74
rect -240 40 1960 70
rect -240 30 80 40
rect -240 -50 -160 30
rect -1590 -150 -160 -50
rect -240 -210 -160 -150
rect -50 -210 80 30
rect 340 -210 1960 40
rect -240 -250 1960 -210
rect 1510 -310 1960 -250
rect -312 -351 -221 -338
rect -312 -416 -299 -351
rect -234 -416 -221 -351
rect -312 -429 -221 -416
rect -299 -455 -234 -429
rect 310 -630 470 -610
rect 310 -720 330 -630
rect -190 -740 330 -720
rect -190 -890 -170 -740
rect -30 -750 330 -740
rect 450 -720 470 -630
rect 450 -750 1960 -720
rect -30 -830 1960 -750
rect -30 -890 330 -830
rect -190 -910 330 -890
rect 310 -950 330 -910
rect 450 -910 1960 -830
rect 450 -950 470 -910
rect 310 -970 470 -950
rect 2290 -1320 2620 -1290
rect 2290 -1350 2320 -1320
rect 480 -1390 2320 -1350
rect 480 -1500 1160 -1390
rect 1270 -1500 1470 -1390
rect 1580 -1500 1710 -1390
rect 1820 -1500 1970 -1390
rect 2080 -1500 2320 -1390
rect 480 -1530 2320 -1500
rect 2290 -1560 2320 -1530
rect 2590 -1560 2620 -1320
rect 2290 -1580 2620 -1560
rect 290 -1870 450 -1850
rect 290 -1970 310 -1870
rect -190 -1990 310 -1970
rect 430 -1970 450 -1870
rect 430 -1990 1500 -1970
rect -190 -2130 -170 -1990
rect -30 -2120 1500 -1990
rect -30 -2130 310 -2120
rect -190 -2150 310 -2130
rect 290 -2240 310 -2150
rect 430 -2150 1500 -2120
rect 430 -2240 450 -2150
rect 290 -2260 450 -2240
rect 2290 -2550 2620 -2520
rect 2290 -2590 2320 -2550
rect 480 -2630 2320 -2590
rect 480 -2740 1540 -2630
rect 1650 -2740 1760 -2630
rect 1870 -2740 2000 -2630
rect 2110 -2740 2320 -2630
rect 480 -2770 2320 -2740
rect 2290 -2790 2320 -2770
rect 2590 -2790 2620 -2550
rect 2290 -2820 2620 -2790
rect 3010 -2990 3210 -2790
rect 310 -3130 470 -3110
rect 310 -3210 330 -3130
rect -190 -3230 330 -3210
rect -190 -3390 -170 -3230
rect -30 -3390 330 -3230
rect -190 -3410 330 -3390
rect 310 -3420 330 -3410
rect 450 -3210 470 -3130
rect 450 -3410 950 -3210
rect 3010 -3390 3210 -3190
rect 450 -3420 470 -3410
rect 310 -3440 470 -3420
rect 2290 -3810 2620 -3780
rect 3010 -3790 3210 -3590
rect 2290 -3850 2320 -3810
rect 480 -3880 2320 -3850
rect 480 -3990 1730 -3880
rect 1840 -3990 1960 -3880
rect 2070 -3990 2320 -3880
rect 480 -4020 2320 -3990
rect 2290 -4050 2320 -4020
rect 2590 -4050 2620 -3810
rect 2290 -4080 2620 -4050
rect 3010 -4190 3210 -3990
rect 300 -4380 460 -4360
rect 300 -4460 320 -4380
rect -190 -4480 320 -4460
rect -190 -4620 -170 -4480
rect -30 -4500 320 -4480
rect 440 -4460 460 -4380
rect 440 -4500 1690 -4460
rect -30 -4560 1690 -4500
rect -30 -4620 320 -4560
rect -190 -4640 320 -4620
rect 300 -4680 320 -4640
rect 440 -4640 1690 -4560
rect 440 -4680 460 -4640
rect 300 -4700 460 -4680
rect 2290 -5030 2620 -5000
rect 2290 -5080 2320 -5030
rect 480 -5110 2320 -5080
rect 480 -5220 1190 -5110
rect 1300 -5220 1490 -5110
rect 1600 -5220 1790 -5110
rect 1900 -5220 2320 -5110
rect 480 -5250 2320 -5220
rect 2290 -5270 2320 -5250
rect 2590 -5270 2620 -5030
rect 2290 -5300 2620 -5270
rect 290 -5550 450 -5530
rect 290 -5670 310 -5550
rect 430 -5670 450 -5550
rect -190 -5690 450 -5670
rect -190 -5780 -170 -5690
rect -30 -5780 1140 -5690
rect -190 -5800 1140 -5780
rect 290 -5920 310 -5800
rect 430 -5870 1140 -5800
rect 430 -5920 450 -5870
rect 290 -5940 450 -5920
rect 2290 -6290 2620 -6260
rect 2290 -6310 2320 -6290
rect 480 -6350 2320 -6310
rect 480 -6460 2030 -6350
rect 2140 -6460 2320 -6350
rect 480 -6490 2320 -6460
rect 2290 -6530 2320 -6490
rect 2590 -6530 2620 -6290
rect 2290 -6560 2620 -6530
rect 290 -6790 430 -6780
rect -190 -6800 430 -6790
rect -190 -6810 300 -6800
rect -190 -6910 -170 -6810
rect -30 -6910 300 -6810
rect -190 -6920 300 -6910
rect 420 -6920 430 -6800
rect -190 -6930 430 -6920
rect 290 -7050 1970 -6930
<< via1 >>
rect -3870 280 -3750 470
rect -3620 280 -3500 470
rect -3370 280 -3250 470
rect -3120 280 -3000 470
rect -2870 280 -2750 470
rect -2620 280 -2500 470
rect -2370 280 -2250 470
rect -2120 280 -2000 470
rect -1870 280 -1750 470
rect -3367 182 -3250 234
rect -1680 180 -1620 240
rect -1417 221 -1339 247
rect -1417 187 -1386 221
rect -1386 187 -1339 221
rect -1417 169 -1339 187
rect -1144 221 -1066 247
rect -1144 187 -1143 221
rect -1143 187 -1109 221
rect -1109 187 -1066 221
rect -1144 169 -1066 187
rect -988 220 -923 247
rect -170 300 -30 420
rect -988 186 -962 220
rect -962 186 -928 220
rect -928 186 -923 220
rect -988 169 -923 186
rect -858 220 -780 247
rect -858 186 -832 220
rect -832 186 -780 220
rect -858 169 -780 186
rect -585 221 -507 234
rect -585 187 -559 221
rect -559 187 -507 221
rect -585 169 -507 187
rect -442 221 -364 234
rect -442 187 -410 221
rect -410 187 -376 221
rect -376 187 -364 221
rect -442 156 -364 187
rect -299 220 -247 234
rect -299 186 -284 220
rect -284 186 -247 220
rect -299 156 -247 186
rect 80 -210 340 40
rect -299 -416 -234 -351
rect -170 -890 -30 -740
rect 2320 -1560 2590 -1320
rect -170 -2130 -30 -1990
rect 2320 -2790 2590 -2550
rect -170 -3390 -30 -3230
rect 2320 -4050 2590 -3810
rect -170 -4620 -30 -4480
rect 2320 -5270 2590 -5030
rect -170 -5780 -30 -5690
rect 2320 -6530 2590 -6290
rect -170 -6910 -30 -6810
<< metal2 >>
rect -3880 470 -3740 480
rect -3880 280 -3870 470
rect -3750 280 -3740 470
rect -3880 -7030 -3740 280
rect -3630 470 -3490 480
rect -3630 280 -3620 470
rect -3500 280 -3490 470
rect -3630 -7030 -3490 280
rect -3380 470 -3240 480
rect -3380 280 -3370 470
rect -3250 280 -3240 470
rect -3380 234 -3240 280
rect -3380 182 -3367 234
rect -3250 182 -3240 234
rect -3380 -7030 -3240 182
rect -3130 470 -2990 480
rect -3130 280 -3120 470
rect -3000 280 -2990 470
rect -3130 -7030 -2990 280
rect -2880 470 -2740 480
rect -2880 280 -2870 470
rect -2750 280 -2740 470
rect -2880 -7030 -2740 280
rect -2630 470 -2490 480
rect -2630 280 -2620 470
rect -2500 280 -2490 470
rect -2630 260 -2490 280
rect -2630 156 -2613 260
rect -2496 156 -2490 260
rect -2630 -7030 -2490 156
rect -2380 470 -2240 480
rect -2380 280 -2370 470
rect -2250 280 -2240 470
rect -2380 78 -2240 280
rect -2380 0 -2366 78
rect -2249 0 -2240 78
rect -2380 -7030 -2240 0
rect -2130 470 -1990 480
rect -2130 280 -2120 470
rect -2000 280 -1990 470
rect -2130 -7030 -1990 280
rect -1880 470 -1740 480
rect -1880 280 -1870 470
rect -1750 280 -1740 470
rect -180 420 -20 430
rect -1880 -7030 -1740 280
rect -455 390 -351 403
rect -455 325 -442 390
rect -364 325 -351 390
rect -1690 240 -1610 250
rect -1690 180 -1680 240
rect -1620 180 -1610 240
rect -1690 170 -1610 180
rect -1443 247 -1313 260
rect -1690 169 -1612 170
rect -1443 169 -1417 247
rect -1339 169 -1313 247
rect -1443 -260 -1313 169
rect -1157 247 -1027 260
rect -1157 169 -1144 247
rect -1066 169 -1027 247
rect -1157 -110 -1027 169
rect -988 247 -897 260
rect -910 169 -897 247
rect -988 156 -897 169
rect -858 247 -767 260
rect -780 169 -767 247
rect -858 -52 -767 169
rect -728 104 -637 247
rect -598 234 -494 247
rect -598 169 -585 234
rect -507 169 -494 234
rect -598 156 -494 169
rect -728 26 -715 104
rect -650 26 -637 104
rect -728 13 -637 26
rect -1450 -7030 -1310 -260
rect -1170 -7030 -1020 -110
rect -871 -250 -767 -52
rect -585 -180 -494 156
rect -455 234 -351 325
rect -180 300 -170 420
rect -30 300 -20 420
rect -180 290 -20 300
rect -455 156 -442 234
rect -364 156 -351 234
rect -455 143 -351 156
rect -312 234 -221 247
rect -312 156 -299 234
rect -247 156 -221 234
rect -890 -7030 -740 -250
rect -610 -7030 -470 -180
rect -312 -351 -221 156
rect 70 40 350 50
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect -312 -416 -299 -351
rect -234 -416 -221 -351
rect -312 -3090 -221 -416
rect -180 -740 -20 -730
rect -180 -890 -170 -740
rect -30 -890 -20 -740
rect -180 -900 -20 -890
rect 2310 -1320 2600 -1310
rect 2310 -1560 2320 -1320
rect 2590 -1560 2600 -1320
rect 2310 -1570 2600 -1560
rect -180 -1990 -20 -1980
rect -180 -2130 -170 -1990
rect -30 -2130 -20 -1990
rect -180 -2140 -20 -2130
rect 2310 -2550 2600 -2540
rect 2310 -2790 2320 -2550
rect 2590 -2790 2600 -2550
rect 2310 -2800 2600 -2790
rect -312 -3094 -220 -3090
rect -310 -7030 -220 -3094
rect -180 -3230 -20 -3220
rect -180 -3390 -170 -3230
rect -30 -3390 -20 -3230
rect -180 -3400 -20 -3390
rect 2310 -3810 2600 -3800
rect 2310 -4050 2320 -3810
rect 2590 -4050 2600 -3810
rect 2310 -4060 2600 -4050
rect -180 -4480 -20 -4470
rect -180 -4620 -170 -4480
rect -30 -4620 -20 -4480
rect -180 -4630 -20 -4620
rect 2310 -5030 2600 -5020
rect 2310 -5270 2320 -5030
rect 2590 -5270 2600 -5030
rect 2310 -5280 2600 -5270
rect -180 -5690 -20 -5680
rect -180 -5780 -170 -5690
rect -30 -5780 -20 -5690
rect -180 -5790 -20 -5780
rect 2310 -6290 2600 -6280
rect 2310 -6530 2320 -6290
rect 2590 -6530 2600 -6290
rect 2310 -6540 2600 -6530
rect -180 -6810 -20 -6800
rect -180 -6910 -170 -6810
rect -30 -6910 -20 -6810
rect -180 -6920 -20 -6910
<< via2 >>
rect -2613 156 -2496 260
rect -2366 0 -2249 78
rect -1859 338 -1768 403
rect -442 325 -364 390
rect -988 169 -923 247
rect -923 169 -910 247
rect -715 26 -650 104
rect -170 300 -30 420
rect 80 -210 340 40
rect -170 -890 -30 -740
rect 2320 -1560 2590 -1320
rect -170 -2130 -30 -1990
rect 2320 -2790 2590 -2550
rect -170 -3390 -30 -3230
rect 2320 -4050 2590 -3810
rect -170 -4620 -30 -4480
rect 2320 -5270 2590 -5030
rect -170 -5780 -30 -5690
rect 2320 -6530 2590 -6290
rect -170 -6910 -30 -6810
<< metal3 >>
rect -190 430 -10 440
rect -1890 403 -1710 420
rect -1890 338 -1859 403
rect -1768 390 -1710 403
rect -455 390 -351 403
rect -1768 338 -442 390
rect -1890 325 -442 338
rect -364 325 -351 390
rect -1890 320 -351 325
rect -455 312 -351 320
rect -190 290 -180 430
rect -20 290 -10 430
rect -190 280 -10 290
rect -2639 260 -2470 273
rect -2639 156 -2613 260
rect -2496 247 -897 260
rect -2496 169 -988 247
rect -910 169 -897 247
rect -2496 156 -897 169
rect -2639 143 -2470 156
rect -728 104 -637 117
rect -728 91 -715 104
rect -2379 78 -715 91
rect -2379 0 -2366 78
rect -2249 26 -715 78
rect -650 26 -637 104
rect -2249 13 -637 26
rect 70 40 350 50
rect -2249 0 -2236 13
rect -2379 -13 -2236 0
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect -180 -740 -20 -730
rect -180 -890 -170 -740
rect -30 -890 -20 -740
rect -180 -900 -20 -890
rect 2310 -1320 2600 -1310
rect 2310 -1560 2320 -1320
rect 2590 -1560 2600 -1320
rect 2310 -1570 2600 -1560
rect -180 -1990 -20 -1980
rect -180 -2130 -170 -1990
rect -30 -2130 -20 -1990
rect -180 -2140 -20 -2130
rect 2310 -2550 2600 -2540
rect 2310 -2790 2320 -2550
rect 2590 -2790 2600 -2550
rect 2310 -2800 2600 -2790
rect -180 -3230 -20 -3220
rect -180 -3390 -170 -3230
rect -30 -3390 -20 -3230
rect -180 -3400 -20 -3390
rect 2310 -3810 2600 -3800
rect 2310 -4050 2320 -3810
rect 2590 -4050 2600 -3810
rect 2310 -4060 2600 -4050
rect -180 -4480 -20 -4470
rect -180 -4620 -170 -4480
rect -30 -4620 -20 -4480
rect -180 -4630 -20 -4620
rect 2310 -5030 2600 -5020
rect 2310 -5270 2320 -5030
rect 2590 -5270 2600 -5030
rect 2310 -5280 2600 -5270
rect -180 -5690 -20 -5680
rect -180 -5780 -170 -5690
rect -30 -5780 -20 -5690
rect -180 -5790 -20 -5780
rect 2310 -6290 2600 -6280
rect 2310 -6530 2320 -6290
rect 2590 -6530 2600 -6290
rect 2310 -6540 2600 -6530
rect -180 -6810 -20 -6800
rect -180 -6910 -170 -6810
rect -30 -6910 -20 -6810
rect -180 -6920 -20 -6910
<< via3 >>
rect -180 420 -20 430
rect -180 300 -170 420
rect -170 300 -30 420
rect -30 300 -20 420
rect -180 290 -20 300
rect 80 -210 340 40
rect -170 -890 -30 -740
rect 2320 -1560 2590 -1320
rect -170 -2130 -30 -1990
rect 2320 -2790 2590 -2550
rect -170 -3390 -30 -3230
rect 2320 -4050 2590 -3810
rect -170 -4620 -30 -4480
rect 2320 -5270 2590 -5030
rect -170 -5780 -30 -5690
rect 2320 -6530 2590 -6290
rect -170 -6910 -30 -6810
<< metal4 >>
rect -190 430 -10 700
rect -190 290 -180 430
rect -20 290 -10 430
rect -190 -740 -10 290
rect 70 40 350 50
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect -190 -890 -170 -740
rect -30 -890 -10 -740
rect -190 -1990 -10 -890
rect 2310 -1320 2600 -1310
rect 2310 -1560 2320 -1320
rect 2590 -1560 2600 -1320
rect 2310 -1570 2600 -1560
rect -190 -2130 -170 -1990
rect -30 -2130 -10 -1990
rect -190 -3230 -10 -2130
rect 2310 -2550 2600 -2540
rect 2310 -2790 2320 -2550
rect 2590 -2790 2600 -2550
rect 2310 -2800 2600 -2790
rect -190 -3390 -170 -3230
rect -30 -3390 -10 -3230
rect -190 -4480 -10 -3390
rect 2310 -3810 2600 -3800
rect 2310 -4050 2320 -3810
rect 2590 -4050 2600 -3810
rect 2310 -4060 2600 -4050
rect -190 -4620 -170 -4480
rect -30 -4620 -10 -4480
rect -190 -5690 -10 -4620
rect 2310 -5030 2600 -5020
rect 2310 -5270 2320 -5030
rect 2590 -5270 2600 -5030
rect 2310 -5280 2600 -5270
rect -190 -5780 -170 -5690
rect -30 -5780 -10 -5690
rect -190 -6810 -10 -5780
rect 2310 -6290 2600 -6280
rect 2310 -6530 2320 -6290
rect 2590 -6530 2600 -6290
rect 2310 -6540 2600 -6530
rect -190 -6910 -170 -6810
rect -30 -6910 -10 -6810
rect -190 -7030 -10 -6910
<< via4 >>
rect 80 -210 340 40
rect 2320 -1560 2590 -1320
rect 2320 -2790 2590 -2550
rect 2320 -4050 2590 -3810
rect 2320 -5270 2590 -5030
rect 2320 -6530 2590 -6290
<< metal5 >>
rect 2290 70 2620 700
rect -1590 40 2620 70
rect -1590 -210 80 40
rect 340 -210 2620 40
rect -1590 -250 2620 -210
rect 2290 -1320 2620 -250
rect 2290 -1560 2320 -1320
rect 2590 -1560 2620 -1320
rect 2290 -2550 2620 -1560
rect 2290 -2790 2320 -2550
rect 2590 -2790 2620 -2550
rect 2290 -3810 2620 -2790
rect 2290 -4050 2320 -3810
rect 2590 -4050 2620 -3810
rect 2290 -5030 2620 -4050
rect 2290 -5270 2320 -5030
rect 2590 -5270 2620 -5030
rect 2290 -6290 2620 -5270
rect 2290 -6530 2320 -6290
rect 2590 -6530 2620 -6290
rect 2290 -6560 2620 -6530
use sky130_fd_sc_hd__or4_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 488 0 1 -772
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  x2
timestamp 1701704242
transform 1 0 488 0 -1 -858
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 -758 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1040 0 1 -772
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1701704242
transform 1 0 -1034 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1701704242
transform 1 0 -1308 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1701704242
transform 1 0 -1584 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1500 0 1 -772
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1701704242
transform 1 0 -482 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x10
timestamp 1701704242
transform 1 0 488 0 1 -2022
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x11
timestamp 1701704242
transform 1 0 488 0 -1 -2098
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x12
timestamp 1701704242
transform 1 0 488 0 1 -3262
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x13
timestamp 1701704242
transform 1 0 490 0 -1 -3352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x14
timestamp 1701704242
transform 1 0 948 0 -1 -2098
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 488 0 1 -4512
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x16
timestamp 1701704242
transform 1 0 488 0 -1 -4584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  x17
timestamp 1701704242
transform 1 0 1132 0 1 -4512
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x18
timestamp 1701704242
transform 1 0 488 0 1 -5744
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x19
timestamp 1701704242
transform 1 0 488 0 -1 -5818
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 488 0 1 -6982
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x21
timestamp 1701704242
transform 1 0 948 0 1 -6982
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x22
timestamp 1701704242
transform -1 0 1960 0 1 -6982
box -38 -48 590 592
<< labels >>
flabel metal1 -3910 490 -3710 690 0 FreeSans 256 0 0 0 I0
port 3 nsew
flabel metal1 -3660 490 -3460 690 0 FreeSans 256 0 0 0 I1
port 0 nsew
flabel metal1 -3410 490 -3210 690 0 FreeSans 256 0 0 0 I2
port 4 nsew
flabel metal1 -3160 490 -2960 690 0 FreeSans 256 0 0 0 I3
port 2 nsew
flabel metal1 -2910 490 -2710 690 0 FreeSans 256 0 0 0 I4
port 7 nsew
flabel metal1 -2660 490 -2460 690 0 FreeSans 256 0 0 0 I5
port 1 nsew
flabel metal1 -2410 490 -2210 690 0 FreeSans 256 0 0 0 I6
port 5 nsew
flabel metal1 -2160 490 -1960 690 0 FreeSans 256 0 0 0 I7
port 6 nsew
flabel metal1 -1910 490 -1710 690 0 FreeSans 256 0 0 0 EI
port 13 nsew
flabel metal1 3010 -4190 3210 -3990 0 FreeSans 256 0 0 0 A1
port 11 nsew
flabel metal1 3010 -3790 3210 -3590 0 FreeSans 256 0 0 0 A2
port 10 nsew
flabel metal1 3010 -2990 3210 -2790 0 FreeSans 256 0 0 0 EO
port 8 nsew
flabel metal1 3010 -3390 3210 -3190 0 FreeSans 256 0 0 0 GS
port 9 nsew
<< end >>
