magic
tech sky130A
magscale 1 2
timestamp 1713140669
<< pwell >>
rect -325 -460 325 460
<< nmos >>
rect -129 -250 -29 250
rect 29 -250 129 250
<< ndiff >>
rect -187 238 -129 250
rect -187 -238 -175 238
rect -141 -238 -129 238
rect -187 -250 -129 -238
rect -29 238 29 250
rect -29 -238 -17 238
rect 17 -238 29 238
rect -29 -250 29 -238
rect 129 238 187 250
rect 129 -238 141 238
rect 175 -238 187 238
rect 129 -250 187 -238
<< ndiffc >>
rect -175 -238 -141 238
rect -17 -238 17 238
rect 141 -238 175 238
<< psubdiff >>
rect -289 390 -193 424
rect 193 390 289 424
rect -289 328 -255 390
rect 255 328 289 390
rect -289 -390 -255 -328
rect 255 -390 289 -328
rect -289 -424 -193 -390
rect 193 -424 289 -390
<< psubdiffcont >>
rect -193 390 193 424
rect -289 -328 -255 328
rect 255 -328 289 328
rect -193 -424 193 -390
<< poly >>
rect -129 322 -29 338
rect -129 288 -113 322
rect -45 288 -29 322
rect -129 250 -29 288
rect 29 322 129 338
rect 29 288 45 322
rect 113 288 129 322
rect 29 250 129 288
rect -129 -288 -29 -250
rect -129 -322 -113 -288
rect -45 -322 -29 -288
rect -129 -338 -29 -322
rect 29 -288 129 -250
rect 29 -322 45 -288
rect 113 -322 129 -288
rect 29 -338 129 -322
<< polycont >>
rect -113 288 -45 322
rect 45 288 113 322
rect -113 -322 -45 -288
rect 45 -322 113 -288
<< locali >>
rect -289 390 -193 424
rect 193 390 289 424
rect -289 328 -255 390
rect 255 328 289 390
rect -129 288 -113 322
rect -45 288 -29 322
rect 29 288 45 322
rect 113 288 129 322
rect -175 238 -141 254
rect -175 -254 -141 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 141 238 175 254
rect 141 -254 175 -238
rect -129 -322 -113 -288
rect -45 -322 -29 -288
rect 29 -322 45 -288
rect 113 -322 129 -288
rect -289 -390 -255 -328
rect 255 -390 289 -328
rect -289 -424 -193 -390
rect 193 -424 289 -390
<< viali >>
rect -113 288 -45 322
rect 45 288 113 322
rect -175 -238 -141 238
rect -17 -238 17 238
rect 141 -238 175 238
rect -113 -322 -45 -288
rect 45 -322 113 -288
<< metal1 >>
rect -125 322 -33 328
rect -125 288 -113 322
rect -45 288 -33 322
rect -125 282 -33 288
rect 33 322 125 328
rect 33 288 45 322
rect 113 288 125 322
rect 33 282 125 288
rect -181 238 -135 250
rect -181 -238 -175 238
rect -141 -238 -135 238
rect -181 -250 -135 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 135 238 181 250
rect 135 -238 141 238
rect 175 -238 181 238
rect 135 -250 181 -238
rect -125 -288 -33 -282
rect -125 -322 -113 -288
rect -45 -322 -33 -288
rect -125 -328 -33 -322
rect 33 -288 125 -282
rect 33 -322 45 -288
rect 113 -322 125 -288
rect 33 -328 125 -322
<< properties >>
string FIXED_BBOX -272 -407 272 407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
