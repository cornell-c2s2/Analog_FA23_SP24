magic
tech sky130A
magscale 1 2
timestamp 1714792946
<< pwell >>
rect -5086 -18510 5086 18510
<< psubdiff >>
rect -5050 18440 -4954 18474
rect 4954 18440 5050 18474
rect -5050 18378 -5016 18440
rect 5016 18378 5050 18440
rect -5050 -18440 -5016 -18378
rect 5016 -18440 5050 -18378
rect -5050 -18474 -4954 -18440
rect 4954 -18474 5050 -18440
<< psubdiffcont >>
rect -4954 18440 4954 18474
rect -5050 -18378 -5016 18378
rect 5016 -18378 5050 18378
rect -4954 -18474 4954 -18440
<< xpolycontact >>
rect -4920 17912 -3774 18344
rect -4920 16404 -3774 16836
rect -3678 17912 -2532 18344
rect -3678 16404 -2532 16836
rect -2436 17912 -1290 18344
rect -2436 16404 -1290 16836
rect -1194 17912 -48 18344
rect -1194 16404 -48 16836
rect 48 17912 1194 18344
rect 48 16404 1194 16836
rect 1290 17912 2436 18344
rect 1290 16404 2436 16836
rect 2532 17912 3678 18344
rect 2532 16404 3678 16836
rect 3774 17912 4920 18344
rect 3774 16404 4920 16836
rect -4920 15868 -3774 16300
rect -4920 14360 -3774 14792
rect -3678 15868 -2532 16300
rect -3678 14360 -2532 14792
rect -2436 15868 -1290 16300
rect -2436 14360 -1290 14792
rect -1194 15868 -48 16300
rect -1194 14360 -48 14792
rect 48 15868 1194 16300
rect 48 14360 1194 14792
rect 1290 15868 2436 16300
rect 1290 14360 2436 14792
rect 2532 15868 3678 16300
rect 2532 14360 3678 14792
rect 3774 15868 4920 16300
rect 3774 14360 4920 14792
rect -4920 13824 -3774 14256
rect -4920 12316 -3774 12748
rect -3678 13824 -2532 14256
rect -3678 12316 -2532 12748
rect -2436 13824 -1290 14256
rect -2436 12316 -1290 12748
rect -1194 13824 -48 14256
rect -1194 12316 -48 12748
rect 48 13824 1194 14256
rect 48 12316 1194 12748
rect 1290 13824 2436 14256
rect 1290 12316 2436 12748
rect 2532 13824 3678 14256
rect 2532 12316 3678 12748
rect 3774 13824 4920 14256
rect 3774 12316 4920 12748
rect -4920 11780 -3774 12212
rect -4920 10272 -3774 10704
rect -3678 11780 -2532 12212
rect -3678 10272 -2532 10704
rect -2436 11780 -1290 12212
rect -2436 10272 -1290 10704
rect -1194 11780 -48 12212
rect -1194 10272 -48 10704
rect 48 11780 1194 12212
rect 48 10272 1194 10704
rect 1290 11780 2436 12212
rect 1290 10272 2436 10704
rect 2532 11780 3678 12212
rect 2532 10272 3678 10704
rect 3774 11780 4920 12212
rect 3774 10272 4920 10704
rect -4920 9736 -3774 10168
rect -4920 8228 -3774 8660
rect -3678 9736 -2532 10168
rect -3678 8228 -2532 8660
rect -2436 9736 -1290 10168
rect -2436 8228 -1290 8660
rect -1194 9736 -48 10168
rect -1194 8228 -48 8660
rect 48 9736 1194 10168
rect 48 8228 1194 8660
rect 1290 9736 2436 10168
rect 1290 8228 2436 8660
rect 2532 9736 3678 10168
rect 2532 8228 3678 8660
rect 3774 9736 4920 10168
rect 3774 8228 4920 8660
rect -4920 7692 -3774 8124
rect -4920 6184 -3774 6616
rect -3678 7692 -2532 8124
rect -3678 6184 -2532 6616
rect -2436 7692 -1290 8124
rect -2436 6184 -1290 6616
rect -1194 7692 -48 8124
rect -1194 6184 -48 6616
rect 48 7692 1194 8124
rect 48 6184 1194 6616
rect 1290 7692 2436 8124
rect 1290 6184 2436 6616
rect 2532 7692 3678 8124
rect 2532 6184 3678 6616
rect 3774 7692 4920 8124
rect 3774 6184 4920 6616
rect -4920 5648 -3774 6080
rect -4920 4140 -3774 4572
rect -3678 5648 -2532 6080
rect -3678 4140 -2532 4572
rect -2436 5648 -1290 6080
rect -2436 4140 -1290 4572
rect -1194 5648 -48 6080
rect -1194 4140 -48 4572
rect 48 5648 1194 6080
rect 48 4140 1194 4572
rect 1290 5648 2436 6080
rect 1290 4140 2436 4572
rect 2532 5648 3678 6080
rect 2532 4140 3678 4572
rect 3774 5648 4920 6080
rect 3774 4140 4920 4572
rect -4920 3604 -3774 4036
rect -4920 2096 -3774 2528
rect -3678 3604 -2532 4036
rect -3678 2096 -2532 2528
rect -2436 3604 -1290 4036
rect -2436 2096 -1290 2528
rect -1194 3604 -48 4036
rect -1194 2096 -48 2528
rect 48 3604 1194 4036
rect 48 2096 1194 2528
rect 1290 3604 2436 4036
rect 1290 2096 2436 2528
rect 2532 3604 3678 4036
rect 2532 2096 3678 2528
rect 3774 3604 4920 4036
rect 3774 2096 4920 2528
rect -4920 1560 -3774 1992
rect -4920 52 -3774 484
rect -3678 1560 -2532 1992
rect -3678 52 -2532 484
rect -2436 1560 -1290 1992
rect -2436 52 -1290 484
rect -1194 1560 -48 1992
rect -1194 52 -48 484
rect 48 1560 1194 1992
rect 48 52 1194 484
rect 1290 1560 2436 1992
rect 1290 52 2436 484
rect 2532 1560 3678 1992
rect 2532 52 3678 484
rect 3774 1560 4920 1992
rect 3774 52 4920 484
rect -4920 -484 -3774 -52
rect -4920 -1992 -3774 -1560
rect -3678 -484 -2532 -52
rect -3678 -1992 -2532 -1560
rect -2436 -484 -1290 -52
rect -2436 -1992 -1290 -1560
rect -1194 -484 -48 -52
rect -1194 -1992 -48 -1560
rect 48 -484 1194 -52
rect 48 -1992 1194 -1560
rect 1290 -484 2436 -52
rect 1290 -1992 2436 -1560
rect 2532 -484 3678 -52
rect 2532 -1992 3678 -1560
rect 3774 -484 4920 -52
rect 3774 -1992 4920 -1560
rect -4920 -2528 -3774 -2096
rect -4920 -4036 -3774 -3604
rect -3678 -2528 -2532 -2096
rect -3678 -4036 -2532 -3604
rect -2436 -2528 -1290 -2096
rect -2436 -4036 -1290 -3604
rect -1194 -2528 -48 -2096
rect -1194 -4036 -48 -3604
rect 48 -2528 1194 -2096
rect 48 -4036 1194 -3604
rect 1290 -2528 2436 -2096
rect 1290 -4036 2436 -3604
rect 2532 -2528 3678 -2096
rect 2532 -4036 3678 -3604
rect 3774 -2528 4920 -2096
rect 3774 -4036 4920 -3604
rect -4920 -4572 -3774 -4140
rect -4920 -6080 -3774 -5648
rect -3678 -4572 -2532 -4140
rect -3678 -6080 -2532 -5648
rect -2436 -4572 -1290 -4140
rect -2436 -6080 -1290 -5648
rect -1194 -4572 -48 -4140
rect -1194 -6080 -48 -5648
rect 48 -4572 1194 -4140
rect 48 -6080 1194 -5648
rect 1290 -4572 2436 -4140
rect 1290 -6080 2436 -5648
rect 2532 -4572 3678 -4140
rect 2532 -6080 3678 -5648
rect 3774 -4572 4920 -4140
rect 3774 -6080 4920 -5648
rect -4920 -6616 -3774 -6184
rect -4920 -8124 -3774 -7692
rect -3678 -6616 -2532 -6184
rect -3678 -8124 -2532 -7692
rect -2436 -6616 -1290 -6184
rect -2436 -8124 -1290 -7692
rect -1194 -6616 -48 -6184
rect -1194 -8124 -48 -7692
rect 48 -6616 1194 -6184
rect 48 -8124 1194 -7692
rect 1290 -6616 2436 -6184
rect 1290 -8124 2436 -7692
rect 2532 -6616 3678 -6184
rect 2532 -8124 3678 -7692
rect 3774 -6616 4920 -6184
rect 3774 -8124 4920 -7692
rect -4920 -8660 -3774 -8228
rect -4920 -10168 -3774 -9736
rect -3678 -8660 -2532 -8228
rect -3678 -10168 -2532 -9736
rect -2436 -8660 -1290 -8228
rect -2436 -10168 -1290 -9736
rect -1194 -8660 -48 -8228
rect -1194 -10168 -48 -9736
rect 48 -8660 1194 -8228
rect 48 -10168 1194 -9736
rect 1290 -8660 2436 -8228
rect 1290 -10168 2436 -9736
rect 2532 -8660 3678 -8228
rect 2532 -10168 3678 -9736
rect 3774 -8660 4920 -8228
rect 3774 -10168 4920 -9736
rect -4920 -10704 -3774 -10272
rect -4920 -12212 -3774 -11780
rect -3678 -10704 -2532 -10272
rect -3678 -12212 -2532 -11780
rect -2436 -10704 -1290 -10272
rect -2436 -12212 -1290 -11780
rect -1194 -10704 -48 -10272
rect -1194 -12212 -48 -11780
rect 48 -10704 1194 -10272
rect 48 -12212 1194 -11780
rect 1290 -10704 2436 -10272
rect 1290 -12212 2436 -11780
rect 2532 -10704 3678 -10272
rect 2532 -12212 3678 -11780
rect 3774 -10704 4920 -10272
rect 3774 -12212 4920 -11780
rect -4920 -12748 -3774 -12316
rect -4920 -14256 -3774 -13824
rect -3678 -12748 -2532 -12316
rect -3678 -14256 -2532 -13824
rect -2436 -12748 -1290 -12316
rect -2436 -14256 -1290 -13824
rect -1194 -12748 -48 -12316
rect -1194 -14256 -48 -13824
rect 48 -12748 1194 -12316
rect 48 -14256 1194 -13824
rect 1290 -12748 2436 -12316
rect 1290 -14256 2436 -13824
rect 2532 -12748 3678 -12316
rect 2532 -14256 3678 -13824
rect 3774 -12748 4920 -12316
rect 3774 -14256 4920 -13824
rect -4920 -14792 -3774 -14360
rect -4920 -16300 -3774 -15868
rect -3678 -14792 -2532 -14360
rect -3678 -16300 -2532 -15868
rect -2436 -14792 -1290 -14360
rect -2436 -16300 -1290 -15868
rect -1194 -14792 -48 -14360
rect -1194 -16300 -48 -15868
rect 48 -14792 1194 -14360
rect 48 -16300 1194 -15868
rect 1290 -14792 2436 -14360
rect 1290 -16300 2436 -15868
rect 2532 -14792 3678 -14360
rect 2532 -16300 3678 -15868
rect 3774 -14792 4920 -14360
rect 3774 -16300 4920 -15868
rect -4920 -16836 -3774 -16404
rect -4920 -18344 -3774 -17912
rect -3678 -16836 -2532 -16404
rect -3678 -18344 -2532 -17912
rect -2436 -16836 -1290 -16404
rect -2436 -18344 -1290 -17912
rect -1194 -16836 -48 -16404
rect -1194 -18344 -48 -17912
rect 48 -16836 1194 -16404
rect 48 -18344 1194 -17912
rect 1290 -16836 2436 -16404
rect 1290 -18344 2436 -17912
rect 2532 -16836 3678 -16404
rect 2532 -18344 3678 -17912
rect 3774 -16836 4920 -16404
rect 3774 -18344 4920 -17912
<< xpolyres >>
rect -4920 16836 -3774 17912
rect -3678 16836 -2532 17912
rect -2436 16836 -1290 17912
rect -1194 16836 -48 17912
rect 48 16836 1194 17912
rect 1290 16836 2436 17912
rect 2532 16836 3678 17912
rect 3774 16836 4920 17912
rect -4920 14792 -3774 15868
rect -3678 14792 -2532 15868
rect -2436 14792 -1290 15868
rect -1194 14792 -48 15868
rect 48 14792 1194 15868
rect 1290 14792 2436 15868
rect 2532 14792 3678 15868
rect 3774 14792 4920 15868
rect -4920 12748 -3774 13824
rect -3678 12748 -2532 13824
rect -2436 12748 -1290 13824
rect -1194 12748 -48 13824
rect 48 12748 1194 13824
rect 1290 12748 2436 13824
rect 2532 12748 3678 13824
rect 3774 12748 4920 13824
rect -4920 10704 -3774 11780
rect -3678 10704 -2532 11780
rect -2436 10704 -1290 11780
rect -1194 10704 -48 11780
rect 48 10704 1194 11780
rect 1290 10704 2436 11780
rect 2532 10704 3678 11780
rect 3774 10704 4920 11780
rect -4920 8660 -3774 9736
rect -3678 8660 -2532 9736
rect -2436 8660 -1290 9736
rect -1194 8660 -48 9736
rect 48 8660 1194 9736
rect 1290 8660 2436 9736
rect 2532 8660 3678 9736
rect 3774 8660 4920 9736
rect -4920 6616 -3774 7692
rect -3678 6616 -2532 7692
rect -2436 6616 -1290 7692
rect -1194 6616 -48 7692
rect 48 6616 1194 7692
rect 1290 6616 2436 7692
rect 2532 6616 3678 7692
rect 3774 6616 4920 7692
rect -4920 4572 -3774 5648
rect -3678 4572 -2532 5648
rect -2436 4572 -1290 5648
rect -1194 4572 -48 5648
rect 48 4572 1194 5648
rect 1290 4572 2436 5648
rect 2532 4572 3678 5648
rect 3774 4572 4920 5648
rect -4920 2528 -3774 3604
rect -3678 2528 -2532 3604
rect -2436 2528 -1290 3604
rect -1194 2528 -48 3604
rect 48 2528 1194 3604
rect 1290 2528 2436 3604
rect 2532 2528 3678 3604
rect 3774 2528 4920 3604
rect -4920 484 -3774 1560
rect -3678 484 -2532 1560
rect -2436 484 -1290 1560
rect -1194 484 -48 1560
rect 48 484 1194 1560
rect 1290 484 2436 1560
rect 2532 484 3678 1560
rect 3774 484 4920 1560
rect -4920 -1560 -3774 -484
rect -3678 -1560 -2532 -484
rect -2436 -1560 -1290 -484
rect -1194 -1560 -48 -484
rect 48 -1560 1194 -484
rect 1290 -1560 2436 -484
rect 2532 -1560 3678 -484
rect 3774 -1560 4920 -484
rect -4920 -3604 -3774 -2528
rect -3678 -3604 -2532 -2528
rect -2436 -3604 -1290 -2528
rect -1194 -3604 -48 -2528
rect 48 -3604 1194 -2528
rect 1290 -3604 2436 -2528
rect 2532 -3604 3678 -2528
rect 3774 -3604 4920 -2528
rect -4920 -5648 -3774 -4572
rect -3678 -5648 -2532 -4572
rect -2436 -5648 -1290 -4572
rect -1194 -5648 -48 -4572
rect 48 -5648 1194 -4572
rect 1290 -5648 2436 -4572
rect 2532 -5648 3678 -4572
rect 3774 -5648 4920 -4572
rect -4920 -7692 -3774 -6616
rect -3678 -7692 -2532 -6616
rect -2436 -7692 -1290 -6616
rect -1194 -7692 -48 -6616
rect 48 -7692 1194 -6616
rect 1290 -7692 2436 -6616
rect 2532 -7692 3678 -6616
rect 3774 -7692 4920 -6616
rect -4920 -9736 -3774 -8660
rect -3678 -9736 -2532 -8660
rect -2436 -9736 -1290 -8660
rect -1194 -9736 -48 -8660
rect 48 -9736 1194 -8660
rect 1290 -9736 2436 -8660
rect 2532 -9736 3678 -8660
rect 3774 -9736 4920 -8660
rect -4920 -11780 -3774 -10704
rect -3678 -11780 -2532 -10704
rect -2436 -11780 -1290 -10704
rect -1194 -11780 -48 -10704
rect 48 -11780 1194 -10704
rect 1290 -11780 2436 -10704
rect 2532 -11780 3678 -10704
rect 3774 -11780 4920 -10704
rect -4920 -13824 -3774 -12748
rect -3678 -13824 -2532 -12748
rect -2436 -13824 -1290 -12748
rect -1194 -13824 -48 -12748
rect 48 -13824 1194 -12748
rect 1290 -13824 2436 -12748
rect 2532 -13824 3678 -12748
rect 3774 -13824 4920 -12748
rect -4920 -15868 -3774 -14792
rect -3678 -15868 -2532 -14792
rect -2436 -15868 -1290 -14792
rect -1194 -15868 -48 -14792
rect 48 -15868 1194 -14792
rect 1290 -15868 2436 -14792
rect 2532 -15868 3678 -14792
rect 3774 -15868 4920 -14792
rect -4920 -17912 -3774 -16836
rect -3678 -17912 -2532 -16836
rect -2436 -17912 -1290 -16836
rect -1194 -17912 -48 -16836
rect 48 -17912 1194 -16836
rect 1290 -17912 2436 -16836
rect 2532 -17912 3678 -16836
rect 3774 -17912 4920 -16836
<< locali >>
rect -5050 18440 -4954 18474
rect 4954 18440 5050 18474
rect -5050 18378 -5016 18440
rect 5016 18378 5050 18440
rect -5050 -18440 -5016 -18378
rect 5016 -18440 5050 -18378
rect -5050 -18474 -4954 -18440
rect 4954 -18474 5050 -18440
<< viali >>
rect -4904 17929 -3790 18326
rect -3662 17929 -2548 18326
rect -2420 17929 -1306 18326
rect -1178 17929 -64 18326
rect 64 17929 1178 18326
rect 1306 17929 2420 18326
rect 2548 17929 3662 18326
rect 3790 17929 4904 18326
rect -4904 16422 -3790 16819
rect -3662 16422 -2548 16819
rect -2420 16422 -1306 16819
rect -1178 16422 -64 16819
rect 64 16422 1178 16819
rect 1306 16422 2420 16819
rect 2548 16422 3662 16819
rect 3790 16422 4904 16819
rect -4904 15885 -3790 16282
rect -3662 15885 -2548 16282
rect -2420 15885 -1306 16282
rect -1178 15885 -64 16282
rect 64 15885 1178 16282
rect 1306 15885 2420 16282
rect 2548 15885 3662 16282
rect 3790 15885 4904 16282
rect -4904 14378 -3790 14775
rect -3662 14378 -2548 14775
rect -2420 14378 -1306 14775
rect -1178 14378 -64 14775
rect 64 14378 1178 14775
rect 1306 14378 2420 14775
rect 2548 14378 3662 14775
rect 3790 14378 4904 14775
rect -4904 13841 -3790 14238
rect -3662 13841 -2548 14238
rect -2420 13841 -1306 14238
rect -1178 13841 -64 14238
rect 64 13841 1178 14238
rect 1306 13841 2420 14238
rect 2548 13841 3662 14238
rect 3790 13841 4904 14238
rect -4904 12334 -3790 12731
rect -3662 12334 -2548 12731
rect -2420 12334 -1306 12731
rect -1178 12334 -64 12731
rect 64 12334 1178 12731
rect 1306 12334 2420 12731
rect 2548 12334 3662 12731
rect 3790 12334 4904 12731
rect -4904 11797 -3790 12194
rect -3662 11797 -2548 12194
rect -2420 11797 -1306 12194
rect -1178 11797 -64 12194
rect 64 11797 1178 12194
rect 1306 11797 2420 12194
rect 2548 11797 3662 12194
rect 3790 11797 4904 12194
rect -4904 10290 -3790 10687
rect -3662 10290 -2548 10687
rect -2420 10290 -1306 10687
rect -1178 10290 -64 10687
rect 64 10290 1178 10687
rect 1306 10290 2420 10687
rect 2548 10290 3662 10687
rect 3790 10290 4904 10687
rect -4904 9753 -3790 10150
rect -3662 9753 -2548 10150
rect -2420 9753 -1306 10150
rect -1178 9753 -64 10150
rect 64 9753 1178 10150
rect 1306 9753 2420 10150
rect 2548 9753 3662 10150
rect 3790 9753 4904 10150
rect -4904 8246 -3790 8643
rect -3662 8246 -2548 8643
rect -2420 8246 -1306 8643
rect -1178 8246 -64 8643
rect 64 8246 1178 8643
rect 1306 8246 2420 8643
rect 2548 8246 3662 8643
rect 3790 8246 4904 8643
rect -4904 7709 -3790 8106
rect -3662 7709 -2548 8106
rect -2420 7709 -1306 8106
rect -1178 7709 -64 8106
rect 64 7709 1178 8106
rect 1306 7709 2420 8106
rect 2548 7709 3662 8106
rect 3790 7709 4904 8106
rect -4904 6202 -3790 6599
rect -3662 6202 -2548 6599
rect -2420 6202 -1306 6599
rect -1178 6202 -64 6599
rect 64 6202 1178 6599
rect 1306 6202 2420 6599
rect 2548 6202 3662 6599
rect 3790 6202 4904 6599
rect -4904 5665 -3790 6062
rect -3662 5665 -2548 6062
rect -2420 5665 -1306 6062
rect -1178 5665 -64 6062
rect 64 5665 1178 6062
rect 1306 5665 2420 6062
rect 2548 5665 3662 6062
rect 3790 5665 4904 6062
rect -4904 4158 -3790 4555
rect -3662 4158 -2548 4555
rect -2420 4158 -1306 4555
rect -1178 4158 -64 4555
rect 64 4158 1178 4555
rect 1306 4158 2420 4555
rect 2548 4158 3662 4555
rect 3790 4158 4904 4555
rect -4904 3621 -3790 4018
rect -3662 3621 -2548 4018
rect -2420 3621 -1306 4018
rect -1178 3621 -64 4018
rect 64 3621 1178 4018
rect 1306 3621 2420 4018
rect 2548 3621 3662 4018
rect 3790 3621 4904 4018
rect -4904 2114 -3790 2511
rect -3662 2114 -2548 2511
rect -2420 2114 -1306 2511
rect -1178 2114 -64 2511
rect 64 2114 1178 2511
rect 1306 2114 2420 2511
rect 2548 2114 3662 2511
rect 3790 2114 4904 2511
rect -4904 1577 -3790 1974
rect -3662 1577 -2548 1974
rect -2420 1577 -1306 1974
rect -1178 1577 -64 1974
rect 64 1577 1178 1974
rect 1306 1577 2420 1974
rect 2548 1577 3662 1974
rect 3790 1577 4904 1974
rect -4904 70 -3790 467
rect -3662 70 -2548 467
rect -2420 70 -1306 467
rect -1178 70 -64 467
rect 64 70 1178 467
rect 1306 70 2420 467
rect 2548 70 3662 467
rect 3790 70 4904 467
rect -4904 -467 -3790 -70
rect -3662 -467 -2548 -70
rect -2420 -467 -1306 -70
rect -1178 -467 -64 -70
rect 64 -467 1178 -70
rect 1306 -467 2420 -70
rect 2548 -467 3662 -70
rect 3790 -467 4904 -70
rect -4904 -1974 -3790 -1577
rect -3662 -1974 -2548 -1577
rect -2420 -1974 -1306 -1577
rect -1178 -1974 -64 -1577
rect 64 -1974 1178 -1577
rect 1306 -1974 2420 -1577
rect 2548 -1974 3662 -1577
rect 3790 -1974 4904 -1577
rect -4904 -2511 -3790 -2114
rect -3662 -2511 -2548 -2114
rect -2420 -2511 -1306 -2114
rect -1178 -2511 -64 -2114
rect 64 -2511 1178 -2114
rect 1306 -2511 2420 -2114
rect 2548 -2511 3662 -2114
rect 3790 -2511 4904 -2114
rect -4904 -4018 -3790 -3621
rect -3662 -4018 -2548 -3621
rect -2420 -4018 -1306 -3621
rect -1178 -4018 -64 -3621
rect 64 -4018 1178 -3621
rect 1306 -4018 2420 -3621
rect 2548 -4018 3662 -3621
rect 3790 -4018 4904 -3621
rect -4904 -4555 -3790 -4158
rect -3662 -4555 -2548 -4158
rect -2420 -4555 -1306 -4158
rect -1178 -4555 -64 -4158
rect 64 -4555 1178 -4158
rect 1306 -4555 2420 -4158
rect 2548 -4555 3662 -4158
rect 3790 -4555 4904 -4158
rect -4904 -6062 -3790 -5665
rect -3662 -6062 -2548 -5665
rect -2420 -6062 -1306 -5665
rect -1178 -6062 -64 -5665
rect 64 -6062 1178 -5665
rect 1306 -6062 2420 -5665
rect 2548 -6062 3662 -5665
rect 3790 -6062 4904 -5665
rect -4904 -6599 -3790 -6202
rect -3662 -6599 -2548 -6202
rect -2420 -6599 -1306 -6202
rect -1178 -6599 -64 -6202
rect 64 -6599 1178 -6202
rect 1306 -6599 2420 -6202
rect 2548 -6599 3662 -6202
rect 3790 -6599 4904 -6202
rect -4904 -8106 -3790 -7709
rect -3662 -8106 -2548 -7709
rect -2420 -8106 -1306 -7709
rect -1178 -8106 -64 -7709
rect 64 -8106 1178 -7709
rect 1306 -8106 2420 -7709
rect 2548 -8106 3662 -7709
rect 3790 -8106 4904 -7709
rect -4904 -8643 -3790 -8246
rect -3662 -8643 -2548 -8246
rect -2420 -8643 -1306 -8246
rect -1178 -8643 -64 -8246
rect 64 -8643 1178 -8246
rect 1306 -8643 2420 -8246
rect 2548 -8643 3662 -8246
rect 3790 -8643 4904 -8246
rect -4904 -10150 -3790 -9753
rect -3662 -10150 -2548 -9753
rect -2420 -10150 -1306 -9753
rect -1178 -10150 -64 -9753
rect 64 -10150 1178 -9753
rect 1306 -10150 2420 -9753
rect 2548 -10150 3662 -9753
rect 3790 -10150 4904 -9753
rect -4904 -10687 -3790 -10290
rect -3662 -10687 -2548 -10290
rect -2420 -10687 -1306 -10290
rect -1178 -10687 -64 -10290
rect 64 -10687 1178 -10290
rect 1306 -10687 2420 -10290
rect 2548 -10687 3662 -10290
rect 3790 -10687 4904 -10290
rect -4904 -12194 -3790 -11797
rect -3662 -12194 -2548 -11797
rect -2420 -12194 -1306 -11797
rect -1178 -12194 -64 -11797
rect 64 -12194 1178 -11797
rect 1306 -12194 2420 -11797
rect 2548 -12194 3662 -11797
rect 3790 -12194 4904 -11797
rect -4904 -12731 -3790 -12334
rect -3662 -12731 -2548 -12334
rect -2420 -12731 -1306 -12334
rect -1178 -12731 -64 -12334
rect 64 -12731 1178 -12334
rect 1306 -12731 2420 -12334
rect 2548 -12731 3662 -12334
rect 3790 -12731 4904 -12334
rect -4904 -14238 -3790 -13841
rect -3662 -14238 -2548 -13841
rect -2420 -14238 -1306 -13841
rect -1178 -14238 -64 -13841
rect 64 -14238 1178 -13841
rect 1306 -14238 2420 -13841
rect 2548 -14238 3662 -13841
rect 3790 -14238 4904 -13841
rect -4904 -14775 -3790 -14378
rect -3662 -14775 -2548 -14378
rect -2420 -14775 -1306 -14378
rect -1178 -14775 -64 -14378
rect 64 -14775 1178 -14378
rect 1306 -14775 2420 -14378
rect 2548 -14775 3662 -14378
rect 3790 -14775 4904 -14378
rect -4904 -16282 -3790 -15885
rect -3662 -16282 -2548 -15885
rect -2420 -16282 -1306 -15885
rect -1178 -16282 -64 -15885
rect 64 -16282 1178 -15885
rect 1306 -16282 2420 -15885
rect 2548 -16282 3662 -15885
rect 3790 -16282 4904 -15885
rect -4904 -16819 -3790 -16422
rect -3662 -16819 -2548 -16422
rect -2420 -16819 -1306 -16422
rect -1178 -16819 -64 -16422
rect 64 -16819 1178 -16422
rect 1306 -16819 2420 -16422
rect 2548 -16819 3662 -16422
rect 3790 -16819 4904 -16422
rect -4904 -18326 -3790 -17929
rect -3662 -18326 -2548 -17929
rect -2420 -18326 -1306 -17929
rect -1178 -18326 -64 -17929
rect 64 -18326 1178 -17929
rect 1306 -18326 2420 -17929
rect 2548 -18326 3662 -17929
rect 3790 -18326 4904 -17929
<< metal1 >>
rect -4916 18326 -3778 18332
rect -4916 17929 -4904 18326
rect -3790 17929 -3778 18326
rect -4916 17923 -3778 17929
rect -3674 18326 -2536 18332
rect -3674 17929 -3662 18326
rect -2548 17929 -2536 18326
rect -3674 17923 -2536 17929
rect -2432 18326 -1294 18332
rect -2432 17929 -2420 18326
rect -1306 17929 -1294 18326
rect -2432 17923 -1294 17929
rect -1190 18326 -52 18332
rect -1190 17929 -1178 18326
rect -64 17929 -52 18326
rect -1190 17923 -52 17929
rect 52 18326 1190 18332
rect 52 17929 64 18326
rect 1178 17929 1190 18326
rect 52 17923 1190 17929
rect 1294 18326 2432 18332
rect 1294 17929 1306 18326
rect 2420 17929 2432 18326
rect 1294 17923 2432 17929
rect 2536 18326 3674 18332
rect 2536 17929 2548 18326
rect 3662 17929 3674 18326
rect 2536 17923 3674 17929
rect 3778 18326 4916 18332
rect 3778 17929 3790 18326
rect 4904 17929 4916 18326
rect 3778 17923 4916 17929
rect -4916 16819 -3778 16825
rect -4916 16422 -4904 16819
rect -3790 16422 -3778 16819
rect -4916 16416 -3778 16422
rect -3674 16819 -2536 16825
rect -3674 16422 -3662 16819
rect -2548 16422 -2536 16819
rect -3674 16416 -2536 16422
rect -2432 16819 -1294 16825
rect -2432 16422 -2420 16819
rect -1306 16422 -1294 16819
rect -2432 16416 -1294 16422
rect -1190 16819 -52 16825
rect -1190 16422 -1178 16819
rect -64 16422 -52 16819
rect -1190 16416 -52 16422
rect 52 16819 1190 16825
rect 52 16422 64 16819
rect 1178 16422 1190 16819
rect 52 16416 1190 16422
rect 1294 16819 2432 16825
rect 1294 16422 1306 16819
rect 2420 16422 2432 16819
rect 1294 16416 2432 16422
rect 2536 16819 3674 16825
rect 2536 16422 2548 16819
rect 3662 16422 3674 16819
rect 2536 16416 3674 16422
rect 3778 16819 4916 16825
rect 3778 16422 3790 16819
rect 4904 16422 4916 16819
rect 3778 16416 4916 16422
rect -4916 16282 -3778 16288
rect -4916 15885 -4904 16282
rect -3790 15885 -3778 16282
rect -4916 15879 -3778 15885
rect -3674 16282 -2536 16288
rect -3674 15885 -3662 16282
rect -2548 15885 -2536 16282
rect -3674 15879 -2536 15885
rect -2432 16282 -1294 16288
rect -2432 15885 -2420 16282
rect -1306 15885 -1294 16282
rect -2432 15879 -1294 15885
rect -1190 16282 -52 16288
rect -1190 15885 -1178 16282
rect -64 15885 -52 16282
rect -1190 15879 -52 15885
rect 52 16282 1190 16288
rect 52 15885 64 16282
rect 1178 15885 1190 16282
rect 52 15879 1190 15885
rect 1294 16282 2432 16288
rect 1294 15885 1306 16282
rect 2420 15885 2432 16282
rect 1294 15879 2432 15885
rect 2536 16282 3674 16288
rect 2536 15885 2548 16282
rect 3662 15885 3674 16282
rect 2536 15879 3674 15885
rect 3778 16282 4916 16288
rect 3778 15885 3790 16282
rect 4904 15885 4916 16282
rect 3778 15879 4916 15885
rect -4916 14775 -3778 14781
rect -4916 14378 -4904 14775
rect -3790 14378 -3778 14775
rect -4916 14372 -3778 14378
rect -3674 14775 -2536 14781
rect -3674 14378 -3662 14775
rect -2548 14378 -2536 14775
rect -3674 14372 -2536 14378
rect -2432 14775 -1294 14781
rect -2432 14378 -2420 14775
rect -1306 14378 -1294 14775
rect -2432 14372 -1294 14378
rect -1190 14775 -52 14781
rect -1190 14378 -1178 14775
rect -64 14378 -52 14775
rect -1190 14372 -52 14378
rect 52 14775 1190 14781
rect 52 14378 64 14775
rect 1178 14378 1190 14775
rect 52 14372 1190 14378
rect 1294 14775 2432 14781
rect 1294 14378 1306 14775
rect 2420 14378 2432 14775
rect 1294 14372 2432 14378
rect 2536 14775 3674 14781
rect 2536 14378 2548 14775
rect 3662 14378 3674 14775
rect 2536 14372 3674 14378
rect 3778 14775 4916 14781
rect 3778 14378 3790 14775
rect 4904 14378 4916 14775
rect 3778 14372 4916 14378
rect -4916 14238 -3778 14244
rect -4916 13841 -4904 14238
rect -3790 13841 -3778 14238
rect -4916 13835 -3778 13841
rect -3674 14238 -2536 14244
rect -3674 13841 -3662 14238
rect -2548 13841 -2536 14238
rect -3674 13835 -2536 13841
rect -2432 14238 -1294 14244
rect -2432 13841 -2420 14238
rect -1306 13841 -1294 14238
rect -2432 13835 -1294 13841
rect -1190 14238 -52 14244
rect -1190 13841 -1178 14238
rect -64 13841 -52 14238
rect -1190 13835 -52 13841
rect 52 14238 1190 14244
rect 52 13841 64 14238
rect 1178 13841 1190 14238
rect 52 13835 1190 13841
rect 1294 14238 2432 14244
rect 1294 13841 1306 14238
rect 2420 13841 2432 14238
rect 1294 13835 2432 13841
rect 2536 14238 3674 14244
rect 2536 13841 2548 14238
rect 3662 13841 3674 14238
rect 2536 13835 3674 13841
rect 3778 14238 4916 14244
rect 3778 13841 3790 14238
rect 4904 13841 4916 14238
rect 3778 13835 4916 13841
rect -4916 12731 -3778 12737
rect -4916 12334 -4904 12731
rect -3790 12334 -3778 12731
rect -4916 12328 -3778 12334
rect -3674 12731 -2536 12737
rect -3674 12334 -3662 12731
rect -2548 12334 -2536 12731
rect -3674 12328 -2536 12334
rect -2432 12731 -1294 12737
rect -2432 12334 -2420 12731
rect -1306 12334 -1294 12731
rect -2432 12328 -1294 12334
rect -1190 12731 -52 12737
rect -1190 12334 -1178 12731
rect -64 12334 -52 12731
rect -1190 12328 -52 12334
rect 52 12731 1190 12737
rect 52 12334 64 12731
rect 1178 12334 1190 12731
rect 52 12328 1190 12334
rect 1294 12731 2432 12737
rect 1294 12334 1306 12731
rect 2420 12334 2432 12731
rect 1294 12328 2432 12334
rect 2536 12731 3674 12737
rect 2536 12334 2548 12731
rect 3662 12334 3674 12731
rect 2536 12328 3674 12334
rect 3778 12731 4916 12737
rect 3778 12334 3790 12731
rect 4904 12334 4916 12731
rect 3778 12328 4916 12334
rect -4916 12194 -3778 12200
rect -4916 11797 -4904 12194
rect -3790 11797 -3778 12194
rect -4916 11791 -3778 11797
rect -3674 12194 -2536 12200
rect -3674 11797 -3662 12194
rect -2548 11797 -2536 12194
rect -3674 11791 -2536 11797
rect -2432 12194 -1294 12200
rect -2432 11797 -2420 12194
rect -1306 11797 -1294 12194
rect -2432 11791 -1294 11797
rect -1190 12194 -52 12200
rect -1190 11797 -1178 12194
rect -64 11797 -52 12194
rect -1190 11791 -52 11797
rect 52 12194 1190 12200
rect 52 11797 64 12194
rect 1178 11797 1190 12194
rect 52 11791 1190 11797
rect 1294 12194 2432 12200
rect 1294 11797 1306 12194
rect 2420 11797 2432 12194
rect 1294 11791 2432 11797
rect 2536 12194 3674 12200
rect 2536 11797 2548 12194
rect 3662 11797 3674 12194
rect 2536 11791 3674 11797
rect 3778 12194 4916 12200
rect 3778 11797 3790 12194
rect 4904 11797 4916 12194
rect 3778 11791 4916 11797
rect -4916 10687 -3778 10693
rect -4916 10290 -4904 10687
rect -3790 10290 -3778 10687
rect -4916 10284 -3778 10290
rect -3674 10687 -2536 10693
rect -3674 10290 -3662 10687
rect -2548 10290 -2536 10687
rect -3674 10284 -2536 10290
rect -2432 10687 -1294 10693
rect -2432 10290 -2420 10687
rect -1306 10290 -1294 10687
rect -2432 10284 -1294 10290
rect -1190 10687 -52 10693
rect -1190 10290 -1178 10687
rect -64 10290 -52 10687
rect -1190 10284 -52 10290
rect 52 10687 1190 10693
rect 52 10290 64 10687
rect 1178 10290 1190 10687
rect 52 10284 1190 10290
rect 1294 10687 2432 10693
rect 1294 10290 1306 10687
rect 2420 10290 2432 10687
rect 1294 10284 2432 10290
rect 2536 10687 3674 10693
rect 2536 10290 2548 10687
rect 3662 10290 3674 10687
rect 2536 10284 3674 10290
rect 3778 10687 4916 10693
rect 3778 10290 3790 10687
rect 4904 10290 4916 10687
rect 3778 10284 4916 10290
rect -4916 10150 -3778 10156
rect -4916 9753 -4904 10150
rect -3790 9753 -3778 10150
rect -4916 9747 -3778 9753
rect -3674 10150 -2536 10156
rect -3674 9753 -3662 10150
rect -2548 9753 -2536 10150
rect -3674 9747 -2536 9753
rect -2432 10150 -1294 10156
rect -2432 9753 -2420 10150
rect -1306 9753 -1294 10150
rect -2432 9747 -1294 9753
rect -1190 10150 -52 10156
rect -1190 9753 -1178 10150
rect -64 9753 -52 10150
rect -1190 9747 -52 9753
rect 52 10150 1190 10156
rect 52 9753 64 10150
rect 1178 9753 1190 10150
rect 52 9747 1190 9753
rect 1294 10150 2432 10156
rect 1294 9753 1306 10150
rect 2420 9753 2432 10150
rect 1294 9747 2432 9753
rect 2536 10150 3674 10156
rect 2536 9753 2548 10150
rect 3662 9753 3674 10150
rect 2536 9747 3674 9753
rect 3778 10150 4916 10156
rect 3778 9753 3790 10150
rect 4904 9753 4916 10150
rect 3778 9747 4916 9753
rect -4916 8643 -3778 8649
rect -4916 8246 -4904 8643
rect -3790 8246 -3778 8643
rect -4916 8240 -3778 8246
rect -3674 8643 -2536 8649
rect -3674 8246 -3662 8643
rect -2548 8246 -2536 8643
rect -3674 8240 -2536 8246
rect -2432 8643 -1294 8649
rect -2432 8246 -2420 8643
rect -1306 8246 -1294 8643
rect -2432 8240 -1294 8246
rect -1190 8643 -52 8649
rect -1190 8246 -1178 8643
rect -64 8246 -52 8643
rect -1190 8240 -52 8246
rect 52 8643 1190 8649
rect 52 8246 64 8643
rect 1178 8246 1190 8643
rect 52 8240 1190 8246
rect 1294 8643 2432 8649
rect 1294 8246 1306 8643
rect 2420 8246 2432 8643
rect 1294 8240 2432 8246
rect 2536 8643 3674 8649
rect 2536 8246 2548 8643
rect 3662 8246 3674 8643
rect 2536 8240 3674 8246
rect 3778 8643 4916 8649
rect 3778 8246 3790 8643
rect 4904 8246 4916 8643
rect 3778 8240 4916 8246
rect -4916 8106 -3778 8112
rect -4916 7709 -4904 8106
rect -3790 7709 -3778 8106
rect -4916 7703 -3778 7709
rect -3674 8106 -2536 8112
rect -3674 7709 -3662 8106
rect -2548 7709 -2536 8106
rect -3674 7703 -2536 7709
rect -2432 8106 -1294 8112
rect -2432 7709 -2420 8106
rect -1306 7709 -1294 8106
rect -2432 7703 -1294 7709
rect -1190 8106 -52 8112
rect -1190 7709 -1178 8106
rect -64 7709 -52 8106
rect -1190 7703 -52 7709
rect 52 8106 1190 8112
rect 52 7709 64 8106
rect 1178 7709 1190 8106
rect 52 7703 1190 7709
rect 1294 8106 2432 8112
rect 1294 7709 1306 8106
rect 2420 7709 2432 8106
rect 1294 7703 2432 7709
rect 2536 8106 3674 8112
rect 2536 7709 2548 8106
rect 3662 7709 3674 8106
rect 2536 7703 3674 7709
rect 3778 8106 4916 8112
rect 3778 7709 3790 8106
rect 4904 7709 4916 8106
rect 3778 7703 4916 7709
rect -4916 6599 -3778 6605
rect -4916 6202 -4904 6599
rect -3790 6202 -3778 6599
rect -4916 6196 -3778 6202
rect -3674 6599 -2536 6605
rect -3674 6202 -3662 6599
rect -2548 6202 -2536 6599
rect -3674 6196 -2536 6202
rect -2432 6599 -1294 6605
rect -2432 6202 -2420 6599
rect -1306 6202 -1294 6599
rect -2432 6196 -1294 6202
rect -1190 6599 -52 6605
rect -1190 6202 -1178 6599
rect -64 6202 -52 6599
rect -1190 6196 -52 6202
rect 52 6599 1190 6605
rect 52 6202 64 6599
rect 1178 6202 1190 6599
rect 52 6196 1190 6202
rect 1294 6599 2432 6605
rect 1294 6202 1306 6599
rect 2420 6202 2432 6599
rect 1294 6196 2432 6202
rect 2536 6599 3674 6605
rect 2536 6202 2548 6599
rect 3662 6202 3674 6599
rect 2536 6196 3674 6202
rect 3778 6599 4916 6605
rect 3778 6202 3790 6599
rect 4904 6202 4916 6599
rect 3778 6196 4916 6202
rect -4916 6062 -3778 6068
rect -4916 5665 -4904 6062
rect -3790 5665 -3778 6062
rect -4916 5659 -3778 5665
rect -3674 6062 -2536 6068
rect -3674 5665 -3662 6062
rect -2548 5665 -2536 6062
rect -3674 5659 -2536 5665
rect -2432 6062 -1294 6068
rect -2432 5665 -2420 6062
rect -1306 5665 -1294 6062
rect -2432 5659 -1294 5665
rect -1190 6062 -52 6068
rect -1190 5665 -1178 6062
rect -64 5665 -52 6062
rect -1190 5659 -52 5665
rect 52 6062 1190 6068
rect 52 5665 64 6062
rect 1178 5665 1190 6062
rect 52 5659 1190 5665
rect 1294 6062 2432 6068
rect 1294 5665 1306 6062
rect 2420 5665 2432 6062
rect 1294 5659 2432 5665
rect 2536 6062 3674 6068
rect 2536 5665 2548 6062
rect 3662 5665 3674 6062
rect 2536 5659 3674 5665
rect 3778 6062 4916 6068
rect 3778 5665 3790 6062
rect 4904 5665 4916 6062
rect 3778 5659 4916 5665
rect -4916 4555 -3778 4561
rect -4916 4158 -4904 4555
rect -3790 4158 -3778 4555
rect -4916 4152 -3778 4158
rect -3674 4555 -2536 4561
rect -3674 4158 -3662 4555
rect -2548 4158 -2536 4555
rect -3674 4152 -2536 4158
rect -2432 4555 -1294 4561
rect -2432 4158 -2420 4555
rect -1306 4158 -1294 4555
rect -2432 4152 -1294 4158
rect -1190 4555 -52 4561
rect -1190 4158 -1178 4555
rect -64 4158 -52 4555
rect -1190 4152 -52 4158
rect 52 4555 1190 4561
rect 52 4158 64 4555
rect 1178 4158 1190 4555
rect 52 4152 1190 4158
rect 1294 4555 2432 4561
rect 1294 4158 1306 4555
rect 2420 4158 2432 4555
rect 1294 4152 2432 4158
rect 2536 4555 3674 4561
rect 2536 4158 2548 4555
rect 3662 4158 3674 4555
rect 2536 4152 3674 4158
rect 3778 4555 4916 4561
rect 3778 4158 3790 4555
rect 4904 4158 4916 4555
rect 3778 4152 4916 4158
rect -4916 4018 -3778 4024
rect -4916 3621 -4904 4018
rect -3790 3621 -3778 4018
rect -4916 3615 -3778 3621
rect -3674 4018 -2536 4024
rect -3674 3621 -3662 4018
rect -2548 3621 -2536 4018
rect -3674 3615 -2536 3621
rect -2432 4018 -1294 4024
rect -2432 3621 -2420 4018
rect -1306 3621 -1294 4018
rect -2432 3615 -1294 3621
rect -1190 4018 -52 4024
rect -1190 3621 -1178 4018
rect -64 3621 -52 4018
rect -1190 3615 -52 3621
rect 52 4018 1190 4024
rect 52 3621 64 4018
rect 1178 3621 1190 4018
rect 52 3615 1190 3621
rect 1294 4018 2432 4024
rect 1294 3621 1306 4018
rect 2420 3621 2432 4018
rect 1294 3615 2432 3621
rect 2536 4018 3674 4024
rect 2536 3621 2548 4018
rect 3662 3621 3674 4018
rect 2536 3615 3674 3621
rect 3778 4018 4916 4024
rect 3778 3621 3790 4018
rect 4904 3621 4916 4018
rect 3778 3615 4916 3621
rect -4916 2511 -3778 2517
rect -4916 2114 -4904 2511
rect -3790 2114 -3778 2511
rect -4916 2108 -3778 2114
rect -3674 2511 -2536 2517
rect -3674 2114 -3662 2511
rect -2548 2114 -2536 2511
rect -3674 2108 -2536 2114
rect -2432 2511 -1294 2517
rect -2432 2114 -2420 2511
rect -1306 2114 -1294 2511
rect -2432 2108 -1294 2114
rect -1190 2511 -52 2517
rect -1190 2114 -1178 2511
rect -64 2114 -52 2511
rect -1190 2108 -52 2114
rect 52 2511 1190 2517
rect 52 2114 64 2511
rect 1178 2114 1190 2511
rect 52 2108 1190 2114
rect 1294 2511 2432 2517
rect 1294 2114 1306 2511
rect 2420 2114 2432 2511
rect 1294 2108 2432 2114
rect 2536 2511 3674 2517
rect 2536 2114 2548 2511
rect 3662 2114 3674 2511
rect 2536 2108 3674 2114
rect 3778 2511 4916 2517
rect 3778 2114 3790 2511
rect 4904 2114 4916 2511
rect 3778 2108 4916 2114
rect -4916 1974 -3778 1980
rect -4916 1577 -4904 1974
rect -3790 1577 -3778 1974
rect -4916 1571 -3778 1577
rect -3674 1974 -2536 1980
rect -3674 1577 -3662 1974
rect -2548 1577 -2536 1974
rect -3674 1571 -2536 1577
rect -2432 1974 -1294 1980
rect -2432 1577 -2420 1974
rect -1306 1577 -1294 1974
rect -2432 1571 -1294 1577
rect -1190 1974 -52 1980
rect -1190 1577 -1178 1974
rect -64 1577 -52 1974
rect -1190 1571 -52 1577
rect 52 1974 1190 1980
rect 52 1577 64 1974
rect 1178 1577 1190 1974
rect 52 1571 1190 1577
rect 1294 1974 2432 1980
rect 1294 1577 1306 1974
rect 2420 1577 2432 1974
rect 1294 1571 2432 1577
rect 2536 1974 3674 1980
rect 2536 1577 2548 1974
rect 3662 1577 3674 1974
rect 2536 1571 3674 1577
rect 3778 1974 4916 1980
rect 3778 1577 3790 1974
rect 4904 1577 4916 1974
rect 3778 1571 4916 1577
rect -4916 467 -3778 473
rect -4916 70 -4904 467
rect -3790 70 -3778 467
rect -4916 64 -3778 70
rect -3674 467 -2536 473
rect -3674 70 -3662 467
rect -2548 70 -2536 467
rect -3674 64 -2536 70
rect -2432 467 -1294 473
rect -2432 70 -2420 467
rect -1306 70 -1294 467
rect -2432 64 -1294 70
rect -1190 467 -52 473
rect -1190 70 -1178 467
rect -64 70 -52 467
rect -1190 64 -52 70
rect 52 467 1190 473
rect 52 70 64 467
rect 1178 70 1190 467
rect 52 64 1190 70
rect 1294 467 2432 473
rect 1294 70 1306 467
rect 2420 70 2432 467
rect 1294 64 2432 70
rect 2536 467 3674 473
rect 2536 70 2548 467
rect 3662 70 3674 467
rect 2536 64 3674 70
rect 3778 467 4916 473
rect 3778 70 3790 467
rect 4904 70 4916 467
rect 3778 64 4916 70
rect -4916 -70 -3778 -64
rect -4916 -467 -4904 -70
rect -3790 -467 -3778 -70
rect -4916 -473 -3778 -467
rect -3674 -70 -2536 -64
rect -3674 -467 -3662 -70
rect -2548 -467 -2536 -70
rect -3674 -473 -2536 -467
rect -2432 -70 -1294 -64
rect -2432 -467 -2420 -70
rect -1306 -467 -1294 -70
rect -2432 -473 -1294 -467
rect -1190 -70 -52 -64
rect -1190 -467 -1178 -70
rect -64 -467 -52 -70
rect -1190 -473 -52 -467
rect 52 -70 1190 -64
rect 52 -467 64 -70
rect 1178 -467 1190 -70
rect 52 -473 1190 -467
rect 1294 -70 2432 -64
rect 1294 -467 1306 -70
rect 2420 -467 2432 -70
rect 1294 -473 2432 -467
rect 2536 -70 3674 -64
rect 2536 -467 2548 -70
rect 3662 -467 3674 -70
rect 2536 -473 3674 -467
rect 3778 -70 4916 -64
rect 3778 -467 3790 -70
rect 4904 -467 4916 -70
rect 3778 -473 4916 -467
rect -4916 -1577 -3778 -1571
rect -4916 -1974 -4904 -1577
rect -3790 -1974 -3778 -1577
rect -4916 -1980 -3778 -1974
rect -3674 -1577 -2536 -1571
rect -3674 -1974 -3662 -1577
rect -2548 -1974 -2536 -1577
rect -3674 -1980 -2536 -1974
rect -2432 -1577 -1294 -1571
rect -2432 -1974 -2420 -1577
rect -1306 -1974 -1294 -1577
rect -2432 -1980 -1294 -1974
rect -1190 -1577 -52 -1571
rect -1190 -1974 -1178 -1577
rect -64 -1974 -52 -1577
rect -1190 -1980 -52 -1974
rect 52 -1577 1190 -1571
rect 52 -1974 64 -1577
rect 1178 -1974 1190 -1577
rect 52 -1980 1190 -1974
rect 1294 -1577 2432 -1571
rect 1294 -1974 1306 -1577
rect 2420 -1974 2432 -1577
rect 1294 -1980 2432 -1974
rect 2536 -1577 3674 -1571
rect 2536 -1974 2548 -1577
rect 3662 -1974 3674 -1577
rect 2536 -1980 3674 -1974
rect 3778 -1577 4916 -1571
rect 3778 -1974 3790 -1577
rect 4904 -1974 4916 -1577
rect 3778 -1980 4916 -1974
rect -4916 -2114 -3778 -2108
rect -4916 -2511 -4904 -2114
rect -3790 -2511 -3778 -2114
rect -4916 -2517 -3778 -2511
rect -3674 -2114 -2536 -2108
rect -3674 -2511 -3662 -2114
rect -2548 -2511 -2536 -2114
rect -3674 -2517 -2536 -2511
rect -2432 -2114 -1294 -2108
rect -2432 -2511 -2420 -2114
rect -1306 -2511 -1294 -2114
rect -2432 -2517 -1294 -2511
rect -1190 -2114 -52 -2108
rect -1190 -2511 -1178 -2114
rect -64 -2511 -52 -2114
rect -1190 -2517 -52 -2511
rect 52 -2114 1190 -2108
rect 52 -2511 64 -2114
rect 1178 -2511 1190 -2114
rect 52 -2517 1190 -2511
rect 1294 -2114 2432 -2108
rect 1294 -2511 1306 -2114
rect 2420 -2511 2432 -2114
rect 1294 -2517 2432 -2511
rect 2536 -2114 3674 -2108
rect 2536 -2511 2548 -2114
rect 3662 -2511 3674 -2114
rect 2536 -2517 3674 -2511
rect 3778 -2114 4916 -2108
rect 3778 -2511 3790 -2114
rect 4904 -2511 4916 -2114
rect 3778 -2517 4916 -2511
rect -4916 -3621 -3778 -3615
rect -4916 -4018 -4904 -3621
rect -3790 -4018 -3778 -3621
rect -4916 -4024 -3778 -4018
rect -3674 -3621 -2536 -3615
rect -3674 -4018 -3662 -3621
rect -2548 -4018 -2536 -3621
rect -3674 -4024 -2536 -4018
rect -2432 -3621 -1294 -3615
rect -2432 -4018 -2420 -3621
rect -1306 -4018 -1294 -3621
rect -2432 -4024 -1294 -4018
rect -1190 -3621 -52 -3615
rect -1190 -4018 -1178 -3621
rect -64 -4018 -52 -3621
rect -1190 -4024 -52 -4018
rect 52 -3621 1190 -3615
rect 52 -4018 64 -3621
rect 1178 -4018 1190 -3621
rect 52 -4024 1190 -4018
rect 1294 -3621 2432 -3615
rect 1294 -4018 1306 -3621
rect 2420 -4018 2432 -3621
rect 1294 -4024 2432 -4018
rect 2536 -3621 3674 -3615
rect 2536 -4018 2548 -3621
rect 3662 -4018 3674 -3621
rect 2536 -4024 3674 -4018
rect 3778 -3621 4916 -3615
rect 3778 -4018 3790 -3621
rect 4904 -4018 4916 -3621
rect 3778 -4024 4916 -4018
rect -4916 -4158 -3778 -4152
rect -4916 -4555 -4904 -4158
rect -3790 -4555 -3778 -4158
rect -4916 -4561 -3778 -4555
rect -3674 -4158 -2536 -4152
rect -3674 -4555 -3662 -4158
rect -2548 -4555 -2536 -4158
rect -3674 -4561 -2536 -4555
rect -2432 -4158 -1294 -4152
rect -2432 -4555 -2420 -4158
rect -1306 -4555 -1294 -4158
rect -2432 -4561 -1294 -4555
rect -1190 -4158 -52 -4152
rect -1190 -4555 -1178 -4158
rect -64 -4555 -52 -4158
rect -1190 -4561 -52 -4555
rect 52 -4158 1190 -4152
rect 52 -4555 64 -4158
rect 1178 -4555 1190 -4158
rect 52 -4561 1190 -4555
rect 1294 -4158 2432 -4152
rect 1294 -4555 1306 -4158
rect 2420 -4555 2432 -4158
rect 1294 -4561 2432 -4555
rect 2536 -4158 3674 -4152
rect 2536 -4555 2548 -4158
rect 3662 -4555 3674 -4158
rect 2536 -4561 3674 -4555
rect 3778 -4158 4916 -4152
rect 3778 -4555 3790 -4158
rect 4904 -4555 4916 -4158
rect 3778 -4561 4916 -4555
rect -4916 -5665 -3778 -5659
rect -4916 -6062 -4904 -5665
rect -3790 -6062 -3778 -5665
rect -4916 -6068 -3778 -6062
rect -3674 -5665 -2536 -5659
rect -3674 -6062 -3662 -5665
rect -2548 -6062 -2536 -5665
rect -3674 -6068 -2536 -6062
rect -2432 -5665 -1294 -5659
rect -2432 -6062 -2420 -5665
rect -1306 -6062 -1294 -5665
rect -2432 -6068 -1294 -6062
rect -1190 -5665 -52 -5659
rect -1190 -6062 -1178 -5665
rect -64 -6062 -52 -5665
rect -1190 -6068 -52 -6062
rect 52 -5665 1190 -5659
rect 52 -6062 64 -5665
rect 1178 -6062 1190 -5665
rect 52 -6068 1190 -6062
rect 1294 -5665 2432 -5659
rect 1294 -6062 1306 -5665
rect 2420 -6062 2432 -5665
rect 1294 -6068 2432 -6062
rect 2536 -5665 3674 -5659
rect 2536 -6062 2548 -5665
rect 3662 -6062 3674 -5665
rect 2536 -6068 3674 -6062
rect 3778 -5665 4916 -5659
rect 3778 -6062 3790 -5665
rect 4904 -6062 4916 -5665
rect 3778 -6068 4916 -6062
rect -4916 -6202 -3778 -6196
rect -4916 -6599 -4904 -6202
rect -3790 -6599 -3778 -6202
rect -4916 -6605 -3778 -6599
rect -3674 -6202 -2536 -6196
rect -3674 -6599 -3662 -6202
rect -2548 -6599 -2536 -6202
rect -3674 -6605 -2536 -6599
rect -2432 -6202 -1294 -6196
rect -2432 -6599 -2420 -6202
rect -1306 -6599 -1294 -6202
rect -2432 -6605 -1294 -6599
rect -1190 -6202 -52 -6196
rect -1190 -6599 -1178 -6202
rect -64 -6599 -52 -6202
rect -1190 -6605 -52 -6599
rect 52 -6202 1190 -6196
rect 52 -6599 64 -6202
rect 1178 -6599 1190 -6202
rect 52 -6605 1190 -6599
rect 1294 -6202 2432 -6196
rect 1294 -6599 1306 -6202
rect 2420 -6599 2432 -6202
rect 1294 -6605 2432 -6599
rect 2536 -6202 3674 -6196
rect 2536 -6599 2548 -6202
rect 3662 -6599 3674 -6202
rect 2536 -6605 3674 -6599
rect 3778 -6202 4916 -6196
rect 3778 -6599 3790 -6202
rect 4904 -6599 4916 -6202
rect 3778 -6605 4916 -6599
rect -4916 -7709 -3778 -7703
rect -4916 -8106 -4904 -7709
rect -3790 -8106 -3778 -7709
rect -4916 -8112 -3778 -8106
rect -3674 -7709 -2536 -7703
rect -3674 -8106 -3662 -7709
rect -2548 -8106 -2536 -7709
rect -3674 -8112 -2536 -8106
rect -2432 -7709 -1294 -7703
rect -2432 -8106 -2420 -7709
rect -1306 -8106 -1294 -7709
rect -2432 -8112 -1294 -8106
rect -1190 -7709 -52 -7703
rect -1190 -8106 -1178 -7709
rect -64 -8106 -52 -7709
rect -1190 -8112 -52 -8106
rect 52 -7709 1190 -7703
rect 52 -8106 64 -7709
rect 1178 -8106 1190 -7709
rect 52 -8112 1190 -8106
rect 1294 -7709 2432 -7703
rect 1294 -8106 1306 -7709
rect 2420 -8106 2432 -7709
rect 1294 -8112 2432 -8106
rect 2536 -7709 3674 -7703
rect 2536 -8106 2548 -7709
rect 3662 -8106 3674 -7709
rect 2536 -8112 3674 -8106
rect 3778 -7709 4916 -7703
rect 3778 -8106 3790 -7709
rect 4904 -8106 4916 -7709
rect 3778 -8112 4916 -8106
rect -4916 -8246 -3778 -8240
rect -4916 -8643 -4904 -8246
rect -3790 -8643 -3778 -8246
rect -4916 -8649 -3778 -8643
rect -3674 -8246 -2536 -8240
rect -3674 -8643 -3662 -8246
rect -2548 -8643 -2536 -8246
rect -3674 -8649 -2536 -8643
rect -2432 -8246 -1294 -8240
rect -2432 -8643 -2420 -8246
rect -1306 -8643 -1294 -8246
rect -2432 -8649 -1294 -8643
rect -1190 -8246 -52 -8240
rect -1190 -8643 -1178 -8246
rect -64 -8643 -52 -8246
rect -1190 -8649 -52 -8643
rect 52 -8246 1190 -8240
rect 52 -8643 64 -8246
rect 1178 -8643 1190 -8246
rect 52 -8649 1190 -8643
rect 1294 -8246 2432 -8240
rect 1294 -8643 1306 -8246
rect 2420 -8643 2432 -8246
rect 1294 -8649 2432 -8643
rect 2536 -8246 3674 -8240
rect 2536 -8643 2548 -8246
rect 3662 -8643 3674 -8246
rect 2536 -8649 3674 -8643
rect 3778 -8246 4916 -8240
rect 3778 -8643 3790 -8246
rect 4904 -8643 4916 -8246
rect 3778 -8649 4916 -8643
rect -4916 -9753 -3778 -9747
rect -4916 -10150 -4904 -9753
rect -3790 -10150 -3778 -9753
rect -4916 -10156 -3778 -10150
rect -3674 -9753 -2536 -9747
rect -3674 -10150 -3662 -9753
rect -2548 -10150 -2536 -9753
rect -3674 -10156 -2536 -10150
rect -2432 -9753 -1294 -9747
rect -2432 -10150 -2420 -9753
rect -1306 -10150 -1294 -9753
rect -2432 -10156 -1294 -10150
rect -1190 -9753 -52 -9747
rect -1190 -10150 -1178 -9753
rect -64 -10150 -52 -9753
rect -1190 -10156 -52 -10150
rect 52 -9753 1190 -9747
rect 52 -10150 64 -9753
rect 1178 -10150 1190 -9753
rect 52 -10156 1190 -10150
rect 1294 -9753 2432 -9747
rect 1294 -10150 1306 -9753
rect 2420 -10150 2432 -9753
rect 1294 -10156 2432 -10150
rect 2536 -9753 3674 -9747
rect 2536 -10150 2548 -9753
rect 3662 -10150 3674 -9753
rect 2536 -10156 3674 -10150
rect 3778 -9753 4916 -9747
rect 3778 -10150 3790 -9753
rect 4904 -10150 4916 -9753
rect 3778 -10156 4916 -10150
rect -4916 -10290 -3778 -10284
rect -4916 -10687 -4904 -10290
rect -3790 -10687 -3778 -10290
rect -4916 -10693 -3778 -10687
rect -3674 -10290 -2536 -10284
rect -3674 -10687 -3662 -10290
rect -2548 -10687 -2536 -10290
rect -3674 -10693 -2536 -10687
rect -2432 -10290 -1294 -10284
rect -2432 -10687 -2420 -10290
rect -1306 -10687 -1294 -10290
rect -2432 -10693 -1294 -10687
rect -1190 -10290 -52 -10284
rect -1190 -10687 -1178 -10290
rect -64 -10687 -52 -10290
rect -1190 -10693 -52 -10687
rect 52 -10290 1190 -10284
rect 52 -10687 64 -10290
rect 1178 -10687 1190 -10290
rect 52 -10693 1190 -10687
rect 1294 -10290 2432 -10284
rect 1294 -10687 1306 -10290
rect 2420 -10687 2432 -10290
rect 1294 -10693 2432 -10687
rect 2536 -10290 3674 -10284
rect 2536 -10687 2548 -10290
rect 3662 -10687 3674 -10290
rect 2536 -10693 3674 -10687
rect 3778 -10290 4916 -10284
rect 3778 -10687 3790 -10290
rect 4904 -10687 4916 -10290
rect 3778 -10693 4916 -10687
rect -4916 -11797 -3778 -11791
rect -4916 -12194 -4904 -11797
rect -3790 -12194 -3778 -11797
rect -4916 -12200 -3778 -12194
rect -3674 -11797 -2536 -11791
rect -3674 -12194 -3662 -11797
rect -2548 -12194 -2536 -11797
rect -3674 -12200 -2536 -12194
rect -2432 -11797 -1294 -11791
rect -2432 -12194 -2420 -11797
rect -1306 -12194 -1294 -11797
rect -2432 -12200 -1294 -12194
rect -1190 -11797 -52 -11791
rect -1190 -12194 -1178 -11797
rect -64 -12194 -52 -11797
rect -1190 -12200 -52 -12194
rect 52 -11797 1190 -11791
rect 52 -12194 64 -11797
rect 1178 -12194 1190 -11797
rect 52 -12200 1190 -12194
rect 1294 -11797 2432 -11791
rect 1294 -12194 1306 -11797
rect 2420 -12194 2432 -11797
rect 1294 -12200 2432 -12194
rect 2536 -11797 3674 -11791
rect 2536 -12194 2548 -11797
rect 3662 -12194 3674 -11797
rect 2536 -12200 3674 -12194
rect 3778 -11797 4916 -11791
rect 3778 -12194 3790 -11797
rect 4904 -12194 4916 -11797
rect 3778 -12200 4916 -12194
rect -4916 -12334 -3778 -12328
rect -4916 -12731 -4904 -12334
rect -3790 -12731 -3778 -12334
rect -4916 -12737 -3778 -12731
rect -3674 -12334 -2536 -12328
rect -3674 -12731 -3662 -12334
rect -2548 -12731 -2536 -12334
rect -3674 -12737 -2536 -12731
rect -2432 -12334 -1294 -12328
rect -2432 -12731 -2420 -12334
rect -1306 -12731 -1294 -12334
rect -2432 -12737 -1294 -12731
rect -1190 -12334 -52 -12328
rect -1190 -12731 -1178 -12334
rect -64 -12731 -52 -12334
rect -1190 -12737 -52 -12731
rect 52 -12334 1190 -12328
rect 52 -12731 64 -12334
rect 1178 -12731 1190 -12334
rect 52 -12737 1190 -12731
rect 1294 -12334 2432 -12328
rect 1294 -12731 1306 -12334
rect 2420 -12731 2432 -12334
rect 1294 -12737 2432 -12731
rect 2536 -12334 3674 -12328
rect 2536 -12731 2548 -12334
rect 3662 -12731 3674 -12334
rect 2536 -12737 3674 -12731
rect 3778 -12334 4916 -12328
rect 3778 -12731 3790 -12334
rect 4904 -12731 4916 -12334
rect 3778 -12737 4916 -12731
rect -4916 -13841 -3778 -13835
rect -4916 -14238 -4904 -13841
rect -3790 -14238 -3778 -13841
rect -4916 -14244 -3778 -14238
rect -3674 -13841 -2536 -13835
rect -3674 -14238 -3662 -13841
rect -2548 -14238 -2536 -13841
rect -3674 -14244 -2536 -14238
rect -2432 -13841 -1294 -13835
rect -2432 -14238 -2420 -13841
rect -1306 -14238 -1294 -13841
rect -2432 -14244 -1294 -14238
rect -1190 -13841 -52 -13835
rect -1190 -14238 -1178 -13841
rect -64 -14238 -52 -13841
rect -1190 -14244 -52 -14238
rect 52 -13841 1190 -13835
rect 52 -14238 64 -13841
rect 1178 -14238 1190 -13841
rect 52 -14244 1190 -14238
rect 1294 -13841 2432 -13835
rect 1294 -14238 1306 -13841
rect 2420 -14238 2432 -13841
rect 1294 -14244 2432 -14238
rect 2536 -13841 3674 -13835
rect 2536 -14238 2548 -13841
rect 3662 -14238 3674 -13841
rect 2536 -14244 3674 -14238
rect 3778 -13841 4916 -13835
rect 3778 -14238 3790 -13841
rect 4904 -14238 4916 -13841
rect 3778 -14244 4916 -14238
rect -4916 -14378 -3778 -14372
rect -4916 -14775 -4904 -14378
rect -3790 -14775 -3778 -14378
rect -4916 -14781 -3778 -14775
rect -3674 -14378 -2536 -14372
rect -3674 -14775 -3662 -14378
rect -2548 -14775 -2536 -14378
rect -3674 -14781 -2536 -14775
rect -2432 -14378 -1294 -14372
rect -2432 -14775 -2420 -14378
rect -1306 -14775 -1294 -14378
rect -2432 -14781 -1294 -14775
rect -1190 -14378 -52 -14372
rect -1190 -14775 -1178 -14378
rect -64 -14775 -52 -14378
rect -1190 -14781 -52 -14775
rect 52 -14378 1190 -14372
rect 52 -14775 64 -14378
rect 1178 -14775 1190 -14378
rect 52 -14781 1190 -14775
rect 1294 -14378 2432 -14372
rect 1294 -14775 1306 -14378
rect 2420 -14775 2432 -14378
rect 1294 -14781 2432 -14775
rect 2536 -14378 3674 -14372
rect 2536 -14775 2548 -14378
rect 3662 -14775 3674 -14378
rect 2536 -14781 3674 -14775
rect 3778 -14378 4916 -14372
rect 3778 -14775 3790 -14378
rect 4904 -14775 4916 -14378
rect 3778 -14781 4916 -14775
rect -4916 -15885 -3778 -15879
rect -4916 -16282 -4904 -15885
rect -3790 -16282 -3778 -15885
rect -4916 -16288 -3778 -16282
rect -3674 -15885 -2536 -15879
rect -3674 -16282 -3662 -15885
rect -2548 -16282 -2536 -15885
rect -3674 -16288 -2536 -16282
rect -2432 -15885 -1294 -15879
rect -2432 -16282 -2420 -15885
rect -1306 -16282 -1294 -15885
rect -2432 -16288 -1294 -16282
rect -1190 -15885 -52 -15879
rect -1190 -16282 -1178 -15885
rect -64 -16282 -52 -15885
rect -1190 -16288 -52 -16282
rect 52 -15885 1190 -15879
rect 52 -16282 64 -15885
rect 1178 -16282 1190 -15885
rect 52 -16288 1190 -16282
rect 1294 -15885 2432 -15879
rect 1294 -16282 1306 -15885
rect 2420 -16282 2432 -15885
rect 1294 -16288 2432 -16282
rect 2536 -15885 3674 -15879
rect 2536 -16282 2548 -15885
rect 3662 -16282 3674 -15885
rect 2536 -16288 3674 -16282
rect 3778 -15885 4916 -15879
rect 3778 -16282 3790 -15885
rect 4904 -16282 4916 -15885
rect 3778 -16288 4916 -16282
rect -4916 -16422 -3778 -16416
rect -4916 -16819 -4904 -16422
rect -3790 -16819 -3778 -16422
rect -4916 -16825 -3778 -16819
rect -3674 -16422 -2536 -16416
rect -3674 -16819 -3662 -16422
rect -2548 -16819 -2536 -16422
rect -3674 -16825 -2536 -16819
rect -2432 -16422 -1294 -16416
rect -2432 -16819 -2420 -16422
rect -1306 -16819 -1294 -16422
rect -2432 -16825 -1294 -16819
rect -1190 -16422 -52 -16416
rect -1190 -16819 -1178 -16422
rect -64 -16819 -52 -16422
rect -1190 -16825 -52 -16819
rect 52 -16422 1190 -16416
rect 52 -16819 64 -16422
rect 1178 -16819 1190 -16422
rect 52 -16825 1190 -16819
rect 1294 -16422 2432 -16416
rect 1294 -16819 1306 -16422
rect 2420 -16819 2432 -16422
rect 1294 -16825 2432 -16819
rect 2536 -16422 3674 -16416
rect 2536 -16819 2548 -16422
rect 3662 -16819 3674 -16422
rect 2536 -16825 3674 -16819
rect 3778 -16422 4916 -16416
rect 3778 -16819 3790 -16422
rect 4904 -16819 4916 -16422
rect 3778 -16825 4916 -16819
rect -4916 -17929 -3778 -17923
rect -4916 -18326 -4904 -17929
rect -3790 -18326 -3778 -17929
rect -4916 -18332 -3778 -18326
rect -3674 -17929 -2536 -17923
rect -3674 -18326 -3662 -17929
rect -2548 -18326 -2536 -17929
rect -3674 -18332 -2536 -18326
rect -2432 -17929 -1294 -17923
rect -2432 -18326 -2420 -17929
rect -1306 -18326 -1294 -17929
rect -2432 -18332 -1294 -18326
rect -1190 -17929 -52 -17923
rect -1190 -18326 -1178 -17929
rect -64 -18326 -52 -17929
rect -1190 -18332 -52 -18326
rect 52 -17929 1190 -17923
rect 52 -18326 64 -17929
rect 1178 -18326 1190 -17929
rect 52 -18332 1190 -18326
rect 1294 -17929 2432 -17923
rect 1294 -18326 1306 -17929
rect 2420 -18326 2432 -17929
rect 1294 -18332 2432 -18326
rect 2536 -17929 3674 -17923
rect 2536 -18326 2548 -17929
rect 3662 -18326 3674 -17929
rect 2536 -18332 3674 -18326
rect 3778 -17929 4916 -17923
rect 3778 -18326 3790 -17929
rect 4904 -18326 4916 -17929
rect 3778 -18332 4916 -18326
<< properties >>
string FIXED_BBOX -5033 -18457 5033 18457
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 5.542 m 18 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 2.0k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
