magic
tech sky130A
magscale 1 2
timestamp 1683296730
<< nwell >>
rect -100 -1800 1790 1140
<< pwell >>
rect -2660 -20100 4370 -5290
<< psubdiff >>
rect -2610 -5920 -2370 -5896
rect -2610 -6184 -2370 -6160
rect 4090 -5920 4330 -5896
rect 4090 -6184 4330 -6160
rect -2610 -7640 -2370 -7616
rect -2610 -7904 -2370 -7880
rect 4090 -7640 4330 -7616
rect 4090 -7904 4330 -7880
rect -2610 -9360 -2370 -9336
rect -2610 -9624 -2370 -9600
rect 4090 -9360 4330 -9336
rect 4090 -9624 4330 -9600
rect -2610 -10840 -2370 -10816
rect -2610 -11104 -2370 -11080
rect 4090 -10840 4330 -10816
rect 4090 -11104 4330 -11080
rect -2610 -12560 -2370 -12536
rect -2610 -12824 -2370 -12800
rect 4090 -12560 4330 -12536
rect 4090 -12824 4330 -12800
rect -2610 -14160 -2370 -14136
rect -2610 -14424 -2370 -14400
rect 4090 -14160 4330 -14136
rect 4090 -14424 4330 -14400
rect -2610 -15880 -2370 -15856
rect -2610 -16144 -2370 -16120
rect 4090 -15880 4330 -15856
rect 4090 -16144 4330 -16120
rect -2610 -17480 -2370 -17456
rect -2610 -17744 -2370 -17720
rect 4090 -17480 4330 -17456
rect 4090 -17744 4330 -17720
rect -2610 -19200 -2370 -19176
rect -2610 -19464 -2370 -19440
rect 4090 -19200 4330 -19176
rect 4090 -19464 4330 -19440
<< psubdiffcont >>
rect -2610 -6160 -2370 -5920
rect 4090 -6160 4330 -5920
rect -2610 -7880 -2370 -7640
rect 4090 -7880 4330 -7640
rect -2610 -9600 -2370 -9360
rect 4090 -9600 4330 -9360
rect -2610 -11080 -2370 -10840
rect 4090 -11080 4330 -10840
rect -2610 -12800 -2370 -12560
rect 4090 -12800 4330 -12560
rect -2610 -14400 -2370 -14160
rect 4090 -14400 4330 -14160
rect -2610 -16120 -2370 -15880
rect 4090 -16120 4330 -15880
rect -2610 -17720 -2370 -17480
rect 4090 -17720 4330 -17480
rect -2610 -19440 -2370 -19200
rect 4090 -19440 4330 -19200
<< locali >>
rect -2610 -5920 -2370 -5904
rect -2610 -6176 -2370 -6160
rect 4090 -5920 4330 -5904
rect 4090 -6176 4330 -6160
rect -2610 -7640 -2370 -7624
rect -2610 -7896 -2370 -7880
rect 4090 -7640 4330 -7624
rect 4090 -7896 4330 -7880
rect -2610 -9360 -2370 -9344
rect -2610 -9616 -2370 -9600
rect 4090 -9360 4330 -9344
rect 4090 -9616 4330 -9600
rect -2610 -10840 -2370 -10824
rect -2610 -11096 -2370 -11080
rect 4090 -10840 4330 -10824
rect 4090 -11096 4330 -11080
rect -2610 -12560 -2370 -12544
rect -2610 -12816 -2370 -12800
rect 4090 -12560 4330 -12544
rect 4090 -12816 4330 -12800
rect -2610 -14160 -2370 -14144
rect -2610 -14416 -2370 -14400
rect 4090 -14160 4330 -14144
rect 4090 -14416 4330 -14400
rect -2610 -15880 -2370 -15864
rect -2610 -16136 -2370 -16120
rect 4090 -15880 4330 -15864
rect 4090 -16136 4330 -16120
rect -2610 -17480 -2370 -17464
rect -2610 -17736 -2370 -17720
rect 4090 -17480 4330 -17464
rect 4090 -17736 4330 -17720
rect -2610 -19200 -2370 -19184
rect -2610 -19456 -2370 -19440
rect 4090 -19200 4330 -19184
rect 4090 -19456 4330 -19440
<< viali >>
rect -70 300 -30 530
rect 1710 300 1750 530
rect -70 -1210 -30 -980
rect 1710 -1210 1750 -980
rect 530 -2550 570 -2320
rect 1080 -2550 1120 -2320
rect 150 -3360 240 -3270
rect 1410 -3350 1490 -3270
rect 690 -3620 930 -3580
rect 690 -3800 930 -3760
rect 690 -5120 930 -5080
rect -2610 -6160 -2370 -5920
rect 4090 -6160 4330 -5920
rect -2610 -7880 -2370 -7640
rect 4090 -7880 4330 -7640
rect -2610 -9600 -2370 -9360
rect 4090 -9600 4330 -9360
rect -2610 -11080 -2370 -10840
rect 4090 -11080 4330 -10840
rect -2610 -12800 -2370 -12560
rect 4090 -12800 4330 -12560
rect -2610 -14400 -2370 -14160
rect 4090 -14400 4330 -14160
rect -2610 -16120 -2370 -15880
rect 4090 -16120 4330 -15880
rect -2610 -17720 -2370 -17480
rect 4090 -17720 4330 -17480
rect -2610 -19440 -2370 -19200
rect 4090 -19440 4330 -19200
<< metal1 >>
rect -210 960 1890 1010
rect -210 -120 -140 960
rect 20 620 30 700
rect 110 620 120 700
rect 530 620 540 700
rect 620 620 630 700
rect 1050 620 1060 700
rect 1140 620 1150 700
rect 1570 620 1580 700
rect 1660 620 1670 700
rect -80 530 90 550
rect -80 300 -70 530
rect -30 300 90 530
rect -80 280 90 300
rect 1590 530 1760 550
rect 1590 300 1710 530
rect 1750 300 1760 530
rect 1590 280 1760 300
rect 270 140 280 220
rect 360 140 370 220
rect 790 140 800 220
rect 880 140 890 220
rect 1310 140 1320 220
rect 1400 140 1410 220
rect 1820 -120 1890 960
rect -210 -130 1890 -120
rect -210 -170 110 -130
rect 100 -200 110 -170
rect 180 -170 810 -130
rect 180 -200 190 -170
rect 800 -200 810 -170
rect 880 -170 1500 -130
rect 880 -200 890 -170
rect 1490 -200 1500 -170
rect 1570 -170 1890 -130
rect 1570 -200 1580 -170
rect 100 -490 110 -460
rect 90 -530 110 -490
rect 180 -490 190 -460
rect 800 -490 810 -460
rect 180 -530 810 -490
rect 880 -490 890 -460
rect 1490 -490 1500 -460
rect 880 -530 1500 -490
rect 1570 -490 1580 -460
rect 1570 -530 1590 -490
rect 90 -540 1590 -530
rect 300 -700 350 -540
rect 820 -700 870 -540
rect 1330 -700 1380 -540
rect 20 -840 30 -760
rect 110 -840 120 -760
rect 530 -840 540 -760
rect 620 -840 630 -760
rect 1050 -840 1060 -760
rect 1140 -840 1150 -760
rect 1570 -840 1580 -760
rect 1660 -840 1670 -760
rect -240 -980 -20 -960
rect -240 -1060 -180 -980
rect -100 -1060 -70 -980
rect -240 -1120 -70 -1060
rect -240 -1200 -180 -1120
rect -100 -1200 -70 -1120
rect -240 -1210 -70 -1200
rect -30 -1210 -20 -980
rect -240 -1220 -20 -1210
rect 1700 -980 1920 -960
rect 1700 -1210 1710 -980
rect 1750 -1060 1780 -980
rect 1860 -1060 1920 -980
rect 1750 -1120 1920 -1060
rect 1750 -1200 1780 -1120
rect 1860 -1200 1920 -1120
rect 1750 -1210 1920 -1200
rect 1700 -1220 1920 -1210
rect -76 -1222 -24 -1220
rect 1704 -1222 1756 -1220
rect 300 -1620 350 -1460
rect 820 -1620 870 -1450
rect 1330 -1620 1380 -1460
rect -20 -1630 1670 -1620
rect -20 -1730 0 -1630
rect 100 -1670 790 -1630
rect 100 -1730 120 -1670
rect 780 -1700 790 -1670
rect 860 -1670 1550 -1630
rect 860 -1700 870 -1670
rect -20 -1740 120 -1730
rect 1530 -1730 1550 -1670
rect 1650 -1730 1670 -1630
rect 1530 -1740 1670 -1730
rect 780 -2110 790 -2070
rect 640 -2140 790 -2110
rect 860 -2110 870 -2070
rect 860 -2140 1010 -2110
rect 640 -2160 1010 -2140
rect 524 -2320 576 -2308
rect 524 -2380 530 -2320
rect 570 -2380 576 -2320
rect 640 -2350 690 -2160
rect 960 -2350 1010 -2160
rect 1074 -2320 1126 -2308
rect 1074 -2370 1080 -2320
rect 1120 -2370 1126 -2320
rect 450 -2500 460 -2380
rect 580 -2500 590 -2380
rect 1070 -2490 1080 -2370
rect 1200 -2490 1210 -2370
rect 524 -2550 530 -2500
rect 570 -2550 576 -2500
rect 524 -2562 576 -2550
rect 780 -2610 790 -2540
rect 860 -2610 870 -2540
rect 1074 -2550 1080 -2490
rect 1120 -2550 1126 -2490
rect 1074 -2562 1126 -2550
rect 640 -2720 690 -2680
rect 960 -2720 1010 -2680
rect 640 -2770 1010 -2720
rect 270 -3150 280 -3070
rect 360 -3110 370 -3070
rect 780 -3110 790 -3070
rect 360 -3140 790 -3110
rect 860 -3110 870 -3070
rect 1310 -3110 1320 -3070
rect 860 -3140 1320 -3110
rect 360 -3150 1320 -3140
rect 1400 -3150 1410 -3070
rect 270 -3160 1410 -3150
rect 540 -3200 590 -3160
rect 1060 -3190 1110 -3160
rect 130 -3270 360 -3260
rect 1320 -3270 1510 -3260
rect 130 -3360 150 -3270
rect 240 -3360 260 -3270
rect 350 -3360 360 -3270
rect 770 -3360 780 -3270
rect 870 -3360 880 -3270
rect 1280 -3360 1290 -3270
rect 1380 -3350 1410 -3270
rect 1490 -3350 1510 -3270
rect 1380 -3360 1510 -3350
rect 130 -3370 360 -3360
rect 540 -3470 590 -3430
rect 1060 -3470 1110 -3430
rect 330 -3480 1310 -3470
rect 330 -3520 410 -3480
rect 400 -3540 410 -3520
rect 470 -3520 1180 -3480
rect 470 -3540 480 -3520
rect 1170 -3540 1180 -3520
rect 1240 -3520 1310 -3480
rect 1240 -3540 1250 -3520
rect 670 -3580 950 -3570
rect 670 -3620 690 -3580
rect 930 -3620 950 -3580
rect 670 -3650 950 -3620
rect 670 -3740 770 -3650
rect 860 -3740 950 -3650
rect 670 -3760 950 -3740
rect 670 -3800 690 -3760
rect 930 -3800 950 -3760
rect 670 -3810 950 -3800
rect 400 -3860 410 -3840
rect -90 -3900 410 -3860
rect 470 -3860 480 -3840
rect 1170 -3860 1180 -3840
rect 470 -3900 1180 -3860
rect 1240 -3860 1250 -3840
rect 1240 -3900 1740 -3860
rect -90 -3910 1740 -3900
rect -90 -4970 -30 -3910
rect 10 -4270 20 -4210
rect 80 -4270 90 -4210
rect 530 -4270 540 -4210
rect 600 -4270 610 -4210
rect 1040 -4270 1050 -4210
rect 1110 -4270 1120 -4210
rect 1560 -4270 1570 -4210
rect 1630 -4270 1640 -4210
rect 270 -4680 280 -4620
rect 340 -4680 350 -4620
rect 790 -4680 800 -4620
rect 860 -4680 870 -4620
rect 1300 -4680 1310 -4620
rect 1370 -4680 1380 -4620
rect 1680 -4970 1740 -3910
rect -90 -5020 1740 -4970
rect 670 -5080 950 -5070
rect 670 -5120 690 -5080
rect 930 -5120 950 -5080
rect 670 -5180 770 -5120
rect 860 -5180 950 -5120
rect 670 -5190 950 -5180
rect -1220 -5370 3150 -5350
rect -1220 -5430 280 -5370
rect 340 -5430 1310 -5370
rect 1370 -5430 3150 -5370
rect -1220 -5540 3150 -5430
rect -1220 -5600 280 -5540
rect 340 -5600 1310 -5540
rect 1370 -5600 3150 -5540
rect -1220 -5710 3150 -5600
rect -1220 -5770 280 -5710
rect 340 -5770 1310 -5710
rect 1370 -5770 3150 -5710
rect -1220 -5790 3150 -5770
rect -2622 -5920 -2358 -5914
rect -2622 -6160 -2610 -5920
rect -2370 -6160 -2358 -5920
rect -2622 -6166 -2358 -6160
rect 4078 -5920 4342 -5914
rect 4078 -6160 4090 -5920
rect 4330 -6160 4342 -5920
rect 4078 -6166 4342 -6160
rect -2622 -7640 -2358 -7634
rect -2622 -7880 -2610 -7640
rect -2370 -7880 -2358 -7640
rect -2622 -7886 -2358 -7880
rect 4078 -7640 4342 -7634
rect 4078 -7880 4090 -7640
rect 4330 -7880 4342 -7640
rect 4078 -7886 4342 -7880
rect -2622 -9360 -2358 -9354
rect -2622 -9600 -2610 -9360
rect -2370 -9600 -2358 -9360
rect -2622 -9606 -2358 -9600
rect 4078 -9360 4342 -9354
rect 4078 -9600 4090 -9360
rect 4330 -9600 4342 -9360
rect 4078 -9606 4342 -9600
rect -2622 -10840 -2358 -10834
rect -2622 -11080 -2610 -10840
rect -2370 -11080 -2358 -10840
rect -2622 -11086 -2358 -11080
rect 4078 -10840 4342 -10834
rect 4078 -11080 4090 -10840
rect 4330 -11080 4342 -10840
rect 4078 -11086 4342 -11080
rect -2622 -12560 -2358 -12554
rect -2622 -12800 -2610 -12560
rect -2370 -12800 -2358 -12560
rect -2622 -12806 -2358 -12800
rect 4078 -12560 4342 -12554
rect 4078 -12800 4090 -12560
rect 4330 -12800 4342 -12560
rect 4078 -12806 4342 -12800
rect -2622 -14160 -2358 -14154
rect -2622 -14400 -2610 -14160
rect -2370 -14400 -2358 -14160
rect -2622 -14406 -2358 -14400
rect 4078 -14160 4342 -14154
rect 4078 -14400 4090 -14160
rect 4330 -14400 4342 -14160
rect 4078 -14406 4342 -14400
rect -2622 -15880 -2358 -15874
rect -2622 -16120 -2610 -15880
rect -2370 -16120 -2358 -15880
rect -2622 -16126 -2358 -16120
rect 4078 -15880 4342 -15874
rect 4078 -16120 4090 -15880
rect 4330 -16120 4342 -15880
rect 4078 -16126 4342 -16120
rect -2622 -17480 -2358 -17474
rect -2622 -17720 -2610 -17480
rect -2370 -17720 -2358 -17480
rect -2622 -17726 -2358 -17720
rect 4078 -17480 4342 -17474
rect 4078 -17720 4090 -17480
rect 4330 -17720 4342 -17480
rect 4078 -17726 4342 -17720
rect -2622 -19200 -2358 -19194
rect -2622 -19440 -2610 -19200
rect -2370 -19440 -2358 -19200
rect -2622 -19446 -2358 -19440
rect 4078 -19200 4342 -19194
rect 4078 -19440 4090 -19200
rect 4330 -19440 4342 -19200
rect 4078 -19446 4342 -19440
rect -2630 -19680 4350 -19580
rect -2630 -19920 -2610 -19680
rect -2370 -19920 4090 -19680
rect 4330 -19920 4350 -19680
rect -2630 -20020 4350 -19920
<< via1 >>
rect 30 620 110 700
rect 540 620 620 700
rect 1060 620 1140 700
rect 1580 620 1660 700
rect 280 140 360 220
rect 800 140 880 220
rect 1320 140 1400 220
rect 110 -200 180 -130
rect 810 -200 880 -130
rect 1500 -200 1570 -130
rect 110 -530 180 -460
rect 810 -530 880 -460
rect 1500 -530 1570 -460
rect 30 -840 110 -760
rect 540 -840 620 -760
rect 1060 -840 1140 -760
rect 1580 -840 1660 -760
rect -180 -1060 -100 -980
rect -180 -1200 -100 -1120
rect 1780 -1060 1860 -980
rect 1780 -1200 1860 -1120
rect 0 -1730 100 -1630
rect 790 -1700 860 -1630
rect 1550 -1730 1650 -1630
rect 790 -2140 860 -2070
rect 460 -2500 530 -2380
rect 530 -2500 570 -2380
rect 570 -2500 580 -2380
rect 1080 -2490 1120 -2370
rect 1120 -2490 1200 -2370
rect 790 -2610 860 -2540
rect 280 -3150 360 -3070
rect 790 -3140 860 -3070
rect 1320 -3150 1400 -3070
rect 260 -3360 350 -3270
rect 780 -3360 870 -3270
rect 1290 -3360 1380 -3270
rect 410 -3540 470 -3480
rect 1180 -3540 1240 -3480
rect 770 -3740 860 -3650
rect 410 -3900 470 -3840
rect 1180 -3900 1240 -3840
rect 20 -4270 80 -4210
rect 540 -4270 600 -4210
rect 1050 -4270 1110 -4210
rect 1570 -4270 1630 -4210
rect 280 -4680 340 -4620
rect 800 -4680 860 -4620
rect 1310 -4680 1370 -4620
rect 770 -5120 860 -5090
rect 770 -5180 860 -5120
rect 280 -5430 340 -5370
rect 1310 -5430 1370 -5370
rect 280 -5600 340 -5540
rect 1310 -5600 1370 -5540
rect 280 -5770 340 -5710
rect 1310 -5770 1370 -5710
rect -2610 -6160 -2370 -5920
rect 4090 -6160 4330 -5920
rect -2610 -7880 -2370 -7640
rect 4090 -7880 4330 -7640
rect -2610 -9600 -2370 -9360
rect 4090 -9600 4330 -9360
rect -2610 -11080 -2370 -10840
rect 4090 -11080 4330 -10840
rect -2610 -12800 -2370 -12560
rect 4090 -12800 4330 -12560
rect -2610 -14400 -2370 -14160
rect 4090 -14400 4330 -14160
rect -2610 -16120 -2370 -15880
rect 4090 -16120 4330 -15880
rect -2610 -17720 -2370 -17480
rect 4090 -17720 4330 -17480
rect -2610 -19440 -2370 -19200
rect 4090 -19440 4330 -19200
rect -2610 -19920 -2370 -19680
rect 4090 -19920 4330 -19680
<< metal2 >>
rect 30 700 110 710
rect 30 610 110 620
rect 540 700 620 710
rect 540 610 620 620
rect 1060 700 1140 710
rect 1060 610 1140 620
rect 1580 700 1660 710
rect 1580 610 1660 620
rect 270 220 370 230
rect 270 140 280 220
rect 360 140 370 220
rect 90 -130 200 -120
rect 90 -200 110 -130
rect 180 -200 200 -130
rect 90 -460 200 -200
rect 90 -530 110 -460
rect 180 -530 200 -460
rect 90 -540 200 -530
rect 30 -760 110 -750
rect 30 -850 110 -840
rect -180 -980 -100 -970
rect -180 -1070 -100 -1060
rect -180 -1120 -100 -1110
rect -180 -1210 -100 -1200
rect -20 -1630 120 -1620
rect -20 -1730 0 -1630
rect 100 -1730 120 -1630
rect -20 -4210 120 -1730
rect 270 -3070 370 140
rect 800 220 880 230
rect 800 130 880 140
rect 1310 220 1410 230
rect 1310 140 1320 220
rect 1400 140 1410 220
rect 790 -130 900 -120
rect 790 -200 810 -130
rect 880 -200 900 -130
rect 790 -460 900 -200
rect 790 -530 810 -460
rect 880 -530 900 -460
rect 790 -540 900 -530
rect 540 -760 620 -750
rect 540 -850 620 -840
rect 1060 -760 1140 -750
rect 1060 -850 1140 -840
rect 780 -1630 870 -1620
rect 780 -1700 790 -1630
rect 860 -1700 870 -1630
rect 780 -2070 870 -1700
rect 780 -2140 790 -2070
rect 860 -2140 870 -2070
rect 780 -2150 870 -2140
rect 1080 -2370 1200 -2360
rect 460 -2380 580 -2370
rect 1080 -2500 1200 -2490
rect 460 -2510 580 -2500
rect 270 -3150 280 -3070
rect 360 -3150 370 -3070
rect 780 -2540 870 -2530
rect 780 -2610 790 -2540
rect 860 -2610 870 -2540
rect 780 -3070 870 -2610
rect 780 -3110 790 -3070
rect 860 -3110 870 -3070
rect 1310 -3070 1410 140
rect 1480 -130 1590 -120
rect 1480 -200 1500 -130
rect 1570 -200 1590 -130
rect 1480 -460 1590 -200
rect 1480 -530 1500 -460
rect 1570 -530 1590 -460
rect 1480 -540 1590 -530
rect 1580 -760 1660 -750
rect 1580 -850 1660 -840
rect 1780 -980 1860 -970
rect 1780 -1070 1860 -1060
rect 1780 -1120 1860 -1110
rect 1780 -1210 1860 -1200
rect 790 -3150 860 -3140
rect 1310 -3150 1320 -3070
rect 1400 -3150 1410 -3070
rect 270 -3160 370 -3150
rect 1310 -3160 1410 -3150
rect 1530 -1630 1670 -1620
rect 1530 -1730 1550 -1630
rect 1650 -1730 1670 -1630
rect 260 -3270 350 -3260
rect 260 -3370 350 -3360
rect 780 -3270 870 -3260
rect 780 -3370 870 -3360
rect 1290 -3270 1380 -3260
rect 1290 -3370 1380 -3360
rect 400 -3480 480 -3470
rect 400 -3540 410 -3480
rect 470 -3540 480 -3480
rect 400 -3840 480 -3540
rect 1170 -3480 1250 -3470
rect 1170 -3540 1180 -3480
rect 1240 -3540 1250 -3480
rect 770 -3650 860 -3640
rect 770 -3750 860 -3740
rect 400 -3900 410 -3840
rect 470 -3900 480 -3840
rect 400 -3910 480 -3900
rect 1170 -3840 1250 -3540
rect 1170 -3900 1180 -3840
rect 1240 -3900 1250 -3840
rect 1170 -3910 1250 -3900
rect -20 -4270 20 -4210
rect 80 -4270 120 -4210
rect -20 -4280 120 -4270
rect 540 -4210 600 -4200
rect 540 -4280 600 -4270
rect 1050 -4210 1110 -4200
rect 1050 -4280 1110 -4270
rect 1530 -4210 1670 -1730
rect 1530 -4270 1570 -4210
rect 1630 -4270 1670 -4210
rect 1530 -4280 1670 -4270
rect 260 -4620 360 -4610
rect 260 -4680 280 -4620
rect 340 -4680 360 -4620
rect 260 -5370 360 -4680
rect 800 -4620 860 -4610
rect 800 -4690 860 -4680
rect 1290 -4620 1390 -4610
rect 1290 -4680 1310 -4620
rect 1370 -4680 1390 -4620
rect 770 -5090 860 -5080
rect 770 -5190 860 -5180
rect 260 -5430 280 -5370
rect 340 -5430 360 -5370
rect 260 -5540 360 -5430
rect 260 -5600 280 -5540
rect 340 -5600 360 -5540
rect 260 -5710 360 -5600
rect 260 -5770 280 -5710
rect 340 -5770 360 -5710
rect 260 -5790 360 -5770
rect 1290 -5370 1390 -4680
rect 1290 -5430 1310 -5370
rect 1370 -5430 1390 -5370
rect 1290 -5540 1390 -5430
rect 1290 -5600 1310 -5540
rect 1370 -5600 1390 -5540
rect 1290 -5710 1390 -5600
rect 1290 -5770 1310 -5710
rect 1370 -5770 1390 -5710
rect 1290 -5790 1390 -5770
rect -2630 -5920 -2350 -5880
rect -2630 -6160 -2610 -5920
rect -2370 -6160 -2350 -5920
rect -2630 -7640 -2350 -6160
rect -2630 -7880 -2610 -7640
rect -2370 -7880 -2350 -7640
rect -2630 -9360 -2350 -7880
rect -2630 -9600 -2610 -9360
rect -2370 -9600 -2350 -9360
rect -2630 -10840 -2350 -9600
rect -2630 -11080 -2610 -10840
rect -2370 -11080 -2350 -10840
rect -2630 -12560 -2350 -11080
rect -2630 -12800 -2610 -12560
rect -2370 -12800 -2350 -12560
rect -2630 -14160 -2350 -12800
rect -2630 -14400 -2610 -14160
rect -2370 -14400 -2350 -14160
rect -2630 -15880 -2350 -14400
rect -2630 -16120 -2610 -15880
rect -2370 -16120 -2350 -15880
rect -2630 -17480 -2350 -16120
rect -2630 -17720 -2610 -17480
rect -2370 -17720 -2350 -17480
rect -2630 -19200 -2350 -17720
rect -2630 -19440 -2610 -19200
rect -2370 -19440 -2350 -19200
rect -2630 -19680 -2350 -19440
rect -2630 -19920 -2610 -19680
rect -2370 -19920 -2350 -19680
rect -2630 -20020 -2350 -19920
rect 4070 -5920 4350 -5880
rect 4070 -6160 4090 -5920
rect 4330 -6160 4350 -5920
rect 4070 -7640 4350 -6160
rect 4070 -7880 4090 -7640
rect 4330 -7880 4350 -7640
rect 4070 -9360 4350 -7880
rect 4070 -9600 4090 -9360
rect 4330 -9600 4350 -9360
rect 4070 -10840 4350 -9600
rect 4070 -11080 4090 -10840
rect 4330 -11080 4350 -10840
rect 4070 -12560 4350 -11080
rect 4070 -12800 4090 -12560
rect 4330 -12800 4350 -12560
rect 4070 -14160 4350 -12800
rect 4070 -14400 4090 -14160
rect 4330 -14400 4350 -14160
rect 4070 -15880 4350 -14400
rect 4070 -16120 4090 -15880
rect 4330 -16120 4350 -15880
rect 4070 -17480 4350 -16120
rect 4070 -17720 4090 -17480
rect 4330 -17720 4350 -17480
rect 4070 -19200 4350 -17720
rect 4070 -19440 4090 -19200
rect 4330 -19440 4350 -19200
rect 4070 -19680 4350 -19440
rect 4070 -19920 4090 -19680
rect 4330 -19920 4350 -19680
rect 4070 -20020 4350 -19920
<< via2 >>
rect 30 620 110 700
rect 540 620 620 700
rect 1060 620 1140 700
rect 1580 620 1660 700
rect 280 140 360 220
rect 30 -840 110 -760
rect -180 -1060 -100 -980
rect -180 -1200 -100 -1120
rect 800 140 880 220
rect 1320 140 1400 220
rect 540 -840 620 -760
rect 1060 -840 1140 -760
rect 460 -2500 580 -2380
rect 1080 -2490 1200 -2370
rect 1580 -840 1660 -760
rect 1780 -1060 1860 -980
rect 1780 -1200 1860 -1120
rect 260 -3360 350 -3270
rect 780 -3360 870 -3270
rect 1290 -3360 1380 -3270
rect 770 -3740 860 -3650
rect 20 -4270 80 -4210
rect 540 -4270 600 -4210
rect 1050 -4270 1110 -4210
rect 1570 -4270 1630 -4210
rect 280 -4680 340 -4620
rect 800 -4680 860 -4620
rect 1310 -4680 1370 -4620
rect 770 -5180 860 -5090
rect -2610 -6160 -2370 -5920
rect -2610 -7880 -2370 -7640
rect -2610 -9600 -2370 -9360
rect -2610 -11080 -2370 -10840
rect -2610 -12800 -2370 -12560
rect -2610 -14400 -2370 -14160
rect -2610 -16120 -2370 -15880
rect -2610 -17720 -2370 -17480
rect -2610 -19440 -2370 -19200
rect 4090 -6160 4330 -5920
rect 4090 -7880 4330 -7640
rect 4090 -9600 4330 -9360
rect 4090 -11080 4330 -10840
rect 4090 -12800 4330 -12560
rect 4090 -14400 4330 -14160
rect 4090 -16120 4330 -15880
rect 4090 -17720 4330 -17480
rect 4090 -19440 4330 -19200
<< metal3 >>
rect -10 600 0 720
rect 120 700 1670 720
rect 120 620 540 700
rect 620 620 1060 700
rect 1140 620 1580 700
rect 1660 620 1670 700
rect 120 600 1670 620
rect 40 220 1640 240
rect 40 140 280 220
rect 360 140 800 220
rect 880 140 1320 220
rect 1400 140 1640 220
rect 40 120 1640 140
rect -240 -760 1920 -740
rect -240 -840 -180 -760
rect -100 -840 30 -760
rect 110 -840 540 -760
rect 620 -840 1060 -760
rect 1140 -840 1580 -760
rect 1660 -840 1780 -760
rect 1860 -840 1920 -760
rect -240 -860 1920 -840
rect -200 -980 -80 -960
rect -200 -1060 -180 -980
rect -100 -1060 -80 -980
rect -200 -1120 -80 -1060
rect -200 -1200 -180 -1120
rect -100 -1200 -80 -1120
rect -200 -1220 -80 -1200
rect 1760 -980 1880 -960
rect 1760 -1060 1780 -980
rect 1860 -1060 1880 -980
rect 1760 -1120 1880 -1060
rect 1760 -1200 1780 -1120
rect 1860 -1200 1880 -1120
rect 1760 -1220 1880 -1200
rect 1070 -2370 1210 -2365
rect 450 -2380 590 -2375
rect 450 -2500 460 -2380
rect 580 -2500 590 -2380
rect 1070 -2490 1080 -2370
rect 1200 -2490 1210 -2370
rect 1070 -2495 1210 -2490
rect 450 -2505 590 -2500
rect 240 -3270 1400 -3250
rect 240 -3360 260 -3270
rect 350 -3360 780 -3270
rect 870 -3360 1290 -3270
rect 1380 -3360 1400 -3270
rect 240 -3380 1400 -3360
rect 760 -3650 870 -3645
rect 760 -3740 770 -3650
rect 860 -3740 870 -3650
rect 760 -3745 870 -3740
rect 10 -4210 1640 -4200
rect 10 -4270 20 -4210
rect 80 -4270 540 -4210
rect 600 -4270 1050 -4210
rect 1110 -4270 1570 -4210
rect 1630 -4270 1640 -4210
rect 10 -4280 1640 -4270
rect 30 -4620 1620 -4610
rect 30 -4680 280 -4620
rect 340 -4680 800 -4620
rect 860 -4680 1310 -4620
rect 1370 -4680 1620 -4620
rect 30 -4690 1620 -4680
rect 760 -5090 870 -5085
rect 760 -5180 770 -5090
rect 860 -5180 870 -5090
rect 760 -5185 870 -5180
rect -2620 -5920 -2360 -5915
rect -2620 -6160 -2610 -5920
rect -2370 -6160 -2360 -5920
rect -2620 -6165 -2360 -6160
rect 4080 -5920 4340 -5915
rect 4080 -6160 4090 -5920
rect 4330 -6160 4340 -5920
rect 4080 -6165 4340 -6160
rect -2620 -7640 -2360 -7635
rect -2620 -7880 -2610 -7640
rect -2370 -7880 -2360 -7640
rect -2620 -7885 -2360 -7880
rect 4080 -7640 4340 -7635
rect 4080 -7880 4090 -7640
rect 4330 -7880 4340 -7640
rect 4080 -7885 4340 -7880
rect -2620 -9360 -2360 -9355
rect -2620 -9600 -2610 -9360
rect -2370 -9600 -2360 -9360
rect -2620 -9605 -2360 -9600
rect 4080 -9360 4340 -9355
rect 4080 -9600 4090 -9360
rect 4330 -9600 4340 -9360
rect 4080 -9605 4340 -9600
rect -2620 -10840 -2360 -10835
rect -2620 -11080 -2610 -10840
rect -2370 -11080 -2360 -10840
rect -2620 -11085 -2360 -11080
rect 4080 -10840 4340 -10835
rect 4080 -11080 4090 -10840
rect 4330 -11080 4340 -10840
rect 4080 -11085 4340 -11080
rect -2620 -12560 -2360 -12555
rect -2620 -12800 -2610 -12560
rect -2370 -12800 -2360 -12560
rect -2620 -12805 -2360 -12800
rect 4080 -12560 4340 -12555
rect 4080 -12800 4090 -12560
rect 4330 -12800 4340 -12560
rect 4080 -12805 4340 -12800
rect -2620 -14160 -2360 -14155
rect -2620 -14400 -2610 -14160
rect -2370 -14400 -2360 -14160
rect -2620 -14405 -2360 -14400
rect 4080 -14160 4340 -14155
rect 4080 -14400 4090 -14160
rect 4330 -14400 4340 -14160
rect 4080 -14405 4340 -14400
rect -2620 -15880 -2360 -15875
rect -2620 -16120 -2610 -15880
rect -2370 -16120 -2360 -15880
rect -2620 -16125 -2360 -16120
rect 4080 -15880 4340 -15875
rect 4080 -16120 4090 -15880
rect 4330 -16120 4340 -15880
rect 4080 -16125 4340 -16120
rect -2620 -17480 -2360 -17475
rect -2620 -17720 -2610 -17480
rect -2370 -17720 -2360 -17480
rect -2620 -17725 -2360 -17720
rect 4080 -17480 4340 -17475
rect 4080 -17720 4090 -17480
rect 4330 -17720 4340 -17480
rect 4080 -17725 4340 -17720
rect -2620 -19200 -2360 -19195
rect -2620 -19440 -2610 -19200
rect -2370 -19440 -2360 -19200
rect -2620 -19445 -2360 -19440
rect 4080 -19200 4340 -19195
rect 4080 -19440 4090 -19200
rect 4330 -19440 4340 -19200
rect 4080 -19445 4340 -19440
<< via3 >>
rect 0 700 120 720
rect 0 620 30 700
rect 30 620 110 700
rect 110 620 120 700
rect 540 620 620 700
rect 1060 620 1140 700
rect 1580 620 1660 700
rect 0 600 120 620
rect -180 -840 -100 -760
rect 1780 -840 1860 -760
rect -180 -1060 -100 -980
rect -180 -1200 -100 -1120
rect 1780 -1060 1860 -980
rect 1780 -1200 1860 -1120
rect 460 -2500 580 -2380
rect 1080 -2490 1200 -2370
rect 780 -3360 870 -3270
rect 770 -3740 860 -3650
rect 770 -5180 860 -5090
rect -2610 -9600 -2370 -9360
rect 4090 -9600 4330 -9360
rect -2610 -12800 -2370 -12560
rect 4090 -12800 4330 -12560
rect -2610 -16120 -2370 -15880
rect 4090 -16120 4330 -15880
<< metal4 >>
rect -240 540 -60 780
rect 1740 540 1920 780
rect -240 -760 -20 540
rect -240 -840 -180 -760
rect -100 -840 -20 -760
rect -240 -980 -20 -840
rect -240 -1060 -180 -980
rect -100 -1060 -20 -980
rect -240 -1120 -20 -1060
rect -240 -1200 -180 -1120
rect -100 -1200 -20 -1120
rect -240 -1220 -20 -1200
rect 1700 -760 1920 540
rect 1700 -840 1780 -760
rect 1860 -840 1920 -760
rect 1700 -980 1920 -840
rect 1700 -1060 1780 -980
rect 1860 -1060 1920 -980
rect 1700 -1120 1920 -1060
rect 1700 -1200 1780 -1120
rect 1860 -1200 1920 -1120
rect 1700 -1220 1920 -1200
rect 320 -2370 1280 -2200
rect 320 -2380 1080 -2370
rect 320 -2500 460 -2380
rect 580 -2490 1080 -2380
rect 1200 -2490 1280 -2370
rect 580 -2500 1280 -2490
rect 320 -3270 1280 -2500
rect 320 -3360 780 -3270
rect 870 -3360 1280 -3270
rect 320 -3650 1280 -3360
rect 320 -3740 770 -3650
rect 860 -3740 1280 -3650
rect 320 -5090 1280 -3740
rect 320 -5180 770 -5090
rect 860 -5180 1280 -5090
rect 320 -8880 1280 -5180
rect 320 -9120 400 -8880
rect 640 -9120 960 -8880
rect 1200 -9120 1280 -8880
rect -2611 -9360 -2369 -9359
rect -2611 -9600 -2610 -9360
rect -2370 -9600 -2369 -9360
rect -2611 -9601 -2369 -9600
rect 320 -9360 1280 -9120
rect 320 -9600 400 -9360
rect 640 -9600 960 -9360
rect 1200 -9600 1280 -9360
rect 320 -9840 1280 -9600
rect 4089 -9360 4331 -9359
rect 4089 -9600 4090 -9360
rect 4330 -9600 4331 -9360
rect 4089 -9601 4331 -9600
rect 320 -10080 400 -9840
rect 640 -10080 960 -9840
rect 1200 -10080 1280 -9840
rect 320 -12080 1280 -10080
rect 320 -12320 400 -12080
rect 640 -12320 960 -12080
rect 1200 -12320 1280 -12080
rect -2611 -12560 -2369 -12559
rect -2611 -12800 -2610 -12560
rect -2370 -12800 -2369 -12560
rect -2611 -12801 -2369 -12800
rect 320 -12560 1280 -12320
rect 320 -12800 400 -12560
rect 640 -12800 960 -12560
rect 1200 -12800 1280 -12560
rect 320 -13040 1280 -12800
rect 4089 -12560 4331 -12559
rect 4089 -12800 4090 -12560
rect 4330 -12800 4331 -12560
rect 4089 -12801 4331 -12800
rect 320 -13280 400 -13040
rect 640 -13280 960 -13040
rect 1200 -13280 1280 -13040
rect 320 -15400 1280 -13280
rect 320 -15640 400 -15400
rect 640 -15640 960 -15400
rect 1200 -15640 1280 -15400
rect -2611 -15880 -2369 -15879
rect -2611 -16120 -2610 -15880
rect -2370 -16120 -2369 -15880
rect -2611 -16121 -2369 -16120
rect 320 -15880 1280 -15640
rect 320 -16120 400 -15880
rect 640 -16120 960 -15880
rect 1200 -16120 1280 -15880
rect 320 -16360 1280 -16120
rect 4089 -15880 4331 -15879
rect 4089 -16120 4090 -15880
rect 4330 -16120 4331 -15880
rect 4089 -16121 4331 -16120
rect 320 -16600 400 -16360
rect 640 -16600 960 -16360
rect 1200 -16600 1280 -16360
rect 320 -16680 1280 -16600
<< via4 >>
rect -60 720 180 780
rect -60 600 0 720
rect 0 600 120 720
rect 120 600 180 720
rect -60 540 180 600
rect 460 700 700 780
rect 460 620 540 700
rect 540 620 620 700
rect 620 620 700 700
rect 460 540 700 620
rect 980 700 1220 780
rect 980 620 1060 700
rect 1060 620 1140 700
rect 1140 620 1220 700
rect 980 540 1220 620
rect 1500 700 1740 780
rect 1500 620 1580 700
rect 1580 620 1660 700
rect 1660 620 1740 700
rect 1500 540 1740 620
rect 400 -9120 640 -8880
rect 960 -9120 1200 -8880
rect -2610 -9600 -2370 -9360
rect 400 -9600 640 -9360
rect 960 -9600 1200 -9360
rect 4090 -9600 4330 -9360
rect 400 -10080 640 -9840
rect 960 -10080 1200 -9840
rect 400 -12320 640 -12080
rect 960 -12320 1200 -12080
rect -2610 -12800 -2370 -12560
rect 400 -12800 640 -12560
rect 960 -12800 1200 -12560
rect 4090 -12800 4330 -12560
rect 400 -13280 640 -13040
rect 960 -13280 1200 -13040
rect 400 -15640 640 -15400
rect 960 -15640 1200 -15400
rect -2610 -16120 -2370 -15880
rect 400 -16120 640 -15880
rect 960 -16120 1200 -15880
rect 4090 -16120 4330 -15880
rect 400 -16600 640 -16360
rect 960 -16600 1200 -16360
<< metal5 >>
rect -320 780 2040 1120
rect -320 540 -60 780
rect 180 540 460 780
rect 700 540 980 780
rect 1220 540 1500 780
rect 1740 540 2040 780
rect -320 480 2040 540
rect -2690 -8880 4420 -8790
rect -2690 -9120 400 -8880
rect 640 -9120 960 -8880
rect 1200 -9120 4420 -8880
rect -2690 -9360 4420 -9120
rect -2690 -9600 -2610 -9360
rect -2370 -9600 400 -9360
rect 640 -9600 960 -9360
rect 1200 -9600 4090 -9360
rect 4330 -9600 4420 -9360
rect -2690 -9840 4420 -9600
rect -2690 -10080 400 -9840
rect 640 -10080 960 -9840
rect 1200 -10080 4420 -9840
rect -2690 -10160 4420 -10080
rect -2700 -12080 4410 -12000
rect -2700 -12320 400 -12080
rect 640 -12320 960 -12080
rect 1200 -12320 4410 -12080
rect -2700 -12560 4410 -12320
rect -2700 -12800 -2610 -12560
rect -2370 -12800 400 -12560
rect 640 -12800 960 -12560
rect 1200 -12800 4090 -12560
rect 4330 -12800 4410 -12560
rect -2700 -13040 4410 -12800
rect -2700 -13280 400 -13040
rect 640 -13280 960 -13040
rect 1200 -13280 4410 -13040
rect -2700 -13370 4410 -13280
rect -2690 -15400 4410 -15320
rect -2690 -15640 400 -15400
rect 640 -15640 960 -15400
rect 1200 -15640 4410 -15400
rect -2690 -15880 4410 -15640
rect -2690 -16120 -2610 -15880
rect -2370 -16120 400 -15880
rect 640 -16120 960 -15880
rect 1200 -16120 4090 -15880
rect 4330 -16120 4410 -15880
rect -2690 -16360 4410 -16120
rect -2690 -16600 400 -16360
rect 640 -16600 960 -16360
rect 1200 -16600 4410 -16360
rect -2690 -16680 4410 -16600
use sky130_fd_pr__nfet_01v8_A5635U  sky130_fd_pr__nfet_01v8_A5635U_0
timestamp 1682745745
transform 1 0 823 0 1 -3315
box -683 -335 683 335
use sky130_fd_pr__nfet_01v8_GLZPWL  sky130_fd_pr__nfet_01v8_GLZPWL_0
timestamp 1682745745
transform 1 0 826 0 1 -4440
box -941 -710 941 710
use sky130_fd_pr__nfet_01v8_H7FLKU  sky130_fd_pr__nfet_01v8_H7FLKU_0
timestamp 1682745745
transform 1 0 825 0 1 -2440
box -325 -460 325 460
use sky130_fd_pr__pfet_01v8_LK874N  sky130_fd_pr__pfet_01v8_LK874N_0
timestamp 1682745745
transform 1 0 841 0 1 419
box -941 -719 941 719
use sky130_fd_pr__pfet_01v8_LK874N  sky130_fd_pr__pfet_01v8_LK874N_1
timestamp 1682745745
transform 1 0 841 0 1 -1081
box -941 -719 941 719
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_0
timestamp 1677346452
transform 1 0 1575 0 1 -12688
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_1
timestamp 1677346452
transform 1 0 35 0 1 -12688
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_2
timestamp 1677346452
transform 1 0 -1515 0 1 -12688
box -575 -7332 575 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_3
timestamp 1677346452
transform 1 0 3125 0 1 -12688
box -575 -7332 575 7332
<< labels >>
rlabel metal5 -438 -12860 -438 -12860 1 VSS
port 1 n
rlabel metal3 582 184 582 184 1 Vout
port 2 n
rlabel metal5 290 1000 290 1000 1 VDD
port 3 n
<< end >>
