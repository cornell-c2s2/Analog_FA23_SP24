magic
tech sky130A
magscale 1 2
timestamp 1713414733
<< error_s >>
rect 15660 -2540 16100 -2110
rect 10670 -9901 19302 -9580
rect 11973 -10115 11996 -9985
rect 12026 -10115 12080 -9985
rect 12110 -10115 12164 -9985
rect 12194 -10115 12248 -9985
rect 12278 -10115 12332 -9985
rect 12362 -10115 12416 -9985
rect 12446 -10115 12500 -9985
rect 12530 -10115 12584 -9985
rect 12614 -10115 12668 -9985
rect 12698 -10115 12752 -9985
rect 12782 -10115 12836 -9985
rect 12866 -10115 12920 -9985
rect 12950 -10115 13004 -9985
rect 13034 -10115 13088 -9985
rect 13118 -10115 13172 -9985
rect 13202 -10115 13256 -9985
rect 13286 -10115 13338 -9985
rect 13416 -10115 13468 -9985
rect 13498 -10115 13552 -9985
rect 13582 -10115 13636 -9985
rect 13666 -10115 13720 -9985
rect 13750 -10115 13804 -9985
rect 13834 -10115 13888 -9985
rect 13918 -10115 13972 -9985
rect 14002 -10115 14056 -9985
rect 14086 -10115 14140 -9985
rect 14170 -10115 14224 -9985
rect 14254 -10115 14308 -9985
rect 14338 -10115 14392 -9985
rect 14422 -10115 14476 -9985
rect 14506 -10115 14560 -9985
rect 14590 -10115 14644 -9985
rect 14674 -10115 14728 -9985
rect 14758 -10115 14810 -9985
rect 14888 -10115 14940 -9985
rect 14970 -10115 15024 -9985
rect 15054 -10115 15108 -9985
rect 15138 -10115 15192 -9985
rect 15222 -10115 15276 -9985
rect 15306 -10115 15360 -9985
rect 15390 -10115 15444 -9985
rect 15474 -10115 15528 -9985
rect 15558 -10115 15612 -9985
rect 15642 -10115 15696 -9985
rect 15726 -10115 15780 -9985
rect 15810 -10115 15864 -9985
rect 15894 -10115 15948 -9985
rect 15978 -10115 16032 -9985
rect 16062 -10115 16116 -9985
rect 16146 -10115 16200 -9985
rect 16230 -10115 16282 -9985
rect 16360 -10115 16412 -9985
rect 16442 -10115 16496 -9985
rect 16526 -10115 16580 -9985
rect 16610 -10115 16664 -9985
rect 16694 -10115 16748 -9985
rect 16778 -10115 16832 -9985
rect 16862 -10115 16916 -9985
rect 16946 -10115 17000 -9985
rect 17030 -10115 17084 -9985
rect 17114 -10115 17168 -9985
rect 17198 -10115 17252 -9985
rect 17282 -10115 17336 -9985
rect 17366 -10115 17420 -9985
rect 17450 -10115 17504 -9985
rect 17534 -10115 17588 -9985
rect 17618 -10115 17672 -9985
rect 17702 -10115 17754 -9985
rect 10670 -11551 19302 -11230
rect 10945 -11681 10997 -11635
rect 10764 -11765 10816 -11681
rect 10846 -11765 10900 -11681
rect 10930 -11765 10997 -11681
rect 11027 -11765 11079 -11635
rect 11236 -11765 11288 -11635
rect 11318 -11765 11370 -11635
rect 11481 -11765 11533 -11635
rect 11563 -11765 11617 -11635
rect 11647 -11765 11701 -11635
rect 11731 -11765 11785 -11635
rect 11815 -11765 11867 -11635
rect 11944 -11765 11996 -11635
rect 12026 -11765 12080 -11635
rect 12110 -11765 12164 -11635
rect 12194 -11765 12248 -11635
rect 12278 -11765 12332 -11635
rect 12362 -11765 12416 -11635
rect 12446 -11765 12500 -11635
rect 12530 -11765 12584 -11635
rect 12614 -11765 12668 -11635
rect 12698 -11765 12752 -11635
rect 12782 -11765 12836 -11635
rect 12866 -11765 12920 -11635
rect 12950 -11765 13004 -11635
rect 13034 -11765 13088 -11635
rect 13118 -11765 13172 -11635
rect 13202 -11765 13256 -11635
rect 13286 -11765 13338 -11635
rect 13416 -11765 13468 -11635
rect 13498 -11765 13552 -11635
rect 13582 -11765 13636 -11635
rect 13666 -11765 13720 -11635
rect 13750 -11765 13804 -11635
rect 13834 -11765 13888 -11635
rect 13918 -11765 13972 -11635
rect 14002 -11765 14056 -11635
rect 14086 -11765 14140 -11635
rect 14170 -11765 14224 -11635
rect 14254 -11765 14308 -11635
rect 14338 -11765 14392 -11635
rect 14422 -11765 14476 -11635
rect 14506 -11765 14560 -11635
rect 14590 -11765 14644 -11635
rect 14674 -11765 14728 -11635
rect 14758 -11765 14810 -11635
rect 14888 -11765 14940 -11635
rect 14970 -11765 15024 -11635
rect 15054 -11765 15108 -11635
rect 15138 -11765 15192 -11635
rect 15222 -11765 15276 -11635
rect 15306 -11765 15360 -11635
rect 15390 -11765 15444 -11635
rect 15474 -11765 15528 -11635
rect 15558 -11765 15612 -11635
rect 15642 -11765 15696 -11635
rect 15726 -11765 15780 -11635
rect 15810 -11765 15864 -11635
rect 15894 -11765 15948 -11635
rect 15978 -11765 16032 -11635
rect 16062 -11765 16116 -11635
rect 16146 -11765 16200 -11635
rect 16230 -11765 16282 -11635
rect 16360 -11765 16412 -11635
rect 16442 -11765 16496 -11635
rect 16526 -11765 16580 -11635
rect 16610 -11765 16664 -11635
rect 16694 -11765 16748 -11635
rect 16778 -11765 16832 -11635
rect 16862 -11765 16916 -11635
rect 16946 -11765 17000 -11635
rect 17030 -11765 17084 -11635
rect 17114 -11765 17168 -11635
rect 17198 -11765 17252 -11635
rect 17282 -11765 17336 -11635
rect 17366 -11765 17420 -11635
rect 17450 -11765 17504 -11635
rect 17534 -11765 17588 -11635
rect 17618 -11765 17672 -11635
rect 17702 -11765 17754 -11635
rect 17832 -11765 17884 -11635
rect 17914 -11765 17968 -11635
rect 17998 -11765 18052 -11635
rect 18082 -11765 18136 -11635
rect 18166 -11765 18220 -11635
rect 18250 -11765 18304 -11635
rect 18334 -11765 18388 -11635
rect 18418 -11765 18472 -11635
rect 18502 -11765 18556 -11635
rect 18586 -11765 18640 -11635
rect 18670 -11765 18724 -11635
rect 18754 -11765 18808 -11635
rect 18838 -11765 18892 -11635
rect 18922 -11765 18976 -11635
rect 19006 -11765 19060 -11635
rect 19090 -11765 19144 -11635
rect 19174 -11765 19226 -11635
<< nwell >>
rect 12570 -540 13530 350
rect 8560 -1270 16750 -540
rect 8610 -2410 8980 -1850
rect 15660 -2540 16100 -2110
rect 10660 -7770 19310 -7210
<< pwell >>
rect 8600 -1810 16750 -1310
rect 10870 -2160 11510 -1810
rect 15670 -1850 16710 -1810
rect 16350 -2140 16710 -1850
rect 10660 -8280 19310 -7810
<< pdiff >>
rect 10640 -1190 10700 -1140
<< psubdiff >>
rect 10360 -1640 10530 -1610
rect 9460 -1670 9630 -1640
rect 9460 -1780 9490 -1670
rect 9600 -1780 9630 -1670
rect 10360 -1750 10390 -1640
rect 10500 -1750 10530 -1640
rect 10360 -1780 10530 -1750
rect 11620 -1650 11790 -1620
rect 11620 -1760 11650 -1650
rect 11760 -1760 11790 -1650
rect 9460 -1810 9630 -1780
rect 11620 -1790 11790 -1760
rect 13030 -1640 13200 -1610
rect 13030 -1750 13060 -1640
rect 13170 -1750 13200 -1640
rect 13030 -1780 13200 -1750
rect 14190 -1650 14360 -1620
rect 14190 -1760 14220 -1650
rect 14330 -1760 14360 -1650
rect 14190 -1790 14360 -1760
rect 15260 -1640 15430 -1610
rect 15260 -1750 15290 -1640
rect 15400 -1750 15430 -1640
rect 15260 -1780 15430 -1750
rect 16370 -1630 16540 -1600
rect 16370 -1740 16400 -1630
rect 16510 -1740 16540 -1630
rect 16370 -1770 16540 -1740
rect 11350 -8110 11520 -8080
rect 11350 -8220 11380 -8110
rect 11490 -8220 11520 -8110
rect 11350 -8250 11520 -8220
rect 12990 -8120 13160 -8090
rect 12990 -8230 13020 -8120
rect 13130 -8230 13160 -8120
rect 12990 -8260 13160 -8230
rect 14400 -8110 14570 -8080
rect 14400 -8220 14430 -8110
rect 14540 -8220 14570 -8110
rect 14400 -8250 14570 -8220
rect 15780 -8110 15950 -8080
rect 15780 -8220 15810 -8110
rect 15920 -8220 15950 -8110
rect 15780 -8250 15950 -8220
rect 17320 -8120 17490 -8090
rect 17320 -8230 17350 -8120
rect 17460 -8230 17490 -8120
rect 17320 -8260 17490 -8230
rect 18600 -8120 18770 -8090
rect 18600 -8230 18630 -8120
rect 18740 -8230 18770 -8120
rect 18600 -8260 18770 -8230
<< nsubdiff >>
rect 8760 -690 8940 -660
rect 8760 -800 8790 -690
rect 8900 -800 8940 -690
rect 8760 -830 8940 -800
rect 9370 -690 9550 -660
rect 9370 -800 9410 -690
rect 9520 -800 9550 -690
rect 9370 -830 9550 -800
rect 9980 -700 10160 -670
rect 9980 -810 10010 -700
rect 10120 -810 10160 -700
rect 9980 -840 10160 -810
rect 10630 -710 10810 -680
rect 10630 -820 10660 -710
rect 10770 -820 10810 -710
rect 10630 -850 10810 -820
rect 11340 -700 11520 -670
rect 11340 -810 11380 -700
rect 11490 -810 11520 -700
rect 11340 -840 11520 -810
rect 12060 -700 12240 -670
rect 12060 -810 12090 -700
rect 12200 -810 12240 -700
rect 12060 -840 12240 -810
rect 13710 -720 13890 -690
rect 13710 -830 13750 -720
rect 13860 -830 13890 -720
rect 13710 -860 13890 -830
rect 15150 -730 15330 -700
rect 15150 -840 15190 -730
rect 15300 -840 15330 -730
rect 15150 -870 15330 -840
rect 8720 -2230 8890 -2200
rect 8720 -2340 8750 -2230
rect 8860 -2340 8890 -2230
rect 8720 -2370 8890 -2340
rect 11320 -7280 11490 -7250
rect 11320 -7390 11350 -7280
rect 11460 -7390 11490 -7280
rect 11320 -7420 11490 -7390
rect 13020 -7280 13190 -7250
rect 13020 -7390 13050 -7280
rect 13160 -7390 13190 -7280
rect 13020 -7420 13190 -7390
rect 14400 -7280 14570 -7250
rect 14400 -7390 14430 -7280
rect 14540 -7390 14570 -7280
rect 14400 -7420 14570 -7390
rect 15690 -7280 15860 -7250
rect 15690 -7390 15720 -7280
rect 15830 -7390 15860 -7280
rect 15690 -7420 15860 -7390
rect 17210 -7280 17380 -7250
rect 17210 -7390 17240 -7280
rect 17350 -7390 17380 -7280
rect 17210 -7420 17380 -7390
rect 18620 -7280 18790 -7250
rect 18620 -7390 18650 -7280
rect 18760 -7390 18790 -7280
rect 18620 -7420 18790 -7390
<< psubdiffcont >>
rect 9490 -1780 9600 -1670
rect 10390 -1750 10500 -1640
rect 11650 -1760 11760 -1650
rect 13060 -1750 13170 -1640
rect 14220 -1760 14330 -1650
rect 15290 -1750 15400 -1640
rect 16400 -1740 16510 -1630
rect 11380 -8220 11490 -8110
rect 13020 -8230 13130 -8120
rect 14430 -8220 14540 -8110
rect 15810 -8220 15920 -8110
rect 17350 -8230 17460 -8120
rect 18630 -8230 18740 -8120
<< nsubdiffcont >>
rect 8790 -800 8900 -690
rect 9410 -800 9520 -690
rect 10010 -810 10120 -700
rect 10660 -820 10770 -710
rect 11380 -810 11490 -700
rect 12090 -810 12200 -700
rect 13750 -830 13860 -720
rect 15190 -840 15300 -730
rect 8750 -2340 8860 -2230
rect 11350 -7390 11460 -7280
rect 13050 -7390 13160 -7280
rect 14430 -7390 14540 -7280
rect 15720 -7390 15830 -7280
rect 17240 -7390 17350 -7280
rect 18650 -7390 18760 -7280
<< locali >>
rect 10650 -1110 10690 -1100
rect 10640 -1150 10650 -1140
rect 10690 -1150 10700 -1140
rect 10640 -1190 10700 -1150
rect 8330 -1220 8620 -1200
rect 8330 -1380 8350 -1220
rect 8510 -1260 8620 -1220
rect 8780 -1260 8820 -1250
rect 9270 -1260 9320 -1250
rect 8510 -1270 8680 -1260
rect 8510 -1300 8730 -1270
rect 8510 -1380 8620 -1300
rect 8780 -1310 8980 -1260
rect 9270 -1310 9430 -1260
rect 8330 -1400 8620 -1380
rect 8330 -1670 8600 -1650
rect 8330 -1830 8350 -1670
rect 8510 -1820 8600 -1670
rect 8510 -1830 8780 -1820
rect 8330 -1860 8780 -1830
rect 11090 -7760 11190 -7740
rect 11090 -7800 11290 -7760
rect 11090 -7820 11190 -7800
rect 11340 -7810 11510 -7760
rect 11830 -7810 11970 -7760
<< viali >>
rect 8760 -690 8940 -660
rect 8760 -800 8790 -690
rect 8790 -800 8900 -690
rect 8900 -800 8940 -690
rect 8760 -830 8940 -800
rect 9370 -690 9550 -660
rect 9370 -800 9410 -690
rect 9410 -800 9520 -690
rect 9520 -800 9550 -690
rect 9370 -830 9550 -800
rect 9980 -700 10160 -670
rect 9980 -810 10010 -700
rect 10010 -810 10120 -700
rect 10120 -810 10160 -700
rect 9980 -840 10160 -810
rect 10630 -710 10810 -680
rect 10630 -820 10660 -710
rect 10660 -820 10770 -710
rect 10770 -820 10810 -710
rect 10630 -850 10810 -820
rect 11340 -700 11520 -670
rect 11340 -810 11380 -700
rect 11380 -810 11490 -700
rect 11490 -810 11520 -700
rect 11340 -840 11520 -810
rect 12060 -700 12240 -670
rect 12060 -810 12090 -700
rect 12090 -810 12200 -700
rect 12200 -810 12240 -700
rect 12060 -840 12240 -810
rect 13710 -720 13890 -690
rect 13710 -830 13750 -720
rect 13750 -830 13860 -720
rect 13860 -830 13890 -720
rect 13710 -860 13890 -830
rect 15150 -730 15330 -700
rect 15150 -840 15190 -730
rect 15190 -840 15300 -730
rect 15300 -840 15330 -730
rect 15150 -870 15330 -840
rect 10650 -1150 10690 -1110
rect 8350 -1380 8510 -1220
rect 10650 -1230 10690 -1190
rect 10650 -1310 10690 -1270
rect 11238 -1304 11643 -1264
rect 10650 -1400 10690 -1360
rect 12120 -1400 12160 -1130
rect 12740 -1307 13110 -1267
rect 13600 -1410 13640 -1140
rect 14199 -1304 14569 -1264
rect 15070 -1380 15110 -1110
rect 15339 -1305 15619 -1265
rect 16540 -1400 16580 -1130
rect 10360 -1640 10530 -1610
rect 8350 -1830 8510 -1670
rect 9460 -1670 9630 -1640
rect 9460 -1780 9490 -1670
rect 9490 -1780 9600 -1670
rect 9600 -1780 9630 -1670
rect 10360 -1750 10390 -1640
rect 10390 -1750 10500 -1640
rect 10500 -1750 10530 -1640
rect 10360 -1780 10530 -1750
rect 11620 -1650 11790 -1620
rect 11620 -1760 11650 -1650
rect 11650 -1760 11760 -1650
rect 11760 -1760 11790 -1650
rect 9460 -1810 9630 -1780
rect 11620 -1790 11790 -1760
rect 13030 -1640 13200 -1610
rect 13030 -1750 13060 -1640
rect 13060 -1750 13170 -1640
rect 13170 -1750 13200 -1640
rect 13030 -1780 13200 -1750
rect 14190 -1650 14360 -1620
rect 14190 -1760 14220 -1650
rect 14220 -1760 14330 -1650
rect 14330 -1760 14360 -1650
rect 14190 -1790 14360 -1760
rect 15260 -1640 15430 -1610
rect 15260 -1750 15290 -1640
rect 15290 -1750 15400 -1640
rect 15400 -1750 15430 -1640
rect 15260 -1780 15430 -1750
rect 16370 -1630 16540 -1600
rect 16370 -1740 16400 -1630
rect 16400 -1740 16510 -1630
rect 16510 -1740 16540 -1630
rect 16370 -1770 16540 -1740
rect 8810 -2030 8860 -1920
rect 8720 -2230 8890 -2200
rect 8720 -2340 8750 -2230
rect 8750 -2340 8860 -2230
rect 8860 -2340 8890 -2230
rect 8720 -2370 8890 -2340
rect 11320 -7280 11490 -7250
rect 11320 -7390 11350 -7280
rect 11350 -7390 11460 -7280
rect 11460 -7390 11490 -7280
rect 11320 -7420 11490 -7390
rect 13020 -7280 13190 -7250
rect 13020 -7390 13050 -7280
rect 13050 -7390 13160 -7280
rect 13160 -7390 13190 -7280
rect 13020 -7420 13190 -7390
rect 14400 -7280 14570 -7250
rect 14400 -7390 14430 -7280
rect 14430 -7390 14540 -7280
rect 14540 -7390 14570 -7280
rect 14400 -7420 14570 -7390
rect 15690 -7280 15860 -7250
rect 15690 -7390 15720 -7280
rect 15720 -7390 15830 -7280
rect 15830 -7390 15860 -7280
rect 15690 -7420 15860 -7390
rect 17210 -7280 17380 -7250
rect 17210 -7390 17240 -7280
rect 17240 -7390 17350 -7280
rect 17350 -7390 17380 -7280
rect 17210 -7420 17380 -7390
rect 18620 -7280 18790 -7250
rect 18620 -7390 18650 -7280
rect 18650 -7390 18760 -7280
rect 18760 -7390 18790 -7280
rect 18620 -7420 18790 -7390
rect 13200 -7860 13250 -7690
rect 13480 -7801 14341 -7767
rect 14680 -7860 14730 -7670
rect 14914 -7800 15775 -7766
rect 16150 -7860 16200 -7680
rect 16393 -7800 17254 -7766
rect 17620 -7870 17670 -7680
rect 17850 -7769 18617 -7767
rect 17848 -7803 18618 -7769
rect 19090 -7870 19140 -7680
rect 11350 -8110 11520 -8080
rect 11350 -8220 11380 -8110
rect 11380 -8220 11490 -8110
rect 11490 -8220 11520 -8110
rect 11350 -8250 11520 -8220
rect 12990 -8120 13160 -8090
rect 12990 -8230 13020 -8120
rect 13020 -8230 13130 -8120
rect 13130 -8230 13160 -8120
rect 12990 -8260 13160 -8230
rect 14400 -8110 14570 -8080
rect 14400 -8220 14430 -8110
rect 14430 -8220 14540 -8110
rect 14540 -8220 14570 -8110
rect 14400 -8250 14570 -8220
rect 15780 -8110 15950 -8080
rect 15780 -8220 15810 -8110
rect 15810 -8220 15920 -8110
rect 15920 -8220 15950 -8110
rect 15780 -8250 15950 -8220
rect 17320 -8120 17490 -8090
rect 17320 -8230 17350 -8120
rect 17350 -8230 17460 -8120
rect 17460 -8230 17490 -8120
rect 17320 -8260 17490 -8230
rect 18600 -8120 18770 -8090
rect 18600 -8230 18630 -8120
rect 18630 -8230 18740 -8120
rect 18740 -8230 18770 -8120
rect 18600 -8260 18770 -8230
<< metal1 >>
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 15750 -560 16020 -260
rect 480 -610 920 -600
rect 480 -790 690 -610
rect 910 -790 920 -610
rect 480 -800 920 -790
rect 8600 -660 16020 -560
rect 8600 -830 8760 -660
rect 8940 -830 9370 -660
rect 9550 -670 16020 -660
rect 9550 -830 9980 -670
rect 8600 -840 9980 -830
rect 10160 -680 11340 -670
rect 10160 -840 10630 -680
rect 8600 -850 10630 -840
rect 10810 -840 11340 -680
rect 11520 -840 12060 -670
rect 12240 -690 16020 -670
rect 16460 -690 16710 -260
rect 12240 -840 13710 -690
rect 10810 -850 13710 -840
rect 8600 -860 13710 -850
rect 13890 -700 16710 -690
rect 13890 -860 15150 -700
rect 8600 -870 15150 -860
rect 15330 -870 16710 -700
rect 480 -940 920 -930
rect 480 -1120 690 -940
rect 910 -1120 920 -940
rect 8600 -1030 16710 -870
rect 480 -1130 920 -1120
rect 10630 -1110 10780 -1100
rect 15040 -1110 15140 -1100
rect 10630 -1400 10650 -1110
rect 10690 -1140 10780 -1110
rect 10760 -1390 10780 -1140
rect 12090 -1120 12190 -1110
rect 11220 -1250 11660 -1240
rect 11220 -1264 11240 -1250
rect 11640 -1264 11660 -1250
rect 11220 -1304 11238 -1264
rect 11643 -1304 11660 -1264
rect 11220 -1320 11240 -1304
rect 11640 -1320 11660 -1304
rect 11220 -1330 11660 -1320
rect 10690 -1400 10780 -1390
rect 480 -1430 920 -1420
rect 10630 -1430 10780 -1400
rect 12090 -1410 12100 -1120
rect 12180 -1410 12190 -1120
rect 13570 -1130 13670 -1110
rect 12720 -1250 13130 -1240
rect 12720 -1320 12740 -1250
rect 13110 -1320 13130 -1250
rect 12720 -1330 13130 -1320
rect 12090 -1420 12190 -1410
rect 13570 -1420 13580 -1130
rect 13660 -1420 13670 -1130
rect 14180 -1250 14590 -1240
rect 14180 -1320 14190 -1250
rect 14580 -1320 14590 -1250
rect 14180 -1330 14590 -1320
rect 15040 -1380 15050 -1110
rect 15130 -1380 15140 -1110
rect 16510 -1120 16610 -1110
rect 15310 -1250 15640 -1240
rect 15310 -1320 15320 -1250
rect 15630 -1320 15640 -1250
rect 15310 -1330 15640 -1320
rect 15040 -1390 15140 -1380
rect 16510 -1410 16520 -1120
rect 16600 -1410 16610 -1120
rect 13570 -1430 13670 -1420
rect 480 -1610 690 -1430
rect 910 -1610 920 -1430
rect 17570 -1450 17980 -1420
rect 480 -1620 920 -1610
rect 8600 -1600 16710 -1470
rect 8600 -1610 16370 -1600
rect 8600 -1640 10360 -1610
rect 8600 -1650 9460 -1640
rect 480 -1710 920 -1700
rect 480 -1890 690 -1710
rect 910 -1890 920 -1710
rect 9350 -1810 9460 -1650
rect 9630 -1780 10360 -1640
rect 10530 -1620 13030 -1610
rect 10530 -1700 11620 -1620
rect 10530 -1780 11020 -1700
rect 9630 -1810 11020 -1780
rect 9350 -1850 11020 -1810
rect 480 -1900 920 -1890
rect 8380 -1920 8870 -1900
rect 8380 -1990 8810 -1920
rect 7640 -2000 8810 -1990
rect 480 -2170 920 -2160
rect 480 -2350 690 -2170
rect 910 -2350 920 -2170
rect 7640 -2240 7650 -2000
rect 7780 -2030 8810 -2000
rect 8860 -2030 8870 -1920
rect 7780 -2050 8870 -2030
rect 10870 -2050 11020 -1850
rect 11380 -1790 11620 -1700
rect 11790 -1780 13030 -1620
rect 13200 -1620 15260 -1610
rect 13200 -1780 14190 -1620
rect 11790 -1790 14190 -1780
rect 14360 -1780 15260 -1620
rect 15430 -1770 16370 -1610
rect 16540 -1770 16710 -1600
rect 15430 -1780 16710 -1770
rect 14360 -1790 16710 -1780
rect 11380 -1850 16710 -1790
rect 11380 -2050 11510 -1850
rect 7780 -2240 8560 -2050
rect 7640 -2250 8560 -2240
rect 8600 -2120 9470 -2090
rect 8600 -2200 9010 -2120
rect 480 -2360 920 -2350
rect 8600 -2370 8720 -2200
rect 8890 -2370 9010 -2200
rect 8600 -2380 9010 -2370
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16710 -1850
rect 17570 -1830 17600 -1450
rect 17950 -1530 17980 -1450
rect 17950 -1730 18180 -1530
rect 17950 -1830 17980 -1730
rect 17570 -1860 17980 -1830
rect 8600 -2410 9470 -2380
rect 480 -2530 920 -2520
rect 480 -2710 690 -2530
rect 910 -2710 920 -2530
rect 480 -2720 920 -2710
rect 15390 -2540 15660 -2110
rect 16100 -2140 16710 -2110
rect 16100 -2540 16350 -2140
rect 15390 -2760 16350 -2540
rect 480 -2930 920 -2920
rect 480 -3110 690 -2930
rect 910 -3110 920 -2930
rect 480 -3120 920 -3110
rect 480 -3380 920 -3370
rect 480 -3560 690 -3380
rect 910 -3560 920 -3380
rect 480 -3570 920 -3560
rect 480 -3750 920 -3740
rect 480 -3930 690 -3750
rect 910 -3930 920 -3750
rect 480 -3940 920 -3930
rect 11090 -5210 11290 -5010
rect 11670 -5150 11870 -4950
rect 12130 -5190 12330 -4990
rect 10660 -6610 19310 -6580
rect 10660 -7180 10690 -6610
rect 19280 -7180 19310 -6610
rect 10660 -7250 19310 -7180
rect 10660 -7420 11320 -7250
rect 11490 -7420 13020 -7250
rect 13190 -7420 14400 -7250
rect 14570 -7420 15690 -7250
rect 15860 -7420 17210 -7250
rect 17380 -7420 18620 -7250
rect 18790 -7420 19310 -7250
rect 10660 -7530 19310 -7420
rect 14660 -7660 14750 -7650
rect 13180 -7680 13270 -7670
rect 13180 -7870 13190 -7680
rect 13260 -7870 13270 -7680
rect 13450 -7740 14360 -7730
rect 13450 -7820 13460 -7740
rect 14350 -7820 14360 -7740
rect 13450 -7830 14360 -7820
rect 13180 -7880 13270 -7870
rect 14660 -7870 14670 -7660
rect 14740 -7870 14750 -7660
rect 16130 -7670 16220 -7660
rect 14900 -7740 15800 -7730
rect 14900 -7820 14910 -7740
rect 15790 -7820 15800 -7740
rect 14900 -7830 15800 -7820
rect 14660 -7880 14750 -7870
rect 16130 -7870 16140 -7670
rect 16210 -7870 16220 -7670
rect 17600 -7670 17690 -7660
rect 16370 -7750 17270 -7740
rect 16370 -7820 16380 -7750
rect 17260 -7820 17270 -7750
rect 16370 -7830 17270 -7820
rect 16130 -7880 16220 -7870
rect 17600 -7880 17610 -7670
rect 17680 -7880 17690 -7670
rect 19070 -7670 19160 -7660
rect 17840 -7749 18640 -7740
rect 17840 -7767 17852 -7749
rect 17840 -7769 17850 -7767
rect 17840 -7803 17848 -7769
rect 17840 -7821 17852 -7803
rect 18632 -7821 18640 -7749
rect 17840 -7830 18640 -7821
rect 17600 -7890 17690 -7880
rect 19070 -7880 19080 -7670
rect 19150 -7880 19160 -7670
rect 19070 -7890 19160 -7880
rect 10660 -8080 19310 -7970
rect 10660 -8250 11350 -8080
rect 11520 -8090 14400 -8080
rect 11520 -8250 12990 -8090
rect 10660 -8260 12990 -8250
rect 13160 -8250 14400 -8090
rect 14570 -8250 15780 -8080
rect 15950 -8090 19310 -8080
rect 15950 -8250 17320 -8090
rect 13160 -8260 17320 -8250
rect 17490 -8260 18600 -8090
rect 18770 -8260 19310 -8090
rect 10660 -8310 19310 -8260
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8950 920 -8770
rect 10660 -8880 10690 -8310
rect 19280 -8880 19310 -8310
rect 10660 -8910 19310 -8880
rect 680 -8960 920 -8950
rect 470 -9100 920 -9090
rect 470 -9280 690 -9100
rect 910 -9280 920 -9100
rect 470 -9290 920 -9280
rect 470 -9590 920 -9580
rect 470 -9770 690 -9590
rect 910 -9770 920 -9590
rect 470 -9780 920 -9770
rect 470 -9870 920 -9860
rect 470 -10050 690 -9870
rect 910 -10050 920 -9870
rect 470 -10060 920 -10050
rect 470 -10330 920 -10320
rect 470 -10510 690 -10330
rect 910 -10510 920 -10330
rect 470 -10520 920 -10510
rect 470 -10690 920 -10680
rect 470 -10870 690 -10690
rect 910 -10870 920 -10690
rect 470 -10880 920 -10870
rect 470 -11090 920 -11080
rect 470 -11270 690 -11090
rect 910 -11270 920 -11090
rect 470 -11280 920 -11270
rect 470 -11540 920 -11530
rect 470 -11720 690 -11540
rect 910 -11720 920 -11540
rect 470 -11730 920 -11720
rect 480 -11910 920 -11900
rect 480 -12090 690 -11910
rect 910 -12090 920 -11910
rect 480 -12100 920 -12090
<< via1 >>
rect 12830 -350 13270 80
rect 690 -790 910 -610
rect 16020 -690 16460 -260
rect 690 -1120 910 -940
rect 10650 -1150 10690 -1140
rect 10690 -1150 10760 -1140
rect 10650 -1190 10760 -1150
rect 10650 -1230 10690 -1190
rect 10690 -1230 10760 -1190
rect 10650 -1270 10760 -1230
rect 10650 -1310 10690 -1270
rect 10690 -1310 10760 -1270
rect 10650 -1360 10760 -1310
rect 10650 -1390 10690 -1360
rect 10690 -1390 10760 -1360
rect 11240 -1264 11640 -1250
rect 11240 -1304 11640 -1264
rect 11240 -1320 11640 -1304
rect 12100 -1130 12180 -1120
rect 12100 -1400 12120 -1130
rect 12120 -1400 12160 -1130
rect 12160 -1400 12180 -1130
rect 12100 -1410 12180 -1400
rect 12740 -1267 13110 -1250
rect 12740 -1307 13110 -1267
rect 12740 -1320 13110 -1307
rect 13580 -1140 13660 -1130
rect 13580 -1410 13600 -1140
rect 13600 -1410 13640 -1140
rect 13640 -1410 13660 -1140
rect 13580 -1420 13660 -1410
rect 14190 -1264 14580 -1250
rect 14190 -1304 14199 -1264
rect 14199 -1304 14569 -1264
rect 14569 -1304 14580 -1264
rect 14190 -1320 14580 -1304
rect 15050 -1380 15070 -1110
rect 15070 -1380 15110 -1110
rect 15110 -1380 15130 -1110
rect 15320 -1265 15630 -1250
rect 15320 -1305 15339 -1265
rect 15339 -1305 15619 -1265
rect 15619 -1305 15630 -1265
rect 15320 -1320 15630 -1305
rect 16520 -1130 16600 -1120
rect 16520 -1400 16540 -1130
rect 16540 -1400 16580 -1130
rect 16580 -1400 16600 -1130
rect 16520 -1410 16600 -1400
rect 690 -1610 910 -1430
rect 690 -1890 910 -1710
rect 690 -2350 910 -2170
rect 7650 -2240 7780 -2000
rect 11020 -2050 11380 -1700
rect 9010 -2380 9440 -2120
rect 17600 -1830 17950 -1450
rect 690 -2710 910 -2530
rect 15660 -2540 16100 -2110
rect 690 -3110 910 -2930
rect 690 -3560 910 -3380
rect 690 -3930 910 -3750
rect 10690 -7180 19280 -6610
rect 13190 -7690 13260 -7680
rect 13190 -7860 13200 -7690
rect 13200 -7860 13250 -7690
rect 13250 -7860 13260 -7690
rect 13190 -7870 13260 -7860
rect 13460 -7767 14350 -7740
rect 13460 -7801 13480 -7767
rect 13480 -7801 14341 -7767
rect 14341 -7801 14350 -7767
rect 13460 -7820 14350 -7801
rect 14670 -7670 14740 -7660
rect 14670 -7860 14680 -7670
rect 14680 -7860 14730 -7670
rect 14730 -7860 14740 -7670
rect 14670 -7870 14740 -7860
rect 14910 -7766 15790 -7740
rect 14910 -7800 14914 -7766
rect 14914 -7800 15775 -7766
rect 15775 -7800 15790 -7766
rect 14910 -7820 15790 -7800
rect 16140 -7680 16210 -7670
rect 16140 -7860 16150 -7680
rect 16150 -7860 16200 -7680
rect 16200 -7860 16210 -7680
rect 16140 -7870 16210 -7860
rect 16380 -7766 17260 -7750
rect 16380 -7800 16393 -7766
rect 16393 -7800 17254 -7766
rect 17254 -7800 17260 -7766
rect 16380 -7820 17260 -7800
rect 17610 -7680 17680 -7670
rect 17610 -7870 17620 -7680
rect 17620 -7870 17670 -7680
rect 17670 -7870 17680 -7680
rect 17610 -7880 17680 -7870
rect 17852 -7767 18632 -7749
rect 17852 -7769 18617 -7767
rect 18617 -7769 18632 -7767
rect 17852 -7803 18618 -7769
rect 18618 -7803 18632 -7769
rect 17852 -7821 18632 -7803
rect 19080 -7680 19150 -7670
rect 19080 -7870 19090 -7680
rect 19090 -7870 19140 -7680
rect 19140 -7870 19150 -7680
rect 19080 -7880 19150 -7870
rect 690 -8950 910 -8770
rect 10690 -8880 19280 -8310
rect 690 -9280 910 -9100
rect 690 -9770 910 -9590
rect 690 -10050 910 -9870
rect 690 -10510 910 -10330
rect 690 -10870 910 -10690
rect 690 -11270 910 -11090
rect 690 -11720 910 -11540
rect 690 -12090 910 -11910
<< metal2 >>
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 680 -610 920 -600
rect 680 -790 690 -610
rect 910 -790 920 -610
rect 15750 -690 16020 -260
rect 16460 -690 16710 -260
rect 680 -800 920 -790
rect 10630 -880 10780 -860
rect 680 -940 920 -930
rect 680 -1120 690 -940
rect 910 -1120 920 -940
rect 10630 -970 10650 -880
rect 10760 -970 10780 -880
rect 680 -1130 920 -1120
rect 10630 -1140 10780 -970
rect 680 -1430 920 -1420
rect 680 -1610 690 -1430
rect 910 -1610 920 -1430
rect 680 -1620 920 -1610
rect 680 -1710 920 -1700
rect 680 -1890 690 -1710
rect 910 -1890 920 -1710
rect 680 -1900 920 -1890
rect 680 -2170 920 -2160
rect 680 -2350 690 -2170
rect 910 -2350 920 -2170
rect 680 -2360 920 -2350
rect 680 -2530 920 -2520
rect 680 -2710 690 -2530
rect 910 -2710 920 -2530
rect 680 -2720 920 -2710
rect 680 -2930 920 -2920
rect 680 -3110 690 -2930
rect 910 -3110 920 -2930
rect 680 -3120 920 -3110
rect 680 -3380 920 -3370
rect 680 -3560 690 -3380
rect 910 -3560 920 -3380
rect 680 -3570 920 -3560
rect 680 -3750 920 -3740
rect 680 -3930 690 -3750
rect 910 -3930 920 -3750
rect 680 -3940 920 -3930
rect 1080 -3770 1220 -1150
rect 10630 -1390 10650 -1140
rect 10760 -1390 10780 -1140
rect 11220 -880 11630 -860
rect 11220 -950 11240 -880
rect 11610 -950 11630 -880
rect 11220 -1240 11630 -950
rect 12720 -870 13130 -860
rect 12720 -940 12740 -870
rect 13110 -940 13130 -870
rect 12090 -1120 12190 -1110
rect 11220 -1250 11660 -1240
rect 11220 -1320 11240 -1250
rect 11640 -1320 11660 -1250
rect 11220 -1330 11660 -1320
rect 10630 -1430 10780 -1390
rect 12090 -1410 12100 -1120
rect 12180 -1410 12190 -1120
rect 12720 -1250 13130 -940
rect 14180 -870 14590 -860
rect 14180 -940 14200 -870
rect 14570 -940 14590 -870
rect 12720 -1320 12740 -1250
rect 13110 -1320 13130 -1250
rect 12720 -1330 13130 -1320
rect 13570 -1130 13670 -1110
rect 12090 -1570 12190 -1410
rect 10870 -1700 11510 -1570
rect 12090 -1680 12100 -1570
rect 12180 -1680 12190 -1570
rect 12090 -1690 12190 -1680
rect 13570 -1420 13580 -1130
rect 13660 -1420 13670 -1130
rect 14180 -1250 14590 -940
rect 15310 -870 15640 -860
rect 15310 -940 15330 -870
rect 15620 -940 15640 -870
rect 15750 -920 16710 -690
rect 14180 -1320 14190 -1250
rect 14580 -1320 14590 -1250
rect 14180 -1330 14590 -1320
rect 15040 -1110 15140 -1100
rect 13570 -1570 13670 -1420
rect 13570 -1680 13580 -1570
rect 13660 -1680 13670 -1570
rect 13570 -1690 13670 -1680
rect 15040 -1380 15050 -1110
rect 15130 -1380 15140 -1110
rect 15310 -1250 15640 -940
rect 15310 -1320 15320 -1250
rect 15630 -1320 15640 -1250
rect 15310 -1330 15640 -1320
rect 16510 -1120 16610 -1110
rect 15040 -1570 15140 -1380
rect 15040 -1680 15050 -1570
rect 15130 -1680 15140 -1570
rect 15040 -1690 15140 -1680
rect 16510 -1410 16520 -1120
rect 16600 -1410 16610 -1120
rect 16510 -1570 16610 -1410
rect 16510 -1680 16520 -1570
rect 16600 -1680 16610 -1570
rect 16510 -1690 16610 -1680
rect 17570 -1450 17980 -1420
rect 7600 -2000 7790 -1990
rect 7600 -2240 7650 -2000
rect 7780 -2240 7790 -2000
rect 10870 -2050 11020 -1700
rect 11380 -2050 11510 -1700
rect 17570 -1830 17600 -1450
rect 17950 -1830 17980 -1450
rect 1080 -3910 1090 -3770
rect 1210 -3910 1220 -3770
rect 1080 -3940 1220 -3910
rect 7600 -8060 7790 -2240
rect 8980 -2120 9470 -2090
rect 8980 -2380 9010 -2120
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16350 -1850
rect 17570 -1860 17980 -1830
rect 8980 -2410 9470 -2380
rect 15390 -2540 15660 -2110
rect 16100 -2540 16350 -2110
rect 15390 -2760 16350 -2540
rect 10660 -6610 19310 -6580
rect 10660 -7180 10690 -6610
rect 19280 -7180 19310 -6610
rect 10660 -7210 19310 -7180
rect 13180 -7320 13270 -7310
rect 13180 -7410 13190 -7320
rect 13260 -7410 13270 -7320
rect 13180 -7680 13270 -7410
rect 13180 -7870 13190 -7680
rect 13260 -7870 13270 -7680
rect 13450 -7320 14360 -7310
rect 13450 -7410 13460 -7320
rect 14350 -7410 14360 -7320
rect 13450 -7740 14360 -7410
rect 14900 -7320 15800 -7310
rect 14900 -7410 14910 -7320
rect 15790 -7410 15800 -7320
rect 13450 -7820 13460 -7740
rect 14350 -7820 14360 -7740
rect 13450 -7830 14360 -7820
rect 14660 -7660 14750 -7650
rect 13180 -7880 13270 -7870
rect 14660 -7870 14670 -7660
rect 14740 -7870 14750 -7660
rect 14900 -7740 15800 -7410
rect 16370 -7320 17270 -7310
rect 16370 -7410 16380 -7320
rect 17260 -7410 17270 -7320
rect 14900 -7820 14910 -7740
rect 15790 -7820 15800 -7740
rect 14900 -7830 15800 -7820
rect 16130 -7670 16220 -7660
rect 7600 -8180 7610 -8060
rect 7780 -8180 7790 -8060
rect 7600 -8190 7790 -8180
rect 14660 -8100 14750 -7870
rect 14660 -8180 14670 -8100
rect 14740 -8180 14750 -8100
rect 14660 -8190 14750 -8180
rect 16130 -7870 16140 -7670
rect 16210 -7870 16220 -7670
rect 16370 -7750 17270 -7410
rect 17840 -7320 18640 -7310
rect 17840 -7410 17850 -7320
rect 18630 -7410 18640 -7320
rect 16370 -7820 16380 -7750
rect 17260 -7820 17270 -7750
rect 16370 -7830 17270 -7820
rect 17610 -7670 17690 -7660
rect 16130 -8100 16220 -7870
rect 16130 -8180 16140 -8100
rect 16210 -8180 16220 -8100
rect 16130 -8190 16220 -8180
rect 17680 -7880 17690 -7670
rect 17840 -7749 18640 -7410
rect 17840 -7821 17852 -7749
rect 18632 -7821 18640 -7749
rect 17840 -7831 18640 -7821
rect 19070 -7670 19160 -7660
rect 17610 -8100 17690 -7880
rect 17610 -8180 17620 -8100
rect 17680 -8180 17690 -8100
rect 17610 -8190 17690 -8180
rect 19070 -7880 19080 -7670
rect 19150 -7880 19160 -7670
rect 19070 -8100 19160 -7880
rect 19070 -8180 19080 -8100
rect 19150 -8180 19160 -8100
rect 19070 -8190 19160 -8180
rect 10660 -8310 19310 -8280
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8950 920 -8770
rect 10660 -8880 10690 -8310
rect 19280 -8880 19310 -8310
rect 10660 -8910 19310 -8880
rect 680 -8960 920 -8950
rect 680 -9100 920 -9090
rect 680 -9280 690 -9100
rect 910 -9280 920 -9100
rect 680 -9290 920 -9280
rect 680 -9590 920 -9580
rect 680 -9770 690 -9590
rect 910 -9770 920 -9590
rect 680 -9780 920 -9770
rect 680 -9870 920 -9860
rect 680 -10050 690 -9870
rect 910 -10050 920 -9870
rect 680 -10060 920 -10050
rect 680 -10330 920 -10320
rect 680 -10510 690 -10330
rect 910 -10510 920 -10330
rect 680 -10520 920 -10510
rect 680 -10690 920 -10680
rect 680 -10870 690 -10690
rect 910 -10870 920 -10690
rect 680 -10880 920 -10870
rect 680 -11090 920 -11080
rect 680 -11270 690 -11090
rect 910 -11270 920 -11090
rect 680 -11280 920 -11270
rect 680 -11540 920 -11530
rect 680 -11720 690 -11540
rect 910 -11720 920 -11540
rect 680 -11730 920 -11720
rect 680 -11910 920 -11900
rect 680 -12090 690 -11910
rect 910 -12090 920 -11910
rect 680 -12100 920 -12090
rect 1080 -11930 1220 -9310
rect 1080 -12070 1090 -11930
rect 1210 -12070 1220 -11930
rect 1080 -12100 1220 -12070
<< via2 >>
rect 12830 -350 13270 80
rect 690 -790 910 -610
rect 16020 -690 16460 -260
rect 3090 -890 3210 -790
rect 690 -1120 910 -940
rect 10650 -970 10760 -880
rect 2840 -1090 2960 -970
rect 690 -1610 910 -1430
rect 690 -1890 910 -1710
rect 690 -2350 910 -2170
rect 690 -2710 910 -2530
rect 690 -3110 910 -2930
rect 690 -3560 910 -3380
rect 690 -3930 910 -3750
rect 11240 -950 11610 -880
rect 12740 -940 13110 -870
rect 14200 -940 14570 -870
rect 2590 -1590 2710 -1450
rect 12100 -1680 12180 -1570
rect 15330 -940 15620 -870
rect 13580 -1680 13660 -1570
rect 15050 -1680 15130 -1570
rect 16520 -1680 16600 -1570
rect 2340 -1870 2460 -1730
rect 11020 -2050 11380 -1700
rect 17600 -1830 17950 -1450
rect 1840 -2690 1960 -2550
rect 1590 -3090 1710 -2960
rect 1340 -3540 1460 -3400
rect 1090 -3910 1210 -3770
rect 9010 -2380 9440 -2120
rect 15660 -2540 16100 -2110
rect 10690 -7180 19280 -6610
rect 13190 -7410 13260 -7320
rect 13460 -7410 14350 -7320
rect 14910 -7410 15790 -7320
rect 16380 -7410 17260 -7320
rect 7610 -8180 7780 -8060
rect 14670 -8180 14740 -8100
rect 17850 -7410 18630 -7320
rect 16140 -8180 16210 -8100
rect 17620 -8180 17680 -8100
rect 19080 -8180 19150 -8100
rect 690 -8950 910 -8770
rect 10690 -8880 19280 -8310
rect 3090 -9050 3210 -8950
rect 690 -9280 910 -9100
rect 2840 -9250 2960 -9130
rect 690 -9770 910 -9590
rect 690 -10050 910 -9870
rect 690 -10510 910 -10330
rect 690 -10870 910 -10690
rect 690 -11270 910 -11090
rect 690 -11720 910 -11540
rect 690 -12090 910 -11910
rect 2590 -9750 2710 -9610
rect 1840 -10850 1960 -10710
rect 1590 -11250 1710 -11110
rect 1340 -11700 1460 -11560
rect 1090 -12070 1210 -11930
<< metal3 >>
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 680 -610 920 -600
rect 680 -790 690 -610
rect 910 -620 920 -610
rect 910 -780 1240 -620
rect 15750 -690 16020 -260
rect 16460 -690 16710 -260
rect 910 -790 920 -780
rect 680 -800 920 -790
rect 1080 -790 3220 -780
rect 1080 -890 3090 -790
rect 3210 -890 3220 -790
rect 1080 -900 3220 -890
rect 10630 -870 15640 -860
rect 10630 -880 12740 -870
rect 680 -940 920 -930
rect 680 -1120 690 -940
rect 910 -960 920 -940
rect 910 -970 2970 -960
rect 910 -1090 2840 -970
rect 2960 -1090 2970 -970
rect 10630 -970 10650 -880
rect 10760 -950 11240 -880
rect 11610 -940 12740 -880
rect 13110 -940 14200 -870
rect 14570 -940 15330 -870
rect 15620 -940 15640 -870
rect 15750 -920 16710 -690
rect 11610 -950 15640 -940
rect 10760 -960 15640 -950
rect 10760 -970 10780 -960
rect 10630 -990 10780 -970
rect 910 -1100 2970 -1090
rect 910 -1120 920 -1100
rect 680 -1130 920 -1120
rect 680 -1430 920 -1420
rect 680 -1610 690 -1430
rect 910 -1440 920 -1430
rect 910 -1450 2720 -1440
rect 910 -1590 2590 -1450
rect 2710 -1590 2720 -1450
rect 17570 -1450 17980 -1420
rect 17570 -1560 17600 -1450
rect 12090 -1570 17600 -1560
rect 910 -1600 2720 -1590
rect 910 -1610 920 -1600
rect 680 -1620 920 -1610
rect 10870 -1700 11510 -1570
rect 12090 -1680 12100 -1570
rect 12180 -1680 13580 -1570
rect 13660 -1680 15050 -1570
rect 15130 -1680 16520 -1570
rect 16600 -1680 17600 -1570
rect 12090 -1690 17600 -1680
rect 680 -1710 920 -1700
rect 680 -1890 690 -1710
rect 910 -1720 920 -1710
rect 910 -1730 2470 -1720
rect 910 -1870 2340 -1730
rect 2460 -1870 2470 -1730
rect 910 -1880 2470 -1870
rect 910 -1890 920 -1880
rect 680 -1900 920 -1890
rect 10870 -2050 11020 -1700
rect 11380 -2050 11510 -1700
rect 17570 -1830 17600 -1690
rect 17950 -1830 17980 -1450
rect 8980 -2120 9470 -2090
rect 680 -2170 920 -2160
rect 680 -2350 690 -2170
rect 910 -2180 920 -2170
rect 910 -2340 2220 -2180
rect 910 -2350 920 -2340
rect 680 -2360 920 -2350
rect 8980 -2380 9010 -2120
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16350 -1850
rect 17570 -1860 17980 -1830
rect 8980 -2410 9470 -2380
rect 680 -2530 920 -2520
rect 680 -2710 690 -2530
rect 910 -2540 920 -2530
rect 15390 -2540 15660 -2110
rect 16100 -2540 16350 -2110
rect 910 -2550 1970 -2540
rect 910 -2690 1840 -2550
rect 1960 -2690 1970 -2550
rect 910 -2700 1970 -2690
rect 910 -2710 920 -2700
rect 680 -2720 920 -2710
rect 15390 -2760 16350 -2540
rect 680 -2930 920 -2920
rect 680 -3110 690 -2930
rect 910 -2950 920 -2930
rect 910 -2960 1720 -2950
rect 910 -3090 1590 -2960
rect 1710 -3090 1720 -2960
rect 910 -3100 1720 -3090
rect 910 -3110 920 -3100
rect 680 -3120 920 -3110
rect 680 -3380 920 -3370
rect 680 -3560 690 -3380
rect 910 -3390 920 -3380
rect 910 -3400 1470 -3390
rect 910 -3540 1340 -3400
rect 1460 -3540 1470 -3400
rect 910 -3550 1470 -3540
rect 910 -3560 920 -3550
rect 680 -3570 920 -3560
rect 680 -3750 920 -3740
rect 680 -3930 690 -3750
rect 910 -3760 920 -3750
rect 910 -3770 1220 -3760
rect 910 -3910 1090 -3770
rect 1210 -3910 1220 -3770
rect 910 -3920 1220 -3910
rect 910 -3930 920 -3920
rect 680 -3940 920 -3930
rect 10660 -6610 19310 -6580
rect 10660 -7180 10690 -6610
rect 19280 -7180 19310 -6610
rect 10660 -7210 19310 -7180
rect 13180 -7320 18640 -7310
rect 13180 -7410 13190 -7320
rect 13260 -7410 13460 -7320
rect 14350 -7410 14910 -7320
rect 15790 -7410 16380 -7320
rect 17260 -7410 17850 -7320
rect 18630 -7410 18640 -7320
rect 13180 -7420 18640 -7410
rect 6630 -8060 7790 -8050
rect 6630 -8180 7610 -8060
rect 7780 -8180 7790 -8060
rect 6630 -8190 7790 -8180
rect 14660 -8100 19620 -8090
rect 14660 -8180 14670 -8100
rect 14740 -8180 16140 -8100
rect 16210 -8180 17620 -8100
rect 17680 -8180 19080 -8100
rect 19150 -8180 19620 -8100
rect 14660 -8190 19620 -8180
rect 10660 -8310 19310 -8280
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8780 920 -8770
rect 910 -8940 1240 -8780
rect 10660 -8880 10690 -8310
rect 19280 -8880 19310 -8310
rect 10660 -8910 19310 -8880
rect 910 -8950 920 -8940
rect 680 -8960 920 -8950
rect 1080 -8950 3220 -8940
rect 1080 -9050 3090 -8950
rect 3210 -9050 3220 -8950
rect 1080 -9060 3220 -9050
rect 680 -9100 920 -9090
rect 680 -9280 690 -9100
rect 910 -9120 920 -9100
rect 910 -9130 2970 -9120
rect 910 -9250 2840 -9130
rect 2960 -9250 2970 -9130
rect 910 -9260 2970 -9250
rect 910 -9280 920 -9260
rect 680 -9290 920 -9280
rect 680 -9590 920 -9580
rect 680 -9770 690 -9590
rect 910 -9600 920 -9590
rect 910 -9610 2720 -9600
rect 910 -9750 2590 -9610
rect 2710 -9750 2720 -9610
rect 910 -9760 2720 -9750
rect 910 -9770 920 -9760
rect 680 -9780 920 -9770
rect 680 -9870 920 -9860
rect 680 -10050 690 -9870
rect 910 -9880 920 -9870
rect 910 -10040 2470 -9880
rect 910 -10050 920 -10040
rect 680 -10060 920 -10050
rect 2250 -10100 2470 -10040
rect 680 -10330 920 -10320
rect 680 -10510 690 -10330
rect 910 -10340 920 -10330
rect 910 -10500 2220 -10340
rect 910 -10510 920 -10500
rect 680 -10520 920 -10510
rect 680 -10690 920 -10680
rect 680 -10870 690 -10690
rect 910 -10700 920 -10690
rect 910 -10710 1970 -10700
rect 910 -10850 1840 -10710
rect 1960 -10850 1970 -10710
rect 910 -10860 1970 -10850
rect 910 -10870 920 -10860
rect 680 -10880 920 -10870
rect 680 -11090 920 -11080
rect 680 -11270 690 -11090
rect 910 -11100 920 -11090
rect 910 -11110 1720 -11100
rect 910 -11250 1590 -11110
rect 1710 -11250 1720 -11110
rect 910 -11260 1720 -11250
rect 910 -11270 920 -11260
rect 680 -11280 920 -11270
rect 680 -11540 920 -11530
rect 680 -11720 690 -11540
rect 910 -11550 920 -11540
rect 910 -11560 1470 -11550
rect 910 -11700 1340 -11560
rect 1460 -11700 1470 -11560
rect 910 -11710 1470 -11700
rect 910 -11720 920 -11710
rect 680 -11730 920 -11720
rect 680 -11910 920 -11900
rect 680 -12090 690 -11910
rect 910 -11920 920 -11910
rect 910 -11930 1220 -11920
rect 910 -12070 1090 -11930
rect 1210 -12070 1220 -11930
rect 910 -12080 1220 -12070
rect 910 -12090 920 -12080
rect 680 -12100 920 -12090
<< via3 >>
rect 12830 -350 13270 80
rect 16020 -690 16460 -260
rect 11020 -2050 11380 -1700
rect 9010 -2380 9440 -2120
rect 15660 -2540 16100 -2110
rect 10690 -7180 19280 -6610
rect 10690 -8880 19280 -8310
<< metal4 >>
rect 4140 -500 8590 300
rect 4140 -15670 4950 -500
rect 7640 -1470 8590 -500
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 15750 -690 16020 -260
rect 16460 -690 16710 -260
rect 15750 -920 16710 -690
rect 7640 -1700 17310 -1470
rect 7640 -1850 11020 -1700
rect 7640 -15750 8590 -1850
rect 10870 -2050 11020 -1850
rect 11380 -1850 17310 -1700
rect 11380 -2050 11510 -1850
rect 8980 -2120 9470 -2090
rect 8980 -2380 9010 -2120
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16960 -1850
rect 8980 -2410 9470 -2380
rect 15390 -2540 15660 -2110
rect 16100 -2200 16960 -2110
rect 16100 -2540 16350 -2200
rect 15390 -2760 16350 -2540
rect 10660 -6610 19310 -6580
rect 10660 -7180 10690 -6610
rect 19280 -7180 19310 -6610
rect 10660 -7210 19310 -7180
rect 10660 -8310 19310 -8280
rect 10660 -8880 10690 -8310
rect 19280 -8880 19310 -8310
rect 10660 -8910 19310 -8880
<< via4 >>
rect 12830 -350 13270 80
rect 16020 -690 16460 -260
rect 9010 -2380 9440 -2120
rect 15660 -2540 16100 -2110
rect 10690 -7180 19280 -6610
<< metal5 >>
rect 12570 80 13530 350
rect 12570 10 12830 80
rect 7160 -350 12830 10
rect 13270 10 13530 80
rect 13270 -260 17310 10
rect 13270 -350 16020 -260
rect 7160 -690 16020 -350
rect 16460 -690 17310 -260
rect 7160 -1130 17310 -690
rect 7160 -1760 8400 -1130
rect 7160 -2110 17310 -1760
rect 7160 -2120 15660 -2110
rect 7160 -2380 9010 -2120
rect 9440 -2200 15660 -2120
rect 9440 -2380 9470 -2200
rect 7160 -2410 9470 -2380
rect 7160 -15300 8400 -2410
rect 15390 -2540 15660 -2200
rect 16100 -2200 17310 -2110
rect 16100 -2540 16350 -2200
rect 15390 -2760 16350 -2540
rect 10660 -6610 19310 -6580
rect 10660 -7180 10690 -6610
rect 19280 -7180 19310 -6610
rect 10660 -7210 19310 -7180
use sky130_fd_sc_hd__or2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713414733
transform 1 0 10708 0 1 -10162
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  x2
timestamp 1713414733
transform 1 0 10708 0 1 -11812
box -38 -48 498 592
use 8to3_Priority_Encoder_v0p2p0  x3
timestamp 1713414733
transform 1 0 4960 0 1 -8740
box -3910 -7130 3570 700
use sky130_fd_sc_hd__inv_16  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713414733
transform 1 0 12288 0 1 -1522
box -38 -48 1510 592
use 8to3_Priority_Encoder_v0p2p0  x5
timestamp 1713414733
transform 1 0 4960 0 1 -700
box -3910 -7130 3570 700
use sky130_fd_sc_hd__inv_16  x6
timestamp 1713414733
transform 1 0 10816 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713414733
transform 1 0 8658 0 -1 -1598
box -38 -48 314 592
use sky130_fd_sc_hd__inv_16  x8
timestamp 1713414733
transform 1 0 13760 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x9
timestamp 1713414733
transform 1 0 15232 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x10
timestamp 1713414733
transform 1 0 13376 0 1 -8022
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  x11
timestamp 1713414733
transform 1 0 10708 0 1 -8022
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x12
timestamp 1713414733
transform 1 0 14848 0 1 -8022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x13
timestamp 1713414733
transform 1 0 16320 0 1 -8022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x14
timestamp 1713414733
transform 1 0 17792 0 1 -8022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x15
timestamp 1713414733
transform 1 0 13376 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x16
timestamp 1713414733
transform 1 0 14848 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x17
timestamp 1713414733
transform 1 0 16320 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x18
timestamp 1713414733
transform 1 0 17792 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x19
timestamp 1713414733
transform 1 0 13376 0 1 -11812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x20
timestamp 1713414733
transform 1 0 11168 0 1 -11812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1713414733
transform 1 0 11444 0 1 -11812
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x22
timestamp 1713414733
transform 1 0 11904 0 1 -11812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x23
timestamp 1713414733
transform 1 0 14848 0 1 -11812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x24
timestamp 1713414733
transform 1 0 16320 0 1 -11812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x25
timestamp 1713414733
transform 1 0 17792 0 1 -11812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x27
timestamp 1713414733
transform 1 0 11168 0 1 -10162
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x28
timestamp 1713414733
transform 1 0 11444 0 1 -10162
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x29
timestamp 1713414733
transform 1 0 11904 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x34
timestamp 1713414733
transform 1 0 11168 0 1 -8022
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x35
timestamp 1713414733
transform 1 0 11444 0 1 -8022
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x36
timestamp 1713414733
transform 1 0 11904 0 1 -8022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x41
timestamp 1713414733
transform 1 0 8608 0 1 -1522
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x42
timestamp 1713414733
transform 1 0 8884 0 1 -1522
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x43
timestamp 1713414733
transform 1 0 9344 0 1 -1522
box -38 -48 1510 592
<< labels >>
flabel metal1 480 -1130 680 -930 0 FreeSans 256 0 0 0 I15
port 2 nsew
flabel metal1 480 -800 680 -600 0 FreeSans 256 0 0 0 EI
port 1 nsew
flabel metal1 480 -1620 680 -1420 0 FreeSans 256 0 0 0 I14
port 3 nsew
flabel metal1 480 -1900 680 -1700 0 FreeSans 256 0 0 0 I13
port 4 nsew
flabel metal1 480 -2360 680 -2160 0 FreeSans 256 0 0 0 I12
port 5 nsew
flabel metal1 480 -2720 680 -2520 0 FreeSans 256 0 0 0 I11
port 6 nsew
flabel metal1 480 -3120 680 -2920 0 FreeSans 256 0 0 0 I10
port 7 nsew
flabel metal1 480 -3570 680 -3370 0 FreeSans 256 0 0 0 I9
port 9 nsew
flabel metal1 480 -3940 680 -3740 0 FreeSans 256 0 0 0 I8
port 10 nsew
flabel metal1 480 -12100 680 -11900 0 FreeSans 256 0 0 0 I0
port 19 nsew
flabel metal1 470 -11730 670 -11530 0 FreeSans 256 0 0 0 I1
port 18 nsew
flabel metal1 470 -11280 670 -11080 0 FreeSans 256 0 0 0 I2
port 17 nsew
flabel metal1 470 -10880 670 -10680 0 FreeSans 256 0 0 0 I3
port 16 nsew
flabel metal1 470 -10520 670 -10320 0 FreeSans 256 0 0 0 I4
port 14 nsew
flabel metal1 470 -10060 670 -9860 0 FreeSans 256 0 0 0 I5
port 13 nsew
flabel metal1 470 -9780 670 -9580 0 FreeSans 256 0 0 0 I6
port 12 nsew
flabel metal1 470 -9290 670 -9090 0 FreeSans 256 0 0 0 I7
port 11 nsew
flabel metal1 17980 -1730 18180 -1530 0 FreeSans 256 0 0 0 A3
port 0 nsew
flabel metal1 11090 -5210 11290 -5010 0 FreeSans 256 0 0 0 A2
port 8 nsew
flabel metal1 11670 -5150 11870 -4950 0 FreeSans 256 0 0 0 A1
port 15 nsew
flabel metal1 12130 -5190 12330 -4990 0 FreeSans 256 0 0 0 A0
port 20 nsew
<< end >>
