magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< pwell >>
rect -5086 -1136 5086 1136
<< psubdiff >>
rect -5050 1066 -4954 1100
rect 4954 1066 5050 1100
rect -5050 1004 -5016 1066
rect 5016 1004 5050 1066
rect -5050 -1066 -5016 -1004
rect 5016 -1066 5050 -1004
rect -5050 -1100 -4954 -1066
rect 4954 -1100 5050 -1066
<< psubdiffcont >>
rect -4954 1066 4954 1100
rect -5050 -1004 -5016 1004
rect 5016 -1004 5050 1004
rect -4954 -1100 4954 -1066
<< xpolycontact >>
rect -4920 538 -3774 970
rect -4920 -970 -3774 -538
rect -3678 538 -2532 970
rect -3678 -970 -2532 -538
rect -2436 538 -1290 970
rect -2436 -970 -1290 -538
rect -1194 538 -48 970
rect -1194 -970 -48 -538
rect 48 538 1194 970
rect 48 -970 1194 -538
rect 1290 538 2436 970
rect 1290 -970 2436 -538
rect 2532 538 3678 970
rect 2532 -970 3678 -538
rect 3774 538 4920 970
rect 3774 -970 4920 -538
<< xpolyres >>
rect -4920 -538 -3774 538
rect -3678 -538 -2532 538
rect -2436 -538 -1290 538
rect -1194 -538 -48 538
rect 48 -538 1194 538
rect 1290 -538 2436 538
rect 2532 -538 3678 538
rect 3774 -538 4920 538
<< locali >>
rect -5050 1066 -4954 1100
rect 4954 1066 5050 1100
rect -5050 1004 -5016 1066
rect 5016 1004 5050 1066
rect -5050 -1066 -5016 -1004
rect 5016 -1066 5050 -1004
rect -5050 -1100 -4954 -1066
rect 4954 -1100 5050 -1066
<< viali >>
rect -4904 555 -3790 952
rect -3662 555 -2548 952
rect -2420 555 -1306 952
rect -1178 555 -64 952
rect 64 555 1178 952
rect 1306 555 2420 952
rect 2548 555 3662 952
rect 3790 555 4904 952
rect -4904 -952 -3790 -555
rect -3662 -952 -2548 -555
rect -2420 -952 -1306 -555
rect -1178 -952 -64 -555
rect 64 -952 1178 -555
rect 1306 -952 2420 -555
rect 2548 -952 3662 -555
rect 3790 -952 4904 -555
<< metal1 >>
rect -4916 952 -3778 958
rect -4916 555 -4904 952
rect -3790 555 -3778 952
rect -4916 549 -3778 555
rect -3674 952 -2536 958
rect -3674 555 -3662 952
rect -2548 555 -2536 952
rect -3674 549 -2536 555
rect -2432 952 -1294 958
rect -2432 555 -2420 952
rect -1306 555 -1294 952
rect -2432 549 -1294 555
rect -1190 952 -52 958
rect -1190 555 -1178 952
rect -64 555 -52 952
rect -1190 549 -52 555
rect 52 952 1190 958
rect 52 555 64 952
rect 1178 555 1190 952
rect 52 549 1190 555
rect 1294 952 2432 958
rect 1294 555 1306 952
rect 2420 555 2432 952
rect 1294 549 2432 555
rect 2536 952 3674 958
rect 2536 555 2548 952
rect 3662 555 3674 952
rect 2536 549 3674 555
rect 3778 952 4916 958
rect 3778 555 3790 952
rect 4904 555 4916 952
rect 3778 549 4916 555
rect -4916 -555 -3778 -549
rect -4916 -952 -4904 -555
rect -3790 -952 -3778 -555
rect -4916 -958 -3778 -952
rect -3674 -555 -2536 -549
rect -3674 -952 -3662 -555
rect -2548 -952 -2536 -555
rect -3674 -958 -2536 -952
rect -2432 -555 -1294 -549
rect -2432 -952 -2420 -555
rect -1306 -952 -1294 -555
rect -2432 -958 -1294 -952
rect -1190 -555 -52 -549
rect -1190 -952 -1178 -555
rect -64 -952 -52 -555
rect -1190 -958 -52 -952
rect 52 -555 1190 -549
rect 52 -952 64 -555
rect 1178 -952 1190 -555
rect 52 -958 1190 -952
rect 1294 -555 2432 -549
rect 1294 -952 1306 -555
rect 2420 -952 2432 -555
rect 1294 -958 2432 -952
rect 2536 -555 3674 -549
rect 2536 -952 2548 -555
rect 3662 -952 3674 -555
rect 2536 -958 3674 -952
rect 3778 -555 4916 -549
rect 3778 -952 3790 -555
rect 4904 -952 4916 -555
rect 3778 -958 4916 -952
<< properties >>
string FIXED_BBOX -5033 -1083 5033 1083
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 5.542 m 1 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 2.0k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
