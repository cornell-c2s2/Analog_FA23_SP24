magic
tech sky130A
magscale 1 2
timestamp 1716326491
<< nwell >>
rect 53860 -2340 55098 -1522
rect 57056 -2024 57406 -1830
rect 57056 -2320 57410 -2024
rect 57058 -2345 57410 -2320
rect 55000 -2638 55630 -2626
rect 55000 -2928 55640 -2638
rect 55000 -3538 55640 -3248
rect 55000 -3550 55630 -3538
rect 56280 -3706 56742 -2468
rect 58894 -2447 59732 -1897
rect 53850 -4656 55088 -3838
rect 58894 -3804 59346 -2447
rect 60405 -3426 61056 -2890
rect 60406 -3570 61056 -3426
rect 57056 -4460 57416 -3840
rect 58894 -4354 59732 -3804
rect 20696 -11875 22260 -7637
rect 53860 -7740 55098 -6922
rect 57056 -7424 57406 -7230
rect 57056 -7720 57410 -7424
rect 57058 -7745 57410 -7720
rect 55000 -8038 55630 -8026
rect 55000 -8328 55640 -8038
rect 55000 -8938 55640 -8648
rect 55000 -8950 55630 -8938
rect 56280 -9106 56742 -7868
rect 58894 -7847 59732 -7297
rect 53850 -10056 55088 -9238
rect 58894 -9204 59346 -7847
rect 60405 -8826 61056 -8290
rect 60406 -8970 61056 -8826
rect 57056 -9860 57416 -9240
rect 58894 -9754 59732 -9204
rect 53860 -13140 55098 -12322
rect 57056 -12824 57406 -12630
rect 57056 -13120 57410 -12824
rect 57058 -13145 57410 -13120
rect 55000 -13438 55630 -13426
rect 55000 -13728 55640 -13438
rect 55000 -14338 55640 -14048
rect 55000 -14350 55630 -14338
rect 56280 -14506 56742 -13268
rect 58894 -13247 59732 -12697
rect 53850 -15456 55088 -14638
rect 58894 -14604 59346 -13247
rect 60405 -14226 61056 -13690
rect 60406 -14370 61056 -14226
rect 57056 -15260 57416 -14640
rect 58894 -15154 59732 -14604
rect 53860 -18540 55098 -17722
rect 57056 -18224 57406 -18030
rect 57056 -18520 57410 -18224
rect 57058 -18545 57410 -18520
rect 55000 -18838 55630 -18826
rect 55000 -19128 55640 -18838
rect 55000 -19738 55640 -19448
rect 55000 -19750 55630 -19738
rect 56280 -19906 56742 -18668
rect 58894 -18647 59732 -18097
rect 53850 -20856 55088 -20038
rect 58894 -20004 59346 -18647
rect 60405 -19626 61056 -19090
rect 60406 -19770 61056 -19626
rect 57056 -20660 57416 -20040
rect 58894 -20554 59732 -20004
rect 53860 -23940 55098 -23122
rect 57056 -23624 57406 -23430
rect 57056 -23920 57410 -23624
rect 57058 -23945 57410 -23920
rect 55000 -24238 55630 -24226
rect 55000 -24528 55640 -24238
rect 55000 -25138 55640 -24848
rect 55000 -25150 55630 -25138
rect 56280 -25306 56742 -24068
rect 58894 -24047 59732 -23497
rect 53850 -26256 55088 -25438
rect 58894 -25404 59346 -24047
rect 60405 -25026 61056 -24490
rect 60406 -25170 61056 -25026
rect 57056 -26060 57416 -25440
rect 58894 -25954 59732 -25404
rect 53860 -29340 55098 -28522
rect 57056 -29024 57406 -28830
rect 57056 -29320 57410 -29024
rect 57058 -29345 57410 -29320
rect 55000 -29638 55630 -29626
rect 55000 -29928 55640 -29638
rect 55000 -30538 55640 -30248
rect 55000 -30550 55630 -30538
rect 56280 -30706 56742 -29468
rect 58894 -29447 59732 -28897
rect 53850 -31656 55088 -30838
rect 58894 -30804 59346 -29447
rect 60405 -30426 61056 -29890
rect 60406 -30570 61056 -30426
rect 57056 -31460 57416 -30840
rect 58894 -31354 59732 -30804
rect 53860 -34740 55098 -33922
rect 57056 -34424 57406 -34230
rect 57056 -34720 57410 -34424
rect 57058 -34745 57410 -34720
rect 55000 -35038 55630 -35026
rect 55000 -35328 55640 -35038
rect 55000 -35938 55640 -35648
rect 55000 -35950 55630 -35938
rect 56280 -36106 56742 -34868
rect 58894 -34847 59732 -34297
rect 53850 -37056 55088 -36238
rect 58894 -36204 59346 -34847
rect 60405 -35826 61056 -35290
rect 60406 -35970 61056 -35826
rect 57056 -36860 57416 -36240
rect 58894 -36754 59732 -36204
rect 75468 -38650 76922 -38649
rect 75460 -39080 79280 -38650
rect 84700 -38670 85660 -37780
rect 53860 -40140 55098 -39322
rect 77540 -39340 79280 -39080
rect 77540 -39341 79088 -39340
rect 80690 -39400 88880 -38670
rect 57056 -39824 57406 -39630
rect 57056 -40120 57410 -39824
rect 57058 -40145 57410 -40120
rect 55000 -40438 55630 -40426
rect 55000 -40728 55640 -40438
rect 55000 -41338 55640 -41048
rect 55000 -41350 55630 -41338
rect 56280 -41506 56742 -40268
rect 58894 -40247 59732 -39697
rect 77540 -39950 78168 -39949
rect 53850 -42456 55088 -41638
rect 58894 -41604 59346 -40247
rect 60405 -41226 61056 -40690
rect 77540 -40600 79280 -39950
rect 80740 -40540 81110 -39980
rect 77540 -41190 78628 -41189
rect 60406 -41370 61056 -41226
rect 57056 -42260 57416 -41640
rect 58894 -42154 59732 -41604
rect 77530 -41840 79280 -41190
rect 77540 -43080 79280 -42440
rect 77540 -43081 78912 -43080
rect 77530 -44320 79280 -43670
rect 82790 -43900 91440 -43340
rect 53860 -45540 55098 -44722
rect 57056 -45224 57406 -45030
rect 57056 -45520 57410 -45224
rect 57058 -45545 57410 -45520
rect 55000 -45838 55630 -45826
rect 55000 -46128 55640 -45838
rect 55000 -46738 55640 -46448
rect 55000 -46750 55630 -46738
rect 56280 -46906 56742 -45668
rect 58894 -45647 59732 -45097
rect 53850 -47856 55088 -47038
rect 58894 -47004 59346 -45647
rect 77530 -45560 79280 -44900
rect 60405 -46626 61056 -46090
rect 60406 -46770 61056 -46626
rect 75468 -46690 76922 -46689
rect 57056 -47660 57416 -47040
rect 58894 -47554 59732 -47004
rect 75460 -47120 79280 -46690
rect 77540 -47380 79280 -47120
rect 77540 -47381 79088 -47380
rect 77540 -47990 78168 -47989
rect 77540 -48640 79280 -47990
rect 82794 -48038 91444 -47478
rect 77540 -49230 78628 -49229
rect 77530 -49880 79280 -49230
rect 53860 -50940 55098 -50122
rect 57056 -50624 57406 -50430
rect 57056 -50920 57410 -50624
rect 57058 -50945 57410 -50920
rect 55000 -51238 55630 -51226
rect 55000 -51528 55640 -51238
rect 55000 -52138 55640 -51848
rect 55000 -52150 55630 -52138
rect 56280 -52306 56742 -51068
rect 58894 -51047 59732 -50497
rect 53850 -53256 55088 -52438
rect 58894 -52404 59346 -51047
rect 77540 -51120 79280 -50480
rect 77540 -51121 78912 -51120
rect 60405 -52026 61056 -51490
rect 82790 -51690 91440 -51130
rect 60406 -52170 61056 -52026
rect 57056 -53060 57416 -52440
rect 58894 -52954 59732 -52404
rect 77530 -52360 79280 -51710
rect 77530 -53600 79280 -52940
rect 53860 -56340 55098 -55522
rect 57056 -56024 57406 -55830
rect 57056 -56320 57410 -56024
rect 57058 -56345 57410 -56320
rect 55000 -56638 55630 -56626
rect 55000 -56928 55640 -56638
rect 55000 -57538 55640 -57248
rect 55000 -57550 55630 -57538
rect 56280 -57706 56742 -56468
rect 58894 -56447 59732 -55897
rect 53850 -58656 55088 -57838
rect 58894 -57804 59346 -56447
rect 60405 -57426 61056 -56890
rect 60406 -57570 61056 -57426
rect 57056 -58460 57416 -57840
rect 58894 -58354 59732 -57804
rect 53860 -61740 55098 -60922
rect 57056 -61424 57406 -61230
rect 57056 -61720 57410 -61424
rect 57058 -61745 57410 -61720
rect 55000 -62038 55630 -62026
rect 55000 -62328 55640 -62038
rect 55000 -62938 55640 -62648
rect 55000 -62950 55630 -62938
rect 56280 -63106 56742 -61868
rect 58894 -61847 59732 -61297
rect 53850 -64056 55088 -63238
rect 58894 -63204 59346 -61847
rect 60405 -62826 61056 -62290
rect 60406 -62970 61056 -62826
rect 57056 -63860 57416 -63240
rect 58894 -63754 59732 -63204
rect 53860 -67140 55098 -66322
rect 57056 -66824 57406 -66630
rect 57056 -67120 57410 -66824
rect 57058 -67145 57410 -67120
rect 55000 -67438 55630 -67426
rect 55000 -67728 55640 -67438
rect 55000 -68338 55640 -68048
rect 55000 -68350 55630 -68338
rect 56280 -68506 56742 -67268
rect 58894 -67247 59732 -66697
rect 53850 -69456 55088 -68638
rect 58894 -68604 59346 -67247
rect 60405 -68226 61056 -67690
rect 60406 -68370 61056 -68226
rect 57056 -69260 57416 -68640
rect 58894 -69154 59732 -68604
rect 53860 -72540 55098 -71722
rect 57056 -72224 57406 -72030
rect 57056 -72520 57410 -72224
rect 57058 -72545 57410 -72520
rect 55000 -72838 55630 -72826
rect 55000 -73128 55640 -72838
rect 55000 -73738 55640 -73448
rect 55000 -73750 55630 -73738
rect 56280 -73906 56742 -72668
rect 58894 -72647 59732 -72097
rect 53850 -74856 55088 -74038
rect 58894 -74004 59346 -72647
rect 60405 -73626 61056 -73090
rect 60406 -73770 61056 -73626
rect 57056 -74660 57416 -74040
rect 58894 -74554 59732 -74004
rect 53860 -77940 55098 -77122
rect 57056 -77624 57406 -77430
rect 57056 -77920 57410 -77624
rect 57058 -77945 57410 -77920
rect 55000 -78238 55630 -78226
rect 55000 -78528 55640 -78238
rect 55000 -79138 55640 -78848
rect 55000 -79150 55630 -79138
rect 56280 -79306 56742 -78068
rect 58894 -78047 59732 -77497
rect 53850 -80256 55088 -79438
rect 58894 -79404 59346 -78047
rect 60405 -79026 61056 -78490
rect 60406 -79170 61056 -79026
rect 57056 -80060 57416 -79440
rect 58894 -79954 59732 -79404
rect 53860 -83340 55098 -82522
rect 57056 -83024 57406 -82830
rect 57056 -83320 57410 -83024
rect 57058 -83345 57410 -83320
rect 55000 -83638 55630 -83626
rect 55000 -83928 55640 -83638
rect 55000 -84538 55640 -84248
rect 55000 -84550 55630 -84538
rect 56280 -84706 56742 -83468
rect 58894 -83447 59732 -82897
rect 53850 -85656 55088 -84838
rect 58894 -84804 59346 -83447
rect 60405 -84426 61056 -83890
rect 60406 -84570 61056 -84426
rect 57056 -85460 57416 -84840
rect 58894 -85354 59732 -84804
<< pwell >>
rect 53314 -2628 53826 -1968
rect 55140 -2458 55562 -2030
rect 55670 -2458 56182 -1918
rect 57097 -2430 57371 -2429
rect 54834 -2626 56182 -2458
rect 54834 -2628 55000 -2626
rect 53314 -2928 55000 -2628
rect 55630 -2638 56182 -2626
rect 55640 -2928 56182 -2638
rect 53314 -3248 56182 -2928
rect 53314 -3546 55000 -3248
rect 55640 -3538 56182 -3248
rect 53314 -4206 53826 -3546
rect 54834 -3550 55000 -3546
rect 55630 -3550 56182 -3538
rect 54834 -3708 56182 -3550
rect 57086 -2810 57376 -2430
rect 59826 -2220 59976 -2130
rect 55130 -4146 55552 -3708
rect 55670 -4252 56182 -3708
rect 57008 -3760 57462 -3318
rect 59736 -2560 60556 -2220
rect 59352 -2666 60556 -2560
rect 59352 -3073 60090 -2666
rect 61106 -2780 61366 -2760
rect 60165 -2957 60347 -2939
rect 60127 -2991 60347 -2957
rect 59351 -3180 60090 -3073
rect 59351 -3590 60089 -3180
rect 60165 -3377 60347 -2991
rect 60196 -3590 60276 -3377
rect 61106 -2900 61386 -2780
rect 61106 -2939 61376 -2900
rect 61105 -2960 61376 -2939
rect 61105 -2991 61325 -2960
rect 61105 -3377 61287 -2991
rect 59351 -3693 60556 -3590
rect 55140 -4830 55698 -4408
rect 59736 -4032 60556 -3693
rect 20120 -12107 20562 -11780
rect 53314 -8028 53826 -7368
rect 55140 -7858 55562 -7430
rect 55670 -7858 56182 -7318
rect 57097 -7830 57371 -7829
rect 54834 -8026 56182 -7858
rect 54834 -8028 55000 -8026
rect 53314 -8328 55000 -8028
rect 55630 -8038 56182 -8026
rect 55640 -8328 56182 -8038
rect 53314 -8648 56182 -8328
rect 53314 -8946 55000 -8648
rect 55640 -8938 56182 -8648
rect 53314 -9606 53826 -8946
rect 54834 -8950 55000 -8946
rect 55630 -8950 56182 -8938
rect 54834 -9108 56182 -8950
rect 57086 -8210 57376 -7830
rect 59826 -7620 59976 -7530
rect 55130 -9546 55552 -9108
rect 55670 -9652 56182 -9108
rect 57008 -9160 57462 -8718
rect 59736 -7960 60556 -7620
rect 59352 -8066 60556 -7960
rect 59352 -8473 60090 -8066
rect 61106 -8180 61366 -8160
rect 60165 -8357 60347 -8339
rect 60127 -8391 60347 -8357
rect 59351 -8580 60090 -8473
rect 59351 -8990 60089 -8580
rect 60165 -8777 60347 -8391
rect 60196 -8990 60276 -8777
rect 61106 -8300 61386 -8180
rect 61106 -8339 61376 -8300
rect 61105 -8360 61376 -8339
rect 61105 -8391 61325 -8360
rect 61105 -8777 61287 -8391
rect 59351 -9093 60556 -8990
rect 55140 -10230 55698 -9808
rect 59736 -9432 60556 -9093
rect 16403 -13327 25441 -12107
rect 16400 -16200 34752 -13350
rect 53314 -13428 53826 -12768
rect 55140 -13258 55562 -12830
rect 55670 -13258 56182 -12718
rect 57097 -13230 57371 -13229
rect 54834 -13426 56182 -13258
rect 54834 -13428 55000 -13426
rect 53314 -13728 55000 -13428
rect 55630 -13438 56182 -13426
rect 55640 -13728 56182 -13438
rect 53314 -14048 56182 -13728
rect 53314 -14346 55000 -14048
rect 55640 -14338 56182 -14048
rect 53314 -15006 53826 -14346
rect 54834 -14350 55000 -14346
rect 55630 -14350 56182 -14338
rect 54834 -14508 56182 -14350
rect 57086 -13610 57376 -13230
rect 59826 -13020 59976 -12930
rect 55130 -14946 55552 -14508
rect 55670 -15052 56182 -14508
rect 57008 -14560 57462 -14118
rect 59736 -13360 60556 -13020
rect 59352 -13466 60556 -13360
rect 59352 -13873 60090 -13466
rect 61106 -13580 61366 -13560
rect 60165 -13757 60347 -13739
rect 60127 -13791 60347 -13757
rect 59351 -13980 60090 -13873
rect 59351 -14390 60089 -13980
rect 60165 -14177 60347 -13791
rect 60196 -14390 60276 -14177
rect 61106 -13700 61386 -13580
rect 61106 -13739 61376 -13700
rect 61105 -13760 61376 -13739
rect 61105 -13791 61325 -13760
rect 61105 -14177 61287 -13791
rect 59351 -14493 60556 -14390
rect 55140 -15630 55698 -15208
rect 59736 -14832 60556 -14493
rect 53314 -18828 53826 -18168
rect 55140 -18658 55562 -18230
rect 55670 -18658 56182 -18118
rect 57097 -18630 57371 -18629
rect 54834 -18826 56182 -18658
rect 54834 -18828 55000 -18826
rect 53314 -19128 55000 -18828
rect 55630 -18838 56182 -18826
rect 55640 -19128 56182 -18838
rect 53314 -19448 56182 -19128
rect 53314 -19746 55000 -19448
rect 55640 -19738 56182 -19448
rect 53314 -20406 53826 -19746
rect 54834 -19750 55000 -19746
rect 55630 -19750 56182 -19738
rect 54834 -19908 56182 -19750
rect 57086 -19010 57376 -18630
rect 59826 -18420 59976 -18330
rect 55130 -20346 55552 -19908
rect 55670 -20452 56182 -19908
rect 57008 -19960 57462 -19518
rect 59736 -18760 60556 -18420
rect 59352 -18866 60556 -18760
rect 59352 -19273 60090 -18866
rect 61106 -18980 61366 -18960
rect 60165 -19157 60347 -19139
rect 60127 -19191 60347 -19157
rect 59351 -19380 60090 -19273
rect 59351 -19790 60089 -19380
rect 60165 -19577 60347 -19191
rect 60196 -19790 60276 -19577
rect 61106 -19100 61386 -18980
rect 61106 -19139 61376 -19100
rect 61105 -19160 61376 -19139
rect 61105 -19191 61325 -19160
rect 61105 -19577 61287 -19191
rect 59351 -19893 60556 -19790
rect 55140 -21030 55698 -20608
rect 59736 -20232 60556 -19893
rect 53314 -24228 53826 -23568
rect 55140 -24058 55562 -23630
rect 55670 -24058 56182 -23518
rect 57097 -24030 57371 -24029
rect 54834 -24226 56182 -24058
rect 54834 -24228 55000 -24226
rect 53314 -24528 55000 -24228
rect 55630 -24238 56182 -24226
rect 55640 -24528 56182 -24238
rect 53314 -24848 56182 -24528
rect 53314 -25146 55000 -24848
rect 55640 -25138 56182 -24848
rect 53314 -25806 53826 -25146
rect 54834 -25150 55000 -25146
rect 55630 -25150 56182 -25138
rect 54834 -25308 56182 -25150
rect 57086 -24410 57376 -24030
rect 59826 -23820 59976 -23730
rect 55130 -25746 55552 -25308
rect 55670 -25852 56182 -25308
rect 57008 -25360 57462 -24918
rect 59736 -24160 60556 -23820
rect 59352 -24266 60556 -24160
rect 59352 -24673 60090 -24266
rect 61106 -24380 61366 -24360
rect 60165 -24557 60347 -24539
rect 60127 -24591 60347 -24557
rect 59351 -24780 60090 -24673
rect 59351 -25190 60089 -24780
rect 60165 -24977 60347 -24591
rect 60196 -25190 60276 -24977
rect 61106 -24500 61386 -24380
rect 61106 -24539 61376 -24500
rect 61105 -24560 61376 -24539
rect 61105 -24591 61325 -24560
rect 61105 -24977 61287 -24591
rect 59351 -25293 60556 -25190
rect 55140 -26430 55698 -26008
rect 59736 -25632 60556 -25293
rect 53314 -29628 53826 -28968
rect 55140 -29458 55562 -29030
rect 55670 -29458 56182 -28918
rect 57097 -29430 57371 -29429
rect 54834 -29626 56182 -29458
rect 54834 -29628 55000 -29626
rect 53314 -29928 55000 -29628
rect 55630 -29638 56182 -29626
rect 55640 -29928 56182 -29638
rect 53314 -30248 56182 -29928
rect 53314 -30546 55000 -30248
rect 55640 -30538 56182 -30248
rect 25702 -31020 35874 -30962
rect 25700 -31180 35874 -31020
rect 25702 -31280 35874 -31180
rect 53314 -31206 53826 -30546
rect 54834 -30550 55000 -30546
rect 55630 -30550 56182 -30538
rect 54834 -30708 56182 -30550
rect 57086 -29810 57376 -29430
rect 59826 -29220 59976 -29130
rect 24540 -32662 35874 -31280
rect 55130 -31146 55552 -30708
rect 55670 -31252 56182 -30708
rect 57008 -30760 57462 -30318
rect 59736 -29560 60556 -29220
rect 59352 -29666 60556 -29560
rect 59352 -30073 60090 -29666
rect 61106 -29780 61366 -29760
rect 60165 -29957 60347 -29939
rect 60127 -29991 60347 -29957
rect 59351 -30180 60090 -30073
rect 59351 -30590 60089 -30180
rect 60165 -30377 60347 -29991
rect 60196 -30590 60276 -30377
rect 61106 -29900 61386 -29780
rect 61106 -29939 61376 -29900
rect 61105 -29960 61376 -29939
rect 61105 -29991 61325 -29960
rect 61105 -30377 61287 -29991
rect 59351 -30693 60556 -30590
rect 55140 -31830 55698 -31408
rect 59736 -31032 60556 -30693
rect 24540 -38962 35872 -32662
rect 53314 -35028 53826 -34368
rect 55140 -34858 55562 -34430
rect 55670 -34858 56182 -34318
rect 57097 -34830 57371 -34829
rect 54834 -35026 56182 -34858
rect 54834 -35028 55000 -35026
rect 53314 -35328 55000 -35028
rect 55630 -35038 56182 -35026
rect 55640 -35328 56182 -35038
rect 53314 -35648 56182 -35328
rect 53314 -35946 55000 -35648
rect 55640 -35938 56182 -35648
rect 53314 -36606 53826 -35946
rect 54834 -35950 55000 -35946
rect 55630 -35950 56182 -35938
rect 54834 -36108 56182 -35950
rect 57086 -35210 57376 -34830
rect 59826 -34620 59976 -34530
rect 55130 -36546 55552 -36108
rect 55670 -36652 56182 -36108
rect 57008 -36160 57462 -35718
rect 59736 -34960 60556 -34620
rect 59352 -35066 60556 -34960
rect 59352 -35473 60090 -35066
rect 61106 -35180 61366 -35160
rect 60165 -35357 60347 -35339
rect 60127 -35391 60347 -35357
rect 59351 -35580 60090 -35473
rect 59351 -35990 60089 -35580
rect 60165 -35777 60347 -35391
rect 60196 -35990 60276 -35777
rect 61106 -35300 61386 -35180
rect 61106 -35339 61376 -35300
rect 61105 -35360 61376 -35339
rect 61105 -35391 61325 -35360
rect 61105 -35777 61287 -35391
rect 59351 -36093 60556 -35990
rect 55140 -37230 55698 -36808
rect 59736 -36432 60556 -36093
rect 75490 -38600 77260 -38330
rect 24540 -40662 35874 -38962
rect 53314 -40428 53826 -39768
rect 77940 -39400 78129 -39399
rect 78398 -39400 78589 -39399
rect 78819 -39400 79009 -39399
rect 55140 -40258 55562 -39830
rect 55670 -40258 56182 -39718
rect 57097 -40230 57371 -40229
rect 54834 -40426 56182 -40258
rect 54834 -40428 55000 -40426
rect 24540 -53352 35872 -40662
rect 53314 -40728 55000 -40428
rect 55630 -40438 56182 -40426
rect 55640 -40728 56182 -40438
rect 53314 -41048 56182 -40728
rect 53314 -41346 55000 -41048
rect 55640 -41338 56182 -41048
rect 53314 -42006 53826 -41346
rect 54834 -41350 55000 -41346
rect 55630 -41350 56182 -41338
rect 54834 -41508 56182 -41350
rect 57086 -40610 57376 -40230
rect 77340 -39850 79030 -39400
rect 77579 -39851 78129 -39850
rect 77940 -39891 78129 -39851
rect 59826 -40020 59976 -39930
rect 80730 -39940 88880 -39440
rect 55130 -41946 55552 -41508
rect 55670 -42052 56182 -41508
rect 57008 -41560 57462 -41118
rect 59736 -40360 60556 -40020
rect 59352 -40466 60556 -40360
rect 59352 -40873 60090 -40466
rect 61106 -40580 61366 -40560
rect 60165 -40757 60347 -40739
rect 60127 -40791 60347 -40757
rect 59351 -40980 60090 -40873
rect 59351 -41390 60089 -40980
rect 60165 -41177 60347 -40791
rect 60196 -41390 60276 -41177
rect 61106 -40700 61386 -40580
rect 83000 -40290 83640 -39940
rect 87800 -39980 88840 -39940
rect 87520 -40220 88840 -39980
rect 77807 -40660 77997 -40649
rect 61106 -40739 61376 -40700
rect 61105 -40760 61376 -40739
rect 61105 -40791 61325 -40760
rect 61105 -41177 61287 -40791
rect 77340 -41110 78590 -40660
rect 87520 -40890 88480 -40220
rect 88690 -40270 88840 -40220
rect 77611 -41113 77997 -41110
rect 77807 -41131 77997 -41113
rect 78400 -41131 78589 -41110
rect 59351 -41493 60556 -41390
rect 55140 -42630 55698 -42208
rect 59736 -41832 60556 -41493
rect 77807 -41900 77997 -41889
rect 77340 -42380 78030 -41900
rect 77809 -42385 77999 -42380
rect 77340 -43140 77750 -43130
rect 77830 -43140 78240 -43130
rect 78310 -43140 78340 -43130
rect 78480 -43140 78520 -43130
rect 78600 -43139 78780 -43130
rect 78600 -43140 78873 -43139
rect 77340 -43620 78880 -43140
rect 53314 -45828 53826 -45168
rect 77340 -44860 78230 -44360
rect 82790 -44410 91440 -43940
rect 55140 -45658 55562 -45230
rect 55670 -45658 56182 -45118
rect 57097 -45630 57371 -45629
rect 54834 -45826 56182 -45658
rect 54834 -45828 55000 -45826
rect 53314 -46128 55000 -45828
rect 55630 -45838 56182 -45826
rect 55640 -46128 56182 -45838
rect 53314 -46448 56182 -46128
rect 53314 -46746 55000 -46448
rect 55640 -46738 56182 -46448
rect 53314 -47406 53826 -46746
rect 54834 -46750 55000 -46746
rect 55630 -46750 56182 -46738
rect 54834 -46908 56182 -46750
rect 57086 -46010 57376 -45630
rect 59826 -45420 59976 -45330
rect 55130 -47346 55552 -46908
rect 55670 -47452 56182 -46908
rect 57008 -46960 57462 -46518
rect 59736 -45760 60556 -45420
rect 59352 -45866 60556 -45760
rect 77340 -45620 78670 -45590
rect 78750 -45620 79060 -45590
rect 77340 -45800 79060 -45620
rect 77607 -45829 77641 -45800
rect 78067 -45829 78101 -45800
rect 78528 -45829 78562 -45800
rect 59352 -46273 60090 -45866
rect 61106 -45980 61366 -45960
rect 60165 -46157 60347 -46139
rect 60127 -46191 60347 -46157
rect 59351 -46380 60090 -46273
rect 59351 -46790 60089 -46380
rect 60165 -46577 60347 -46191
rect 60196 -46790 60276 -46577
rect 61106 -46100 61386 -45980
rect 61106 -46139 61376 -46100
rect 61105 -46160 61376 -46139
rect 61105 -46191 61325 -46160
rect 61105 -46577 61287 -46191
rect 75490 -46640 77260 -46370
rect 59351 -46893 60556 -46790
rect 55140 -48030 55698 -47608
rect 59736 -47232 60556 -46893
rect 77940 -47440 78129 -47439
rect 78398 -47440 78589 -47439
rect 78819 -47440 79009 -47439
rect 77340 -47890 79030 -47440
rect 77579 -47891 78129 -47890
rect 77940 -47931 78129 -47891
rect 82794 -48548 91444 -48078
rect 77807 -48700 77997 -48689
rect 77340 -49150 78590 -48700
rect 77611 -49153 77997 -49150
rect 77807 -49171 77997 -49153
rect 78400 -49171 78589 -49150
rect 77807 -49940 77997 -49929
rect 53314 -51228 53826 -50568
rect 77340 -50420 78030 -49940
rect 77809 -50425 77999 -50420
rect 55140 -51058 55562 -50630
rect 55670 -51058 56182 -50518
rect 57097 -51030 57371 -51029
rect 54834 -51226 56182 -51058
rect 54834 -51228 55000 -51226
rect 53314 -51528 55000 -51228
rect 55630 -51238 56182 -51226
rect 55640 -51528 56182 -51238
rect 53314 -51848 56182 -51528
rect 53314 -52146 55000 -51848
rect 55640 -52138 56182 -51848
rect 53314 -52806 53826 -52146
rect 54834 -52150 55000 -52146
rect 55630 -52150 56182 -52138
rect 54834 -52308 56182 -52150
rect 57086 -51410 57376 -51030
rect 59826 -50820 59976 -50730
rect 55130 -52746 55552 -52308
rect 55670 -52852 56182 -52308
rect 57008 -52360 57462 -51918
rect 59736 -51160 60556 -50820
rect 59352 -51266 60556 -51160
rect 77340 -51180 77750 -51170
rect 77830 -51180 78240 -51170
rect 78310 -51180 78340 -51170
rect 78480 -51180 78520 -51170
rect 78600 -51179 78780 -51170
rect 78600 -51180 78873 -51179
rect 59352 -51673 60090 -51266
rect 61106 -51380 61366 -51360
rect 60165 -51557 60347 -51539
rect 60127 -51591 60347 -51557
rect 59351 -51780 60090 -51673
rect 59351 -52190 60089 -51780
rect 60165 -51977 60347 -51591
rect 60196 -52190 60276 -51977
rect 61106 -51500 61386 -51380
rect 61106 -51539 61376 -51500
rect 61105 -51560 61376 -51539
rect 61105 -51591 61325 -51560
rect 61105 -51977 61287 -51591
rect 77340 -51660 78880 -51180
rect 59351 -52293 60556 -52190
rect 24540 -55052 35874 -53352
rect 55140 -53430 55698 -53008
rect 59736 -52632 60556 -52293
rect 82790 -52200 91440 -51730
rect 77340 -52900 78230 -52400
rect 77340 -53660 78670 -53630
rect 78750 -53660 79060 -53630
rect 77340 -53840 79060 -53660
rect 77607 -53869 77641 -53840
rect 78067 -53869 78101 -53840
rect 78528 -53869 78562 -53840
rect 24540 -57880 35872 -55052
rect 25700 -58250 35872 -57880
rect 53314 -56628 53826 -55968
rect 55140 -56458 55562 -56030
rect 55670 -56458 56182 -55918
rect 57097 -56430 57371 -56429
rect 54834 -56626 56182 -56458
rect 54834 -56628 55000 -56626
rect 53314 -56928 55000 -56628
rect 55630 -56638 56182 -56626
rect 55640 -56928 56182 -56638
rect 53314 -57248 56182 -56928
rect 53314 -57546 55000 -57248
rect 55640 -57538 56182 -57248
rect 53314 -58206 53826 -57546
rect 54834 -57550 55000 -57546
rect 55630 -57550 56182 -57538
rect 54834 -57708 56182 -57550
rect 57086 -56810 57376 -56430
rect 59826 -56220 59976 -56130
rect 55130 -58146 55552 -57708
rect 55670 -58252 56182 -57708
rect 57008 -57760 57462 -57318
rect 59736 -56560 60556 -56220
rect 59352 -56666 60556 -56560
rect 59352 -57073 60090 -56666
rect 61106 -56780 61366 -56760
rect 60165 -56957 60347 -56939
rect 60127 -56991 60347 -56957
rect 59351 -57180 60090 -57073
rect 59351 -57590 60089 -57180
rect 60165 -57377 60347 -56991
rect 60196 -57590 60276 -57377
rect 61106 -56900 61386 -56780
rect 61106 -56939 61376 -56900
rect 61105 -56960 61376 -56939
rect 61105 -56991 61325 -56960
rect 61105 -57377 61287 -56991
rect 59351 -57693 60556 -57590
rect 55140 -58830 55698 -58408
rect 59736 -58032 60556 -57693
rect 53314 -62028 53826 -61368
rect 55140 -61858 55562 -61430
rect 55670 -61858 56182 -61318
rect 57097 -61830 57371 -61829
rect 54834 -62026 56182 -61858
rect 54834 -62028 55000 -62026
rect 53314 -62328 55000 -62028
rect 55630 -62038 56182 -62026
rect 55640 -62328 56182 -62038
rect 53314 -62648 56182 -62328
rect 53314 -62946 55000 -62648
rect 55640 -62938 56182 -62648
rect 53314 -63606 53826 -62946
rect 54834 -62950 55000 -62946
rect 55630 -62950 56182 -62938
rect 54834 -63108 56182 -62950
rect 57086 -62210 57376 -61830
rect 59826 -61620 59976 -61530
rect 55130 -63546 55552 -63108
rect 55670 -63652 56182 -63108
rect 57008 -63160 57462 -62718
rect 59736 -61960 60556 -61620
rect 59352 -62066 60556 -61960
rect 59352 -62473 60090 -62066
rect 61106 -62180 61366 -62160
rect 60165 -62357 60347 -62339
rect 60127 -62391 60347 -62357
rect 59351 -62580 60090 -62473
rect 59351 -62990 60089 -62580
rect 60165 -62777 60347 -62391
rect 60196 -62990 60276 -62777
rect 61106 -62300 61386 -62180
rect 61106 -62339 61376 -62300
rect 61105 -62360 61376 -62339
rect 61105 -62391 61325 -62360
rect 61105 -62777 61287 -62391
rect 59351 -63093 60556 -62990
rect 55140 -64230 55698 -63808
rect 59736 -63432 60556 -63093
rect 53314 -67428 53826 -66768
rect 55140 -67258 55562 -66830
rect 55670 -67258 56182 -66718
rect 57097 -67230 57371 -67229
rect 54834 -67426 56182 -67258
rect 54834 -67428 55000 -67426
rect 53314 -67728 55000 -67428
rect 55630 -67438 56182 -67426
rect 55640 -67728 56182 -67438
rect 53314 -68048 56182 -67728
rect 53314 -68346 55000 -68048
rect 55640 -68338 56182 -68048
rect 53314 -69006 53826 -68346
rect 54834 -68350 55000 -68346
rect 55630 -68350 56182 -68338
rect 54834 -68508 56182 -68350
rect 57086 -67610 57376 -67230
rect 59826 -67020 59976 -66930
rect 55130 -68946 55552 -68508
rect 55670 -69052 56182 -68508
rect 57008 -68560 57462 -68118
rect 59736 -67360 60556 -67020
rect 59352 -67466 60556 -67360
rect 59352 -67873 60090 -67466
rect 61106 -67580 61366 -67560
rect 60165 -67757 60347 -67739
rect 60127 -67791 60347 -67757
rect 59351 -67980 60090 -67873
rect 59351 -68390 60089 -67980
rect 60165 -68177 60347 -67791
rect 60196 -68390 60276 -68177
rect 61106 -67700 61386 -67580
rect 61106 -67739 61376 -67700
rect 61105 -67760 61376 -67739
rect 61105 -67791 61325 -67760
rect 61105 -68177 61287 -67791
rect 59351 -68493 60556 -68390
rect 55140 -69630 55698 -69208
rect 59736 -68832 60556 -68493
rect 53314 -72828 53826 -72168
rect 55140 -72658 55562 -72230
rect 55670 -72658 56182 -72118
rect 57097 -72630 57371 -72629
rect 54834 -72826 56182 -72658
rect 54834 -72828 55000 -72826
rect 53314 -73128 55000 -72828
rect 55630 -72838 56182 -72826
rect 55640 -73128 56182 -72838
rect 53314 -73448 56182 -73128
rect 53314 -73746 55000 -73448
rect 55640 -73738 56182 -73448
rect 53314 -74406 53826 -73746
rect 54834 -73750 55000 -73746
rect 55630 -73750 56182 -73738
rect 54834 -73908 56182 -73750
rect 57086 -73010 57376 -72630
rect 59826 -72420 59976 -72330
rect 55130 -74346 55552 -73908
rect 55670 -74452 56182 -73908
rect 57008 -73960 57462 -73518
rect 59736 -72760 60556 -72420
rect 59352 -72866 60556 -72760
rect 59352 -73273 60090 -72866
rect 61106 -72980 61366 -72960
rect 60165 -73157 60347 -73139
rect 60127 -73191 60347 -73157
rect 59351 -73380 60090 -73273
rect 59351 -73790 60089 -73380
rect 60165 -73577 60347 -73191
rect 60196 -73790 60276 -73577
rect 61106 -73100 61386 -72980
rect 61106 -73139 61376 -73100
rect 61105 -73160 61376 -73139
rect 61105 -73191 61325 -73160
rect 61105 -73577 61287 -73191
rect 59351 -73893 60556 -73790
rect 55140 -75030 55698 -74608
rect 59736 -74232 60556 -73893
rect 53314 -78228 53826 -77568
rect 55140 -78058 55562 -77630
rect 55670 -78058 56182 -77518
rect 57097 -78030 57371 -78029
rect 54834 -78226 56182 -78058
rect 54834 -78228 55000 -78226
rect 53314 -78528 55000 -78228
rect 55630 -78238 56182 -78226
rect 55640 -78528 56182 -78238
rect 53314 -78848 56182 -78528
rect 53314 -79146 55000 -78848
rect 55640 -79138 56182 -78848
rect 53314 -79806 53826 -79146
rect 54834 -79150 55000 -79146
rect 55630 -79150 56182 -79138
rect 54834 -79308 56182 -79150
rect 57086 -78410 57376 -78030
rect 59826 -77820 59976 -77730
rect 55130 -79746 55552 -79308
rect 55670 -79852 56182 -79308
rect 57008 -79360 57462 -78918
rect 59736 -78160 60556 -77820
rect 59352 -78266 60556 -78160
rect 59352 -78673 60090 -78266
rect 61106 -78380 61366 -78360
rect 60165 -78557 60347 -78539
rect 60127 -78591 60347 -78557
rect 59351 -78780 60090 -78673
rect 59351 -79190 60089 -78780
rect 60165 -78977 60347 -78591
rect 60196 -79190 60276 -78977
rect 61106 -78500 61386 -78380
rect 61106 -78539 61376 -78500
rect 61105 -78560 61376 -78539
rect 61105 -78591 61325 -78560
rect 61105 -78977 61287 -78591
rect 59351 -79293 60556 -79190
rect 55140 -80430 55698 -80008
rect 59736 -79632 60556 -79293
rect 53314 -83628 53826 -82968
rect 55140 -83458 55562 -83030
rect 55670 -83458 56182 -82918
rect 57097 -83430 57371 -83429
rect 54834 -83626 56182 -83458
rect 54834 -83628 55000 -83626
rect 53314 -83928 55000 -83628
rect 55630 -83638 56182 -83626
rect 55640 -83928 56182 -83638
rect 53314 -84248 56182 -83928
rect 53314 -84546 55000 -84248
rect 55640 -84538 56182 -84248
rect 53314 -85206 53826 -84546
rect 54834 -84550 55000 -84546
rect 55630 -84550 56182 -84538
rect 54834 -84708 56182 -84550
rect 57086 -83810 57376 -83430
rect 59826 -83220 59976 -83130
rect 55130 -85146 55552 -84708
rect 55670 -85252 56182 -84708
rect 57008 -84760 57462 -84318
rect 59736 -83560 60556 -83220
rect 59352 -83666 60556 -83560
rect 59352 -84073 60090 -83666
rect 61106 -83780 61366 -83760
rect 60165 -83957 60347 -83939
rect 60127 -83991 60347 -83957
rect 59351 -84180 60090 -84073
rect 59351 -84590 60089 -84180
rect 60165 -84377 60347 -83991
rect 60196 -84590 60276 -84377
rect 61106 -83900 61386 -83780
rect 61106 -83939 61376 -83900
rect 61105 -83960 61376 -83939
rect 61105 -83991 61325 -83960
rect 61105 -84377 61287 -83991
rect 59351 -84693 60556 -84590
rect 55140 -85830 55698 -85408
rect 59736 -85032 60556 -84693
<< nmos >>
rect 59946 -2470 60346 -2420
rect 59548 -2970 59578 -2770
rect 59864 -2970 59894 -2770
rect 59547 -3483 59577 -3283
rect 59863 -3483 59893 -3283
rect 59946 -3836 60346 -3786
rect 59946 -7870 60346 -7820
rect 59548 -8370 59578 -8170
rect 59864 -8370 59894 -8170
rect 59547 -8883 59577 -8683
rect 59863 -8883 59893 -8683
rect 59946 -9236 60346 -9186
rect 59946 -13270 60346 -13220
rect 59548 -13770 59578 -13570
rect 59864 -13770 59894 -13570
rect 59547 -14283 59577 -14083
rect 59863 -14283 59893 -14083
rect 59946 -14636 60346 -14586
rect 59946 -18670 60346 -18620
rect 59548 -19170 59578 -18970
rect 59864 -19170 59894 -18970
rect 59547 -19683 59577 -19483
rect 59863 -19683 59893 -19483
rect 59946 -20036 60346 -19986
rect 59946 -24070 60346 -24020
rect 59548 -24570 59578 -24370
rect 59864 -24570 59894 -24370
rect 59547 -25083 59577 -24883
rect 59863 -25083 59893 -24883
rect 59946 -25436 60346 -25386
rect 59946 -29470 60346 -29420
rect 59548 -29970 59578 -29770
rect 59864 -29970 59894 -29770
rect 59547 -30483 59577 -30283
rect 59863 -30483 59893 -30283
rect 59946 -30836 60346 -30786
rect 59946 -34870 60346 -34820
rect 59548 -35370 59578 -35170
rect 59864 -35370 59894 -35170
rect 59547 -35883 59577 -35683
rect 59863 -35883 59893 -35683
rect 59946 -36236 60346 -36186
rect 59946 -40270 60346 -40220
rect 59548 -40770 59578 -40570
rect 59864 -40770 59894 -40570
rect 59547 -41283 59577 -41083
rect 59863 -41283 59893 -41083
rect 59946 -41636 60346 -41586
rect 59946 -45670 60346 -45620
rect 59548 -46170 59578 -45970
rect 59864 -46170 59894 -45970
rect 59547 -46683 59577 -46483
rect 59863 -46683 59893 -46483
rect 59946 -47036 60346 -46986
rect 59946 -51070 60346 -51020
rect 59548 -51570 59578 -51370
rect 59864 -51570 59894 -51370
rect 59547 -52083 59577 -51883
rect 59863 -52083 59893 -51883
rect 59946 -52436 60346 -52386
rect 59946 -56470 60346 -56420
rect 59548 -56970 59578 -56770
rect 59864 -56970 59894 -56770
rect 59547 -57483 59577 -57283
rect 59863 -57483 59893 -57283
rect 59946 -57836 60346 -57786
rect 59946 -61870 60346 -61820
rect 59548 -62370 59578 -62170
rect 59864 -62370 59894 -62170
rect 59547 -62883 59577 -62683
rect 59863 -62883 59893 -62683
rect 59946 -63236 60346 -63186
rect 59946 -67270 60346 -67220
rect 59548 -67770 59578 -67570
rect 59864 -67770 59894 -67570
rect 59547 -68283 59577 -68083
rect 59863 -68283 59893 -68083
rect 59946 -68636 60346 -68586
rect 59946 -72670 60346 -72620
rect 59548 -73170 59578 -72970
rect 59864 -73170 59894 -72970
rect 59547 -73683 59577 -73483
rect 59863 -73683 59893 -73483
rect 59946 -74036 60346 -73986
rect 59946 -78070 60346 -78020
rect 59548 -78570 59578 -78370
rect 59864 -78570 59894 -78370
rect 59547 -79083 59577 -78883
rect 59863 -79083 59893 -78883
rect 59946 -79436 60346 -79386
rect 59946 -83470 60346 -83420
rect 59548 -83970 59578 -83770
rect 59864 -83970 59894 -83770
rect 59547 -84483 59577 -84283
rect 59863 -84483 59893 -84283
rect 59946 -84836 60346 -84786
<< scnmos >>
rect 57175 -2559 57205 -2455
rect 57263 -2559 57293 -2455
rect 60191 -3047 60321 -3017
rect 61131 -3047 61261 -3017
rect 57175 -3733 57205 -3629
rect 57263 -3733 57293 -3629
rect 60191 -3131 60321 -3101
rect 61131 -3131 61261 -3101
rect 60191 -3215 60321 -3185
rect 61131 -3215 61261 -3185
rect 60191 -3299 60321 -3269
rect 61131 -3299 61261 -3269
rect 57175 -7959 57205 -7855
rect 57263 -7959 57293 -7855
rect 60191 -8447 60321 -8417
rect 61131 -8447 61261 -8417
rect 57175 -9133 57205 -9029
rect 57263 -9133 57293 -9029
rect 60191 -8531 60321 -8501
rect 61131 -8531 61261 -8501
rect 60191 -8615 60321 -8585
rect 61131 -8615 61261 -8585
rect 60191 -8699 60321 -8669
rect 61131 -8699 61261 -8669
rect 57175 -13359 57205 -13255
rect 57263 -13359 57293 -13255
rect 60191 -13847 60321 -13817
rect 61131 -13847 61261 -13817
rect 57175 -14533 57205 -14429
rect 57263 -14533 57293 -14429
rect 60191 -13931 60321 -13901
rect 61131 -13931 61261 -13901
rect 60191 -14015 60321 -13985
rect 61131 -14015 61261 -13985
rect 60191 -14099 60321 -14069
rect 61131 -14099 61261 -14069
rect 57175 -18759 57205 -18655
rect 57263 -18759 57293 -18655
rect 60191 -19247 60321 -19217
rect 61131 -19247 61261 -19217
rect 57175 -19933 57205 -19829
rect 57263 -19933 57293 -19829
rect 60191 -19331 60321 -19301
rect 61131 -19331 61261 -19301
rect 60191 -19415 60321 -19385
rect 61131 -19415 61261 -19385
rect 60191 -19499 60321 -19469
rect 61131 -19499 61261 -19469
rect 57175 -24159 57205 -24055
rect 57263 -24159 57293 -24055
rect 60191 -24647 60321 -24617
rect 61131 -24647 61261 -24617
rect 57175 -25333 57205 -25229
rect 57263 -25333 57293 -25229
rect 60191 -24731 60321 -24701
rect 61131 -24731 61261 -24701
rect 60191 -24815 60321 -24785
rect 61131 -24815 61261 -24785
rect 60191 -24899 60321 -24869
rect 61131 -24899 61261 -24869
rect 57175 -29559 57205 -29455
rect 57263 -29559 57293 -29455
rect 60191 -30047 60321 -30017
rect 61131 -30047 61261 -30017
rect 57175 -30733 57205 -30629
rect 57263 -30733 57293 -30629
rect 60191 -30131 60321 -30101
rect 61131 -30131 61261 -30101
rect 60191 -30215 60321 -30185
rect 61131 -30215 61261 -30185
rect 60191 -30299 60321 -30269
rect 61131 -30299 61261 -30269
rect 57175 -34959 57205 -34855
rect 57263 -34959 57293 -34855
rect 60191 -35447 60321 -35417
rect 61131 -35447 61261 -35417
rect 57175 -36133 57205 -36029
rect 57263 -36133 57293 -36029
rect 60191 -35531 60321 -35501
rect 61131 -35531 61261 -35501
rect 60191 -35615 60321 -35585
rect 61131 -35615 61261 -35585
rect 60191 -35699 60321 -35669
rect 61131 -35699 61261 -35669
rect 75626 -38565 75656 -38435
rect 75902 -38565 75932 -38435
rect 76176 -38565 76206 -38435
rect 76452 -38565 76482 -38435
rect 76728 -38565 76758 -38435
rect 77657 -39549 77687 -39465
rect 77753 -39549 77783 -39465
rect 77837 -39549 77867 -39465
rect 77921 -39549 77951 -39465
rect 78019 -39555 78049 -39425
rect 78211 -39549 78241 -39465
rect 78295 -39549 78325 -39465
rect 78379 -39549 78409 -39465
rect 78477 -39555 78507 -39425
rect 78705 -39527 78735 -39443
rect 78789 -39527 78819 -39443
rect 78897 -39555 78927 -39425
rect 80858 -39605 80888 -39475
rect 81103 -39605 81133 -39475
rect 81187 -39605 81217 -39475
rect 81271 -39605 81301 -39475
rect 81355 -39605 81385 -39475
rect 81566 -39605 81596 -39475
rect 81650 -39605 81680 -39475
rect 81734 -39605 81764 -39475
rect 81818 -39605 81848 -39475
rect 81902 -39605 81932 -39475
rect 81986 -39605 82016 -39475
rect 82070 -39605 82100 -39475
rect 82154 -39605 82184 -39475
rect 82238 -39605 82268 -39475
rect 82322 -39605 82352 -39475
rect 82406 -39605 82436 -39475
rect 82490 -39605 82520 -39475
rect 82574 -39605 82604 -39475
rect 82658 -39605 82688 -39475
rect 82742 -39605 82772 -39475
rect 82826 -39605 82856 -39475
rect 83038 -39605 83068 -39475
rect 83122 -39605 83152 -39475
rect 83206 -39605 83236 -39475
rect 83290 -39605 83320 -39475
rect 83374 -39605 83404 -39475
rect 83458 -39605 83488 -39475
rect 83542 -39605 83572 -39475
rect 83626 -39605 83656 -39475
rect 83710 -39605 83740 -39475
rect 83794 -39605 83824 -39475
rect 83878 -39605 83908 -39475
rect 83962 -39605 83992 -39475
rect 84046 -39605 84076 -39475
rect 84130 -39605 84160 -39475
rect 84214 -39605 84244 -39475
rect 84298 -39605 84328 -39475
rect 84510 -39605 84540 -39475
rect 84594 -39605 84624 -39475
rect 84678 -39605 84708 -39475
rect 84762 -39605 84792 -39475
rect 84846 -39605 84876 -39475
rect 84930 -39605 84960 -39475
rect 85014 -39605 85044 -39475
rect 85098 -39605 85128 -39475
rect 85182 -39605 85212 -39475
rect 85266 -39605 85296 -39475
rect 85350 -39605 85380 -39475
rect 85434 -39605 85464 -39475
rect 85518 -39605 85548 -39475
rect 85602 -39605 85632 -39475
rect 85686 -39605 85716 -39475
rect 85770 -39605 85800 -39475
rect 85982 -39605 86012 -39475
rect 86066 -39605 86096 -39475
rect 86150 -39605 86180 -39475
rect 86234 -39605 86264 -39475
rect 86318 -39605 86348 -39475
rect 86402 -39605 86432 -39475
rect 86486 -39605 86516 -39475
rect 86570 -39605 86600 -39475
rect 86654 -39605 86684 -39475
rect 86738 -39605 86768 -39475
rect 86822 -39605 86852 -39475
rect 86906 -39605 86936 -39475
rect 86990 -39605 87020 -39475
rect 87074 -39605 87104 -39475
rect 87158 -39605 87188 -39475
rect 87242 -39605 87272 -39475
rect 87454 -39605 87484 -39475
rect 87538 -39605 87568 -39475
rect 87622 -39605 87652 -39475
rect 87706 -39605 87736 -39475
rect 87790 -39605 87820 -39475
rect 87874 -39605 87904 -39475
rect 87958 -39605 87988 -39475
rect 88042 -39605 88072 -39475
rect 88126 -39605 88156 -39475
rect 88210 -39605 88240 -39475
rect 88294 -39605 88324 -39475
rect 88378 -39605 88408 -39475
rect 88462 -39605 88492 -39475
rect 88546 -39605 88576 -39475
rect 88630 -39605 88660 -39475
rect 88714 -39605 88744 -39475
rect 77657 -39825 77687 -39741
rect 77753 -39825 77783 -39741
rect 77837 -39825 77867 -39741
rect 77921 -39825 77951 -39741
rect 78019 -39865 78049 -39735
rect 80908 -39905 80938 -39775
rect 57175 -40359 57205 -40255
rect 57263 -40359 57293 -40255
rect 77693 -40777 77723 -40693
rect 77777 -40777 77807 -40693
rect 60191 -40847 60321 -40817
rect 61131 -40847 61261 -40817
rect 77885 -40805 77915 -40675
rect 57175 -41533 57205 -41429
rect 57263 -41533 57293 -41429
rect 60191 -40931 60321 -40901
rect 61131 -40931 61261 -40901
rect 60191 -41015 60321 -40985
rect 61131 -41015 61261 -40985
rect 60191 -41099 60321 -41069
rect 61131 -41099 61261 -41069
rect 77693 -41087 77723 -41003
rect 77777 -41087 77807 -41003
rect 77885 -41105 77915 -40975
rect 78117 -41065 78147 -40981
rect 78213 -41065 78243 -40981
rect 78297 -41065 78327 -40981
rect 78381 -41065 78411 -40981
rect 78479 -41105 78509 -40975
rect 77693 -42017 77723 -41933
rect 77777 -42017 77807 -41933
rect 77885 -42045 77915 -41915
rect 77695 -42341 77725 -42257
rect 77779 -42341 77809 -42257
rect 77887 -42359 77917 -42229
rect 77657 -43295 77687 -43211
rect 77745 -43295 77775 -43211
rect 77851 -43295 77881 -43211
rect 77947 -43295 77977 -43211
rect 78113 -43295 78143 -43165
rect 78401 -43289 78431 -43205
rect 78497 -43289 78527 -43205
rect 78581 -43289 78611 -43205
rect 78665 -43289 78695 -43205
rect 78763 -43295 78793 -43165
rect 77657 -43545 77687 -43461
rect 77745 -43545 77775 -43461
rect 77851 -43545 77881 -43461
rect 77947 -43545 77977 -43461
rect 78113 -43591 78143 -43461
rect 82946 -44105 82976 -44021
rect 83030 -44105 83060 -44021
rect 83127 -44105 83157 -43975
rect 83418 -44105 83448 -43975
rect 83663 -44105 83693 -43975
rect 83747 -44105 83777 -43975
rect 83831 -44105 83861 -43975
rect 83915 -44105 83945 -43975
rect 84126 -44105 84156 -43975
rect 84210 -44105 84240 -43975
rect 84294 -44105 84324 -43975
rect 84378 -44105 84408 -43975
rect 84462 -44105 84492 -43975
rect 84546 -44105 84576 -43975
rect 84630 -44105 84660 -43975
rect 84714 -44105 84744 -43975
rect 84798 -44105 84828 -43975
rect 84882 -44105 84912 -43975
rect 84966 -44105 84996 -43975
rect 85050 -44105 85080 -43975
rect 85134 -44105 85164 -43975
rect 85218 -44105 85248 -43975
rect 85302 -44105 85332 -43975
rect 85386 -44105 85416 -43975
rect 85598 -44105 85628 -43975
rect 85682 -44105 85712 -43975
rect 85766 -44105 85796 -43975
rect 85850 -44105 85880 -43975
rect 85934 -44105 85964 -43975
rect 86018 -44105 86048 -43975
rect 86102 -44105 86132 -43975
rect 86186 -44105 86216 -43975
rect 86270 -44105 86300 -43975
rect 86354 -44105 86384 -43975
rect 86438 -44105 86468 -43975
rect 86522 -44105 86552 -43975
rect 86606 -44105 86636 -43975
rect 86690 -44105 86720 -43975
rect 86774 -44105 86804 -43975
rect 86858 -44105 86888 -43975
rect 87070 -44105 87100 -43975
rect 87154 -44105 87184 -43975
rect 87238 -44105 87268 -43975
rect 87322 -44105 87352 -43975
rect 87406 -44105 87436 -43975
rect 87490 -44105 87520 -43975
rect 87574 -44105 87604 -43975
rect 87658 -44105 87688 -43975
rect 87742 -44105 87772 -43975
rect 87826 -44105 87856 -43975
rect 87910 -44105 87940 -43975
rect 87994 -44105 88024 -43975
rect 88078 -44105 88108 -43975
rect 88162 -44105 88192 -43975
rect 88246 -44105 88276 -43975
rect 88330 -44105 88360 -43975
rect 88542 -44105 88572 -43975
rect 88626 -44105 88656 -43975
rect 88710 -44105 88740 -43975
rect 88794 -44105 88824 -43975
rect 88878 -44105 88908 -43975
rect 88962 -44105 88992 -43975
rect 89046 -44105 89076 -43975
rect 89130 -44105 89160 -43975
rect 89214 -44105 89244 -43975
rect 89298 -44105 89328 -43975
rect 89382 -44105 89412 -43975
rect 89466 -44105 89496 -43975
rect 89550 -44105 89580 -43975
rect 89634 -44105 89664 -43975
rect 89718 -44105 89748 -43975
rect 89802 -44105 89832 -43975
rect 90014 -44105 90044 -43975
rect 90098 -44105 90128 -43975
rect 90182 -44105 90212 -43975
rect 90266 -44105 90296 -43975
rect 90350 -44105 90380 -43975
rect 90434 -44105 90464 -43975
rect 90518 -44105 90548 -43975
rect 90602 -44105 90632 -43975
rect 90686 -44105 90716 -43975
rect 90770 -44105 90800 -43975
rect 90854 -44105 90884 -43975
rect 90938 -44105 90968 -43975
rect 91022 -44105 91052 -43975
rect 91106 -44105 91136 -43975
rect 91190 -44105 91220 -43975
rect 91274 -44105 91304 -43975
rect 77657 -44527 77687 -44443
rect 77745 -44527 77775 -44443
rect 77851 -44527 77881 -44443
rect 77947 -44527 77977 -44443
rect 78113 -44527 78143 -44397
rect 77657 -44779 77687 -44695
rect 77745 -44779 77775 -44695
rect 77851 -44779 77881 -44695
rect 77947 -44779 77977 -44695
rect 78113 -44825 78143 -44695
rect 57175 -45759 57205 -45655
rect 57263 -45759 57293 -45655
rect 77657 -45765 77687 -45681
rect 77729 -45765 77759 -45681
rect 77801 -45765 77831 -45681
rect 77929 -45765 77959 -45635
rect 78153 -45737 78183 -45653
rect 78237 -45737 78267 -45653
rect 78345 -45765 78375 -45635
rect 78577 -45759 78607 -45675
rect 78673 -45759 78703 -45675
rect 78757 -45759 78787 -45675
rect 78841 -45759 78871 -45675
rect 78939 -45765 78969 -45635
rect 60191 -46247 60321 -46217
rect 61131 -46247 61261 -46217
rect 57175 -46933 57205 -46829
rect 57263 -46933 57293 -46829
rect 60191 -46331 60321 -46301
rect 61131 -46331 61261 -46301
rect 60191 -46415 60321 -46385
rect 61131 -46415 61261 -46385
rect 60191 -46499 60321 -46469
rect 61131 -46499 61261 -46469
rect 75626 -46605 75656 -46475
rect 75902 -46605 75932 -46475
rect 76176 -46605 76206 -46475
rect 76452 -46605 76482 -46475
rect 76728 -46605 76758 -46475
rect 77657 -47589 77687 -47505
rect 77753 -47589 77783 -47505
rect 77837 -47589 77867 -47505
rect 77921 -47589 77951 -47505
rect 78019 -47595 78049 -47465
rect 78211 -47589 78241 -47505
rect 78295 -47589 78325 -47505
rect 78379 -47589 78409 -47505
rect 78477 -47595 78507 -47465
rect 78705 -47567 78735 -47483
rect 78789 -47567 78819 -47483
rect 78897 -47595 78927 -47465
rect 77657 -47865 77687 -47781
rect 77753 -47865 77783 -47781
rect 77837 -47865 77867 -47781
rect 77921 -47865 77951 -47781
rect 78019 -47905 78049 -47775
rect 82946 -48245 82976 -48161
rect 83030 -48245 83060 -48161
rect 83127 -48245 83157 -48115
rect 83418 -48245 83448 -48115
rect 83663 -48245 83693 -48115
rect 83747 -48245 83777 -48115
rect 83831 -48245 83861 -48115
rect 83915 -48245 83945 -48115
rect 84126 -48245 84156 -48115
rect 84210 -48245 84240 -48115
rect 84294 -48245 84324 -48115
rect 84378 -48245 84408 -48115
rect 84462 -48245 84492 -48115
rect 84546 -48245 84576 -48115
rect 84630 -48245 84660 -48115
rect 84714 -48245 84744 -48115
rect 84798 -48245 84828 -48115
rect 84882 -48245 84912 -48115
rect 84966 -48245 84996 -48115
rect 85050 -48245 85080 -48115
rect 85134 -48245 85164 -48115
rect 85218 -48245 85248 -48115
rect 85302 -48245 85332 -48115
rect 85386 -48245 85416 -48115
rect 85598 -48245 85628 -48115
rect 85682 -48245 85712 -48115
rect 85766 -48245 85796 -48115
rect 85850 -48245 85880 -48115
rect 85934 -48245 85964 -48115
rect 86018 -48245 86048 -48115
rect 86102 -48245 86132 -48115
rect 86186 -48245 86216 -48115
rect 86270 -48245 86300 -48115
rect 86354 -48245 86384 -48115
rect 86438 -48245 86468 -48115
rect 86522 -48245 86552 -48115
rect 86606 -48245 86636 -48115
rect 86690 -48245 86720 -48115
rect 86774 -48245 86804 -48115
rect 86858 -48245 86888 -48115
rect 87070 -48245 87100 -48115
rect 87154 -48245 87184 -48115
rect 87238 -48245 87268 -48115
rect 87322 -48245 87352 -48115
rect 87406 -48245 87436 -48115
rect 87490 -48245 87520 -48115
rect 87574 -48245 87604 -48115
rect 87658 -48245 87688 -48115
rect 87742 -48245 87772 -48115
rect 87826 -48245 87856 -48115
rect 87910 -48245 87940 -48115
rect 87994 -48245 88024 -48115
rect 88078 -48245 88108 -48115
rect 88162 -48245 88192 -48115
rect 88246 -48245 88276 -48115
rect 88330 -48245 88360 -48115
rect 88542 -48245 88572 -48115
rect 88626 -48245 88656 -48115
rect 88710 -48245 88740 -48115
rect 88794 -48245 88824 -48115
rect 88878 -48245 88908 -48115
rect 88962 -48245 88992 -48115
rect 89046 -48245 89076 -48115
rect 89130 -48245 89160 -48115
rect 89214 -48245 89244 -48115
rect 89298 -48245 89328 -48115
rect 89382 -48245 89412 -48115
rect 89466 -48245 89496 -48115
rect 89550 -48245 89580 -48115
rect 89634 -48245 89664 -48115
rect 89718 -48245 89748 -48115
rect 89802 -48245 89832 -48115
rect 90014 -48245 90044 -48115
rect 90098 -48245 90128 -48115
rect 90182 -48245 90212 -48115
rect 90266 -48245 90296 -48115
rect 90350 -48245 90380 -48115
rect 90434 -48245 90464 -48115
rect 90518 -48245 90548 -48115
rect 90602 -48245 90632 -48115
rect 90686 -48245 90716 -48115
rect 90770 -48245 90800 -48115
rect 90854 -48245 90884 -48115
rect 90938 -48245 90968 -48115
rect 91022 -48245 91052 -48115
rect 91106 -48245 91136 -48115
rect 91190 -48245 91220 -48115
rect 91274 -48245 91304 -48115
rect 77693 -48817 77723 -48733
rect 77777 -48817 77807 -48733
rect 77885 -48845 77915 -48715
rect 77693 -49127 77723 -49043
rect 77777 -49127 77807 -49043
rect 77885 -49145 77915 -49015
rect 78117 -49105 78147 -49021
rect 78213 -49105 78243 -49021
rect 78297 -49105 78327 -49021
rect 78381 -49105 78411 -49021
rect 78479 -49145 78509 -49015
rect 77693 -50057 77723 -49973
rect 77777 -50057 77807 -49973
rect 77885 -50085 77915 -49955
rect 77695 -50381 77725 -50297
rect 77779 -50381 77809 -50297
rect 77887 -50399 77917 -50269
rect 57175 -51159 57205 -51055
rect 57263 -51159 57293 -51055
rect 77657 -51335 77687 -51251
rect 77745 -51335 77775 -51251
rect 77851 -51335 77881 -51251
rect 77947 -51335 77977 -51251
rect 78113 -51335 78143 -51205
rect 78401 -51329 78431 -51245
rect 78497 -51329 78527 -51245
rect 78581 -51329 78611 -51245
rect 78665 -51329 78695 -51245
rect 78763 -51335 78793 -51205
rect 77657 -51585 77687 -51501
rect 77745 -51585 77775 -51501
rect 77851 -51585 77881 -51501
rect 77947 -51585 77977 -51501
rect 60191 -51647 60321 -51617
rect 61131 -51647 61261 -51617
rect 57175 -52333 57205 -52229
rect 57263 -52333 57293 -52229
rect 60191 -51731 60321 -51701
rect 61131 -51731 61261 -51701
rect 78113 -51631 78143 -51501
rect 60191 -51815 60321 -51785
rect 61131 -51815 61261 -51785
rect 60191 -51899 60321 -51869
rect 61131 -51899 61261 -51869
rect 82946 -51895 82976 -51811
rect 83030 -51895 83060 -51811
rect 83127 -51895 83157 -51765
rect 83418 -51895 83448 -51765
rect 83663 -51895 83693 -51765
rect 83747 -51895 83777 -51765
rect 83831 -51895 83861 -51765
rect 83915 -51895 83945 -51765
rect 84126 -51895 84156 -51765
rect 84210 -51895 84240 -51765
rect 84294 -51895 84324 -51765
rect 84378 -51895 84408 -51765
rect 84462 -51895 84492 -51765
rect 84546 -51895 84576 -51765
rect 84630 -51895 84660 -51765
rect 84714 -51895 84744 -51765
rect 84798 -51895 84828 -51765
rect 84882 -51895 84912 -51765
rect 84966 -51895 84996 -51765
rect 85050 -51895 85080 -51765
rect 85134 -51895 85164 -51765
rect 85218 -51895 85248 -51765
rect 85302 -51895 85332 -51765
rect 85386 -51895 85416 -51765
rect 85598 -51895 85628 -51765
rect 85682 -51895 85712 -51765
rect 85766 -51895 85796 -51765
rect 85850 -51895 85880 -51765
rect 85934 -51895 85964 -51765
rect 86018 -51895 86048 -51765
rect 86102 -51895 86132 -51765
rect 86186 -51895 86216 -51765
rect 86270 -51895 86300 -51765
rect 86354 -51895 86384 -51765
rect 86438 -51895 86468 -51765
rect 86522 -51895 86552 -51765
rect 86606 -51895 86636 -51765
rect 86690 -51895 86720 -51765
rect 86774 -51895 86804 -51765
rect 86858 -51895 86888 -51765
rect 87070 -51895 87100 -51765
rect 87154 -51895 87184 -51765
rect 87238 -51895 87268 -51765
rect 87322 -51895 87352 -51765
rect 87406 -51895 87436 -51765
rect 87490 -51895 87520 -51765
rect 87574 -51895 87604 -51765
rect 87658 -51895 87688 -51765
rect 87742 -51895 87772 -51765
rect 87826 -51895 87856 -51765
rect 87910 -51895 87940 -51765
rect 87994 -51895 88024 -51765
rect 88078 -51895 88108 -51765
rect 88162 -51895 88192 -51765
rect 88246 -51895 88276 -51765
rect 88330 -51895 88360 -51765
rect 88542 -51895 88572 -51765
rect 88626 -51895 88656 -51765
rect 88710 -51895 88740 -51765
rect 88794 -51895 88824 -51765
rect 88878 -51895 88908 -51765
rect 88962 -51895 88992 -51765
rect 89046 -51895 89076 -51765
rect 89130 -51895 89160 -51765
rect 89214 -51895 89244 -51765
rect 89298 -51895 89328 -51765
rect 89382 -51895 89412 -51765
rect 89466 -51895 89496 -51765
rect 89550 -51895 89580 -51765
rect 89634 -51895 89664 -51765
rect 89718 -51895 89748 -51765
rect 89802 -51895 89832 -51765
rect 90014 -51895 90044 -51765
rect 90098 -51895 90128 -51765
rect 90182 -51895 90212 -51765
rect 90266 -51895 90296 -51765
rect 90350 -51895 90380 -51765
rect 90434 -51895 90464 -51765
rect 90518 -51895 90548 -51765
rect 90602 -51895 90632 -51765
rect 90686 -51895 90716 -51765
rect 90770 -51895 90800 -51765
rect 90854 -51895 90884 -51765
rect 90938 -51895 90968 -51765
rect 91022 -51895 91052 -51765
rect 91106 -51895 91136 -51765
rect 91190 -51895 91220 -51765
rect 91274 -51895 91304 -51765
rect 77657 -52567 77687 -52483
rect 77745 -52567 77775 -52483
rect 77851 -52567 77881 -52483
rect 77947 -52567 77977 -52483
rect 78113 -52567 78143 -52437
rect 77657 -52819 77687 -52735
rect 77745 -52819 77775 -52735
rect 77851 -52819 77881 -52735
rect 77947 -52819 77977 -52735
rect 78113 -52865 78143 -52735
rect 77657 -53805 77687 -53721
rect 77729 -53805 77759 -53721
rect 77801 -53805 77831 -53721
rect 77929 -53805 77959 -53675
rect 78153 -53777 78183 -53693
rect 78237 -53777 78267 -53693
rect 78345 -53805 78375 -53675
rect 78577 -53799 78607 -53715
rect 78673 -53799 78703 -53715
rect 78757 -53799 78787 -53715
rect 78841 -53799 78871 -53715
rect 78939 -53805 78969 -53675
rect 57175 -56559 57205 -56455
rect 57263 -56559 57293 -56455
rect 60191 -57047 60321 -57017
rect 61131 -57047 61261 -57017
rect 57175 -57733 57205 -57629
rect 57263 -57733 57293 -57629
rect 60191 -57131 60321 -57101
rect 61131 -57131 61261 -57101
rect 60191 -57215 60321 -57185
rect 61131 -57215 61261 -57185
rect 60191 -57299 60321 -57269
rect 61131 -57299 61261 -57269
rect 57175 -61959 57205 -61855
rect 57263 -61959 57293 -61855
rect 60191 -62447 60321 -62417
rect 61131 -62447 61261 -62417
rect 57175 -63133 57205 -63029
rect 57263 -63133 57293 -63029
rect 60191 -62531 60321 -62501
rect 61131 -62531 61261 -62501
rect 60191 -62615 60321 -62585
rect 61131 -62615 61261 -62585
rect 60191 -62699 60321 -62669
rect 61131 -62699 61261 -62669
rect 57175 -67359 57205 -67255
rect 57263 -67359 57293 -67255
rect 60191 -67847 60321 -67817
rect 61131 -67847 61261 -67817
rect 57175 -68533 57205 -68429
rect 57263 -68533 57293 -68429
rect 60191 -67931 60321 -67901
rect 61131 -67931 61261 -67901
rect 60191 -68015 60321 -67985
rect 61131 -68015 61261 -67985
rect 60191 -68099 60321 -68069
rect 61131 -68099 61261 -68069
rect 57175 -72759 57205 -72655
rect 57263 -72759 57293 -72655
rect 60191 -73247 60321 -73217
rect 61131 -73247 61261 -73217
rect 57175 -73933 57205 -73829
rect 57263 -73933 57293 -73829
rect 60191 -73331 60321 -73301
rect 61131 -73331 61261 -73301
rect 60191 -73415 60321 -73385
rect 61131 -73415 61261 -73385
rect 60191 -73499 60321 -73469
rect 61131 -73499 61261 -73469
rect 57175 -78159 57205 -78055
rect 57263 -78159 57293 -78055
rect 60191 -78647 60321 -78617
rect 61131 -78647 61261 -78617
rect 57175 -79333 57205 -79229
rect 57263 -79333 57293 -79229
rect 60191 -78731 60321 -78701
rect 61131 -78731 61261 -78701
rect 60191 -78815 60321 -78785
rect 61131 -78815 61261 -78785
rect 60191 -78899 60321 -78869
rect 61131 -78899 61261 -78869
rect 57175 -83559 57205 -83455
rect 57263 -83559 57293 -83455
rect 60191 -84047 60321 -84017
rect 61131 -84047 61261 -84017
rect 57175 -84733 57205 -84629
rect 57263 -84733 57293 -84629
rect 60191 -84131 60321 -84101
rect 61131 -84131 61261 -84101
rect 60191 -84215 60321 -84185
rect 61131 -84215 61261 -84185
rect 60191 -84299 60321 -84269
rect 61131 -84299 61261 -84269
<< pmos >>
rect 59113 -2143 59513 -2093
rect 59113 -2251 59513 -2201
rect 59090 -2959 59150 -2559
rect 59090 -3689 59150 -3289
rect 59113 -4050 59513 -4000
rect 59113 -4158 59513 -4108
rect 59113 -7543 59513 -7493
rect 59113 -7651 59513 -7601
rect 59090 -8359 59150 -7959
rect 59090 -9089 59150 -8689
rect 59113 -9450 59513 -9400
rect 59113 -9558 59513 -9508
rect 59113 -12943 59513 -12893
rect 59113 -13051 59513 -13001
rect 59090 -13759 59150 -13359
rect 59090 -14489 59150 -14089
rect 59113 -14850 59513 -14800
rect 59113 -14958 59513 -14908
rect 59113 -18343 59513 -18293
rect 59113 -18451 59513 -18401
rect 59090 -19159 59150 -18759
rect 59090 -19889 59150 -19489
rect 59113 -20250 59513 -20200
rect 59113 -20358 59513 -20308
rect 59113 -23743 59513 -23693
rect 59113 -23851 59513 -23801
rect 59090 -24559 59150 -24159
rect 59090 -25289 59150 -24889
rect 59113 -25650 59513 -25600
rect 59113 -25758 59513 -25708
rect 59113 -29143 59513 -29093
rect 59113 -29251 59513 -29201
rect 59090 -29959 59150 -29559
rect 59090 -30689 59150 -30289
rect 59113 -31050 59513 -31000
rect 59113 -31158 59513 -31108
rect 59113 -34543 59513 -34493
rect 59113 -34651 59513 -34601
rect 59090 -35359 59150 -34959
rect 59090 -36089 59150 -35689
rect 59113 -36450 59513 -36400
rect 59113 -36558 59513 -36508
rect 59113 -39943 59513 -39893
rect 59113 -40051 59513 -40001
rect 59090 -40759 59150 -40359
rect 59090 -41489 59150 -41089
rect 59113 -41850 59513 -41800
rect 59113 -41958 59513 -41908
rect 59113 -45343 59513 -45293
rect 59113 -45451 59513 -45401
rect 59090 -46159 59150 -45759
rect 59090 -46889 59150 -46489
rect 59113 -47250 59513 -47200
rect 59113 -47358 59513 -47308
rect 59113 -50743 59513 -50693
rect 59113 -50851 59513 -50801
rect 59090 -51559 59150 -51159
rect 59090 -52289 59150 -51889
rect 59113 -52650 59513 -52600
rect 59113 -52758 59513 -52708
rect 59113 -56143 59513 -56093
rect 59113 -56251 59513 -56201
rect 59090 -56959 59150 -56559
rect 59090 -57689 59150 -57289
rect 59113 -58050 59513 -58000
rect 59113 -58158 59513 -58108
rect 59113 -61543 59513 -61493
rect 59113 -61651 59513 -61601
rect 59090 -62359 59150 -61959
rect 59090 -63089 59150 -62689
rect 59113 -63450 59513 -63400
rect 59113 -63558 59513 -63508
rect 59113 -66943 59513 -66893
rect 59113 -67051 59513 -67001
rect 59090 -67759 59150 -67359
rect 59090 -68489 59150 -68089
rect 59113 -68850 59513 -68800
rect 59113 -68958 59513 -68908
rect 59113 -72343 59513 -72293
rect 59113 -72451 59513 -72401
rect 59090 -73159 59150 -72759
rect 59090 -73889 59150 -73489
rect 59113 -74250 59513 -74200
rect 59113 -74358 59513 -74308
rect 59113 -77743 59513 -77693
rect 59113 -77851 59513 -77801
rect 59090 -78559 59150 -78159
rect 59090 -79289 59150 -78889
rect 59113 -79650 59513 -79600
rect 59113 -79758 59513 -79708
rect 59113 -83143 59513 -83093
rect 59113 -83251 59513 -83201
rect 59090 -83959 59150 -83559
rect 59090 -84689 59150 -84289
rect 59113 -85050 59513 -85000
rect 59113 -85158 59513 -85108
<< scpmoshvt >>
rect 57175 -2267 57205 -2109
rect 57263 -2267 57293 -2109
rect 60441 -3047 60641 -3017
rect 60811 -3047 61011 -3017
rect 60441 -3131 60641 -3101
rect 60811 -3131 61011 -3101
rect 60441 -3215 60641 -3185
rect 60811 -3215 61011 -3185
rect 60441 -3299 60641 -3269
rect 60811 -3299 61011 -3269
rect 57175 -4079 57205 -3921
rect 57263 -4079 57293 -3921
rect 57175 -7667 57205 -7509
rect 57263 -7667 57293 -7509
rect 60441 -8447 60641 -8417
rect 60811 -8447 61011 -8417
rect 60441 -8531 60641 -8501
rect 60811 -8531 61011 -8501
rect 60441 -8615 60641 -8585
rect 60811 -8615 61011 -8585
rect 60441 -8699 60641 -8669
rect 60811 -8699 61011 -8669
rect 57175 -9479 57205 -9321
rect 57263 -9479 57293 -9321
rect 57175 -13067 57205 -12909
rect 57263 -13067 57293 -12909
rect 60441 -13847 60641 -13817
rect 60811 -13847 61011 -13817
rect 60441 -13931 60641 -13901
rect 60811 -13931 61011 -13901
rect 60441 -14015 60641 -13985
rect 60811 -14015 61011 -13985
rect 60441 -14099 60641 -14069
rect 60811 -14099 61011 -14069
rect 57175 -14879 57205 -14721
rect 57263 -14879 57293 -14721
rect 57175 -18467 57205 -18309
rect 57263 -18467 57293 -18309
rect 60441 -19247 60641 -19217
rect 60811 -19247 61011 -19217
rect 60441 -19331 60641 -19301
rect 60811 -19331 61011 -19301
rect 60441 -19415 60641 -19385
rect 60811 -19415 61011 -19385
rect 60441 -19499 60641 -19469
rect 60811 -19499 61011 -19469
rect 57175 -20279 57205 -20121
rect 57263 -20279 57293 -20121
rect 57175 -23867 57205 -23709
rect 57263 -23867 57293 -23709
rect 60441 -24647 60641 -24617
rect 60811 -24647 61011 -24617
rect 60441 -24731 60641 -24701
rect 60811 -24731 61011 -24701
rect 60441 -24815 60641 -24785
rect 60811 -24815 61011 -24785
rect 60441 -24899 60641 -24869
rect 60811 -24899 61011 -24869
rect 57175 -25679 57205 -25521
rect 57263 -25679 57293 -25521
rect 57175 -29267 57205 -29109
rect 57263 -29267 57293 -29109
rect 60441 -30047 60641 -30017
rect 60811 -30047 61011 -30017
rect 60441 -30131 60641 -30101
rect 60811 -30131 61011 -30101
rect 60441 -30215 60641 -30185
rect 60811 -30215 61011 -30185
rect 60441 -30299 60641 -30269
rect 60811 -30299 61011 -30269
rect 57175 -31079 57205 -30921
rect 57263 -31079 57293 -30921
rect 57175 -34667 57205 -34509
rect 57263 -34667 57293 -34509
rect 60441 -35447 60641 -35417
rect 60811 -35447 61011 -35417
rect 60441 -35531 60641 -35501
rect 60811 -35531 61011 -35501
rect 60441 -35615 60641 -35585
rect 60811 -35615 61011 -35585
rect 60441 -35699 60641 -35669
rect 60811 -35699 61011 -35669
rect 57175 -36479 57205 -36321
rect 57263 -36479 57293 -36321
rect 75626 -38885 75656 -38685
rect 75902 -38885 75932 -38685
rect 76176 -38885 76206 -38685
rect 76452 -38885 76482 -38685
rect 76728 -38885 76758 -38685
rect 77657 -39305 77687 -39221
rect 77753 -39305 77783 -39221
rect 77825 -39305 77855 -39221
rect 77921 -39305 77951 -39221
rect 78019 -39305 78049 -39105
rect 78211 -39305 78241 -39221
rect 78283 -39305 78313 -39221
rect 78379 -39305 78409 -39221
rect 78477 -39305 78507 -39105
rect 78705 -39231 78735 -39147
rect 78789 -39231 78819 -39147
rect 78897 -39305 78927 -39105
rect 80858 -39355 80888 -39155
rect 81103 -39355 81133 -39155
rect 81187 -39355 81217 -39155
rect 81271 -39355 81301 -39155
rect 81355 -39355 81385 -39155
rect 81566 -39355 81596 -39155
rect 81650 -39355 81680 -39155
rect 81734 -39355 81764 -39155
rect 81818 -39355 81848 -39155
rect 81902 -39355 81932 -39155
rect 81986 -39355 82016 -39155
rect 82070 -39355 82100 -39155
rect 82154 -39355 82184 -39155
rect 82238 -39355 82268 -39155
rect 82322 -39355 82352 -39155
rect 82406 -39355 82436 -39155
rect 82490 -39355 82520 -39155
rect 82574 -39355 82604 -39155
rect 82658 -39355 82688 -39155
rect 82742 -39355 82772 -39155
rect 82826 -39355 82856 -39155
rect 83038 -39355 83068 -39155
rect 83122 -39355 83152 -39155
rect 83206 -39355 83236 -39155
rect 83290 -39355 83320 -39155
rect 83374 -39355 83404 -39155
rect 83458 -39355 83488 -39155
rect 83542 -39355 83572 -39155
rect 83626 -39355 83656 -39155
rect 83710 -39355 83740 -39155
rect 83794 -39355 83824 -39155
rect 83878 -39355 83908 -39155
rect 83962 -39355 83992 -39155
rect 84046 -39355 84076 -39155
rect 84130 -39355 84160 -39155
rect 84214 -39355 84244 -39155
rect 84298 -39355 84328 -39155
rect 84510 -39355 84540 -39155
rect 84594 -39355 84624 -39155
rect 84678 -39355 84708 -39155
rect 84762 -39355 84792 -39155
rect 84846 -39355 84876 -39155
rect 84930 -39355 84960 -39155
rect 85014 -39355 85044 -39155
rect 85098 -39355 85128 -39155
rect 85182 -39355 85212 -39155
rect 85266 -39355 85296 -39155
rect 85350 -39355 85380 -39155
rect 85434 -39355 85464 -39155
rect 85518 -39355 85548 -39155
rect 85602 -39355 85632 -39155
rect 85686 -39355 85716 -39155
rect 85770 -39355 85800 -39155
rect 85982 -39355 86012 -39155
rect 86066 -39355 86096 -39155
rect 86150 -39355 86180 -39155
rect 86234 -39355 86264 -39155
rect 86318 -39355 86348 -39155
rect 86402 -39355 86432 -39155
rect 86486 -39355 86516 -39155
rect 86570 -39355 86600 -39155
rect 86654 -39355 86684 -39155
rect 86738 -39355 86768 -39155
rect 86822 -39355 86852 -39155
rect 86906 -39355 86936 -39155
rect 86990 -39355 87020 -39155
rect 87074 -39355 87104 -39155
rect 87158 -39355 87188 -39155
rect 87242 -39355 87272 -39155
rect 87454 -39355 87484 -39155
rect 87538 -39355 87568 -39155
rect 87622 -39355 87652 -39155
rect 87706 -39355 87736 -39155
rect 87790 -39355 87820 -39155
rect 87874 -39355 87904 -39155
rect 87958 -39355 87988 -39155
rect 88042 -39355 88072 -39155
rect 88126 -39355 88156 -39155
rect 88210 -39355 88240 -39155
rect 88294 -39355 88324 -39155
rect 88378 -39355 88408 -39155
rect 88462 -39355 88492 -39155
rect 88546 -39355 88576 -39155
rect 88630 -39355 88660 -39155
rect 88714 -39355 88744 -39155
rect 57175 -40067 57205 -39909
rect 57263 -40067 57293 -39909
rect 77657 -40069 77687 -39985
rect 77753 -40069 77783 -39985
rect 77825 -40069 77855 -39985
rect 77921 -40069 77951 -39985
rect 78019 -40185 78049 -39985
rect 80908 -40225 80938 -40025
rect 77693 -40481 77723 -40397
rect 77777 -40481 77807 -40397
rect 77885 -40555 77915 -40355
rect 60441 -40847 60641 -40817
rect 60811 -40847 61011 -40817
rect 60441 -40931 60641 -40901
rect 60811 -40931 61011 -40901
rect 60441 -41015 60641 -40985
rect 60811 -41015 61011 -40985
rect 60441 -41099 60641 -41069
rect 60811 -41099 61011 -41069
rect 77693 -41383 77723 -41299
rect 77777 -41383 77807 -41299
rect 77885 -41425 77915 -41225
rect 78117 -41309 78147 -41225
rect 78213 -41309 78243 -41225
rect 78285 -41309 78315 -41225
rect 78381 -41309 78411 -41225
rect 78479 -41425 78509 -41225
rect 57175 -41879 57205 -41721
rect 57263 -41879 57293 -41721
rect 77693 -41721 77723 -41637
rect 77777 -41721 77807 -41637
rect 77885 -41795 77915 -41595
rect 77695 -42637 77725 -42553
rect 77779 -42637 77809 -42553
rect 77887 -42679 77917 -42479
rect 77657 -42929 77687 -42845
rect 77757 -42929 77787 -42845
rect 77861 -42929 77891 -42845
rect 77947 -42929 77977 -42845
rect 78113 -43045 78143 -42845
rect 78401 -43045 78431 -42961
rect 78497 -43045 78527 -42961
rect 78569 -43045 78599 -42961
rect 78665 -43045 78695 -42961
rect 78763 -43045 78793 -42845
rect 77657 -43911 77687 -43827
rect 77757 -43911 77787 -43827
rect 77861 -43911 77891 -43827
rect 77947 -43911 77977 -43827
rect 78113 -43911 78143 -43711
rect 82958 -43855 82988 -43771
rect 83030 -43855 83060 -43771
rect 83127 -43855 83157 -43655
rect 83418 -43855 83448 -43655
rect 83663 -43855 83693 -43655
rect 83747 -43855 83777 -43655
rect 83831 -43855 83861 -43655
rect 83915 -43855 83945 -43655
rect 84126 -43855 84156 -43655
rect 84210 -43855 84240 -43655
rect 84294 -43855 84324 -43655
rect 84378 -43855 84408 -43655
rect 84462 -43855 84492 -43655
rect 84546 -43855 84576 -43655
rect 84630 -43855 84660 -43655
rect 84714 -43855 84744 -43655
rect 84798 -43855 84828 -43655
rect 84882 -43855 84912 -43655
rect 84966 -43855 84996 -43655
rect 85050 -43855 85080 -43655
rect 85134 -43855 85164 -43655
rect 85218 -43855 85248 -43655
rect 85302 -43855 85332 -43655
rect 85386 -43855 85416 -43655
rect 85598 -43855 85628 -43655
rect 85682 -43855 85712 -43655
rect 85766 -43855 85796 -43655
rect 85850 -43855 85880 -43655
rect 85934 -43855 85964 -43655
rect 86018 -43855 86048 -43655
rect 86102 -43855 86132 -43655
rect 86186 -43855 86216 -43655
rect 86270 -43855 86300 -43655
rect 86354 -43855 86384 -43655
rect 86438 -43855 86468 -43655
rect 86522 -43855 86552 -43655
rect 86606 -43855 86636 -43655
rect 86690 -43855 86720 -43655
rect 86774 -43855 86804 -43655
rect 86858 -43855 86888 -43655
rect 87070 -43855 87100 -43655
rect 87154 -43855 87184 -43655
rect 87238 -43855 87268 -43655
rect 87322 -43855 87352 -43655
rect 87406 -43855 87436 -43655
rect 87490 -43855 87520 -43655
rect 87574 -43855 87604 -43655
rect 87658 -43855 87688 -43655
rect 87742 -43855 87772 -43655
rect 87826 -43855 87856 -43655
rect 87910 -43855 87940 -43655
rect 87994 -43855 88024 -43655
rect 88078 -43855 88108 -43655
rect 88162 -43855 88192 -43655
rect 88246 -43855 88276 -43655
rect 88330 -43855 88360 -43655
rect 88542 -43855 88572 -43655
rect 88626 -43855 88656 -43655
rect 88710 -43855 88740 -43655
rect 88794 -43855 88824 -43655
rect 88878 -43855 88908 -43655
rect 88962 -43855 88992 -43655
rect 89046 -43855 89076 -43655
rect 89130 -43855 89160 -43655
rect 89214 -43855 89244 -43655
rect 89298 -43855 89328 -43655
rect 89382 -43855 89412 -43655
rect 89466 -43855 89496 -43655
rect 89550 -43855 89580 -43655
rect 89634 -43855 89664 -43655
rect 89718 -43855 89748 -43655
rect 89802 -43855 89832 -43655
rect 90014 -43855 90044 -43655
rect 90098 -43855 90128 -43655
rect 90182 -43855 90212 -43655
rect 90266 -43855 90296 -43655
rect 90350 -43855 90380 -43655
rect 90434 -43855 90464 -43655
rect 90518 -43855 90548 -43655
rect 90602 -43855 90632 -43655
rect 90686 -43855 90716 -43655
rect 90770 -43855 90800 -43655
rect 90854 -43855 90884 -43655
rect 90938 -43855 90968 -43655
rect 91022 -43855 91052 -43655
rect 91106 -43855 91136 -43655
rect 91190 -43855 91220 -43655
rect 91274 -43855 91304 -43655
rect 77657 -44161 77687 -44077
rect 77757 -44161 77787 -44077
rect 77861 -44161 77891 -44077
rect 77947 -44161 77977 -44077
rect 78113 -44277 78143 -44077
rect 77657 -45145 77687 -45061
rect 77757 -45145 77787 -45061
rect 77861 -45145 77891 -45061
rect 77947 -45145 77977 -45061
rect 78113 -45145 78143 -44945
rect 57175 -45467 57205 -45309
rect 57263 -45467 57293 -45309
rect 77657 -45512 77687 -45428
rect 77741 -45512 77771 -45428
rect 77834 -45512 77864 -45428
rect 77929 -45515 77959 -45315
rect 78153 -45441 78183 -45357
rect 78237 -45441 78267 -45357
rect 78345 -45515 78375 -45315
rect 78577 -45515 78607 -45431
rect 78673 -45515 78703 -45431
rect 78745 -45515 78775 -45431
rect 78841 -45515 78871 -45431
rect 78939 -45515 78969 -45315
rect 60441 -46247 60641 -46217
rect 60811 -46247 61011 -46217
rect 60441 -46331 60641 -46301
rect 60811 -46331 61011 -46301
rect 60441 -46415 60641 -46385
rect 60811 -46415 61011 -46385
rect 60441 -46499 60641 -46469
rect 60811 -46499 61011 -46469
rect 57175 -47279 57205 -47121
rect 57263 -47279 57293 -47121
rect 75626 -46925 75656 -46725
rect 75902 -46925 75932 -46725
rect 76176 -46925 76206 -46725
rect 76452 -46925 76482 -46725
rect 76728 -46925 76758 -46725
rect 77657 -47345 77687 -47261
rect 77753 -47345 77783 -47261
rect 77825 -47345 77855 -47261
rect 77921 -47345 77951 -47261
rect 78019 -47345 78049 -47145
rect 78211 -47345 78241 -47261
rect 78283 -47345 78313 -47261
rect 78379 -47345 78409 -47261
rect 78477 -47345 78507 -47145
rect 78705 -47271 78735 -47187
rect 78789 -47271 78819 -47187
rect 78897 -47345 78927 -47145
rect 82958 -47995 82988 -47911
rect 83030 -47995 83060 -47911
rect 83127 -47995 83157 -47795
rect 83418 -47995 83448 -47795
rect 83663 -47995 83693 -47795
rect 83747 -47995 83777 -47795
rect 83831 -47995 83861 -47795
rect 83915 -47995 83945 -47795
rect 84126 -47995 84156 -47795
rect 84210 -47995 84240 -47795
rect 84294 -47995 84324 -47795
rect 84378 -47995 84408 -47795
rect 84462 -47995 84492 -47795
rect 84546 -47995 84576 -47795
rect 84630 -47995 84660 -47795
rect 84714 -47995 84744 -47795
rect 84798 -47995 84828 -47795
rect 84882 -47995 84912 -47795
rect 84966 -47995 84996 -47795
rect 85050 -47995 85080 -47795
rect 85134 -47995 85164 -47795
rect 85218 -47995 85248 -47795
rect 85302 -47995 85332 -47795
rect 85386 -47995 85416 -47795
rect 85598 -47995 85628 -47795
rect 85682 -47995 85712 -47795
rect 85766 -47995 85796 -47795
rect 85850 -47995 85880 -47795
rect 85934 -47995 85964 -47795
rect 86018 -47995 86048 -47795
rect 86102 -47995 86132 -47795
rect 86186 -47995 86216 -47795
rect 86270 -47995 86300 -47795
rect 86354 -47995 86384 -47795
rect 86438 -47995 86468 -47795
rect 86522 -47995 86552 -47795
rect 86606 -47995 86636 -47795
rect 86690 -47995 86720 -47795
rect 86774 -47995 86804 -47795
rect 86858 -47995 86888 -47795
rect 87070 -47995 87100 -47795
rect 87154 -47995 87184 -47795
rect 87238 -47995 87268 -47795
rect 87322 -47995 87352 -47795
rect 87406 -47995 87436 -47795
rect 87490 -47995 87520 -47795
rect 87574 -47995 87604 -47795
rect 87658 -47995 87688 -47795
rect 87742 -47995 87772 -47795
rect 87826 -47995 87856 -47795
rect 87910 -47995 87940 -47795
rect 87994 -47995 88024 -47795
rect 88078 -47995 88108 -47795
rect 88162 -47995 88192 -47795
rect 88246 -47995 88276 -47795
rect 88330 -47995 88360 -47795
rect 88542 -47995 88572 -47795
rect 88626 -47995 88656 -47795
rect 88710 -47995 88740 -47795
rect 88794 -47995 88824 -47795
rect 88878 -47995 88908 -47795
rect 88962 -47995 88992 -47795
rect 89046 -47995 89076 -47795
rect 89130 -47995 89160 -47795
rect 89214 -47995 89244 -47795
rect 89298 -47995 89328 -47795
rect 89382 -47995 89412 -47795
rect 89466 -47995 89496 -47795
rect 89550 -47995 89580 -47795
rect 89634 -47995 89664 -47795
rect 89718 -47995 89748 -47795
rect 89802 -47995 89832 -47795
rect 90014 -47995 90044 -47795
rect 90098 -47995 90128 -47795
rect 90182 -47995 90212 -47795
rect 90266 -47995 90296 -47795
rect 90350 -47995 90380 -47795
rect 90434 -47995 90464 -47795
rect 90518 -47995 90548 -47795
rect 90602 -47995 90632 -47795
rect 90686 -47995 90716 -47795
rect 90770 -47995 90800 -47795
rect 90854 -47995 90884 -47795
rect 90938 -47995 90968 -47795
rect 91022 -47995 91052 -47795
rect 91106 -47995 91136 -47795
rect 91190 -47995 91220 -47795
rect 91274 -47995 91304 -47795
rect 77657 -48109 77687 -48025
rect 77753 -48109 77783 -48025
rect 77825 -48109 77855 -48025
rect 77921 -48109 77951 -48025
rect 78019 -48225 78049 -48025
rect 77693 -48521 77723 -48437
rect 77777 -48521 77807 -48437
rect 77885 -48595 77915 -48395
rect 77693 -49423 77723 -49339
rect 77777 -49423 77807 -49339
rect 77885 -49465 77915 -49265
rect 78117 -49349 78147 -49265
rect 78213 -49349 78243 -49265
rect 78285 -49349 78315 -49265
rect 78381 -49349 78411 -49265
rect 78479 -49465 78509 -49265
rect 77693 -49761 77723 -49677
rect 77777 -49761 77807 -49677
rect 77885 -49835 77915 -49635
rect 57175 -50867 57205 -50709
rect 57263 -50867 57293 -50709
rect 77695 -50677 77725 -50593
rect 77779 -50677 77809 -50593
rect 77887 -50719 77917 -50519
rect 77657 -50969 77687 -50885
rect 77757 -50969 77787 -50885
rect 77861 -50969 77891 -50885
rect 77947 -50969 77977 -50885
rect 78113 -51085 78143 -50885
rect 78401 -51085 78431 -51001
rect 78497 -51085 78527 -51001
rect 78569 -51085 78599 -51001
rect 78665 -51085 78695 -51001
rect 78763 -51085 78793 -50885
rect 60441 -51647 60641 -51617
rect 60811 -51647 61011 -51617
rect 60441 -51731 60641 -51701
rect 60811 -51731 61011 -51701
rect 82958 -51645 82988 -51561
rect 83030 -51645 83060 -51561
rect 83127 -51645 83157 -51445
rect 83418 -51645 83448 -51445
rect 83663 -51645 83693 -51445
rect 83747 -51645 83777 -51445
rect 83831 -51645 83861 -51445
rect 83915 -51645 83945 -51445
rect 84126 -51645 84156 -51445
rect 84210 -51645 84240 -51445
rect 84294 -51645 84324 -51445
rect 84378 -51645 84408 -51445
rect 84462 -51645 84492 -51445
rect 84546 -51645 84576 -51445
rect 84630 -51645 84660 -51445
rect 84714 -51645 84744 -51445
rect 84798 -51645 84828 -51445
rect 84882 -51645 84912 -51445
rect 84966 -51645 84996 -51445
rect 85050 -51645 85080 -51445
rect 85134 -51645 85164 -51445
rect 85218 -51645 85248 -51445
rect 85302 -51645 85332 -51445
rect 85386 -51645 85416 -51445
rect 85598 -51645 85628 -51445
rect 85682 -51645 85712 -51445
rect 85766 -51645 85796 -51445
rect 85850 -51645 85880 -51445
rect 85934 -51645 85964 -51445
rect 86018 -51645 86048 -51445
rect 86102 -51645 86132 -51445
rect 86186 -51645 86216 -51445
rect 86270 -51645 86300 -51445
rect 86354 -51645 86384 -51445
rect 86438 -51645 86468 -51445
rect 86522 -51645 86552 -51445
rect 86606 -51645 86636 -51445
rect 86690 -51645 86720 -51445
rect 86774 -51645 86804 -51445
rect 86858 -51645 86888 -51445
rect 87070 -51645 87100 -51445
rect 87154 -51645 87184 -51445
rect 87238 -51645 87268 -51445
rect 87322 -51645 87352 -51445
rect 87406 -51645 87436 -51445
rect 87490 -51645 87520 -51445
rect 87574 -51645 87604 -51445
rect 87658 -51645 87688 -51445
rect 87742 -51645 87772 -51445
rect 87826 -51645 87856 -51445
rect 87910 -51645 87940 -51445
rect 87994 -51645 88024 -51445
rect 88078 -51645 88108 -51445
rect 88162 -51645 88192 -51445
rect 88246 -51645 88276 -51445
rect 88330 -51645 88360 -51445
rect 88542 -51645 88572 -51445
rect 88626 -51645 88656 -51445
rect 88710 -51645 88740 -51445
rect 88794 -51645 88824 -51445
rect 88878 -51645 88908 -51445
rect 88962 -51645 88992 -51445
rect 89046 -51645 89076 -51445
rect 89130 -51645 89160 -51445
rect 89214 -51645 89244 -51445
rect 89298 -51645 89328 -51445
rect 89382 -51645 89412 -51445
rect 89466 -51645 89496 -51445
rect 89550 -51645 89580 -51445
rect 89634 -51645 89664 -51445
rect 89718 -51645 89748 -51445
rect 89802 -51645 89832 -51445
rect 90014 -51645 90044 -51445
rect 90098 -51645 90128 -51445
rect 90182 -51645 90212 -51445
rect 90266 -51645 90296 -51445
rect 90350 -51645 90380 -51445
rect 90434 -51645 90464 -51445
rect 90518 -51645 90548 -51445
rect 90602 -51645 90632 -51445
rect 90686 -51645 90716 -51445
rect 90770 -51645 90800 -51445
rect 90854 -51645 90884 -51445
rect 90938 -51645 90968 -51445
rect 91022 -51645 91052 -51445
rect 91106 -51645 91136 -51445
rect 91190 -51645 91220 -51445
rect 91274 -51645 91304 -51445
rect 60441 -51815 60641 -51785
rect 60811 -51815 61011 -51785
rect 60441 -51899 60641 -51869
rect 60811 -51899 61011 -51869
rect 77657 -51951 77687 -51867
rect 77757 -51951 77787 -51867
rect 77861 -51951 77891 -51867
rect 77947 -51951 77977 -51867
rect 78113 -51951 78143 -51751
rect 77657 -52201 77687 -52117
rect 77757 -52201 77787 -52117
rect 77861 -52201 77891 -52117
rect 77947 -52201 77977 -52117
rect 57175 -52679 57205 -52521
rect 57263 -52679 57293 -52521
rect 78113 -52317 78143 -52117
rect 77657 -53185 77687 -53101
rect 77757 -53185 77787 -53101
rect 77861 -53185 77891 -53101
rect 77947 -53185 77977 -53101
rect 78113 -53185 78143 -52985
rect 77657 -53552 77687 -53468
rect 77741 -53552 77771 -53468
rect 77834 -53552 77864 -53468
rect 77929 -53555 77959 -53355
rect 78153 -53481 78183 -53397
rect 78237 -53481 78267 -53397
rect 78345 -53555 78375 -53355
rect 78577 -53555 78607 -53471
rect 78673 -53555 78703 -53471
rect 78745 -53555 78775 -53471
rect 78841 -53555 78871 -53471
rect 78939 -53555 78969 -53355
rect 57175 -56267 57205 -56109
rect 57263 -56267 57293 -56109
rect 60441 -57047 60641 -57017
rect 60811 -57047 61011 -57017
rect 60441 -57131 60641 -57101
rect 60811 -57131 61011 -57101
rect 60441 -57215 60641 -57185
rect 60811 -57215 61011 -57185
rect 60441 -57299 60641 -57269
rect 60811 -57299 61011 -57269
rect 57175 -58079 57205 -57921
rect 57263 -58079 57293 -57921
rect 57175 -61667 57205 -61509
rect 57263 -61667 57293 -61509
rect 60441 -62447 60641 -62417
rect 60811 -62447 61011 -62417
rect 60441 -62531 60641 -62501
rect 60811 -62531 61011 -62501
rect 60441 -62615 60641 -62585
rect 60811 -62615 61011 -62585
rect 60441 -62699 60641 -62669
rect 60811 -62699 61011 -62669
rect 57175 -63479 57205 -63321
rect 57263 -63479 57293 -63321
rect 57175 -67067 57205 -66909
rect 57263 -67067 57293 -66909
rect 60441 -67847 60641 -67817
rect 60811 -67847 61011 -67817
rect 60441 -67931 60641 -67901
rect 60811 -67931 61011 -67901
rect 60441 -68015 60641 -67985
rect 60811 -68015 61011 -67985
rect 60441 -68099 60641 -68069
rect 60811 -68099 61011 -68069
rect 57175 -68879 57205 -68721
rect 57263 -68879 57293 -68721
rect 57175 -72467 57205 -72309
rect 57263 -72467 57293 -72309
rect 60441 -73247 60641 -73217
rect 60811 -73247 61011 -73217
rect 60441 -73331 60641 -73301
rect 60811 -73331 61011 -73301
rect 60441 -73415 60641 -73385
rect 60811 -73415 61011 -73385
rect 60441 -73499 60641 -73469
rect 60811 -73499 61011 -73469
rect 57175 -74279 57205 -74121
rect 57263 -74279 57293 -74121
rect 57175 -77867 57205 -77709
rect 57263 -77867 57293 -77709
rect 60441 -78647 60641 -78617
rect 60811 -78647 61011 -78617
rect 60441 -78731 60641 -78701
rect 60811 -78731 61011 -78701
rect 60441 -78815 60641 -78785
rect 60811 -78815 61011 -78785
rect 60441 -78899 60641 -78869
rect 60811 -78899 61011 -78869
rect 57175 -79679 57205 -79521
rect 57263 -79679 57293 -79521
rect 57175 -83267 57205 -83109
rect 57263 -83267 57293 -83109
rect 60441 -84047 60641 -84017
rect 60811 -84047 61011 -84017
rect 60441 -84131 60641 -84101
rect 60811 -84131 61011 -84101
rect 60441 -84215 60641 -84185
rect 60811 -84215 61011 -84185
rect 60441 -84299 60641 -84269
rect 60811 -84299 61011 -84269
rect 57175 -85079 57205 -84921
rect 57263 -85079 57293 -84921
<< varactor >>
rect 55118 -2795 55518 -2759
rect 55118 -3417 55518 -3381
rect 55118 -8195 55518 -8159
rect 55118 -8817 55518 -8781
rect 55118 -13595 55518 -13559
rect 55118 -14217 55518 -14181
rect 55118 -18995 55518 -18959
rect 55118 -19617 55518 -19581
rect 55118 -24395 55518 -24359
rect 55118 -25017 55518 -24981
rect 55118 -29795 55518 -29759
rect 55118 -30417 55518 -30381
rect 55118 -35195 55518 -35159
rect 55118 -35817 55518 -35781
rect 55118 -40595 55518 -40559
rect 55118 -41217 55518 -41181
rect 55118 -45995 55518 -45959
rect 55118 -46617 55518 -46581
rect 55118 -51395 55518 -51359
rect 55118 -52017 55518 -51981
rect 55118 -56795 55518 -56759
rect 55118 -57417 55518 -57381
rect 55118 -62195 55518 -62159
rect 55118 -62817 55518 -62781
rect 55118 -67595 55518 -67559
rect 55118 -68217 55518 -68181
rect 55118 -72995 55518 -72959
rect 55118 -73617 55518 -73581
rect 55118 -78395 55518 -78359
rect 55118 -79017 55518 -78981
rect 55118 -83795 55518 -83759
rect 55118 -84417 55518 -84381
<< pmoslvt >>
rect 54079 -1788 54879 -1718
rect 54079 -2144 54879 -2074
rect 54069 -4104 54869 -4034
rect 56476 -3487 56546 -2687
rect 54069 -4460 54869 -4390
rect 54079 -7188 54879 -7118
rect 20892 -11656 21092 -7856
rect 21378 -11656 21578 -7856
rect 21864 -11656 22064 -7856
rect 54079 -7544 54879 -7474
rect 54069 -9504 54869 -9434
rect 56476 -8887 56546 -8087
rect 54069 -9860 54869 -9790
rect 54079 -12588 54879 -12518
rect 54079 -12944 54879 -12874
rect 54069 -14904 54869 -14834
rect 56476 -14287 56546 -13487
rect 54069 -15260 54869 -15190
rect 54079 -17988 54879 -17918
rect 54079 -18344 54879 -18274
rect 54069 -20304 54869 -20234
rect 56476 -19687 56546 -18887
rect 54069 -20660 54869 -20590
rect 54079 -23388 54879 -23318
rect 54079 -23744 54879 -23674
rect 54069 -25704 54869 -25634
rect 56476 -25087 56546 -24287
rect 54069 -26060 54869 -25990
rect 54079 -28788 54879 -28718
rect 54079 -29144 54879 -29074
rect 54069 -31104 54869 -31034
rect 56476 -30487 56546 -29687
rect 54069 -31460 54869 -31390
rect 54079 -34188 54879 -34118
rect 54079 -34544 54879 -34474
rect 54069 -36504 54869 -36434
rect 56476 -35887 56546 -35087
rect 54069 -36860 54869 -36790
rect 54079 -39588 54879 -39518
rect 54079 -39944 54879 -39874
rect 54069 -41904 54869 -41834
rect 56476 -41287 56546 -40487
rect 54069 -42260 54869 -42190
rect 54079 -44988 54879 -44918
rect 54079 -45344 54879 -45274
rect 54069 -47304 54869 -47234
rect 56476 -46687 56546 -45887
rect 54069 -47660 54869 -47590
rect 54079 -50388 54879 -50318
rect 54079 -50744 54879 -50674
rect 54069 -52704 54869 -52634
rect 56476 -52087 56546 -51287
rect 54069 -53060 54869 -52990
rect 54079 -55788 54879 -55718
rect 54079 -56144 54879 -56074
rect 54069 -58104 54869 -58034
rect 56476 -57487 56546 -56687
rect 54069 -58460 54869 -58390
rect 54079 -61188 54879 -61118
rect 54079 -61544 54879 -61474
rect 54069 -63504 54869 -63434
rect 56476 -62887 56546 -62087
rect 54069 -63860 54869 -63790
rect 54079 -66588 54879 -66518
rect 54079 -66944 54879 -66874
rect 54069 -68904 54869 -68834
rect 56476 -68287 56546 -67487
rect 54069 -69260 54869 -69190
rect 54079 -71988 54879 -71918
rect 54079 -72344 54879 -72274
rect 54069 -74304 54869 -74234
rect 56476 -73687 56546 -72887
rect 54069 -74660 54869 -74590
rect 54079 -77388 54879 -77318
rect 54079 -77744 54879 -77674
rect 54069 -79704 54869 -79634
rect 56476 -79087 56546 -78287
rect 54069 -80060 54869 -79990
rect 54079 -82788 54879 -82718
rect 54079 -83144 54879 -83074
rect 54069 -85104 54869 -85034
rect 56476 -84487 56546 -83687
rect 54069 -85460 54869 -85390
<< nmoslvt >>
rect 53510 -2978 53630 -2178
rect 55336 -2440 55366 -2240
rect 53930 -2944 54730 -2824
rect 55866 -2928 55986 -2128
rect 53510 -3996 53630 -3196
rect 53930 -3350 54730 -3230
rect 55326 -3936 55356 -3736
rect 55866 -4042 55986 -3242
rect 55288 -4634 55488 -4604
rect 53510 -8378 53630 -7578
rect 55336 -7840 55366 -7640
rect 53930 -8344 54730 -8224
rect 55866 -8328 55986 -7528
rect 53510 -9396 53630 -8596
rect 53930 -8750 54730 -8630
rect 55326 -9336 55356 -9136
rect 55866 -9442 55986 -8642
rect 55288 -10034 55488 -10004
rect 20268 -12006 20352 -11976
rect 16599 -13117 16719 -12317
rect 17005 -13117 17125 -12317
rect 17411 -13117 17531 -12317
rect 17817 -13117 17937 -12317
rect 18223 -13117 18343 -12317
rect 18629 -13117 18749 -12317
rect 19035 -13117 19155 -12317
rect 19441 -13117 19561 -12317
rect 19847 -13117 19967 -12317
rect 20253 -13117 20373 -12317
rect 20659 -13117 20779 -12317
rect 21065 -13117 21185 -12317
rect 21471 -13117 21591 -12317
rect 21877 -13117 21997 -12317
rect 22283 -13117 22403 -12317
rect 22689 -13117 22809 -12317
rect 23095 -13117 23215 -12317
rect 23501 -13117 23621 -12317
rect 23907 -13117 24027 -12317
rect 24313 -13117 24433 -12317
rect 24719 -13117 24839 -12317
rect 25125 -13117 25245 -12317
rect 53510 -13778 53630 -12978
rect 55336 -13240 55366 -13040
rect 53930 -13744 54730 -13624
rect 55866 -13728 55986 -12928
rect 53510 -14796 53630 -13996
rect 53930 -14150 54730 -14030
rect 55326 -14736 55356 -14536
rect 55866 -14842 55986 -14042
rect 55288 -15434 55488 -15404
rect 53510 -19178 53630 -18378
rect 55336 -18640 55366 -18440
rect 53930 -19144 54730 -19024
rect 55866 -19128 55986 -18328
rect 53510 -20196 53630 -19396
rect 53930 -19550 54730 -19430
rect 55326 -20136 55356 -19936
rect 55866 -20242 55986 -19442
rect 55288 -20834 55488 -20804
rect 53510 -24578 53630 -23778
rect 55336 -24040 55366 -23840
rect 53930 -24544 54730 -24424
rect 55866 -24528 55986 -23728
rect 53510 -25596 53630 -24796
rect 53930 -24950 54730 -24830
rect 55326 -25536 55356 -25336
rect 55866 -25642 55986 -24842
rect 55288 -26234 55488 -26204
rect 53510 -29978 53630 -29178
rect 55336 -29440 55366 -29240
rect 53930 -29944 54730 -29824
rect 55866 -29928 55986 -29128
rect 53510 -30996 53630 -30196
rect 53930 -30350 54730 -30230
rect 55326 -30936 55356 -30736
rect 55866 -31042 55986 -30242
rect 55288 -31634 55488 -31604
rect 53510 -35378 53630 -34578
rect 55336 -34840 55366 -34640
rect 53930 -35344 54730 -35224
rect 55866 -35328 55986 -34528
rect 53510 -36396 53630 -35596
rect 53930 -35750 54730 -35630
rect 55326 -36336 55356 -36136
rect 55866 -36442 55986 -35642
rect 55288 -37034 55488 -37004
rect 53510 -40778 53630 -39978
rect 55336 -40240 55366 -40040
rect 53930 -40744 54730 -40624
rect 55866 -40728 55986 -39928
rect 53510 -41796 53630 -40996
rect 53930 -41150 54730 -41030
rect 55326 -41736 55356 -41536
rect 55866 -41842 55986 -41042
rect 55288 -42434 55488 -42404
rect 53510 -46178 53630 -45378
rect 55336 -45640 55366 -45440
rect 53930 -46144 54730 -46024
rect 55866 -46128 55986 -45328
rect 53510 -47196 53630 -46396
rect 53930 -46550 54730 -46430
rect 55326 -47136 55356 -46936
rect 55866 -47242 55986 -46442
rect 55288 -47834 55488 -47804
rect 53510 -51578 53630 -50778
rect 55336 -51040 55366 -50840
rect 53930 -51544 54730 -51424
rect 55866 -51528 55986 -50728
rect 53510 -52596 53630 -51796
rect 53930 -51950 54730 -51830
rect 55326 -52536 55356 -52336
rect 55866 -52642 55986 -51842
rect 55288 -53234 55488 -53204
rect 53510 -56978 53630 -56178
rect 55336 -56440 55366 -56240
rect 53930 -56944 54730 -56824
rect 55866 -56928 55986 -56128
rect 53510 -57996 53630 -57196
rect 53930 -57350 54730 -57230
rect 55326 -57936 55356 -57736
rect 55866 -58042 55986 -57242
rect 55288 -58634 55488 -58604
rect 53510 -62378 53630 -61578
rect 55336 -61840 55366 -61640
rect 53930 -62344 54730 -62224
rect 55866 -62328 55986 -61528
rect 53510 -63396 53630 -62596
rect 53930 -62750 54730 -62630
rect 55326 -63336 55356 -63136
rect 55866 -63442 55986 -62642
rect 55288 -64034 55488 -64004
rect 53510 -67778 53630 -66978
rect 55336 -67240 55366 -67040
rect 53930 -67744 54730 -67624
rect 55866 -67728 55986 -66928
rect 53510 -68796 53630 -67996
rect 53930 -68150 54730 -68030
rect 55326 -68736 55356 -68536
rect 55866 -68842 55986 -68042
rect 55288 -69434 55488 -69404
rect 53510 -73178 53630 -72378
rect 55336 -72640 55366 -72440
rect 53930 -73144 54730 -73024
rect 55866 -73128 55986 -72328
rect 53510 -74196 53630 -73396
rect 53930 -73550 54730 -73430
rect 55326 -74136 55356 -73936
rect 55866 -74242 55986 -73442
rect 55288 -74834 55488 -74804
rect 53510 -78578 53630 -77778
rect 55336 -78040 55366 -77840
rect 53930 -78544 54730 -78424
rect 55866 -78528 55986 -77728
rect 53510 -79596 53630 -78796
rect 53930 -78950 54730 -78830
rect 55326 -79536 55356 -79336
rect 55866 -79642 55986 -78842
rect 55288 -80234 55488 -80204
rect 53510 -83978 53630 -83178
rect 55336 -83440 55366 -83240
rect 53930 -83944 54730 -83824
rect 55866 -83928 55986 -83128
rect 53510 -84996 53630 -84196
rect 53930 -84350 54730 -84230
rect 55326 -84936 55356 -84736
rect 55866 -85042 55986 -84242
rect 55288 -85634 55488 -85604
<< ndiff >>
rect 53452 -2190 53510 -2178
rect 53452 -2966 53464 -2190
rect 53498 -2966 53510 -2190
rect 53452 -2978 53510 -2966
rect 53630 -2190 53688 -2178
rect 53630 -2966 53642 -2190
rect 53676 -2966 53688 -2190
rect 53630 -2978 53688 -2966
rect 55278 -2252 55336 -2240
rect 55278 -2428 55290 -2252
rect 55324 -2428 55336 -2252
rect 55278 -2440 55336 -2428
rect 55366 -2252 55424 -2240
rect 55366 -2428 55378 -2252
rect 55412 -2428 55424 -2252
rect 55366 -2440 55424 -2428
rect 53930 -2778 54730 -2766
rect 53930 -2812 53942 -2778
rect 54718 -2812 54730 -2778
rect 53930 -2824 54730 -2812
rect 53930 -2956 54730 -2944
rect 53930 -2990 53942 -2956
rect 54718 -2990 54730 -2956
rect 53930 -3002 54730 -2990
rect 55808 -2140 55866 -2128
rect 55808 -2916 55820 -2140
rect 55854 -2916 55866 -2140
rect 55808 -2928 55866 -2916
rect 55986 -2140 56044 -2128
rect 55986 -2916 55998 -2140
rect 56032 -2916 56044 -2140
rect 55986 -2928 56044 -2916
rect 57123 -2500 57175 -2455
rect 53452 -3208 53510 -3196
rect 53452 -3984 53464 -3208
rect 53498 -3984 53510 -3208
rect 53452 -3996 53510 -3984
rect 53630 -3208 53688 -3196
rect 53630 -3984 53642 -3208
rect 53676 -3984 53688 -3208
rect 53630 -3996 53688 -3984
rect 53930 -3184 54730 -3172
rect 53930 -3218 53942 -3184
rect 54718 -3218 54730 -3184
rect 53930 -3230 54730 -3218
rect 53930 -3362 54730 -3350
rect 53930 -3396 53942 -3362
rect 54718 -3396 54730 -3362
rect 53930 -3408 54730 -3396
rect 55268 -3748 55326 -3736
rect 55268 -3924 55280 -3748
rect 55314 -3924 55326 -3748
rect 55268 -3936 55326 -3924
rect 55356 -3748 55414 -3736
rect 55356 -3924 55368 -3748
rect 55402 -3924 55414 -3748
rect 55356 -3936 55414 -3924
rect 55808 -3254 55866 -3242
rect 55808 -4030 55820 -3254
rect 55854 -4030 55866 -3254
rect 55808 -4042 55866 -4030
rect 55986 -3254 56044 -3242
rect 55986 -4030 55998 -3254
rect 56032 -4030 56044 -3254
rect 55986 -4042 56044 -4030
rect 57123 -2534 57131 -2500
rect 57165 -2534 57175 -2500
rect 57123 -2559 57175 -2534
rect 57205 -2513 57263 -2455
rect 57205 -2547 57217 -2513
rect 57251 -2547 57263 -2513
rect 57205 -2559 57263 -2547
rect 57293 -2483 57345 -2455
rect 57293 -2517 57303 -2483
rect 57337 -2517 57345 -2483
rect 57293 -2559 57345 -2517
rect 59946 -2374 60346 -2362
rect 59946 -2408 59958 -2374
rect 60334 -2408 60346 -2374
rect 59946 -2420 60346 -2408
rect 59946 -2482 60346 -2470
rect 59946 -2516 59958 -2482
rect 60334 -2516 60346 -2482
rect 59946 -2528 60346 -2516
rect 59490 -2782 59548 -2770
rect 59490 -2850 59502 -2782
rect 59476 -2920 59502 -2850
rect 59490 -2958 59502 -2920
rect 59536 -2958 59548 -2782
rect 59490 -2970 59548 -2958
rect 59578 -2782 59636 -2770
rect 59578 -2958 59590 -2782
rect 59624 -2958 59636 -2782
rect 59578 -2970 59636 -2958
rect 59806 -2782 59864 -2770
rect 59806 -2958 59818 -2782
rect 59852 -2958 59864 -2782
rect 59806 -2970 59864 -2958
rect 59894 -2782 59952 -2770
rect 59894 -2958 59906 -2782
rect 59940 -2958 59952 -2782
rect 59894 -2970 59952 -2958
rect 60191 -2973 60321 -2965
rect 60191 -3007 60203 -2973
rect 60237 -3007 60321 -2973
rect 60191 -3017 60321 -3007
rect 61131 -2973 61261 -2965
rect 61131 -3007 61215 -2973
rect 61249 -3007 61261 -2973
rect 61131 -3017 61261 -3007
rect 60191 -3057 60321 -3047
rect 60191 -3091 60211 -3057
rect 60245 -3091 60321 -3057
rect 60191 -3101 60321 -3091
rect 61131 -3057 61261 -3047
rect 61131 -3091 61207 -3057
rect 61241 -3091 61261 -3057
rect 61131 -3101 61261 -3091
rect 57123 -3654 57175 -3629
rect 57123 -3688 57131 -3654
rect 57165 -3688 57175 -3654
rect 57123 -3733 57175 -3688
rect 57205 -3641 57263 -3629
rect 57205 -3675 57217 -3641
rect 57251 -3675 57263 -3641
rect 57205 -3733 57263 -3675
rect 57293 -3671 57345 -3629
rect 57293 -3705 57303 -3671
rect 57337 -3705 57345 -3671
rect 57293 -3733 57345 -3705
rect 60191 -3141 60321 -3131
rect 59489 -3295 59547 -3283
rect 59489 -3471 59501 -3295
rect 59535 -3471 59547 -3295
rect 59489 -3483 59547 -3471
rect 59577 -3295 59635 -3283
rect 59577 -3471 59589 -3295
rect 59623 -3471 59635 -3295
rect 59577 -3483 59635 -3471
rect 60191 -3175 60203 -3141
rect 60237 -3175 60321 -3141
rect 60191 -3185 60321 -3175
rect 61131 -3141 61261 -3131
rect 61131 -3175 61215 -3141
rect 61249 -3175 61261 -3141
rect 61131 -3185 61261 -3175
rect 59805 -3295 59863 -3283
rect 59805 -3471 59817 -3295
rect 59851 -3471 59863 -3295
rect 59805 -3483 59863 -3471
rect 59893 -3295 59951 -3283
rect 59893 -3471 59905 -3295
rect 59939 -3471 59951 -3295
rect 59893 -3483 59951 -3471
rect 60191 -3225 60321 -3215
rect 60191 -3259 60211 -3225
rect 60245 -3259 60321 -3225
rect 60191 -3269 60321 -3259
rect 61131 -3225 61261 -3215
rect 61131 -3259 61207 -3225
rect 61241 -3259 61261 -3225
rect 61131 -3269 61261 -3259
rect 60191 -3309 60321 -3299
rect 60191 -3343 60204 -3309
rect 60238 -3343 60321 -3309
rect 60191 -3351 60321 -3343
rect 61131 -3309 61261 -3299
rect 61131 -3343 61214 -3309
rect 61248 -3343 61261 -3309
rect 61131 -3351 61261 -3343
rect 59946 -3740 60346 -3728
rect 59946 -3774 59958 -3740
rect 60334 -3774 60346 -3740
rect 59946 -3786 60346 -3774
rect 59946 -3848 60346 -3836
rect 59946 -3882 59958 -3848
rect 60334 -3882 60346 -3848
rect 59946 -3894 60346 -3882
rect 55288 -4558 55488 -4546
rect 55288 -4592 55300 -4558
rect 55476 -4592 55488 -4558
rect 55288 -4604 55488 -4592
rect 55288 -4646 55488 -4634
rect 55288 -4680 55300 -4646
rect 55476 -4680 55488 -4646
rect 55288 -4692 55488 -4680
rect 53452 -7590 53510 -7578
rect 53452 -8366 53464 -7590
rect 53498 -8366 53510 -7590
rect 53452 -8378 53510 -8366
rect 53630 -7590 53688 -7578
rect 53630 -8366 53642 -7590
rect 53676 -8366 53688 -7590
rect 53630 -8378 53688 -8366
rect 55278 -7652 55336 -7640
rect 55278 -7828 55290 -7652
rect 55324 -7828 55336 -7652
rect 55278 -7840 55336 -7828
rect 55366 -7652 55424 -7640
rect 55366 -7828 55378 -7652
rect 55412 -7828 55424 -7652
rect 55366 -7840 55424 -7828
rect 53930 -8178 54730 -8166
rect 53930 -8212 53942 -8178
rect 54718 -8212 54730 -8178
rect 53930 -8224 54730 -8212
rect 53930 -8356 54730 -8344
rect 53930 -8390 53942 -8356
rect 54718 -8390 54730 -8356
rect 53930 -8402 54730 -8390
rect 55808 -7540 55866 -7528
rect 55808 -8316 55820 -7540
rect 55854 -8316 55866 -7540
rect 55808 -8328 55866 -8316
rect 55986 -7540 56044 -7528
rect 55986 -8316 55998 -7540
rect 56032 -8316 56044 -7540
rect 55986 -8328 56044 -8316
rect 57123 -7900 57175 -7855
rect 53452 -8608 53510 -8596
rect 53452 -9384 53464 -8608
rect 53498 -9384 53510 -8608
rect 53452 -9396 53510 -9384
rect 53630 -8608 53688 -8596
rect 53630 -9384 53642 -8608
rect 53676 -9384 53688 -8608
rect 53630 -9396 53688 -9384
rect 53930 -8584 54730 -8572
rect 53930 -8618 53942 -8584
rect 54718 -8618 54730 -8584
rect 53930 -8630 54730 -8618
rect 53930 -8762 54730 -8750
rect 53930 -8796 53942 -8762
rect 54718 -8796 54730 -8762
rect 53930 -8808 54730 -8796
rect 55268 -9148 55326 -9136
rect 55268 -9324 55280 -9148
rect 55314 -9324 55326 -9148
rect 55268 -9336 55326 -9324
rect 55356 -9148 55414 -9136
rect 55356 -9324 55368 -9148
rect 55402 -9324 55414 -9148
rect 55356 -9336 55414 -9324
rect 55808 -8654 55866 -8642
rect 55808 -9430 55820 -8654
rect 55854 -9430 55866 -8654
rect 55808 -9442 55866 -9430
rect 55986 -8654 56044 -8642
rect 55986 -9430 55998 -8654
rect 56032 -9430 56044 -8654
rect 55986 -9442 56044 -9430
rect 57123 -7934 57131 -7900
rect 57165 -7934 57175 -7900
rect 57123 -7959 57175 -7934
rect 57205 -7913 57263 -7855
rect 57205 -7947 57217 -7913
rect 57251 -7947 57263 -7913
rect 57205 -7959 57263 -7947
rect 57293 -7883 57345 -7855
rect 57293 -7917 57303 -7883
rect 57337 -7917 57345 -7883
rect 57293 -7959 57345 -7917
rect 59946 -7774 60346 -7762
rect 59946 -7808 59958 -7774
rect 60334 -7808 60346 -7774
rect 59946 -7820 60346 -7808
rect 59946 -7882 60346 -7870
rect 59946 -7916 59958 -7882
rect 60334 -7916 60346 -7882
rect 59946 -7928 60346 -7916
rect 59490 -8182 59548 -8170
rect 59490 -8250 59502 -8182
rect 59476 -8320 59502 -8250
rect 59490 -8358 59502 -8320
rect 59536 -8358 59548 -8182
rect 59490 -8370 59548 -8358
rect 59578 -8182 59636 -8170
rect 59578 -8358 59590 -8182
rect 59624 -8358 59636 -8182
rect 59578 -8370 59636 -8358
rect 59806 -8182 59864 -8170
rect 59806 -8358 59818 -8182
rect 59852 -8358 59864 -8182
rect 59806 -8370 59864 -8358
rect 59894 -8182 59952 -8170
rect 59894 -8358 59906 -8182
rect 59940 -8358 59952 -8182
rect 59894 -8370 59952 -8358
rect 60191 -8373 60321 -8365
rect 60191 -8407 60203 -8373
rect 60237 -8407 60321 -8373
rect 60191 -8417 60321 -8407
rect 61131 -8373 61261 -8365
rect 61131 -8407 61215 -8373
rect 61249 -8407 61261 -8373
rect 61131 -8417 61261 -8407
rect 60191 -8457 60321 -8447
rect 60191 -8491 60211 -8457
rect 60245 -8491 60321 -8457
rect 60191 -8501 60321 -8491
rect 61131 -8457 61261 -8447
rect 61131 -8491 61207 -8457
rect 61241 -8491 61261 -8457
rect 61131 -8501 61261 -8491
rect 57123 -9054 57175 -9029
rect 57123 -9088 57131 -9054
rect 57165 -9088 57175 -9054
rect 57123 -9133 57175 -9088
rect 57205 -9041 57263 -9029
rect 57205 -9075 57217 -9041
rect 57251 -9075 57263 -9041
rect 57205 -9133 57263 -9075
rect 57293 -9071 57345 -9029
rect 57293 -9105 57303 -9071
rect 57337 -9105 57345 -9071
rect 57293 -9133 57345 -9105
rect 60191 -8541 60321 -8531
rect 59489 -8695 59547 -8683
rect 59489 -8871 59501 -8695
rect 59535 -8871 59547 -8695
rect 59489 -8883 59547 -8871
rect 59577 -8695 59635 -8683
rect 59577 -8871 59589 -8695
rect 59623 -8871 59635 -8695
rect 59577 -8883 59635 -8871
rect 60191 -8575 60203 -8541
rect 60237 -8575 60321 -8541
rect 60191 -8585 60321 -8575
rect 61131 -8541 61261 -8531
rect 61131 -8575 61215 -8541
rect 61249 -8575 61261 -8541
rect 61131 -8585 61261 -8575
rect 59805 -8695 59863 -8683
rect 59805 -8871 59817 -8695
rect 59851 -8871 59863 -8695
rect 59805 -8883 59863 -8871
rect 59893 -8695 59951 -8683
rect 59893 -8871 59905 -8695
rect 59939 -8871 59951 -8695
rect 59893 -8883 59951 -8871
rect 60191 -8625 60321 -8615
rect 60191 -8659 60211 -8625
rect 60245 -8659 60321 -8625
rect 60191 -8669 60321 -8659
rect 61131 -8625 61261 -8615
rect 61131 -8659 61207 -8625
rect 61241 -8659 61261 -8625
rect 61131 -8669 61261 -8659
rect 60191 -8709 60321 -8699
rect 60191 -8743 60204 -8709
rect 60238 -8743 60321 -8709
rect 60191 -8751 60321 -8743
rect 61131 -8709 61261 -8699
rect 61131 -8743 61214 -8709
rect 61248 -8743 61261 -8709
rect 61131 -8751 61261 -8743
rect 59946 -9140 60346 -9128
rect 59946 -9174 59958 -9140
rect 60334 -9174 60346 -9140
rect 59946 -9186 60346 -9174
rect 59946 -9248 60346 -9236
rect 59946 -9282 59958 -9248
rect 60334 -9282 60346 -9248
rect 59946 -9294 60346 -9282
rect 55288 -9958 55488 -9946
rect 55288 -9992 55300 -9958
rect 55476 -9992 55488 -9958
rect 55288 -10004 55488 -9992
rect 55288 -10046 55488 -10034
rect 55288 -10080 55300 -10046
rect 55476 -10080 55488 -10046
rect 55288 -10092 55488 -10080
rect 20268 -11930 20352 -11918
rect 20268 -11964 20280 -11930
rect 20340 -11964 20352 -11930
rect 20268 -11976 20352 -11964
rect 20268 -12018 20352 -12006
rect 20268 -12052 20280 -12018
rect 20340 -12052 20352 -12018
rect 20268 -12064 20352 -12052
rect 16541 -12329 16599 -12317
rect 16541 -13105 16553 -12329
rect 16587 -13105 16599 -12329
rect 16541 -13117 16599 -13105
rect 16719 -12329 16777 -12317
rect 16719 -13105 16731 -12329
rect 16765 -13105 16777 -12329
rect 16719 -13117 16777 -13105
rect 16947 -12329 17005 -12317
rect 16947 -13105 16959 -12329
rect 16993 -13105 17005 -12329
rect 16947 -13117 17005 -13105
rect 17125 -12329 17183 -12317
rect 17125 -13105 17137 -12329
rect 17171 -13105 17183 -12329
rect 17125 -13117 17183 -13105
rect 17353 -12329 17411 -12317
rect 17353 -13105 17365 -12329
rect 17399 -13105 17411 -12329
rect 17353 -13117 17411 -13105
rect 17531 -12329 17589 -12317
rect 17531 -13105 17543 -12329
rect 17577 -13105 17589 -12329
rect 17531 -13117 17589 -13105
rect 17759 -12329 17817 -12317
rect 17759 -13105 17771 -12329
rect 17805 -13105 17817 -12329
rect 17759 -13117 17817 -13105
rect 17937 -12329 17995 -12317
rect 17937 -13105 17949 -12329
rect 17983 -13105 17995 -12329
rect 17937 -13117 17995 -13105
rect 18165 -12329 18223 -12317
rect 18165 -13105 18177 -12329
rect 18211 -13105 18223 -12329
rect 18165 -13117 18223 -13105
rect 18343 -12329 18401 -12317
rect 18343 -13105 18355 -12329
rect 18389 -13105 18401 -12329
rect 18343 -13117 18401 -13105
rect 18571 -12329 18629 -12317
rect 18571 -13105 18583 -12329
rect 18617 -13105 18629 -12329
rect 18571 -13117 18629 -13105
rect 18749 -12329 18807 -12317
rect 18749 -13105 18761 -12329
rect 18795 -13105 18807 -12329
rect 18749 -13117 18807 -13105
rect 18977 -12329 19035 -12317
rect 18977 -13105 18989 -12329
rect 19023 -13105 19035 -12329
rect 18977 -13117 19035 -13105
rect 19155 -12329 19213 -12317
rect 19155 -13105 19167 -12329
rect 19201 -13105 19213 -12329
rect 19155 -13117 19213 -13105
rect 19383 -12329 19441 -12317
rect 19383 -13105 19395 -12329
rect 19429 -13105 19441 -12329
rect 19383 -13117 19441 -13105
rect 19561 -12329 19619 -12317
rect 19561 -13105 19573 -12329
rect 19607 -13105 19619 -12329
rect 19561 -13117 19619 -13105
rect 19789 -12329 19847 -12317
rect 19789 -13105 19801 -12329
rect 19835 -13105 19847 -12329
rect 19789 -13117 19847 -13105
rect 19967 -12329 20025 -12317
rect 19967 -13105 19979 -12329
rect 20013 -13105 20025 -12329
rect 19967 -13117 20025 -13105
rect 20195 -12329 20253 -12317
rect 20195 -13105 20207 -12329
rect 20241 -13105 20253 -12329
rect 20195 -13117 20253 -13105
rect 20373 -12329 20431 -12317
rect 20373 -13105 20385 -12329
rect 20419 -13105 20431 -12329
rect 20373 -13117 20431 -13105
rect 20601 -12329 20659 -12317
rect 20601 -13105 20613 -12329
rect 20647 -13105 20659 -12329
rect 20601 -13117 20659 -13105
rect 20779 -12329 20837 -12317
rect 20779 -13105 20791 -12329
rect 20825 -13105 20837 -12329
rect 20779 -13117 20837 -13105
rect 21007 -12329 21065 -12317
rect 21007 -13105 21019 -12329
rect 21053 -13105 21065 -12329
rect 21007 -13117 21065 -13105
rect 21185 -12329 21243 -12317
rect 21185 -13105 21197 -12329
rect 21231 -13105 21243 -12329
rect 21185 -13117 21243 -13105
rect 21413 -12329 21471 -12317
rect 21413 -13105 21425 -12329
rect 21459 -13105 21471 -12329
rect 21413 -13117 21471 -13105
rect 21591 -12329 21649 -12317
rect 21591 -13105 21603 -12329
rect 21637 -13105 21649 -12329
rect 21591 -13117 21649 -13105
rect 21819 -12329 21877 -12317
rect 21819 -13105 21831 -12329
rect 21865 -13105 21877 -12329
rect 21819 -13117 21877 -13105
rect 21997 -12329 22055 -12317
rect 21997 -13105 22009 -12329
rect 22043 -13105 22055 -12329
rect 21997 -13117 22055 -13105
rect 22225 -12329 22283 -12317
rect 22225 -13105 22237 -12329
rect 22271 -13105 22283 -12329
rect 22225 -13117 22283 -13105
rect 22403 -12329 22461 -12317
rect 22403 -13105 22415 -12329
rect 22449 -13105 22461 -12329
rect 22403 -13117 22461 -13105
rect 22631 -12329 22689 -12317
rect 22631 -13105 22643 -12329
rect 22677 -13105 22689 -12329
rect 22631 -13117 22689 -13105
rect 22809 -12329 22867 -12317
rect 22809 -13105 22821 -12329
rect 22855 -13105 22867 -12329
rect 22809 -13117 22867 -13105
rect 23037 -12329 23095 -12317
rect 23037 -13105 23049 -12329
rect 23083 -13105 23095 -12329
rect 23037 -13117 23095 -13105
rect 23215 -12329 23273 -12317
rect 23215 -13105 23227 -12329
rect 23261 -13105 23273 -12329
rect 23215 -13117 23273 -13105
rect 23443 -12329 23501 -12317
rect 23443 -13105 23455 -12329
rect 23489 -13105 23501 -12329
rect 23443 -13117 23501 -13105
rect 23621 -12329 23679 -12317
rect 23621 -13105 23633 -12329
rect 23667 -13105 23679 -12329
rect 23621 -13117 23679 -13105
rect 23849 -12329 23907 -12317
rect 23849 -13105 23861 -12329
rect 23895 -13105 23907 -12329
rect 23849 -13117 23907 -13105
rect 24027 -12329 24085 -12317
rect 24027 -13105 24039 -12329
rect 24073 -13105 24085 -12329
rect 24027 -13117 24085 -13105
rect 24255 -12329 24313 -12317
rect 24255 -13105 24267 -12329
rect 24301 -13105 24313 -12329
rect 24255 -13117 24313 -13105
rect 24433 -12329 24491 -12317
rect 24433 -13105 24445 -12329
rect 24479 -13105 24491 -12329
rect 24433 -13117 24491 -13105
rect 24661 -12329 24719 -12317
rect 24661 -13105 24673 -12329
rect 24707 -13105 24719 -12329
rect 24661 -13117 24719 -13105
rect 24839 -12329 24897 -12317
rect 24839 -13105 24851 -12329
rect 24885 -13105 24897 -12329
rect 24839 -13117 24897 -13105
rect 25067 -12329 25125 -12317
rect 25067 -13105 25079 -12329
rect 25113 -13105 25125 -12329
rect 25067 -13117 25125 -13105
rect 25245 -12329 25303 -12317
rect 25245 -13105 25257 -12329
rect 25291 -13105 25303 -12329
rect 25245 -13117 25303 -13105
rect 53452 -12990 53510 -12978
rect 53452 -13766 53464 -12990
rect 53498 -13766 53510 -12990
rect 53452 -13778 53510 -13766
rect 53630 -12990 53688 -12978
rect 53630 -13766 53642 -12990
rect 53676 -13766 53688 -12990
rect 53630 -13778 53688 -13766
rect 55278 -13052 55336 -13040
rect 55278 -13228 55290 -13052
rect 55324 -13228 55336 -13052
rect 55278 -13240 55336 -13228
rect 55366 -13052 55424 -13040
rect 55366 -13228 55378 -13052
rect 55412 -13228 55424 -13052
rect 55366 -13240 55424 -13228
rect 53930 -13578 54730 -13566
rect 53930 -13612 53942 -13578
rect 54718 -13612 54730 -13578
rect 53930 -13624 54730 -13612
rect 53930 -13756 54730 -13744
rect 53930 -13790 53942 -13756
rect 54718 -13790 54730 -13756
rect 53930 -13802 54730 -13790
rect 55808 -12940 55866 -12928
rect 55808 -13716 55820 -12940
rect 55854 -13716 55866 -12940
rect 55808 -13728 55866 -13716
rect 55986 -12940 56044 -12928
rect 55986 -13716 55998 -12940
rect 56032 -13716 56044 -12940
rect 55986 -13728 56044 -13716
rect 57123 -13300 57175 -13255
rect 53452 -14008 53510 -13996
rect 53452 -14784 53464 -14008
rect 53498 -14784 53510 -14008
rect 53452 -14796 53510 -14784
rect 53630 -14008 53688 -13996
rect 53630 -14784 53642 -14008
rect 53676 -14784 53688 -14008
rect 53630 -14796 53688 -14784
rect 53930 -13984 54730 -13972
rect 53930 -14018 53942 -13984
rect 54718 -14018 54730 -13984
rect 53930 -14030 54730 -14018
rect 53930 -14162 54730 -14150
rect 53930 -14196 53942 -14162
rect 54718 -14196 54730 -14162
rect 53930 -14208 54730 -14196
rect 55268 -14548 55326 -14536
rect 55268 -14724 55280 -14548
rect 55314 -14724 55326 -14548
rect 55268 -14736 55326 -14724
rect 55356 -14548 55414 -14536
rect 55356 -14724 55368 -14548
rect 55402 -14724 55414 -14548
rect 55356 -14736 55414 -14724
rect 55808 -14054 55866 -14042
rect 55808 -14830 55820 -14054
rect 55854 -14830 55866 -14054
rect 55808 -14842 55866 -14830
rect 55986 -14054 56044 -14042
rect 55986 -14830 55998 -14054
rect 56032 -14830 56044 -14054
rect 55986 -14842 56044 -14830
rect 57123 -13334 57131 -13300
rect 57165 -13334 57175 -13300
rect 57123 -13359 57175 -13334
rect 57205 -13313 57263 -13255
rect 57205 -13347 57217 -13313
rect 57251 -13347 57263 -13313
rect 57205 -13359 57263 -13347
rect 57293 -13283 57345 -13255
rect 57293 -13317 57303 -13283
rect 57337 -13317 57345 -13283
rect 57293 -13359 57345 -13317
rect 59946 -13174 60346 -13162
rect 59946 -13208 59958 -13174
rect 60334 -13208 60346 -13174
rect 59946 -13220 60346 -13208
rect 59946 -13282 60346 -13270
rect 59946 -13316 59958 -13282
rect 60334 -13316 60346 -13282
rect 59946 -13328 60346 -13316
rect 59490 -13582 59548 -13570
rect 59490 -13650 59502 -13582
rect 59476 -13720 59502 -13650
rect 59490 -13758 59502 -13720
rect 59536 -13758 59548 -13582
rect 59490 -13770 59548 -13758
rect 59578 -13582 59636 -13570
rect 59578 -13758 59590 -13582
rect 59624 -13758 59636 -13582
rect 59578 -13770 59636 -13758
rect 59806 -13582 59864 -13570
rect 59806 -13758 59818 -13582
rect 59852 -13758 59864 -13582
rect 59806 -13770 59864 -13758
rect 59894 -13582 59952 -13570
rect 59894 -13758 59906 -13582
rect 59940 -13758 59952 -13582
rect 59894 -13770 59952 -13758
rect 60191 -13773 60321 -13765
rect 60191 -13807 60203 -13773
rect 60237 -13807 60321 -13773
rect 60191 -13817 60321 -13807
rect 61131 -13773 61261 -13765
rect 61131 -13807 61215 -13773
rect 61249 -13807 61261 -13773
rect 61131 -13817 61261 -13807
rect 60191 -13857 60321 -13847
rect 60191 -13891 60211 -13857
rect 60245 -13891 60321 -13857
rect 60191 -13901 60321 -13891
rect 61131 -13857 61261 -13847
rect 61131 -13891 61207 -13857
rect 61241 -13891 61261 -13857
rect 61131 -13901 61261 -13891
rect 57123 -14454 57175 -14429
rect 57123 -14488 57131 -14454
rect 57165 -14488 57175 -14454
rect 57123 -14533 57175 -14488
rect 57205 -14441 57263 -14429
rect 57205 -14475 57217 -14441
rect 57251 -14475 57263 -14441
rect 57205 -14533 57263 -14475
rect 57293 -14471 57345 -14429
rect 57293 -14505 57303 -14471
rect 57337 -14505 57345 -14471
rect 57293 -14533 57345 -14505
rect 60191 -13941 60321 -13931
rect 59489 -14095 59547 -14083
rect 59489 -14271 59501 -14095
rect 59535 -14271 59547 -14095
rect 59489 -14283 59547 -14271
rect 59577 -14095 59635 -14083
rect 59577 -14271 59589 -14095
rect 59623 -14271 59635 -14095
rect 59577 -14283 59635 -14271
rect 60191 -13975 60203 -13941
rect 60237 -13975 60321 -13941
rect 60191 -13985 60321 -13975
rect 61131 -13941 61261 -13931
rect 61131 -13975 61215 -13941
rect 61249 -13975 61261 -13941
rect 61131 -13985 61261 -13975
rect 59805 -14095 59863 -14083
rect 59805 -14271 59817 -14095
rect 59851 -14271 59863 -14095
rect 59805 -14283 59863 -14271
rect 59893 -14095 59951 -14083
rect 59893 -14271 59905 -14095
rect 59939 -14271 59951 -14095
rect 59893 -14283 59951 -14271
rect 60191 -14025 60321 -14015
rect 60191 -14059 60211 -14025
rect 60245 -14059 60321 -14025
rect 60191 -14069 60321 -14059
rect 61131 -14025 61261 -14015
rect 61131 -14059 61207 -14025
rect 61241 -14059 61261 -14025
rect 61131 -14069 61261 -14059
rect 60191 -14109 60321 -14099
rect 60191 -14143 60204 -14109
rect 60238 -14143 60321 -14109
rect 60191 -14151 60321 -14143
rect 61131 -14109 61261 -14099
rect 61131 -14143 61214 -14109
rect 61248 -14143 61261 -14109
rect 61131 -14151 61261 -14143
rect 59946 -14540 60346 -14528
rect 59946 -14574 59958 -14540
rect 60334 -14574 60346 -14540
rect 59946 -14586 60346 -14574
rect 59946 -14648 60346 -14636
rect 59946 -14682 59958 -14648
rect 60334 -14682 60346 -14648
rect 59946 -14694 60346 -14682
rect 55288 -15358 55488 -15346
rect 55288 -15392 55300 -15358
rect 55476 -15392 55488 -15358
rect 55288 -15404 55488 -15392
rect 55288 -15446 55488 -15434
rect 55288 -15480 55300 -15446
rect 55476 -15480 55488 -15446
rect 55288 -15492 55488 -15480
rect 53452 -18390 53510 -18378
rect 53452 -19166 53464 -18390
rect 53498 -19166 53510 -18390
rect 53452 -19178 53510 -19166
rect 53630 -18390 53688 -18378
rect 53630 -19166 53642 -18390
rect 53676 -19166 53688 -18390
rect 53630 -19178 53688 -19166
rect 55278 -18452 55336 -18440
rect 55278 -18628 55290 -18452
rect 55324 -18628 55336 -18452
rect 55278 -18640 55336 -18628
rect 55366 -18452 55424 -18440
rect 55366 -18628 55378 -18452
rect 55412 -18628 55424 -18452
rect 55366 -18640 55424 -18628
rect 53930 -18978 54730 -18966
rect 53930 -19012 53942 -18978
rect 54718 -19012 54730 -18978
rect 53930 -19024 54730 -19012
rect 53930 -19156 54730 -19144
rect 53930 -19190 53942 -19156
rect 54718 -19190 54730 -19156
rect 53930 -19202 54730 -19190
rect 55808 -18340 55866 -18328
rect 55808 -19116 55820 -18340
rect 55854 -19116 55866 -18340
rect 55808 -19128 55866 -19116
rect 55986 -18340 56044 -18328
rect 55986 -19116 55998 -18340
rect 56032 -19116 56044 -18340
rect 55986 -19128 56044 -19116
rect 57123 -18700 57175 -18655
rect 53452 -19408 53510 -19396
rect 53452 -20184 53464 -19408
rect 53498 -20184 53510 -19408
rect 53452 -20196 53510 -20184
rect 53630 -19408 53688 -19396
rect 53630 -20184 53642 -19408
rect 53676 -20184 53688 -19408
rect 53630 -20196 53688 -20184
rect 53930 -19384 54730 -19372
rect 53930 -19418 53942 -19384
rect 54718 -19418 54730 -19384
rect 53930 -19430 54730 -19418
rect 53930 -19562 54730 -19550
rect 53930 -19596 53942 -19562
rect 54718 -19596 54730 -19562
rect 53930 -19608 54730 -19596
rect 55268 -19948 55326 -19936
rect 55268 -20124 55280 -19948
rect 55314 -20124 55326 -19948
rect 55268 -20136 55326 -20124
rect 55356 -19948 55414 -19936
rect 55356 -20124 55368 -19948
rect 55402 -20124 55414 -19948
rect 55356 -20136 55414 -20124
rect 55808 -19454 55866 -19442
rect 55808 -20230 55820 -19454
rect 55854 -20230 55866 -19454
rect 55808 -20242 55866 -20230
rect 55986 -19454 56044 -19442
rect 55986 -20230 55998 -19454
rect 56032 -20230 56044 -19454
rect 55986 -20242 56044 -20230
rect 57123 -18734 57131 -18700
rect 57165 -18734 57175 -18700
rect 57123 -18759 57175 -18734
rect 57205 -18713 57263 -18655
rect 57205 -18747 57217 -18713
rect 57251 -18747 57263 -18713
rect 57205 -18759 57263 -18747
rect 57293 -18683 57345 -18655
rect 57293 -18717 57303 -18683
rect 57337 -18717 57345 -18683
rect 57293 -18759 57345 -18717
rect 59946 -18574 60346 -18562
rect 59946 -18608 59958 -18574
rect 60334 -18608 60346 -18574
rect 59946 -18620 60346 -18608
rect 59946 -18682 60346 -18670
rect 59946 -18716 59958 -18682
rect 60334 -18716 60346 -18682
rect 59946 -18728 60346 -18716
rect 59490 -18982 59548 -18970
rect 59490 -19050 59502 -18982
rect 59476 -19120 59502 -19050
rect 59490 -19158 59502 -19120
rect 59536 -19158 59548 -18982
rect 59490 -19170 59548 -19158
rect 59578 -18982 59636 -18970
rect 59578 -19158 59590 -18982
rect 59624 -19158 59636 -18982
rect 59578 -19170 59636 -19158
rect 59806 -18982 59864 -18970
rect 59806 -19158 59818 -18982
rect 59852 -19158 59864 -18982
rect 59806 -19170 59864 -19158
rect 59894 -18982 59952 -18970
rect 59894 -19158 59906 -18982
rect 59940 -19158 59952 -18982
rect 59894 -19170 59952 -19158
rect 60191 -19173 60321 -19165
rect 60191 -19207 60203 -19173
rect 60237 -19207 60321 -19173
rect 60191 -19217 60321 -19207
rect 61131 -19173 61261 -19165
rect 61131 -19207 61215 -19173
rect 61249 -19207 61261 -19173
rect 61131 -19217 61261 -19207
rect 60191 -19257 60321 -19247
rect 60191 -19291 60211 -19257
rect 60245 -19291 60321 -19257
rect 60191 -19301 60321 -19291
rect 61131 -19257 61261 -19247
rect 61131 -19291 61207 -19257
rect 61241 -19291 61261 -19257
rect 61131 -19301 61261 -19291
rect 57123 -19854 57175 -19829
rect 57123 -19888 57131 -19854
rect 57165 -19888 57175 -19854
rect 57123 -19933 57175 -19888
rect 57205 -19841 57263 -19829
rect 57205 -19875 57217 -19841
rect 57251 -19875 57263 -19841
rect 57205 -19933 57263 -19875
rect 57293 -19871 57345 -19829
rect 57293 -19905 57303 -19871
rect 57337 -19905 57345 -19871
rect 57293 -19933 57345 -19905
rect 60191 -19341 60321 -19331
rect 59489 -19495 59547 -19483
rect 59489 -19671 59501 -19495
rect 59535 -19671 59547 -19495
rect 59489 -19683 59547 -19671
rect 59577 -19495 59635 -19483
rect 59577 -19671 59589 -19495
rect 59623 -19671 59635 -19495
rect 59577 -19683 59635 -19671
rect 60191 -19375 60203 -19341
rect 60237 -19375 60321 -19341
rect 60191 -19385 60321 -19375
rect 61131 -19341 61261 -19331
rect 61131 -19375 61215 -19341
rect 61249 -19375 61261 -19341
rect 61131 -19385 61261 -19375
rect 59805 -19495 59863 -19483
rect 59805 -19671 59817 -19495
rect 59851 -19671 59863 -19495
rect 59805 -19683 59863 -19671
rect 59893 -19495 59951 -19483
rect 59893 -19671 59905 -19495
rect 59939 -19671 59951 -19495
rect 59893 -19683 59951 -19671
rect 60191 -19425 60321 -19415
rect 60191 -19459 60211 -19425
rect 60245 -19459 60321 -19425
rect 60191 -19469 60321 -19459
rect 61131 -19425 61261 -19415
rect 61131 -19459 61207 -19425
rect 61241 -19459 61261 -19425
rect 61131 -19469 61261 -19459
rect 60191 -19509 60321 -19499
rect 60191 -19543 60204 -19509
rect 60238 -19543 60321 -19509
rect 60191 -19551 60321 -19543
rect 61131 -19509 61261 -19499
rect 61131 -19543 61214 -19509
rect 61248 -19543 61261 -19509
rect 61131 -19551 61261 -19543
rect 59946 -19940 60346 -19928
rect 59946 -19974 59958 -19940
rect 60334 -19974 60346 -19940
rect 59946 -19986 60346 -19974
rect 59946 -20048 60346 -20036
rect 59946 -20082 59958 -20048
rect 60334 -20082 60346 -20048
rect 59946 -20094 60346 -20082
rect 55288 -20758 55488 -20746
rect 55288 -20792 55300 -20758
rect 55476 -20792 55488 -20758
rect 55288 -20804 55488 -20792
rect 55288 -20846 55488 -20834
rect 55288 -20880 55300 -20846
rect 55476 -20880 55488 -20846
rect 55288 -20892 55488 -20880
rect 53452 -23790 53510 -23778
rect 53452 -24566 53464 -23790
rect 53498 -24566 53510 -23790
rect 53452 -24578 53510 -24566
rect 53630 -23790 53688 -23778
rect 53630 -24566 53642 -23790
rect 53676 -24566 53688 -23790
rect 53630 -24578 53688 -24566
rect 55278 -23852 55336 -23840
rect 55278 -24028 55290 -23852
rect 55324 -24028 55336 -23852
rect 55278 -24040 55336 -24028
rect 55366 -23852 55424 -23840
rect 55366 -24028 55378 -23852
rect 55412 -24028 55424 -23852
rect 55366 -24040 55424 -24028
rect 53930 -24378 54730 -24366
rect 53930 -24412 53942 -24378
rect 54718 -24412 54730 -24378
rect 53930 -24424 54730 -24412
rect 53930 -24556 54730 -24544
rect 53930 -24590 53942 -24556
rect 54718 -24590 54730 -24556
rect 53930 -24602 54730 -24590
rect 55808 -23740 55866 -23728
rect 55808 -24516 55820 -23740
rect 55854 -24516 55866 -23740
rect 55808 -24528 55866 -24516
rect 55986 -23740 56044 -23728
rect 55986 -24516 55998 -23740
rect 56032 -24516 56044 -23740
rect 55986 -24528 56044 -24516
rect 57123 -24100 57175 -24055
rect 53452 -24808 53510 -24796
rect 53452 -25584 53464 -24808
rect 53498 -25584 53510 -24808
rect 53452 -25596 53510 -25584
rect 53630 -24808 53688 -24796
rect 53630 -25584 53642 -24808
rect 53676 -25584 53688 -24808
rect 53630 -25596 53688 -25584
rect 53930 -24784 54730 -24772
rect 53930 -24818 53942 -24784
rect 54718 -24818 54730 -24784
rect 53930 -24830 54730 -24818
rect 53930 -24962 54730 -24950
rect 53930 -24996 53942 -24962
rect 54718 -24996 54730 -24962
rect 53930 -25008 54730 -24996
rect 55268 -25348 55326 -25336
rect 55268 -25524 55280 -25348
rect 55314 -25524 55326 -25348
rect 55268 -25536 55326 -25524
rect 55356 -25348 55414 -25336
rect 55356 -25524 55368 -25348
rect 55402 -25524 55414 -25348
rect 55356 -25536 55414 -25524
rect 55808 -24854 55866 -24842
rect 55808 -25630 55820 -24854
rect 55854 -25630 55866 -24854
rect 55808 -25642 55866 -25630
rect 55986 -24854 56044 -24842
rect 55986 -25630 55998 -24854
rect 56032 -25630 56044 -24854
rect 55986 -25642 56044 -25630
rect 57123 -24134 57131 -24100
rect 57165 -24134 57175 -24100
rect 57123 -24159 57175 -24134
rect 57205 -24113 57263 -24055
rect 57205 -24147 57217 -24113
rect 57251 -24147 57263 -24113
rect 57205 -24159 57263 -24147
rect 57293 -24083 57345 -24055
rect 57293 -24117 57303 -24083
rect 57337 -24117 57345 -24083
rect 57293 -24159 57345 -24117
rect 59946 -23974 60346 -23962
rect 59946 -24008 59958 -23974
rect 60334 -24008 60346 -23974
rect 59946 -24020 60346 -24008
rect 59946 -24082 60346 -24070
rect 59946 -24116 59958 -24082
rect 60334 -24116 60346 -24082
rect 59946 -24128 60346 -24116
rect 59490 -24382 59548 -24370
rect 59490 -24450 59502 -24382
rect 59476 -24520 59502 -24450
rect 59490 -24558 59502 -24520
rect 59536 -24558 59548 -24382
rect 59490 -24570 59548 -24558
rect 59578 -24382 59636 -24370
rect 59578 -24558 59590 -24382
rect 59624 -24558 59636 -24382
rect 59578 -24570 59636 -24558
rect 59806 -24382 59864 -24370
rect 59806 -24558 59818 -24382
rect 59852 -24558 59864 -24382
rect 59806 -24570 59864 -24558
rect 59894 -24382 59952 -24370
rect 59894 -24558 59906 -24382
rect 59940 -24558 59952 -24382
rect 59894 -24570 59952 -24558
rect 60191 -24573 60321 -24565
rect 60191 -24607 60203 -24573
rect 60237 -24607 60321 -24573
rect 60191 -24617 60321 -24607
rect 61131 -24573 61261 -24565
rect 61131 -24607 61215 -24573
rect 61249 -24607 61261 -24573
rect 61131 -24617 61261 -24607
rect 60191 -24657 60321 -24647
rect 60191 -24691 60211 -24657
rect 60245 -24691 60321 -24657
rect 60191 -24701 60321 -24691
rect 61131 -24657 61261 -24647
rect 61131 -24691 61207 -24657
rect 61241 -24691 61261 -24657
rect 61131 -24701 61261 -24691
rect 57123 -25254 57175 -25229
rect 57123 -25288 57131 -25254
rect 57165 -25288 57175 -25254
rect 57123 -25333 57175 -25288
rect 57205 -25241 57263 -25229
rect 57205 -25275 57217 -25241
rect 57251 -25275 57263 -25241
rect 57205 -25333 57263 -25275
rect 57293 -25271 57345 -25229
rect 57293 -25305 57303 -25271
rect 57337 -25305 57345 -25271
rect 57293 -25333 57345 -25305
rect 60191 -24741 60321 -24731
rect 59489 -24895 59547 -24883
rect 59489 -25071 59501 -24895
rect 59535 -25071 59547 -24895
rect 59489 -25083 59547 -25071
rect 59577 -24895 59635 -24883
rect 59577 -25071 59589 -24895
rect 59623 -25071 59635 -24895
rect 59577 -25083 59635 -25071
rect 60191 -24775 60203 -24741
rect 60237 -24775 60321 -24741
rect 60191 -24785 60321 -24775
rect 61131 -24741 61261 -24731
rect 61131 -24775 61215 -24741
rect 61249 -24775 61261 -24741
rect 61131 -24785 61261 -24775
rect 59805 -24895 59863 -24883
rect 59805 -25071 59817 -24895
rect 59851 -25071 59863 -24895
rect 59805 -25083 59863 -25071
rect 59893 -24895 59951 -24883
rect 59893 -25071 59905 -24895
rect 59939 -25071 59951 -24895
rect 59893 -25083 59951 -25071
rect 60191 -24825 60321 -24815
rect 60191 -24859 60211 -24825
rect 60245 -24859 60321 -24825
rect 60191 -24869 60321 -24859
rect 61131 -24825 61261 -24815
rect 61131 -24859 61207 -24825
rect 61241 -24859 61261 -24825
rect 61131 -24869 61261 -24859
rect 60191 -24909 60321 -24899
rect 60191 -24943 60204 -24909
rect 60238 -24943 60321 -24909
rect 60191 -24951 60321 -24943
rect 61131 -24909 61261 -24899
rect 61131 -24943 61214 -24909
rect 61248 -24943 61261 -24909
rect 61131 -24951 61261 -24943
rect 59946 -25340 60346 -25328
rect 59946 -25374 59958 -25340
rect 60334 -25374 60346 -25340
rect 59946 -25386 60346 -25374
rect 59946 -25448 60346 -25436
rect 59946 -25482 59958 -25448
rect 60334 -25482 60346 -25448
rect 59946 -25494 60346 -25482
rect 55288 -26158 55488 -26146
rect 55288 -26192 55300 -26158
rect 55476 -26192 55488 -26158
rect 55288 -26204 55488 -26192
rect 55288 -26246 55488 -26234
rect 55288 -26280 55300 -26246
rect 55476 -26280 55488 -26246
rect 55288 -26292 55488 -26280
rect 53452 -29190 53510 -29178
rect 53452 -29966 53464 -29190
rect 53498 -29966 53510 -29190
rect 53452 -29978 53510 -29966
rect 53630 -29190 53688 -29178
rect 53630 -29966 53642 -29190
rect 53676 -29966 53688 -29190
rect 53630 -29978 53688 -29966
rect 55278 -29252 55336 -29240
rect 55278 -29428 55290 -29252
rect 55324 -29428 55336 -29252
rect 55278 -29440 55336 -29428
rect 55366 -29252 55424 -29240
rect 55366 -29428 55378 -29252
rect 55412 -29428 55424 -29252
rect 55366 -29440 55424 -29428
rect 53930 -29778 54730 -29766
rect 53930 -29812 53942 -29778
rect 54718 -29812 54730 -29778
rect 53930 -29824 54730 -29812
rect 53930 -29956 54730 -29944
rect 53930 -29990 53942 -29956
rect 54718 -29990 54730 -29956
rect 53930 -30002 54730 -29990
rect 55808 -29140 55866 -29128
rect 55808 -29916 55820 -29140
rect 55854 -29916 55866 -29140
rect 55808 -29928 55866 -29916
rect 55986 -29140 56044 -29128
rect 55986 -29916 55998 -29140
rect 56032 -29916 56044 -29140
rect 55986 -29928 56044 -29916
rect 57123 -29500 57175 -29455
rect 53452 -30208 53510 -30196
rect 53452 -30984 53464 -30208
rect 53498 -30984 53510 -30208
rect 53452 -30996 53510 -30984
rect 53630 -30208 53688 -30196
rect 53630 -30984 53642 -30208
rect 53676 -30984 53688 -30208
rect 53630 -30996 53688 -30984
rect 53930 -30184 54730 -30172
rect 53930 -30218 53942 -30184
rect 54718 -30218 54730 -30184
rect 53930 -30230 54730 -30218
rect 53930 -30362 54730 -30350
rect 53930 -30396 53942 -30362
rect 54718 -30396 54730 -30362
rect 53930 -30408 54730 -30396
rect 55268 -30748 55326 -30736
rect 55268 -30924 55280 -30748
rect 55314 -30924 55326 -30748
rect 55268 -30936 55326 -30924
rect 55356 -30748 55414 -30736
rect 55356 -30924 55368 -30748
rect 55402 -30924 55414 -30748
rect 55356 -30936 55414 -30924
rect 55808 -30254 55866 -30242
rect 55808 -31030 55820 -30254
rect 55854 -31030 55866 -30254
rect 55808 -31042 55866 -31030
rect 55986 -30254 56044 -30242
rect 55986 -31030 55998 -30254
rect 56032 -31030 56044 -30254
rect 55986 -31042 56044 -31030
rect 57123 -29534 57131 -29500
rect 57165 -29534 57175 -29500
rect 57123 -29559 57175 -29534
rect 57205 -29513 57263 -29455
rect 57205 -29547 57217 -29513
rect 57251 -29547 57263 -29513
rect 57205 -29559 57263 -29547
rect 57293 -29483 57345 -29455
rect 57293 -29517 57303 -29483
rect 57337 -29517 57345 -29483
rect 57293 -29559 57345 -29517
rect 59946 -29374 60346 -29362
rect 59946 -29408 59958 -29374
rect 60334 -29408 60346 -29374
rect 59946 -29420 60346 -29408
rect 59946 -29482 60346 -29470
rect 59946 -29516 59958 -29482
rect 60334 -29516 60346 -29482
rect 59946 -29528 60346 -29516
rect 59490 -29782 59548 -29770
rect 59490 -29850 59502 -29782
rect 59476 -29920 59502 -29850
rect 59490 -29958 59502 -29920
rect 59536 -29958 59548 -29782
rect 59490 -29970 59548 -29958
rect 59578 -29782 59636 -29770
rect 59578 -29958 59590 -29782
rect 59624 -29958 59636 -29782
rect 59578 -29970 59636 -29958
rect 59806 -29782 59864 -29770
rect 59806 -29958 59818 -29782
rect 59852 -29958 59864 -29782
rect 59806 -29970 59864 -29958
rect 59894 -29782 59952 -29770
rect 59894 -29958 59906 -29782
rect 59940 -29958 59952 -29782
rect 59894 -29970 59952 -29958
rect 60191 -29973 60321 -29965
rect 60191 -30007 60203 -29973
rect 60237 -30007 60321 -29973
rect 60191 -30017 60321 -30007
rect 61131 -29973 61261 -29965
rect 61131 -30007 61215 -29973
rect 61249 -30007 61261 -29973
rect 61131 -30017 61261 -30007
rect 60191 -30057 60321 -30047
rect 60191 -30091 60211 -30057
rect 60245 -30091 60321 -30057
rect 60191 -30101 60321 -30091
rect 61131 -30057 61261 -30047
rect 61131 -30091 61207 -30057
rect 61241 -30091 61261 -30057
rect 61131 -30101 61261 -30091
rect 57123 -30654 57175 -30629
rect 57123 -30688 57131 -30654
rect 57165 -30688 57175 -30654
rect 57123 -30733 57175 -30688
rect 57205 -30641 57263 -30629
rect 57205 -30675 57217 -30641
rect 57251 -30675 57263 -30641
rect 57205 -30733 57263 -30675
rect 57293 -30671 57345 -30629
rect 57293 -30705 57303 -30671
rect 57337 -30705 57345 -30671
rect 57293 -30733 57345 -30705
rect 60191 -30141 60321 -30131
rect 59489 -30295 59547 -30283
rect 59489 -30471 59501 -30295
rect 59535 -30471 59547 -30295
rect 59489 -30483 59547 -30471
rect 59577 -30295 59635 -30283
rect 59577 -30471 59589 -30295
rect 59623 -30471 59635 -30295
rect 59577 -30483 59635 -30471
rect 60191 -30175 60203 -30141
rect 60237 -30175 60321 -30141
rect 60191 -30185 60321 -30175
rect 61131 -30141 61261 -30131
rect 61131 -30175 61215 -30141
rect 61249 -30175 61261 -30141
rect 61131 -30185 61261 -30175
rect 59805 -30295 59863 -30283
rect 59805 -30471 59817 -30295
rect 59851 -30471 59863 -30295
rect 59805 -30483 59863 -30471
rect 59893 -30295 59951 -30283
rect 59893 -30471 59905 -30295
rect 59939 -30471 59951 -30295
rect 59893 -30483 59951 -30471
rect 60191 -30225 60321 -30215
rect 60191 -30259 60211 -30225
rect 60245 -30259 60321 -30225
rect 60191 -30269 60321 -30259
rect 61131 -30225 61261 -30215
rect 61131 -30259 61207 -30225
rect 61241 -30259 61261 -30225
rect 61131 -30269 61261 -30259
rect 60191 -30309 60321 -30299
rect 60191 -30343 60204 -30309
rect 60238 -30343 60321 -30309
rect 60191 -30351 60321 -30343
rect 61131 -30309 61261 -30299
rect 61131 -30343 61214 -30309
rect 61248 -30343 61261 -30309
rect 61131 -30351 61261 -30343
rect 59946 -30740 60346 -30728
rect 59946 -30774 59958 -30740
rect 60334 -30774 60346 -30740
rect 59946 -30786 60346 -30774
rect 59946 -30848 60346 -30836
rect 59946 -30882 59958 -30848
rect 60334 -30882 60346 -30848
rect 59946 -30894 60346 -30882
rect 55288 -31558 55488 -31546
rect 55288 -31592 55300 -31558
rect 55476 -31592 55488 -31558
rect 55288 -31604 55488 -31592
rect 55288 -31646 55488 -31634
rect 55288 -31680 55300 -31646
rect 55476 -31680 55488 -31646
rect 55288 -31692 55488 -31680
rect 53452 -34590 53510 -34578
rect 53452 -35366 53464 -34590
rect 53498 -35366 53510 -34590
rect 53452 -35378 53510 -35366
rect 53630 -34590 53688 -34578
rect 53630 -35366 53642 -34590
rect 53676 -35366 53688 -34590
rect 53630 -35378 53688 -35366
rect 55278 -34652 55336 -34640
rect 55278 -34828 55290 -34652
rect 55324 -34828 55336 -34652
rect 55278 -34840 55336 -34828
rect 55366 -34652 55424 -34640
rect 55366 -34828 55378 -34652
rect 55412 -34828 55424 -34652
rect 55366 -34840 55424 -34828
rect 53930 -35178 54730 -35166
rect 53930 -35212 53942 -35178
rect 54718 -35212 54730 -35178
rect 53930 -35224 54730 -35212
rect 53930 -35356 54730 -35344
rect 53930 -35390 53942 -35356
rect 54718 -35390 54730 -35356
rect 53930 -35402 54730 -35390
rect 55808 -34540 55866 -34528
rect 55808 -35316 55820 -34540
rect 55854 -35316 55866 -34540
rect 55808 -35328 55866 -35316
rect 55986 -34540 56044 -34528
rect 55986 -35316 55998 -34540
rect 56032 -35316 56044 -34540
rect 55986 -35328 56044 -35316
rect 57123 -34900 57175 -34855
rect 53452 -35608 53510 -35596
rect 53452 -36384 53464 -35608
rect 53498 -36384 53510 -35608
rect 53452 -36396 53510 -36384
rect 53630 -35608 53688 -35596
rect 53630 -36384 53642 -35608
rect 53676 -36384 53688 -35608
rect 53630 -36396 53688 -36384
rect 53930 -35584 54730 -35572
rect 53930 -35618 53942 -35584
rect 54718 -35618 54730 -35584
rect 53930 -35630 54730 -35618
rect 53930 -35762 54730 -35750
rect 53930 -35796 53942 -35762
rect 54718 -35796 54730 -35762
rect 53930 -35808 54730 -35796
rect 55268 -36148 55326 -36136
rect 55268 -36324 55280 -36148
rect 55314 -36324 55326 -36148
rect 55268 -36336 55326 -36324
rect 55356 -36148 55414 -36136
rect 55356 -36324 55368 -36148
rect 55402 -36324 55414 -36148
rect 55356 -36336 55414 -36324
rect 55808 -35654 55866 -35642
rect 55808 -36430 55820 -35654
rect 55854 -36430 55866 -35654
rect 55808 -36442 55866 -36430
rect 55986 -35654 56044 -35642
rect 55986 -36430 55998 -35654
rect 56032 -36430 56044 -35654
rect 55986 -36442 56044 -36430
rect 57123 -34934 57131 -34900
rect 57165 -34934 57175 -34900
rect 57123 -34959 57175 -34934
rect 57205 -34913 57263 -34855
rect 57205 -34947 57217 -34913
rect 57251 -34947 57263 -34913
rect 57205 -34959 57263 -34947
rect 57293 -34883 57345 -34855
rect 57293 -34917 57303 -34883
rect 57337 -34917 57345 -34883
rect 57293 -34959 57345 -34917
rect 59946 -34774 60346 -34762
rect 59946 -34808 59958 -34774
rect 60334 -34808 60346 -34774
rect 59946 -34820 60346 -34808
rect 59946 -34882 60346 -34870
rect 59946 -34916 59958 -34882
rect 60334 -34916 60346 -34882
rect 59946 -34928 60346 -34916
rect 59490 -35182 59548 -35170
rect 59490 -35250 59502 -35182
rect 59476 -35320 59502 -35250
rect 59490 -35358 59502 -35320
rect 59536 -35358 59548 -35182
rect 59490 -35370 59548 -35358
rect 59578 -35182 59636 -35170
rect 59578 -35358 59590 -35182
rect 59624 -35358 59636 -35182
rect 59578 -35370 59636 -35358
rect 59806 -35182 59864 -35170
rect 59806 -35358 59818 -35182
rect 59852 -35358 59864 -35182
rect 59806 -35370 59864 -35358
rect 59894 -35182 59952 -35170
rect 59894 -35358 59906 -35182
rect 59940 -35358 59952 -35182
rect 59894 -35370 59952 -35358
rect 60191 -35373 60321 -35365
rect 60191 -35407 60203 -35373
rect 60237 -35407 60321 -35373
rect 60191 -35417 60321 -35407
rect 61131 -35373 61261 -35365
rect 61131 -35407 61215 -35373
rect 61249 -35407 61261 -35373
rect 61131 -35417 61261 -35407
rect 60191 -35457 60321 -35447
rect 60191 -35491 60211 -35457
rect 60245 -35491 60321 -35457
rect 60191 -35501 60321 -35491
rect 61131 -35457 61261 -35447
rect 61131 -35491 61207 -35457
rect 61241 -35491 61261 -35457
rect 61131 -35501 61261 -35491
rect 57123 -36054 57175 -36029
rect 57123 -36088 57131 -36054
rect 57165 -36088 57175 -36054
rect 57123 -36133 57175 -36088
rect 57205 -36041 57263 -36029
rect 57205 -36075 57217 -36041
rect 57251 -36075 57263 -36041
rect 57205 -36133 57263 -36075
rect 57293 -36071 57345 -36029
rect 57293 -36105 57303 -36071
rect 57337 -36105 57345 -36071
rect 57293 -36133 57345 -36105
rect 60191 -35541 60321 -35531
rect 59489 -35695 59547 -35683
rect 59489 -35871 59501 -35695
rect 59535 -35871 59547 -35695
rect 59489 -35883 59547 -35871
rect 59577 -35695 59635 -35683
rect 59577 -35871 59589 -35695
rect 59623 -35871 59635 -35695
rect 59577 -35883 59635 -35871
rect 60191 -35575 60203 -35541
rect 60237 -35575 60321 -35541
rect 60191 -35585 60321 -35575
rect 61131 -35541 61261 -35531
rect 61131 -35575 61215 -35541
rect 61249 -35575 61261 -35541
rect 61131 -35585 61261 -35575
rect 59805 -35695 59863 -35683
rect 59805 -35871 59817 -35695
rect 59851 -35871 59863 -35695
rect 59805 -35883 59863 -35871
rect 59893 -35695 59951 -35683
rect 59893 -35871 59905 -35695
rect 59939 -35871 59951 -35695
rect 59893 -35883 59951 -35871
rect 60191 -35625 60321 -35615
rect 60191 -35659 60211 -35625
rect 60245 -35659 60321 -35625
rect 60191 -35669 60321 -35659
rect 61131 -35625 61261 -35615
rect 61131 -35659 61207 -35625
rect 61241 -35659 61261 -35625
rect 61131 -35669 61261 -35659
rect 60191 -35709 60321 -35699
rect 60191 -35743 60204 -35709
rect 60238 -35743 60321 -35709
rect 60191 -35751 60321 -35743
rect 61131 -35709 61261 -35699
rect 61131 -35743 61214 -35709
rect 61248 -35743 61261 -35709
rect 61131 -35751 61261 -35743
rect 59946 -36140 60346 -36128
rect 59946 -36174 59958 -36140
rect 60334 -36174 60346 -36140
rect 59946 -36186 60346 -36174
rect 59946 -36248 60346 -36236
rect 59946 -36282 59958 -36248
rect 60334 -36282 60346 -36248
rect 59946 -36294 60346 -36282
rect 55288 -36958 55488 -36946
rect 55288 -36992 55300 -36958
rect 55476 -36992 55488 -36958
rect 55288 -37004 55488 -36992
rect 55288 -37046 55488 -37034
rect 55288 -37080 55300 -37046
rect 55476 -37080 55488 -37046
rect 55288 -37092 55488 -37080
rect 75574 -38451 75626 -38435
rect 75574 -38485 75582 -38451
rect 75616 -38485 75626 -38451
rect 75574 -38519 75626 -38485
rect 75574 -38553 75582 -38519
rect 75616 -38553 75626 -38519
rect 75574 -38565 75626 -38553
rect 75656 -38451 75708 -38435
rect 75656 -38485 75666 -38451
rect 75700 -38485 75708 -38451
rect 75656 -38519 75708 -38485
rect 75656 -38553 75666 -38519
rect 75700 -38553 75708 -38519
rect 75656 -38565 75708 -38553
rect 75850 -38451 75902 -38435
rect 75850 -38485 75858 -38451
rect 75892 -38485 75902 -38451
rect 75850 -38519 75902 -38485
rect 75850 -38553 75858 -38519
rect 75892 -38553 75902 -38519
rect 75850 -38565 75902 -38553
rect 75932 -38451 75984 -38435
rect 75932 -38485 75942 -38451
rect 75976 -38485 75984 -38451
rect 75932 -38519 75984 -38485
rect 75932 -38553 75942 -38519
rect 75976 -38553 75984 -38519
rect 75932 -38565 75984 -38553
rect 76124 -38451 76176 -38435
rect 76124 -38485 76132 -38451
rect 76166 -38485 76176 -38451
rect 76124 -38519 76176 -38485
rect 76124 -38553 76132 -38519
rect 76166 -38553 76176 -38519
rect 76124 -38565 76176 -38553
rect 76206 -38451 76258 -38435
rect 76206 -38485 76216 -38451
rect 76250 -38485 76258 -38451
rect 76206 -38519 76258 -38485
rect 76206 -38553 76216 -38519
rect 76250 -38553 76258 -38519
rect 76206 -38565 76258 -38553
rect 76400 -38451 76452 -38435
rect 76400 -38485 76408 -38451
rect 76442 -38485 76452 -38451
rect 76400 -38519 76452 -38485
rect 76400 -38553 76408 -38519
rect 76442 -38553 76452 -38519
rect 76400 -38565 76452 -38553
rect 76482 -38451 76534 -38435
rect 76482 -38485 76492 -38451
rect 76526 -38485 76534 -38451
rect 76482 -38519 76534 -38485
rect 76482 -38553 76492 -38519
rect 76526 -38553 76534 -38519
rect 76482 -38565 76534 -38553
rect 76676 -38451 76728 -38435
rect 76676 -38485 76684 -38451
rect 76718 -38485 76728 -38451
rect 76676 -38519 76728 -38485
rect 76676 -38553 76684 -38519
rect 76718 -38553 76728 -38519
rect 76676 -38565 76728 -38553
rect 76758 -38451 76810 -38435
rect 76758 -38485 76768 -38451
rect 76802 -38485 76810 -38451
rect 76758 -38519 76810 -38485
rect 76758 -38553 76768 -38519
rect 76802 -38553 76810 -38519
rect 76758 -38565 76810 -38553
rect 77966 -39465 78019 -39425
rect 77605 -39485 77657 -39465
rect 77605 -39519 77613 -39485
rect 77647 -39519 77657 -39485
rect 77605 -39549 77657 -39519
rect 77687 -39491 77753 -39465
rect 77687 -39525 77703 -39491
rect 77737 -39525 77753 -39491
rect 77687 -39549 77753 -39525
rect 77783 -39505 77837 -39465
rect 77783 -39539 77793 -39505
rect 77827 -39539 77837 -39505
rect 77783 -39549 77837 -39539
rect 77867 -39491 77921 -39465
rect 77867 -39525 77877 -39491
rect 77911 -39525 77921 -39491
rect 77867 -39549 77921 -39525
rect 77951 -39505 78019 -39465
rect 77951 -39539 77971 -39505
rect 78005 -39539 78019 -39505
rect 77951 -39549 78019 -39539
rect 77966 -39555 78019 -39549
rect 78049 -39467 78103 -39425
rect 78424 -39465 78477 -39425
rect 78049 -39501 78059 -39467
rect 78093 -39501 78103 -39467
rect 78049 -39555 78103 -39501
rect 78159 -39491 78211 -39465
rect 78159 -39525 78167 -39491
rect 78201 -39525 78211 -39491
rect 78159 -39549 78211 -39525
rect 78241 -39505 78295 -39465
rect 78241 -39539 78251 -39505
rect 78285 -39539 78295 -39505
rect 78241 -39549 78295 -39539
rect 78325 -39491 78379 -39465
rect 78325 -39525 78335 -39491
rect 78369 -39525 78379 -39491
rect 78325 -39549 78379 -39525
rect 78409 -39505 78477 -39465
rect 78409 -39539 78429 -39505
rect 78463 -39539 78477 -39505
rect 78409 -39549 78477 -39539
rect 78424 -39555 78477 -39549
rect 78507 -39467 78563 -39425
rect 78845 -39443 78897 -39425
rect 78507 -39501 78517 -39467
rect 78551 -39501 78563 -39467
rect 78507 -39555 78563 -39501
rect 78649 -39481 78705 -39443
rect 78649 -39515 78661 -39481
rect 78695 -39515 78705 -39481
rect 78649 -39527 78705 -39515
rect 78735 -39527 78789 -39443
rect 78819 -39509 78897 -39443
rect 78819 -39527 78853 -39509
rect 78845 -39543 78853 -39527
rect 78887 -39543 78897 -39509
rect 78845 -39555 78897 -39543
rect 78927 -39509 78983 -39425
rect 78927 -39543 78937 -39509
rect 78971 -39543 78983 -39509
rect 78927 -39555 78983 -39543
rect 80806 -39487 80858 -39475
rect 80806 -39521 80814 -39487
rect 80848 -39521 80858 -39487
rect 80806 -39555 80858 -39521
rect 80806 -39589 80814 -39555
rect 80848 -39589 80858 -39555
rect 80806 -39605 80858 -39589
rect 80888 -39487 80940 -39475
rect 80888 -39521 80898 -39487
rect 80932 -39521 80940 -39487
rect 80888 -39555 80940 -39521
rect 80888 -39589 80898 -39555
rect 80932 -39589 80940 -39555
rect 80888 -39605 80940 -39589
rect 81051 -39559 81103 -39475
rect 81051 -39593 81059 -39559
rect 81093 -39593 81103 -39559
rect 81051 -39605 81103 -39593
rect 81133 -39551 81187 -39475
rect 81133 -39585 81143 -39551
rect 81177 -39585 81187 -39551
rect 81133 -39605 81187 -39585
rect 81217 -39559 81271 -39475
rect 81217 -39593 81227 -39559
rect 81261 -39593 81271 -39559
rect 81217 -39605 81271 -39593
rect 81301 -39551 81355 -39475
rect 81301 -39585 81311 -39551
rect 81345 -39585 81355 -39551
rect 81301 -39605 81355 -39585
rect 81385 -39558 81437 -39475
rect 81385 -39592 81395 -39558
rect 81429 -39592 81437 -39558
rect 81385 -39605 81437 -39592
rect 81514 -39491 81566 -39475
rect 81514 -39525 81522 -39491
rect 81556 -39525 81566 -39491
rect 81514 -39559 81566 -39525
rect 81514 -39593 81522 -39559
rect 81556 -39593 81566 -39559
rect 81514 -39605 81566 -39593
rect 81596 -39491 81650 -39475
rect 81596 -39525 81606 -39491
rect 81640 -39525 81650 -39491
rect 81596 -39559 81650 -39525
rect 81596 -39593 81606 -39559
rect 81640 -39593 81650 -39559
rect 81596 -39605 81650 -39593
rect 81680 -39559 81734 -39475
rect 81680 -39593 81690 -39559
rect 81724 -39593 81734 -39559
rect 81680 -39605 81734 -39593
rect 81764 -39491 81818 -39475
rect 81764 -39525 81774 -39491
rect 81808 -39525 81818 -39491
rect 81764 -39559 81818 -39525
rect 81764 -39593 81774 -39559
rect 81808 -39593 81818 -39559
rect 81764 -39605 81818 -39593
rect 81848 -39559 81902 -39475
rect 81848 -39593 81858 -39559
rect 81892 -39593 81902 -39559
rect 81848 -39605 81902 -39593
rect 81932 -39491 81986 -39475
rect 81932 -39525 81942 -39491
rect 81976 -39525 81986 -39491
rect 81932 -39559 81986 -39525
rect 81932 -39593 81942 -39559
rect 81976 -39593 81986 -39559
rect 81932 -39605 81986 -39593
rect 82016 -39559 82070 -39475
rect 82016 -39593 82026 -39559
rect 82060 -39593 82070 -39559
rect 82016 -39605 82070 -39593
rect 82100 -39491 82154 -39475
rect 82100 -39525 82110 -39491
rect 82144 -39525 82154 -39491
rect 82100 -39559 82154 -39525
rect 82100 -39593 82110 -39559
rect 82144 -39593 82154 -39559
rect 82100 -39605 82154 -39593
rect 82184 -39559 82238 -39475
rect 82184 -39593 82194 -39559
rect 82228 -39593 82238 -39559
rect 82184 -39605 82238 -39593
rect 82268 -39491 82322 -39475
rect 82268 -39525 82278 -39491
rect 82312 -39525 82322 -39491
rect 82268 -39559 82322 -39525
rect 82268 -39593 82278 -39559
rect 82312 -39593 82322 -39559
rect 82268 -39605 82322 -39593
rect 82352 -39559 82406 -39475
rect 82352 -39593 82362 -39559
rect 82396 -39593 82406 -39559
rect 82352 -39605 82406 -39593
rect 82436 -39491 82490 -39475
rect 82436 -39525 82446 -39491
rect 82480 -39525 82490 -39491
rect 82436 -39559 82490 -39525
rect 82436 -39593 82446 -39559
rect 82480 -39593 82490 -39559
rect 82436 -39605 82490 -39593
rect 82520 -39559 82574 -39475
rect 82520 -39593 82530 -39559
rect 82564 -39593 82574 -39559
rect 82520 -39605 82574 -39593
rect 82604 -39491 82658 -39475
rect 82604 -39525 82614 -39491
rect 82648 -39525 82658 -39491
rect 82604 -39559 82658 -39525
rect 82604 -39593 82614 -39559
rect 82648 -39593 82658 -39559
rect 82604 -39605 82658 -39593
rect 82688 -39559 82742 -39475
rect 82688 -39593 82698 -39559
rect 82732 -39593 82742 -39559
rect 82688 -39605 82742 -39593
rect 82772 -39491 82826 -39475
rect 82772 -39525 82782 -39491
rect 82816 -39525 82826 -39491
rect 82772 -39559 82826 -39525
rect 82772 -39593 82782 -39559
rect 82816 -39593 82826 -39559
rect 82772 -39605 82826 -39593
rect 82856 -39491 82908 -39475
rect 82856 -39525 82866 -39491
rect 82900 -39525 82908 -39491
rect 82856 -39559 82908 -39525
rect 82856 -39593 82866 -39559
rect 82900 -39593 82908 -39559
rect 82856 -39605 82908 -39593
rect 82986 -39491 83038 -39475
rect 82986 -39525 82994 -39491
rect 83028 -39525 83038 -39491
rect 82986 -39559 83038 -39525
rect 82986 -39593 82994 -39559
rect 83028 -39593 83038 -39559
rect 82986 -39605 83038 -39593
rect 83068 -39491 83122 -39475
rect 83068 -39525 83078 -39491
rect 83112 -39525 83122 -39491
rect 83068 -39559 83122 -39525
rect 83068 -39593 83078 -39559
rect 83112 -39593 83122 -39559
rect 83068 -39605 83122 -39593
rect 83152 -39559 83206 -39475
rect 83152 -39593 83162 -39559
rect 83196 -39593 83206 -39559
rect 83152 -39605 83206 -39593
rect 83236 -39491 83290 -39475
rect 83236 -39525 83246 -39491
rect 83280 -39525 83290 -39491
rect 83236 -39559 83290 -39525
rect 83236 -39593 83246 -39559
rect 83280 -39593 83290 -39559
rect 83236 -39605 83290 -39593
rect 83320 -39559 83374 -39475
rect 83320 -39593 83330 -39559
rect 83364 -39593 83374 -39559
rect 83320 -39605 83374 -39593
rect 83404 -39491 83458 -39475
rect 83404 -39525 83414 -39491
rect 83448 -39525 83458 -39491
rect 83404 -39559 83458 -39525
rect 83404 -39593 83414 -39559
rect 83448 -39593 83458 -39559
rect 83404 -39605 83458 -39593
rect 83488 -39559 83542 -39475
rect 83488 -39593 83498 -39559
rect 83532 -39593 83542 -39559
rect 83488 -39605 83542 -39593
rect 83572 -39491 83626 -39475
rect 83572 -39525 83582 -39491
rect 83616 -39525 83626 -39491
rect 83572 -39559 83626 -39525
rect 83572 -39593 83582 -39559
rect 83616 -39593 83626 -39559
rect 83572 -39605 83626 -39593
rect 83656 -39559 83710 -39475
rect 83656 -39593 83666 -39559
rect 83700 -39593 83710 -39559
rect 83656 -39605 83710 -39593
rect 83740 -39491 83794 -39475
rect 83740 -39525 83750 -39491
rect 83784 -39525 83794 -39491
rect 83740 -39559 83794 -39525
rect 83740 -39593 83750 -39559
rect 83784 -39593 83794 -39559
rect 83740 -39605 83794 -39593
rect 83824 -39559 83878 -39475
rect 83824 -39593 83834 -39559
rect 83868 -39593 83878 -39559
rect 83824 -39605 83878 -39593
rect 83908 -39491 83962 -39475
rect 83908 -39525 83918 -39491
rect 83952 -39525 83962 -39491
rect 83908 -39559 83962 -39525
rect 83908 -39593 83918 -39559
rect 83952 -39593 83962 -39559
rect 83908 -39605 83962 -39593
rect 83992 -39559 84046 -39475
rect 83992 -39593 84002 -39559
rect 84036 -39593 84046 -39559
rect 83992 -39605 84046 -39593
rect 84076 -39491 84130 -39475
rect 84076 -39525 84086 -39491
rect 84120 -39525 84130 -39491
rect 84076 -39559 84130 -39525
rect 84076 -39593 84086 -39559
rect 84120 -39593 84130 -39559
rect 84076 -39605 84130 -39593
rect 84160 -39559 84214 -39475
rect 84160 -39593 84170 -39559
rect 84204 -39593 84214 -39559
rect 84160 -39605 84214 -39593
rect 84244 -39491 84298 -39475
rect 84244 -39525 84254 -39491
rect 84288 -39525 84298 -39491
rect 84244 -39559 84298 -39525
rect 84244 -39593 84254 -39559
rect 84288 -39593 84298 -39559
rect 84244 -39605 84298 -39593
rect 84328 -39491 84380 -39475
rect 84328 -39525 84338 -39491
rect 84372 -39525 84380 -39491
rect 84328 -39559 84380 -39525
rect 84328 -39593 84338 -39559
rect 84372 -39593 84380 -39559
rect 84328 -39605 84380 -39593
rect 84458 -39491 84510 -39475
rect 84458 -39525 84466 -39491
rect 84500 -39525 84510 -39491
rect 84458 -39559 84510 -39525
rect 84458 -39593 84466 -39559
rect 84500 -39593 84510 -39559
rect 84458 -39605 84510 -39593
rect 84540 -39491 84594 -39475
rect 84540 -39525 84550 -39491
rect 84584 -39525 84594 -39491
rect 84540 -39559 84594 -39525
rect 84540 -39593 84550 -39559
rect 84584 -39593 84594 -39559
rect 84540 -39605 84594 -39593
rect 84624 -39559 84678 -39475
rect 84624 -39593 84634 -39559
rect 84668 -39593 84678 -39559
rect 84624 -39605 84678 -39593
rect 84708 -39491 84762 -39475
rect 84708 -39525 84718 -39491
rect 84752 -39525 84762 -39491
rect 84708 -39559 84762 -39525
rect 84708 -39593 84718 -39559
rect 84752 -39593 84762 -39559
rect 84708 -39605 84762 -39593
rect 84792 -39559 84846 -39475
rect 84792 -39593 84802 -39559
rect 84836 -39593 84846 -39559
rect 84792 -39605 84846 -39593
rect 84876 -39491 84930 -39475
rect 84876 -39525 84886 -39491
rect 84920 -39525 84930 -39491
rect 84876 -39559 84930 -39525
rect 84876 -39593 84886 -39559
rect 84920 -39593 84930 -39559
rect 84876 -39605 84930 -39593
rect 84960 -39559 85014 -39475
rect 84960 -39593 84970 -39559
rect 85004 -39593 85014 -39559
rect 84960 -39605 85014 -39593
rect 85044 -39491 85098 -39475
rect 85044 -39525 85054 -39491
rect 85088 -39525 85098 -39491
rect 85044 -39559 85098 -39525
rect 85044 -39593 85054 -39559
rect 85088 -39593 85098 -39559
rect 85044 -39605 85098 -39593
rect 85128 -39559 85182 -39475
rect 85128 -39593 85138 -39559
rect 85172 -39593 85182 -39559
rect 85128 -39605 85182 -39593
rect 85212 -39491 85266 -39475
rect 85212 -39525 85222 -39491
rect 85256 -39525 85266 -39491
rect 85212 -39559 85266 -39525
rect 85212 -39593 85222 -39559
rect 85256 -39593 85266 -39559
rect 85212 -39605 85266 -39593
rect 85296 -39559 85350 -39475
rect 85296 -39593 85306 -39559
rect 85340 -39593 85350 -39559
rect 85296 -39605 85350 -39593
rect 85380 -39491 85434 -39475
rect 85380 -39525 85390 -39491
rect 85424 -39525 85434 -39491
rect 85380 -39559 85434 -39525
rect 85380 -39593 85390 -39559
rect 85424 -39593 85434 -39559
rect 85380 -39605 85434 -39593
rect 85464 -39559 85518 -39475
rect 85464 -39593 85474 -39559
rect 85508 -39593 85518 -39559
rect 85464 -39605 85518 -39593
rect 85548 -39491 85602 -39475
rect 85548 -39525 85558 -39491
rect 85592 -39525 85602 -39491
rect 85548 -39559 85602 -39525
rect 85548 -39593 85558 -39559
rect 85592 -39593 85602 -39559
rect 85548 -39605 85602 -39593
rect 85632 -39559 85686 -39475
rect 85632 -39593 85642 -39559
rect 85676 -39593 85686 -39559
rect 85632 -39605 85686 -39593
rect 85716 -39491 85770 -39475
rect 85716 -39525 85726 -39491
rect 85760 -39525 85770 -39491
rect 85716 -39559 85770 -39525
rect 85716 -39593 85726 -39559
rect 85760 -39593 85770 -39559
rect 85716 -39605 85770 -39593
rect 85800 -39491 85852 -39475
rect 85800 -39525 85810 -39491
rect 85844 -39525 85852 -39491
rect 85800 -39559 85852 -39525
rect 85800 -39593 85810 -39559
rect 85844 -39593 85852 -39559
rect 85800 -39605 85852 -39593
rect 85930 -39491 85982 -39475
rect 85930 -39525 85938 -39491
rect 85972 -39525 85982 -39491
rect 85930 -39559 85982 -39525
rect 85930 -39593 85938 -39559
rect 85972 -39593 85982 -39559
rect 85930 -39605 85982 -39593
rect 86012 -39491 86066 -39475
rect 86012 -39525 86022 -39491
rect 86056 -39525 86066 -39491
rect 86012 -39559 86066 -39525
rect 86012 -39593 86022 -39559
rect 86056 -39593 86066 -39559
rect 86012 -39605 86066 -39593
rect 86096 -39559 86150 -39475
rect 86096 -39593 86106 -39559
rect 86140 -39593 86150 -39559
rect 86096 -39605 86150 -39593
rect 86180 -39491 86234 -39475
rect 86180 -39525 86190 -39491
rect 86224 -39525 86234 -39491
rect 86180 -39559 86234 -39525
rect 86180 -39593 86190 -39559
rect 86224 -39593 86234 -39559
rect 86180 -39605 86234 -39593
rect 86264 -39559 86318 -39475
rect 86264 -39593 86274 -39559
rect 86308 -39593 86318 -39559
rect 86264 -39605 86318 -39593
rect 86348 -39491 86402 -39475
rect 86348 -39525 86358 -39491
rect 86392 -39525 86402 -39491
rect 86348 -39559 86402 -39525
rect 86348 -39593 86358 -39559
rect 86392 -39593 86402 -39559
rect 86348 -39605 86402 -39593
rect 86432 -39559 86486 -39475
rect 86432 -39593 86442 -39559
rect 86476 -39593 86486 -39559
rect 86432 -39605 86486 -39593
rect 86516 -39491 86570 -39475
rect 86516 -39525 86526 -39491
rect 86560 -39525 86570 -39491
rect 86516 -39559 86570 -39525
rect 86516 -39593 86526 -39559
rect 86560 -39593 86570 -39559
rect 86516 -39605 86570 -39593
rect 86600 -39559 86654 -39475
rect 86600 -39593 86610 -39559
rect 86644 -39593 86654 -39559
rect 86600 -39605 86654 -39593
rect 86684 -39491 86738 -39475
rect 86684 -39525 86694 -39491
rect 86728 -39525 86738 -39491
rect 86684 -39559 86738 -39525
rect 86684 -39593 86694 -39559
rect 86728 -39593 86738 -39559
rect 86684 -39605 86738 -39593
rect 86768 -39559 86822 -39475
rect 86768 -39593 86778 -39559
rect 86812 -39593 86822 -39559
rect 86768 -39605 86822 -39593
rect 86852 -39491 86906 -39475
rect 86852 -39525 86862 -39491
rect 86896 -39525 86906 -39491
rect 86852 -39559 86906 -39525
rect 86852 -39593 86862 -39559
rect 86896 -39593 86906 -39559
rect 86852 -39605 86906 -39593
rect 86936 -39559 86990 -39475
rect 86936 -39593 86946 -39559
rect 86980 -39593 86990 -39559
rect 86936 -39605 86990 -39593
rect 87020 -39491 87074 -39475
rect 87020 -39525 87030 -39491
rect 87064 -39525 87074 -39491
rect 87020 -39559 87074 -39525
rect 87020 -39593 87030 -39559
rect 87064 -39593 87074 -39559
rect 87020 -39605 87074 -39593
rect 87104 -39559 87158 -39475
rect 87104 -39593 87114 -39559
rect 87148 -39593 87158 -39559
rect 87104 -39605 87158 -39593
rect 87188 -39491 87242 -39475
rect 87188 -39525 87198 -39491
rect 87232 -39525 87242 -39491
rect 87188 -39559 87242 -39525
rect 87188 -39593 87198 -39559
rect 87232 -39593 87242 -39559
rect 87188 -39605 87242 -39593
rect 87272 -39491 87324 -39475
rect 87272 -39525 87282 -39491
rect 87316 -39525 87324 -39491
rect 87272 -39559 87324 -39525
rect 87272 -39593 87282 -39559
rect 87316 -39593 87324 -39559
rect 87272 -39605 87324 -39593
rect 87402 -39491 87454 -39475
rect 87402 -39525 87410 -39491
rect 87444 -39525 87454 -39491
rect 87402 -39559 87454 -39525
rect 87402 -39593 87410 -39559
rect 87444 -39593 87454 -39559
rect 87402 -39605 87454 -39593
rect 87484 -39491 87538 -39475
rect 87484 -39525 87494 -39491
rect 87528 -39525 87538 -39491
rect 87484 -39559 87538 -39525
rect 87484 -39593 87494 -39559
rect 87528 -39593 87538 -39559
rect 87484 -39605 87538 -39593
rect 87568 -39559 87622 -39475
rect 87568 -39593 87578 -39559
rect 87612 -39593 87622 -39559
rect 87568 -39605 87622 -39593
rect 87652 -39491 87706 -39475
rect 87652 -39525 87662 -39491
rect 87696 -39525 87706 -39491
rect 87652 -39559 87706 -39525
rect 87652 -39593 87662 -39559
rect 87696 -39593 87706 -39559
rect 87652 -39605 87706 -39593
rect 87736 -39559 87790 -39475
rect 87736 -39593 87746 -39559
rect 87780 -39593 87790 -39559
rect 87736 -39605 87790 -39593
rect 87820 -39491 87874 -39475
rect 87820 -39525 87830 -39491
rect 87864 -39525 87874 -39491
rect 87820 -39559 87874 -39525
rect 87820 -39593 87830 -39559
rect 87864 -39593 87874 -39559
rect 87820 -39605 87874 -39593
rect 87904 -39559 87958 -39475
rect 87904 -39593 87914 -39559
rect 87948 -39593 87958 -39559
rect 87904 -39605 87958 -39593
rect 87988 -39491 88042 -39475
rect 87988 -39525 87998 -39491
rect 88032 -39525 88042 -39491
rect 87988 -39559 88042 -39525
rect 87988 -39593 87998 -39559
rect 88032 -39593 88042 -39559
rect 87988 -39605 88042 -39593
rect 88072 -39559 88126 -39475
rect 88072 -39593 88082 -39559
rect 88116 -39593 88126 -39559
rect 88072 -39605 88126 -39593
rect 88156 -39491 88210 -39475
rect 88156 -39525 88166 -39491
rect 88200 -39525 88210 -39491
rect 88156 -39559 88210 -39525
rect 88156 -39593 88166 -39559
rect 88200 -39593 88210 -39559
rect 88156 -39605 88210 -39593
rect 88240 -39559 88294 -39475
rect 88240 -39593 88250 -39559
rect 88284 -39593 88294 -39559
rect 88240 -39605 88294 -39593
rect 88324 -39491 88378 -39475
rect 88324 -39525 88334 -39491
rect 88368 -39525 88378 -39491
rect 88324 -39559 88378 -39525
rect 88324 -39593 88334 -39559
rect 88368 -39593 88378 -39559
rect 88324 -39605 88378 -39593
rect 88408 -39559 88462 -39475
rect 88408 -39593 88418 -39559
rect 88452 -39593 88462 -39559
rect 88408 -39605 88462 -39593
rect 88492 -39491 88546 -39475
rect 88492 -39525 88502 -39491
rect 88536 -39525 88546 -39491
rect 88492 -39559 88546 -39525
rect 88492 -39593 88502 -39559
rect 88536 -39593 88546 -39559
rect 88492 -39605 88546 -39593
rect 88576 -39559 88630 -39475
rect 88576 -39593 88586 -39559
rect 88620 -39593 88630 -39559
rect 88576 -39605 88630 -39593
rect 88660 -39491 88714 -39475
rect 88660 -39525 88670 -39491
rect 88704 -39525 88714 -39491
rect 88660 -39559 88714 -39525
rect 88660 -39593 88670 -39559
rect 88704 -39593 88714 -39559
rect 88660 -39605 88714 -39593
rect 88744 -39491 88796 -39475
rect 88744 -39525 88754 -39491
rect 88788 -39525 88796 -39491
rect 88744 -39559 88796 -39525
rect 88744 -39593 88754 -39559
rect 88788 -39593 88796 -39559
rect 88744 -39605 88796 -39593
rect 53452 -39990 53510 -39978
rect 53452 -40766 53464 -39990
rect 53498 -40766 53510 -39990
rect 53452 -40778 53510 -40766
rect 53630 -39990 53688 -39978
rect 53630 -40766 53642 -39990
rect 53676 -40766 53688 -39990
rect 53630 -40778 53688 -40766
rect 55278 -40052 55336 -40040
rect 55278 -40228 55290 -40052
rect 55324 -40228 55336 -40052
rect 55278 -40240 55336 -40228
rect 55366 -40052 55424 -40040
rect 55366 -40228 55378 -40052
rect 55412 -40228 55424 -40052
rect 55366 -40240 55424 -40228
rect 53930 -40578 54730 -40566
rect 53930 -40612 53942 -40578
rect 54718 -40612 54730 -40578
rect 53930 -40624 54730 -40612
rect 53930 -40756 54730 -40744
rect 53930 -40790 53942 -40756
rect 54718 -40790 54730 -40756
rect 53930 -40802 54730 -40790
rect 55808 -39940 55866 -39928
rect 55808 -40716 55820 -39940
rect 55854 -40716 55866 -39940
rect 55808 -40728 55866 -40716
rect 55986 -39940 56044 -39928
rect 55986 -40716 55998 -39940
rect 56032 -40716 56044 -39940
rect 55986 -40728 56044 -40716
rect 77966 -39741 78019 -39735
rect 77605 -39771 77657 -39741
rect 77605 -39805 77613 -39771
rect 77647 -39805 77657 -39771
rect 77605 -39825 77657 -39805
rect 77687 -39765 77753 -39741
rect 77687 -39799 77703 -39765
rect 77737 -39799 77753 -39765
rect 77687 -39825 77753 -39799
rect 77783 -39751 77837 -39741
rect 77783 -39785 77793 -39751
rect 77827 -39785 77837 -39751
rect 77783 -39825 77837 -39785
rect 77867 -39765 77921 -39741
rect 77867 -39799 77877 -39765
rect 77911 -39799 77921 -39765
rect 77867 -39825 77921 -39799
rect 77951 -39751 78019 -39741
rect 77951 -39785 77971 -39751
rect 78005 -39785 78019 -39751
rect 77951 -39825 78019 -39785
rect 77966 -39865 78019 -39825
rect 78049 -39789 78103 -39735
rect 78049 -39823 78059 -39789
rect 78093 -39823 78103 -39789
rect 78049 -39865 78103 -39823
rect 80856 -39791 80908 -39775
rect 80856 -39825 80864 -39791
rect 80898 -39825 80908 -39791
rect 80856 -39859 80908 -39825
rect 80856 -39893 80864 -39859
rect 80898 -39893 80908 -39859
rect 80856 -39905 80908 -39893
rect 80938 -39791 80990 -39775
rect 80938 -39825 80948 -39791
rect 80982 -39825 80990 -39791
rect 80938 -39859 80990 -39825
rect 80938 -39893 80948 -39859
rect 80982 -39893 80990 -39859
rect 80938 -39905 80990 -39893
rect 57123 -40300 57175 -40255
rect 53452 -41008 53510 -40996
rect 53452 -41784 53464 -41008
rect 53498 -41784 53510 -41008
rect 53452 -41796 53510 -41784
rect 53630 -41008 53688 -40996
rect 53630 -41784 53642 -41008
rect 53676 -41784 53688 -41008
rect 53630 -41796 53688 -41784
rect 53930 -40984 54730 -40972
rect 53930 -41018 53942 -40984
rect 54718 -41018 54730 -40984
rect 53930 -41030 54730 -41018
rect 53930 -41162 54730 -41150
rect 53930 -41196 53942 -41162
rect 54718 -41196 54730 -41162
rect 53930 -41208 54730 -41196
rect 55268 -41548 55326 -41536
rect 55268 -41724 55280 -41548
rect 55314 -41724 55326 -41548
rect 55268 -41736 55326 -41724
rect 55356 -41548 55414 -41536
rect 55356 -41724 55368 -41548
rect 55402 -41724 55414 -41548
rect 55356 -41736 55414 -41724
rect 55808 -41054 55866 -41042
rect 55808 -41830 55820 -41054
rect 55854 -41830 55866 -41054
rect 55808 -41842 55866 -41830
rect 55986 -41054 56044 -41042
rect 55986 -41830 55998 -41054
rect 56032 -41830 56044 -41054
rect 55986 -41842 56044 -41830
rect 57123 -40334 57131 -40300
rect 57165 -40334 57175 -40300
rect 57123 -40359 57175 -40334
rect 57205 -40313 57263 -40255
rect 57205 -40347 57217 -40313
rect 57251 -40347 57263 -40313
rect 57205 -40359 57263 -40347
rect 57293 -40283 57345 -40255
rect 57293 -40317 57303 -40283
rect 57337 -40317 57345 -40283
rect 57293 -40359 57345 -40317
rect 59946 -40174 60346 -40162
rect 59946 -40208 59958 -40174
rect 60334 -40208 60346 -40174
rect 59946 -40220 60346 -40208
rect 59946 -40282 60346 -40270
rect 59946 -40316 59958 -40282
rect 60334 -40316 60346 -40282
rect 59946 -40328 60346 -40316
rect 59490 -40582 59548 -40570
rect 59490 -40650 59502 -40582
rect 59476 -40720 59502 -40650
rect 59490 -40758 59502 -40720
rect 59536 -40758 59548 -40582
rect 59490 -40770 59548 -40758
rect 59578 -40582 59636 -40570
rect 59578 -40758 59590 -40582
rect 59624 -40758 59636 -40582
rect 59578 -40770 59636 -40758
rect 59806 -40582 59864 -40570
rect 59806 -40758 59818 -40582
rect 59852 -40758 59864 -40582
rect 59806 -40770 59864 -40758
rect 59894 -40582 59952 -40570
rect 59894 -40758 59906 -40582
rect 59940 -40758 59952 -40582
rect 59894 -40770 59952 -40758
rect 77833 -40693 77885 -40675
rect 60191 -40773 60321 -40765
rect 60191 -40807 60203 -40773
rect 60237 -40807 60321 -40773
rect 60191 -40817 60321 -40807
rect 61131 -40773 61261 -40765
rect 61131 -40807 61215 -40773
rect 61249 -40807 61261 -40773
rect 61131 -40817 61261 -40807
rect 77637 -40731 77693 -40693
rect 77637 -40765 77649 -40731
rect 77683 -40765 77693 -40731
rect 77637 -40777 77693 -40765
rect 77723 -40777 77777 -40693
rect 77807 -40759 77885 -40693
rect 77807 -40777 77841 -40759
rect 77833 -40793 77841 -40777
rect 77875 -40793 77885 -40759
rect 77833 -40805 77885 -40793
rect 77915 -40759 77971 -40675
rect 77915 -40793 77925 -40759
rect 77959 -40793 77971 -40759
rect 77915 -40805 77971 -40793
rect 60191 -40857 60321 -40847
rect 60191 -40891 60211 -40857
rect 60245 -40891 60321 -40857
rect 60191 -40901 60321 -40891
rect 61131 -40857 61261 -40847
rect 61131 -40891 61207 -40857
rect 61241 -40891 61261 -40857
rect 61131 -40901 61261 -40891
rect 57123 -41454 57175 -41429
rect 57123 -41488 57131 -41454
rect 57165 -41488 57175 -41454
rect 57123 -41533 57175 -41488
rect 57205 -41441 57263 -41429
rect 57205 -41475 57217 -41441
rect 57251 -41475 57263 -41441
rect 57205 -41533 57263 -41475
rect 57293 -41471 57345 -41429
rect 57293 -41505 57303 -41471
rect 57337 -41505 57345 -41471
rect 57293 -41533 57345 -41505
rect 60191 -40941 60321 -40931
rect 59489 -41095 59547 -41083
rect 59489 -41271 59501 -41095
rect 59535 -41271 59547 -41095
rect 59489 -41283 59547 -41271
rect 59577 -41095 59635 -41083
rect 59577 -41271 59589 -41095
rect 59623 -41271 59635 -41095
rect 59577 -41283 59635 -41271
rect 60191 -40975 60203 -40941
rect 60237 -40975 60321 -40941
rect 60191 -40985 60321 -40975
rect 61131 -40941 61261 -40931
rect 61131 -40975 61215 -40941
rect 61249 -40975 61261 -40941
rect 61131 -40985 61261 -40975
rect 59805 -41095 59863 -41083
rect 59805 -41271 59817 -41095
rect 59851 -41271 59863 -41095
rect 59805 -41283 59863 -41271
rect 59893 -41095 59951 -41083
rect 59893 -41271 59905 -41095
rect 59939 -41271 59951 -41095
rect 59893 -41283 59951 -41271
rect 60191 -41025 60321 -41015
rect 60191 -41059 60211 -41025
rect 60245 -41059 60321 -41025
rect 60191 -41069 60321 -41059
rect 61131 -41025 61261 -41015
rect 61131 -41059 61207 -41025
rect 61241 -41059 61261 -41025
rect 61131 -41069 61261 -41059
rect 77833 -40987 77885 -40975
rect 77833 -41003 77841 -40987
rect 77637 -41015 77693 -41003
rect 77637 -41049 77649 -41015
rect 77683 -41049 77693 -41015
rect 77637 -41087 77693 -41049
rect 77723 -41087 77777 -41003
rect 77807 -41021 77841 -41003
rect 77875 -41021 77885 -40987
rect 77807 -41087 77885 -41021
rect 60191 -41109 60321 -41099
rect 60191 -41143 60204 -41109
rect 60238 -41143 60321 -41109
rect 60191 -41151 60321 -41143
rect 61131 -41109 61261 -41099
rect 61131 -41143 61214 -41109
rect 61248 -41143 61261 -41109
rect 61131 -41151 61261 -41143
rect 77833 -41105 77885 -41087
rect 77915 -40987 77971 -40975
rect 78426 -40981 78479 -40975
rect 77915 -41021 77925 -40987
rect 77959 -41021 77971 -40987
rect 77915 -41105 77971 -41021
rect 78065 -41011 78117 -40981
rect 78065 -41045 78073 -41011
rect 78107 -41045 78117 -41011
rect 78065 -41065 78117 -41045
rect 78147 -41005 78213 -40981
rect 78147 -41039 78163 -41005
rect 78197 -41039 78213 -41005
rect 78147 -41065 78213 -41039
rect 78243 -40991 78297 -40981
rect 78243 -41025 78253 -40991
rect 78287 -41025 78297 -40991
rect 78243 -41065 78297 -41025
rect 78327 -41005 78381 -40981
rect 78327 -41039 78337 -41005
rect 78371 -41039 78381 -41005
rect 78327 -41065 78381 -41039
rect 78411 -40991 78479 -40981
rect 78411 -41025 78431 -40991
rect 78465 -41025 78479 -40991
rect 78411 -41065 78479 -41025
rect 78426 -41105 78479 -41065
rect 78509 -41029 78563 -40975
rect 78509 -41063 78519 -41029
rect 78553 -41063 78563 -41029
rect 78509 -41105 78563 -41063
rect 59946 -41540 60346 -41528
rect 59946 -41574 59958 -41540
rect 60334 -41574 60346 -41540
rect 59946 -41586 60346 -41574
rect 59946 -41648 60346 -41636
rect 59946 -41682 59958 -41648
rect 60334 -41682 60346 -41648
rect 59946 -41694 60346 -41682
rect 77833 -41933 77885 -41915
rect 77637 -41971 77693 -41933
rect 77637 -42005 77649 -41971
rect 77683 -42005 77693 -41971
rect 77637 -42017 77693 -42005
rect 77723 -42017 77777 -41933
rect 77807 -41999 77885 -41933
rect 77807 -42017 77841 -41999
rect 77833 -42033 77841 -42017
rect 77875 -42033 77885 -41999
rect 77833 -42045 77885 -42033
rect 77915 -41999 77971 -41915
rect 77915 -42033 77925 -41999
rect 77959 -42033 77971 -41999
rect 77915 -42045 77971 -42033
rect 77835 -42241 77887 -42229
rect 77835 -42257 77843 -42241
rect 55288 -42358 55488 -42346
rect 55288 -42392 55300 -42358
rect 55476 -42392 55488 -42358
rect 55288 -42404 55488 -42392
rect 55288 -42446 55488 -42434
rect 55288 -42480 55300 -42446
rect 55476 -42480 55488 -42446
rect 55288 -42492 55488 -42480
rect 77639 -42269 77695 -42257
rect 77639 -42303 77651 -42269
rect 77685 -42303 77695 -42269
rect 77639 -42341 77695 -42303
rect 77725 -42341 77779 -42257
rect 77809 -42275 77843 -42257
rect 77877 -42275 77887 -42241
rect 77809 -42341 77887 -42275
rect 77835 -42359 77887 -42341
rect 77917 -42241 77973 -42229
rect 77917 -42275 77927 -42241
rect 77961 -42275 77973 -42241
rect 77917 -42359 77973 -42275
rect 78020 -43181 78113 -43165
rect 78020 -43211 78054 -43181
rect 77605 -43241 77657 -43211
rect 77605 -43275 77613 -43241
rect 77647 -43275 77657 -43241
rect 77605 -43295 77657 -43275
rect 77687 -43295 77745 -43211
rect 77775 -43295 77851 -43211
rect 77881 -43295 77947 -43211
rect 77977 -43215 78054 -43211
rect 78088 -43215 78113 -43181
rect 77977 -43249 78113 -43215
rect 77977 -43283 78054 -43249
rect 78088 -43283 78113 -43249
rect 77977 -43295 78113 -43283
rect 78143 -43181 78195 -43165
rect 78143 -43215 78153 -43181
rect 78187 -43215 78195 -43181
rect 78710 -43205 78763 -43165
rect 78143 -43249 78195 -43215
rect 78143 -43283 78153 -43249
rect 78187 -43283 78195 -43249
rect 78143 -43295 78195 -43283
rect 78349 -43225 78401 -43205
rect 78349 -43259 78357 -43225
rect 78391 -43259 78401 -43225
rect 78349 -43289 78401 -43259
rect 78431 -43231 78497 -43205
rect 78431 -43265 78447 -43231
rect 78481 -43265 78497 -43231
rect 78431 -43289 78497 -43265
rect 78527 -43245 78581 -43205
rect 78527 -43279 78537 -43245
rect 78571 -43279 78581 -43245
rect 78527 -43289 78581 -43279
rect 78611 -43231 78665 -43205
rect 78611 -43265 78621 -43231
rect 78655 -43265 78665 -43231
rect 78611 -43289 78665 -43265
rect 78695 -43245 78763 -43205
rect 78695 -43279 78715 -43245
rect 78749 -43279 78763 -43245
rect 78695 -43289 78763 -43279
rect 78710 -43295 78763 -43289
rect 78793 -43207 78847 -43165
rect 78793 -43241 78803 -43207
rect 78837 -43241 78847 -43207
rect 78793 -43295 78847 -43241
rect 77605 -43481 77657 -43461
rect 77605 -43515 77613 -43481
rect 77647 -43515 77657 -43481
rect 77605 -43545 77657 -43515
rect 77687 -43545 77745 -43461
rect 77775 -43545 77851 -43461
rect 77881 -43545 77947 -43461
rect 77977 -43473 78113 -43461
rect 77977 -43507 78054 -43473
rect 78088 -43507 78113 -43473
rect 77977 -43541 78113 -43507
rect 77977 -43545 78054 -43541
rect 78020 -43575 78054 -43545
rect 78088 -43575 78113 -43541
rect 78020 -43591 78113 -43575
rect 78143 -43473 78195 -43461
rect 78143 -43507 78153 -43473
rect 78187 -43507 78195 -43473
rect 78143 -43541 78195 -43507
rect 78143 -43575 78153 -43541
rect 78187 -43575 78195 -43541
rect 78143 -43591 78195 -43575
rect 83075 -44021 83127 -43975
rect 82894 -44049 82946 -44021
rect 82894 -44083 82902 -44049
rect 82936 -44083 82946 -44049
rect 82894 -44105 82946 -44083
rect 82976 -44049 83030 -44021
rect 82976 -44083 82986 -44049
rect 83020 -44083 83030 -44049
rect 82976 -44105 83030 -44083
rect 83060 -44049 83127 -44021
rect 83060 -44083 83082 -44049
rect 83116 -44083 83127 -44049
rect 83060 -44105 83127 -44083
rect 83157 -43989 83209 -43975
rect 83157 -44023 83167 -43989
rect 83201 -44023 83209 -43989
rect 83157 -44057 83209 -44023
rect 83157 -44091 83167 -44057
rect 83201 -44091 83209 -44057
rect 83157 -44105 83209 -44091
rect 83366 -43987 83418 -43975
rect 83366 -44021 83374 -43987
rect 83408 -44021 83418 -43987
rect 83366 -44055 83418 -44021
rect 83366 -44089 83374 -44055
rect 83408 -44089 83418 -44055
rect 83366 -44105 83418 -44089
rect 83448 -43987 83500 -43975
rect 83448 -44021 83458 -43987
rect 83492 -44021 83500 -43987
rect 83448 -44055 83500 -44021
rect 83448 -44089 83458 -44055
rect 83492 -44089 83500 -44055
rect 83448 -44105 83500 -44089
rect 83611 -44059 83663 -43975
rect 83611 -44093 83619 -44059
rect 83653 -44093 83663 -44059
rect 83611 -44105 83663 -44093
rect 83693 -44051 83747 -43975
rect 83693 -44085 83703 -44051
rect 83737 -44085 83747 -44051
rect 83693 -44105 83747 -44085
rect 83777 -44059 83831 -43975
rect 83777 -44093 83787 -44059
rect 83821 -44093 83831 -44059
rect 83777 -44105 83831 -44093
rect 83861 -44051 83915 -43975
rect 83861 -44085 83871 -44051
rect 83905 -44085 83915 -44051
rect 83861 -44105 83915 -44085
rect 83945 -44058 83997 -43975
rect 83945 -44092 83955 -44058
rect 83989 -44092 83997 -44058
rect 83945 -44105 83997 -44092
rect 84074 -43991 84126 -43975
rect 84074 -44025 84082 -43991
rect 84116 -44025 84126 -43991
rect 84074 -44059 84126 -44025
rect 84074 -44093 84082 -44059
rect 84116 -44093 84126 -44059
rect 84074 -44105 84126 -44093
rect 84156 -43991 84210 -43975
rect 84156 -44025 84166 -43991
rect 84200 -44025 84210 -43991
rect 84156 -44059 84210 -44025
rect 84156 -44093 84166 -44059
rect 84200 -44093 84210 -44059
rect 84156 -44105 84210 -44093
rect 84240 -44059 84294 -43975
rect 84240 -44093 84250 -44059
rect 84284 -44093 84294 -44059
rect 84240 -44105 84294 -44093
rect 84324 -43991 84378 -43975
rect 84324 -44025 84334 -43991
rect 84368 -44025 84378 -43991
rect 84324 -44059 84378 -44025
rect 84324 -44093 84334 -44059
rect 84368 -44093 84378 -44059
rect 84324 -44105 84378 -44093
rect 84408 -44059 84462 -43975
rect 84408 -44093 84418 -44059
rect 84452 -44093 84462 -44059
rect 84408 -44105 84462 -44093
rect 84492 -43991 84546 -43975
rect 84492 -44025 84502 -43991
rect 84536 -44025 84546 -43991
rect 84492 -44059 84546 -44025
rect 84492 -44093 84502 -44059
rect 84536 -44093 84546 -44059
rect 84492 -44105 84546 -44093
rect 84576 -44059 84630 -43975
rect 84576 -44093 84586 -44059
rect 84620 -44093 84630 -44059
rect 84576 -44105 84630 -44093
rect 84660 -43991 84714 -43975
rect 84660 -44025 84670 -43991
rect 84704 -44025 84714 -43991
rect 84660 -44059 84714 -44025
rect 84660 -44093 84670 -44059
rect 84704 -44093 84714 -44059
rect 84660 -44105 84714 -44093
rect 84744 -44059 84798 -43975
rect 84744 -44093 84754 -44059
rect 84788 -44093 84798 -44059
rect 84744 -44105 84798 -44093
rect 84828 -43991 84882 -43975
rect 84828 -44025 84838 -43991
rect 84872 -44025 84882 -43991
rect 84828 -44059 84882 -44025
rect 84828 -44093 84838 -44059
rect 84872 -44093 84882 -44059
rect 84828 -44105 84882 -44093
rect 84912 -44059 84966 -43975
rect 84912 -44093 84922 -44059
rect 84956 -44093 84966 -44059
rect 84912 -44105 84966 -44093
rect 84996 -43991 85050 -43975
rect 84996 -44025 85006 -43991
rect 85040 -44025 85050 -43991
rect 84996 -44059 85050 -44025
rect 84996 -44093 85006 -44059
rect 85040 -44093 85050 -44059
rect 84996 -44105 85050 -44093
rect 85080 -44059 85134 -43975
rect 85080 -44093 85090 -44059
rect 85124 -44093 85134 -44059
rect 85080 -44105 85134 -44093
rect 85164 -43991 85218 -43975
rect 85164 -44025 85174 -43991
rect 85208 -44025 85218 -43991
rect 85164 -44059 85218 -44025
rect 85164 -44093 85174 -44059
rect 85208 -44093 85218 -44059
rect 85164 -44105 85218 -44093
rect 85248 -44059 85302 -43975
rect 85248 -44093 85258 -44059
rect 85292 -44093 85302 -44059
rect 85248 -44105 85302 -44093
rect 85332 -43991 85386 -43975
rect 85332 -44025 85342 -43991
rect 85376 -44025 85386 -43991
rect 85332 -44059 85386 -44025
rect 85332 -44093 85342 -44059
rect 85376 -44093 85386 -44059
rect 85332 -44105 85386 -44093
rect 85416 -43991 85468 -43975
rect 85416 -44025 85426 -43991
rect 85460 -44025 85468 -43991
rect 85416 -44059 85468 -44025
rect 85416 -44093 85426 -44059
rect 85460 -44093 85468 -44059
rect 85416 -44105 85468 -44093
rect 85546 -43991 85598 -43975
rect 85546 -44025 85554 -43991
rect 85588 -44025 85598 -43991
rect 85546 -44059 85598 -44025
rect 85546 -44093 85554 -44059
rect 85588 -44093 85598 -44059
rect 85546 -44105 85598 -44093
rect 85628 -43991 85682 -43975
rect 85628 -44025 85638 -43991
rect 85672 -44025 85682 -43991
rect 85628 -44059 85682 -44025
rect 85628 -44093 85638 -44059
rect 85672 -44093 85682 -44059
rect 85628 -44105 85682 -44093
rect 85712 -44059 85766 -43975
rect 85712 -44093 85722 -44059
rect 85756 -44093 85766 -44059
rect 85712 -44105 85766 -44093
rect 85796 -43991 85850 -43975
rect 85796 -44025 85806 -43991
rect 85840 -44025 85850 -43991
rect 85796 -44059 85850 -44025
rect 85796 -44093 85806 -44059
rect 85840 -44093 85850 -44059
rect 85796 -44105 85850 -44093
rect 85880 -44059 85934 -43975
rect 85880 -44093 85890 -44059
rect 85924 -44093 85934 -44059
rect 85880 -44105 85934 -44093
rect 85964 -43991 86018 -43975
rect 85964 -44025 85974 -43991
rect 86008 -44025 86018 -43991
rect 85964 -44059 86018 -44025
rect 85964 -44093 85974 -44059
rect 86008 -44093 86018 -44059
rect 85964 -44105 86018 -44093
rect 86048 -44059 86102 -43975
rect 86048 -44093 86058 -44059
rect 86092 -44093 86102 -44059
rect 86048 -44105 86102 -44093
rect 86132 -43991 86186 -43975
rect 86132 -44025 86142 -43991
rect 86176 -44025 86186 -43991
rect 86132 -44059 86186 -44025
rect 86132 -44093 86142 -44059
rect 86176 -44093 86186 -44059
rect 86132 -44105 86186 -44093
rect 86216 -44059 86270 -43975
rect 86216 -44093 86226 -44059
rect 86260 -44093 86270 -44059
rect 86216 -44105 86270 -44093
rect 86300 -43991 86354 -43975
rect 86300 -44025 86310 -43991
rect 86344 -44025 86354 -43991
rect 86300 -44059 86354 -44025
rect 86300 -44093 86310 -44059
rect 86344 -44093 86354 -44059
rect 86300 -44105 86354 -44093
rect 86384 -44059 86438 -43975
rect 86384 -44093 86394 -44059
rect 86428 -44093 86438 -44059
rect 86384 -44105 86438 -44093
rect 86468 -43991 86522 -43975
rect 86468 -44025 86478 -43991
rect 86512 -44025 86522 -43991
rect 86468 -44059 86522 -44025
rect 86468 -44093 86478 -44059
rect 86512 -44093 86522 -44059
rect 86468 -44105 86522 -44093
rect 86552 -44059 86606 -43975
rect 86552 -44093 86562 -44059
rect 86596 -44093 86606 -44059
rect 86552 -44105 86606 -44093
rect 86636 -43991 86690 -43975
rect 86636 -44025 86646 -43991
rect 86680 -44025 86690 -43991
rect 86636 -44059 86690 -44025
rect 86636 -44093 86646 -44059
rect 86680 -44093 86690 -44059
rect 86636 -44105 86690 -44093
rect 86720 -44059 86774 -43975
rect 86720 -44093 86730 -44059
rect 86764 -44093 86774 -44059
rect 86720 -44105 86774 -44093
rect 86804 -43991 86858 -43975
rect 86804 -44025 86814 -43991
rect 86848 -44025 86858 -43991
rect 86804 -44059 86858 -44025
rect 86804 -44093 86814 -44059
rect 86848 -44093 86858 -44059
rect 86804 -44105 86858 -44093
rect 86888 -43991 86940 -43975
rect 86888 -44025 86898 -43991
rect 86932 -44025 86940 -43991
rect 86888 -44059 86940 -44025
rect 86888 -44093 86898 -44059
rect 86932 -44093 86940 -44059
rect 86888 -44105 86940 -44093
rect 87018 -43991 87070 -43975
rect 87018 -44025 87026 -43991
rect 87060 -44025 87070 -43991
rect 87018 -44059 87070 -44025
rect 87018 -44093 87026 -44059
rect 87060 -44093 87070 -44059
rect 87018 -44105 87070 -44093
rect 87100 -43991 87154 -43975
rect 87100 -44025 87110 -43991
rect 87144 -44025 87154 -43991
rect 87100 -44059 87154 -44025
rect 87100 -44093 87110 -44059
rect 87144 -44093 87154 -44059
rect 87100 -44105 87154 -44093
rect 87184 -44059 87238 -43975
rect 87184 -44093 87194 -44059
rect 87228 -44093 87238 -44059
rect 87184 -44105 87238 -44093
rect 87268 -43991 87322 -43975
rect 87268 -44025 87278 -43991
rect 87312 -44025 87322 -43991
rect 87268 -44059 87322 -44025
rect 87268 -44093 87278 -44059
rect 87312 -44093 87322 -44059
rect 87268 -44105 87322 -44093
rect 87352 -44059 87406 -43975
rect 87352 -44093 87362 -44059
rect 87396 -44093 87406 -44059
rect 87352 -44105 87406 -44093
rect 87436 -43991 87490 -43975
rect 87436 -44025 87446 -43991
rect 87480 -44025 87490 -43991
rect 87436 -44059 87490 -44025
rect 87436 -44093 87446 -44059
rect 87480 -44093 87490 -44059
rect 87436 -44105 87490 -44093
rect 87520 -44059 87574 -43975
rect 87520 -44093 87530 -44059
rect 87564 -44093 87574 -44059
rect 87520 -44105 87574 -44093
rect 87604 -43991 87658 -43975
rect 87604 -44025 87614 -43991
rect 87648 -44025 87658 -43991
rect 87604 -44059 87658 -44025
rect 87604 -44093 87614 -44059
rect 87648 -44093 87658 -44059
rect 87604 -44105 87658 -44093
rect 87688 -44059 87742 -43975
rect 87688 -44093 87698 -44059
rect 87732 -44093 87742 -44059
rect 87688 -44105 87742 -44093
rect 87772 -43991 87826 -43975
rect 87772 -44025 87782 -43991
rect 87816 -44025 87826 -43991
rect 87772 -44059 87826 -44025
rect 87772 -44093 87782 -44059
rect 87816 -44093 87826 -44059
rect 87772 -44105 87826 -44093
rect 87856 -44059 87910 -43975
rect 87856 -44093 87866 -44059
rect 87900 -44093 87910 -44059
rect 87856 -44105 87910 -44093
rect 87940 -43991 87994 -43975
rect 87940 -44025 87950 -43991
rect 87984 -44025 87994 -43991
rect 87940 -44059 87994 -44025
rect 87940 -44093 87950 -44059
rect 87984 -44093 87994 -44059
rect 87940 -44105 87994 -44093
rect 88024 -44059 88078 -43975
rect 88024 -44093 88034 -44059
rect 88068 -44093 88078 -44059
rect 88024 -44105 88078 -44093
rect 88108 -43991 88162 -43975
rect 88108 -44025 88118 -43991
rect 88152 -44025 88162 -43991
rect 88108 -44059 88162 -44025
rect 88108 -44093 88118 -44059
rect 88152 -44093 88162 -44059
rect 88108 -44105 88162 -44093
rect 88192 -44059 88246 -43975
rect 88192 -44093 88202 -44059
rect 88236 -44093 88246 -44059
rect 88192 -44105 88246 -44093
rect 88276 -43991 88330 -43975
rect 88276 -44025 88286 -43991
rect 88320 -44025 88330 -43991
rect 88276 -44059 88330 -44025
rect 88276 -44093 88286 -44059
rect 88320 -44093 88330 -44059
rect 88276 -44105 88330 -44093
rect 88360 -43991 88412 -43975
rect 88360 -44025 88370 -43991
rect 88404 -44025 88412 -43991
rect 88360 -44059 88412 -44025
rect 88360 -44093 88370 -44059
rect 88404 -44093 88412 -44059
rect 88360 -44105 88412 -44093
rect 88490 -43991 88542 -43975
rect 88490 -44025 88498 -43991
rect 88532 -44025 88542 -43991
rect 88490 -44059 88542 -44025
rect 88490 -44093 88498 -44059
rect 88532 -44093 88542 -44059
rect 88490 -44105 88542 -44093
rect 88572 -43991 88626 -43975
rect 88572 -44025 88582 -43991
rect 88616 -44025 88626 -43991
rect 88572 -44059 88626 -44025
rect 88572 -44093 88582 -44059
rect 88616 -44093 88626 -44059
rect 88572 -44105 88626 -44093
rect 88656 -44059 88710 -43975
rect 88656 -44093 88666 -44059
rect 88700 -44093 88710 -44059
rect 88656 -44105 88710 -44093
rect 88740 -43991 88794 -43975
rect 88740 -44025 88750 -43991
rect 88784 -44025 88794 -43991
rect 88740 -44059 88794 -44025
rect 88740 -44093 88750 -44059
rect 88784 -44093 88794 -44059
rect 88740 -44105 88794 -44093
rect 88824 -44059 88878 -43975
rect 88824 -44093 88834 -44059
rect 88868 -44093 88878 -44059
rect 88824 -44105 88878 -44093
rect 88908 -43991 88962 -43975
rect 88908 -44025 88918 -43991
rect 88952 -44025 88962 -43991
rect 88908 -44059 88962 -44025
rect 88908 -44093 88918 -44059
rect 88952 -44093 88962 -44059
rect 88908 -44105 88962 -44093
rect 88992 -44059 89046 -43975
rect 88992 -44093 89002 -44059
rect 89036 -44093 89046 -44059
rect 88992 -44105 89046 -44093
rect 89076 -43991 89130 -43975
rect 89076 -44025 89086 -43991
rect 89120 -44025 89130 -43991
rect 89076 -44059 89130 -44025
rect 89076 -44093 89086 -44059
rect 89120 -44093 89130 -44059
rect 89076 -44105 89130 -44093
rect 89160 -44059 89214 -43975
rect 89160 -44093 89170 -44059
rect 89204 -44093 89214 -44059
rect 89160 -44105 89214 -44093
rect 89244 -43991 89298 -43975
rect 89244 -44025 89254 -43991
rect 89288 -44025 89298 -43991
rect 89244 -44059 89298 -44025
rect 89244 -44093 89254 -44059
rect 89288 -44093 89298 -44059
rect 89244 -44105 89298 -44093
rect 89328 -44059 89382 -43975
rect 89328 -44093 89338 -44059
rect 89372 -44093 89382 -44059
rect 89328 -44105 89382 -44093
rect 89412 -43991 89466 -43975
rect 89412 -44025 89422 -43991
rect 89456 -44025 89466 -43991
rect 89412 -44059 89466 -44025
rect 89412 -44093 89422 -44059
rect 89456 -44093 89466 -44059
rect 89412 -44105 89466 -44093
rect 89496 -44059 89550 -43975
rect 89496 -44093 89506 -44059
rect 89540 -44093 89550 -44059
rect 89496 -44105 89550 -44093
rect 89580 -43991 89634 -43975
rect 89580 -44025 89590 -43991
rect 89624 -44025 89634 -43991
rect 89580 -44059 89634 -44025
rect 89580 -44093 89590 -44059
rect 89624 -44093 89634 -44059
rect 89580 -44105 89634 -44093
rect 89664 -44059 89718 -43975
rect 89664 -44093 89674 -44059
rect 89708 -44093 89718 -44059
rect 89664 -44105 89718 -44093
rect 89748 -43991 89802 -43975
rect 89748 -44025 89758 -43991
rect 89792 -44025 89802 -43991
rect 89748 -44059 89802 -44025
rect 89748 -44093 89758 -44059
rect 89792 -44093 89802 -44059
rect 89748 -44105 89802 -44093
rect 89832 -43991 89884 -43975
rect 89832 -44025 89842 -43991
rect 89876 -44025 89884 -43991
rect 89832 -44059 89884 -44025
rect 89832 -44093 89842 -44059
rect 89876 -44093 89884 -44059
rect 89832 -44105 89884 -44093
rect 89962 -43991 90014 -43975
rect 89962 -44025 89970 -43991
rect 90004 -44025 90014 -43991
rect 89962 -44059 90014 -44025
rect 89962 -44093 89970 -44059
rect 90004 -44093 90014 -44059
rect 89962 -44105 90014 -44093
rect 90044 -43991 90098 -43975
rect 90044 -44025 90054 -43991
rect 90088 -44025 90098 -43991
rect 90044 -44059 90098 -44025
rect 90044 -44093 90054 -44059
rect 90088 -44093 90098 -44059
rect 90044 -44105 90098 -44093
rect 90128 -44059 90182 -43975
rect 90128 -44093 90138 -44059
rect 90172 -44093 90182 -44059
rect 90128 -44105 90182 -44093
rect 90212 -43991 90266 -43975
rect 90212 -44025 90222 -43991
rect 90256 -44025 90266 -43991
rect 90212 -44059 90266 -44025
rect 90212 -44093 90222 -44059
rect 90256 -44093 90266 -44059
rect 90212 -44105 90266 -44093
rect 90296 -44059 90350 -43975
rect 90296 -44093 90306 -44059
rect 90340 -44093 90350 -44059
rect 90296 -44105 90350 -44093
rect 90380 -43991 90434 -43975
rect 90380 -44025 90390 -43991
rect 90424 -44025 90434 -43991
rect 90380 -44059 90434 -44025
rect 90380 -44093 90390 -44059
rect 90424 -44093 90434 -44059
rect 90380 -44105 90434 -44093
rect 90464 -44059 90518 -43975
rect 90464 -44093 90474 -44059
rect 90508 -44093 90518 -44059
rect 90464 -44105 90518 -44093
rect 90548 -43991 90602 -43975
rect 90548 -44025 90558 -43991
rect 90592 -44025 90602 -43991
rect 90548 -44059 90602 -44025
rect 90548 -44093 90558 -44059
rect 90592 -44093 90602 -44059
rect 90548 -44105 90602 -44093
rect 90632 -44059 90686 -43975
rect 90632 -44093 90642 -44059
rect 90676 -44093 90686 -44059
rect 90632 -44105 90686 -44093
rect 90716 -43991 90770 -43975
rect 90716 -44025 90726 -43991
rect 90760 -44025 90770 -43991
rect 90716 -44059 90770 -44025
rect 90716 -44093 90726 -44059
rect 90760 -44093 90770 -44059
rect 90716 -44105 90770 -44093
rect 90800 -44059 90854 -43975
rect 90800 -44093 90810 -44059
rect 90844 -44093 90854 -44059
rect 90800 -44105 90854 -44093
rect 90884 -43991 90938 -43975
rect 90884 -44025 90894 -43991
rect 90928 -44025 90938 -43991
rect 90884 -44059 90938 -44025
rect 90884 -44093 90894 -44059
rect 90928 -44093 90938 -44059
rect 90884 -44105 90938 -44093
rect 90968 -44059 91022 -43975
rect 90968 -44093 90978 -44059
rect 91012 -44093 91022 -44059
rect 90968 -44105 91022 -44093
rect 91052 -43991 91106 -43975
rect 91052 -44025 91062 -43991
rect 91096 -44025 91106 -43991
rect 91052 -44059 91106 -44025
rect 91052 -44093 91062 -44059
rect 91096 -44093 91106 -44059
rect 91052 -44105 91106 -44093
rect 91136 -44059 91190 -43975
rect 91136 -44093 91146 -44059
rect 91180 -44093 91190 -44059
rect 91136 -44105 91190 -44093
rect 91220 -43991 91274 -43975
rect 91220 -44025 91230 -43991
rect 91264 -44025 91274 -43991
rect 91220 -44059 91274 -44025
rect 91220 -44093 91230 -44059
rect 91264 -44093 91274 -44059
rect 91220 -44105 91274 -44093
rect 91304 -43991 91356 -43975
rect 91304 -44025 91314 -43991
rect 91348 -44025 91356 -43991
rect 91304 -44059 91356 -44025
rect 91304 -44093 91314 -44059
rect 91348 -44093 91356 -44059
rect 91304 -44105 91356 -44093
rect 78020 -44413 78113 -44397
rect 78020 -44443 78054 -44413
rect 77605 -44473 77657 -44443
rect 77605 -44507 77613 -44473
rect 77647 -44507 77657 -44473
rect 77605 -44527 77657 -44507
rect 77687 -44527 77745 -44443
rect 77775 -44527 77851 -44443
rect 77881 -44527 77947 -44443
rect 77977 -44447 78054 -44443
rect 78088 -44447 78113 -44413
rect 77977 -44481 78113 -44447
rect 77977 -44515 78054 -44481
rect 78088 -44515 78113 -44481
rect 77977 -44527 78113 -44515
rect 78143 -44413 78195 -44397
rect 78143 -44447 78153 -44413
rect 78187 -44447 78195 -44413
rect 78143 -44481 78195 -44447
rect 78143 -44515 78153 -44481
rect 78187 -44515 78195 -44481
rect 78143 -44527 78195 -44515
rect 77605 -44715 77657 -44695
rect 77605 -44749 77613 -44715
rect 77647 -44749 77657 -44715
rect 77605 -44779 77657 -44749
rect 77687 -44779 77745 -44695
rect 77775 -44779 77851 -44695
rect 77881 -44779 77947 -44695
rect 77977 -44707 78113 -44695
rect 77977 -44741 78054 -44707
rect 78088 -44741 78113 -44707
rect 77977 -44775 78113 -44741
rect 77977 -44779 78054 -44775
rect 78020 -44809 78054 -44779
rect 78088 -44809 78113 -44775
rect 78020 -44825 78113 -44809
rect 78143 -44707 78195 -44695
rect 78143 -44741 78153 -44707
rect 78187 -44741 78195 -44707
rect 78143 -44775 78195 -44741
rect 78143 -44809 78153 -44775
rect 78187 -44809 78195 -44775
rect 78143 -44825 78195 -44809
rect 53452 -45390 53510 -45378
rect 53452 -46166 53464 -45390
rect 53498 -46166 53510 -45390
rect 53452 -46178 53510 -46166
rect 53630 -45390 53688 -45378
rect 53630 -46166 53642 -45390
rect 53676 -46166 53688 -45390
rect 53630 -46178 53688 -46166
rect 55278 -45452 55336 -45440
rect 55278 -45628 55290 -45452
rect 55324 -45628 55336 -45452
rect 55278 -45640 55336 -45628
rect 55366 -45452 55424 -45440
rect 55366 -45628 55378 -45452
rect 55412 -45628 55424 -45452
rect 55366 -45640 55424 -45628
rect 53930 -45978 54730 -45966
rect 53930 -46012 53942 -45978
rect 54718 -46012 54730 -45978
rect 53930 -46024 54730 -46012
rect 53930 -46156 54730 -46144
rect 53930 -46190 53942 -46156
rect 54718 -46190 54730 -46156
rect 53930 -46202 54730 -46190
rect 55808 -45340 55866 -45328
rect 55808 -46116 55820 -45340
rect 55854 -46116 55866 -45340
rect 55808 -46128 55866 -46116
rect 55986 -45340 56044 -45328
rect 55986 -46116 55998 -45340
rect 56032 -46116 56044 -45340
rect 55986 -46128 56044 -46116
rect 57123 -45700 57175 -45655
rect 53452 -46408 53510 -46396
rect 53452 -47184 53464 -46408
rect 53498 -47184 53510 -46408
rect 53452 -47196 53510 -47184
rect 53630 -46408 53688 -46396
rect 53630 -47184 53642 -46408
rect 53676 -47184 53688 -46408
rect 53630 -47196 53688 -47184
rect 53930 -46384 54730 -46372
rect 53930 -46418 53942 -46384
rect 54718 -46418 54730 -46384
rect 53930 -46430 54730 -46418
rect 53930 -46562 54730 -46550
rect 53930 -46596 53942 -46562
rect 54718 -46596 54730 -46562
rect 53930 -46608 54730 -46596
rect 55268 -46948 55326 -46936
rect 55268 -47124 55280 -46948
rect 55314 -47124 55326 -46948
rect 55268 -47136 55326 -47124
rect 55356 -46948 55414 -46936
rect 55356 -47124 55368 -46948
rect 55402 -47124 55414 -46948
rect 55356 -47136 55414 -47124
rect 55808 -46454 55866 -46442
rect 55808 -47230 55820 -46454
rect 55854 -47230 55866 -46454
rect 55808 -47242 55866 -47230
rect 55986 -46454 56044 -46442
rect 55986 -47230 55998 -46454
rect 56032 -47230 56044 -46454
rect 55986 -47242 56044 -47230
rect 57123 -45734 57131 -45700
rect 57165 -45734 57175 -45700
rect 57123 -45759 57175 -45734
rect 57205 -45713 57263 -45655
rect 57205 -45747 57217 -45713
rect 57251 -45747 57263 -45713
rect 57205 -45759 57263 -45747
rect 57293 -45683 57345 -45655
rect 57293 -45717 57303 -45683
rect 57337 -45717 57345 -45683
rect 57293 -45759 57345 -45717
rect 59946 -45574 60346 -45562
rect 59946 -45608 59958 -45574
rect 60334 -45608 60346 -45574
rect 59946 -45620 60346 -45608
rect 59946 -45682 60346 -45670
rect 59946 -45716 59958 -45682
rect 60334 -45716 60346 -45682
rect 59946 -45728 60346 -45716
rect 77879 -45681 77929 -45635
rect 77605 -45719 77657 -45681
rect 77605 -45753 77613 -45719
rect 77647 -45753 77657 -45719
rect 77605 -45765 77657 -45753
rect 77687 -45765 77729 -45681
rect 77759 -45765 77801 -45681
rect 77831 -45703 77929 -45681
rect 77831 -45737 77885 -45703
rect 77919 -45737 77929 -45703
rect 77831 -45765 77929 -45737
rect 77959 -45693 78011 -45635
rect 78293 -45653 78345 -45635
rect 77959 -45727 77969 -45693
rect 78003 -45727 78011 -45693
rect 77959 -45765 78011 -45727
rect 78097 -45691 78153 -45653
rect 78097 -45725 78109 -45691
rect 78143 -45725 78153 -45691
rect 78097 -45737 78153 -45725
rect 78183 -45737 78237 -45653
rect 78267 -45719 78345 -45653
rect 78267 -45737 78301 -45719
rect 78293 -45753 78301 -45737
rect 78335 -45753 78345 -45719
rect 78293 -45765 78345 -45753
rect 78375 -45719 78431 -45635
rect 78886 -45675 78939 -45635
rect 78375 -45753 78385 -45719
rect 78419 -45753 78431 -45719
rect 78375 -45765 78431 -45753
rect 78525 -45695 78577 -45675
rect 78525 -45729 78533 -45695
rect 78567 -45729 78577 -45695
rect 78525 -45759 78577 -45729
rect 78607 -45701 78673 -45675
rect 78607 -45735 78623 -45701
rect 78657 -45735 78673 -45701
rect 78607 -45759 78673 -45735
rect 78703 -45715 78757 -45675
rect 78703 -45749 78713 -45715
rect 78747 -45749 78757 -45715
rect 78703 -45759 78757 -45749
rect 78787 -45701 78841 -45675
rect 78787 -45735 78797 -45701
rect 78831 -45735 78841 -45701
rect 78787 -45759 78841 -45735
rect 78871 -45715 78939 -45675
rect 78871 -45749 78891 -45715
rect 78925 -45749 78939 -45715
rect 78871 -45759 78939 -45749
rect 78886 -45765 78939 -45759
rect 78969 -45677 79023 -45635
rect 78969 -45711 78979 -45677
rect 79013 -45711 79023 -45677
rect 78969 -45765 79023 -45711
rect 59490 -45982 59548 -45970
rect 59490 -46050 59502 -45982
rect 59476 -46120 59502 -46050
rect 59490 -46158 59502 -46120
rect 59536 -46158 59548 -45982
rect 59490 -46170 59548 -46158
rect 59578 -45982 59636 -45970
rect 59578 -46158 59590 -45982
rect 59624 -46158 59636 -45982
rect 59578 -46170 59636 -46158
rect 59806 -45982 59864 -45970
rect 59806 -46158 59818 -45982
rect 59852 -46158 59864 -45982
rect 59806 -46170 59864 -46158
rect 59894 -45982 59952 -45970
rect 59894 -46158 59906 -45982
rect 59940 -46158 59952 -45982
rect 59894 -46170 59952 -46158
rect 60191 -46173 60321 -46165
rect 60191 -46207 60203 -46173
rect 60237 -46207 60321 -46173
rect 60191 -46217 60321 -46207
rect 61131 -46173 61261 -46165
rect 61131 -46207 61215 -46173
rect 61249 -46207 61261 -46173
rect 61131 -46217 61261 -46207
rect 60191 -46257 60321 -46247
rect 60191 -46291 60211 -46257
rect 60245 -46291 60321 -46257
rect 60191 -46301 60321 -46291
rect 61131 -46257 61261 -46247
rect 61131 -46291 61207 -46257
rect 61241 -46291 61261 -46257
rect 61131 -46301 61261 -46291
rect 57123 -46854 57175 -46829
rect 57123 -46888 57131 -46854
rect 57165 -46888 57175 -46854
rect 57123 -46933 57175 -46888
rect 57205 -46841 57263 -46829
rect 57205 -46875 57217 -46841
rect 57251 -46875 57263 -46841
rect 57205 -46933 57263 -46875
rect 57293 -46871 57345 -46829
rect 57293 -46905 57303 -46871
rect 57337 -46905 57345 -46871
rect 57293 -46933 57345 -46905
rect 60191 -46341 60321 -46331
rect 59489 -46495 59547 -46483
rect 59489 -46671 59501 -46495
rect 59535 -46671 59547 -46495
rect 59489 -46683 59547 -46671
rect 59577 -46495 59635 -46483
rect 59577 -46671 59589 -46495
rect 59623 -46671 59635 -46495
rect 59577 -46683 59635 -46671
rect 60191 -46375 60203 -46341
rect 60237 -46375 60321 -46341
rect 60191 -46385 60321 -46375
rect 61131 -46341 61261 -46331
rect 61131 -46375 61215 -46341
rect 61249 -46375 61261 -46341
rect 61131 -46385 61261 -46375
rect 59805 -46495 59863 -46483
rect 59805 -46671 59817 -46495
rect 59851 -46671 59863 -46495
rect 59805 -46683 59863 -46671
rect 59893 -46495 59951 -46483
rect 59893 -46671 59905 -46495
rect 59939 -46671 59951 -46495
rect 59893 -46683 59951 -46671
rect 60191 -46425 60321 -46415
rect 60191 -46459 60211 -46425
rect 60245 -46459 60321 -46425
rect 60191 -46469 60321 -46459
rect 61131 -46425 61261 -46415
rect 61131 -46459 61207 -46425
rect 61241 -46459 61261 -46425
rect 61131 -46469 61261 -46459
rect 75574 -46491 75626 -46475
rect 60191 -46509 60321 -46499
rect 60191 -46543 60204 -46509
rect 60238 -46543 60321 -46509
rect 60191 -46551 60321 -46543
rect 61131 -46509 61261 -46499
rect 61131 -46543 61214 -46509
rect 61248 -46543 61261 -46509
rect 61131 -46551 61261 -46543
rect 75574 -46525 75582 -46491
rect 75616 -46525 75626 -46491
rect 75574 -46559 75626 -46525
rect 75574 -46593 75582 -46559
rect 75616 -46593 75626 -46559
rect 75574 -46605 75626 -46593
rect 75656 -46491 75708 -46475
rect 75656 -46525 75666 -46491
rect 75700 -46525 75708 -46491
rect 75656 -46559 75708 -46525
rect 75656 -46593 75666 -46559
rect 75700 -46593 75708 -46559
rect 75656 -46605 75708 -46593
rect 75850 -46491 75902 -46475
rect 75850 -46525 75858 -46491
rect 75892 -46525 75902 -46491
rect 75850 -46559 75902 -46525
rect 75850 -46593 75858 -46559
rect 75892 -46593 75902 -46559
rect 75850 -46605 75902 -46593
rect 75932 -46491 75984 -46475
rect 75932 -46525 75942 -46491
rect 75976 -46525 75984 -46491
rect 75932 -46559 75984 -46525
rect 75932 -46593 75942 -46559
rect 75976 -46593 75984 -46559
rect 75932 -46605 75984 -46593
rect 76124 -46491 76176 -46475
rect 76124 -46525 76132 -46491
rect 76166 -46525 76176 -46491
rect 76124 -46559 76176 -46525
rect 76124 -46593 76132 -46559
rect 76166 -46593 76176 -46559
rect 76124 -46605 76176 -46593
rect 76206 -46491 76258 -46475
rect 76206 -46525 76216 -46491
rect 76250 -46525 76258 -46491
rect 76206 -46559 76258 -46525
rect 76206 -46593 76216 -46559
rect 76250 -46593 76258 -46559
rect 76206 -46605 76258 -46593
rect 76400 -46491 76452 -46475
rect 76400 -46525 76408 -46491
rect 76442 -46525 76452 -46491
rect 76400 -46559 76452 -46525
rect 76400 -46593 76408 -46559
rect 76442 -46593 76452 -46559
rect 76400 -46605 76452 -46593
rect 76482 -46491 76534 -46475
rect 76482 -46525 76492 -46491
rect 76526 -46525 76534 -46491
rect 76482 -46559 76534 -46525
rect 76482 -46593 76492 -46559
rect 76526 -46593 76534 -46559
rect 76482 -46605 76534 -46593
rect 76676 -46491 76728 -46475
rect 76676 -46525 76684 -46491
rect 76718 -46525 76728 -46491
rect 76676 -46559 76728 -46525
rect 76676 -46593 76684 -46559
rect 76718 -46593 76728 -46559
rect 76676 -46605 76728 -46593
rect 76758 -46491 76810 -46475
rect 76758 -46525 76768 -46491
rect 76802 -46525 76810 -46491
rect 76758 -46559 76810 -46525
rect 76758 -46593 76768 -46559
rect 76802 -46593 76810 -46559
rect 76758 -46605 76810 -46593
rect 59946 -46940 60346 -46928
rect 59946 -46974 59958 -46940
rect 60334 -46974 60346 -46940
rect 59946 -46986 60346 -46974
rect 59946 -47048 60346 -47036
rect 59946 -47082 59958 -47048
rect 60334 -47082 60346 -47048
rect 59946 -47094 60346 -47082
rect 77966 -47505 78019 -47465
rect 77605 -47525 77657 -47505
rect 77605 -47559 77613 -47525
rect 77647 -47559 77657 -47525
rect 77605 -47589 77657 -47559
rect 77687 -47531 77753 -47505
rect 77687 -47565 77703 -47531
rect 77737 -47565 77753 -47531
rect 77687 -47589 77753 -47565
rect 77783 -47545 77837 -47505
rect 77783 -47579 77793 -47545
rect 77827 -47579 77837 -47545
rect 77783 -47589 77837 -47579
rect 77867 -47531 77921 -47505
rect 77867 -47565 77877 -47531
rect 77911 -47565 77921 -47531
rect 77867 -47589 77921 -47565
rect 77951 -47545 78019 -47505
rect 77951 -47579 77971 -47545
rect 78005 -47579 78019 -47545
rect 77951 -47589 78019 -47579
rect 77966 -47595 78019 -47589
rect 78049 -47507 78103 -47465
rect 78424 -47505 78477 -47465
rect 78049 -47541 78059 -47507
rect 78093 -47541 78103 -47507
rect 78049 -47595 78103 -47541
rect 78159 -47531 78211 -47505
rect 78159 -47565 78167 -47531
rect 78201 -47565 78211 -47531
rect 78159 -47589 78211 -47565
rect 78241 -47545 78295 -47505
rect 78241 -47579 78251 -47545
rect 78285 -47579 78295 -47545
rect 78241 -47589 78295 -47579
rect 78325 -47531 78379 -47505
rect 78325 -47565 78335 -47531
rect 78369 -47565 78379 -47531
rect 78325 -47589 78379 -47565
rect 78409 -47545 78477 -47505
rect 78409 -47579 78429 -47545
rect 78463 -47579 78477 -47545
rect 78409 -47589 78477 -47579
rect 78424 -47595 78477 -47589
rect 78507 -47507 78563 -47465
rect 78845 -47483 78897 -47465
rect 78507 -47541 78517 -47507
rect 78551 -47541 78563 -47507
rect 78507 -47595 78563 -47541
rect 78649 -47521 78705 -47483
rect 78649 -47555 78661 -47521
rect 78695 -47555 78705 -47521
rect 78649 -47567 78705 -47555
rect 78735 -47567 78789 -47483
rect 78819 -47549 78897 -47483
rect 78819 -47567 78853 -47549
rect 78845 -47583 78853 -47567
rect 78887 -47583 78897 -47549
rect 78845 -47595 78897 -47583
rect 78927 -47549 78983 -47465
rect 78927 -47583 78937 -47549
rect 78971 -47583 78983 -47549
rect 78927 -47595 78983 -47583
rect 55288 -47758 55488 -47746
rect 55288 -47792 55300 -47758
rect 55476 -47792 55488 -47758
rect 55288 -47804 55488 -47792
rect 55288 -47846 55488 -47834
rect 55288 -47880 55300 -47846
rect 55476 -47880 55488 -47846
rect 55288 -47892 55488 -47880
rect 77966 -47781 78019 -47775
rect 77605 -47811 77657 -47781
rect 77605 -47845 77613 -47811
rect 77647 -47845 77657 -47811
rect 77605 -47865 77657 -47845
rect 77687 -47805 77753 -47781
rect 77687 -47839 77703 -47805
rect 77737 -47839 77753 -47805
rect 77687 -47865 77753 -47839
rect 77783 -47791 77837 -47781
rect 77783 -47825 77793 -47791
rect 77827 -47825 77837 -47791
rect 77783 -47865 77837 -47825
rect 77867 -47805 77921 -47781
rect 77867 -47839 77877 -47805
rect 77911 -47839 77921 -47805
rect 77867 -47865 77921 -47839
rect 77951 -47791 78019 -47781
rect 77951 -47825 77971 -47791
rect 78005 -47825 78019 -47791
rect 77951 -47865 78019 -47825
rect 77966 -47905 78019 -47865
rect 78049 -47829 78103 -47775
rect 78049 -47863 78059 -47829
rect 78093 -47863 78103 -47829
rect 78049 -47905 78103 -47863
rect 83075 -48161 83127 -48115
rect 82894 -48189 82946 -48161
rect 82894 -48223 82902 -48189
rect 82936 -48223 82946 -48189
rect 82894 -48245 82946 -48223
rect 82976 -48189 83030 -48161
rect 82976 -48223 82986 -48189
rect 83020 -48223 83030 -48189
rect 82976 -48245 83030 -48223
rect 83060 -48189 83127 -48161
rect 83060 -48223 83082 -48189
rect 83116 -48223 83127 -48189
rect 83060 -48245 83127 -48223
rect 83157 -48129 83209 -48115
rect 83157 -48163 83167 -48129
rect 83201 -48163 83209 -48129
rect 83157 -48197 83209 -48163
rect 83157 -48231 83167 -48197
rect 83201 -48231 83209 -48197
rect 83157 -48245 83209 -48231
rect 83366 -48127 83418 -48115
rect 83366 -48161 83374 -48127
rect 83408 -48161 83418 -48127
rect 83366 -48195 83418 -48161
rect 83366 -48229 83374 -48195
rect 83408 -48229 83418 -48195
rect 83366 -48245 83418 -48229
rect 83448 -48127 83500 -48115
rect 83448 -48161 83458 -48127
rect 83492 -48161 83500 -48127
rect 83448 -48195 83500 -48161
rect 83448 -48229 83458 -48195
rect 83492 -48229 83500 -48195
rect 83448 -48245 83500 -48229
rect 83611 -48199 83663 -48115
rect 83611 -48233 83619 -48199
rect 83653 -48233 83663 -48199
rect 83611 -48245 83663 -48233
rect 83693 -48191 83747 -48115
rect 83693 -48225 83703 -48191
rect 83737 -48225 83747 -48191
rect 83693 -48245 83747 -48225
rect 83777 -48199 83831 -48115
rect 83777 -48233 83787 -48199
rect 83821 -48233 83831 -48199
rect 83777 -48245 83831 -48233
rect 83861 -48191 83915 -48115
rect 83861 -48225 83871 -48191
rect 83905 -48225 83915 -48191
rect 83861 -48245 83915 -48225
rect 83945 -48198 83997 -48115
rect 83945 -48232 83955 -48198
rect 83989 -48232 83997 -48198
rect 83945 -48245 83997 -48232
rect 84074 -48131 84126 -48115
rect 84074 -48165 84082 -48131
rect 84116 -48165 84126 -48131
rect 84074 -48199 84126 -48165
rect 84074 -48233 84082 -48199
rect 84116 -48233 84126 -48199
rect 84074 -48245 84126 -48233
rect 84156 -48131 84210 -48115
rect 84156 -48165 84166 -48131
rect 84200 -48165 84210 -48131
rect 84156 -48199 84210 -48165
rect 84156 -48233 84166 -48199
rect 84200 -48233 84210 -48199
rect 84156 -48245 84210 -48233
rect 84240 -48199 84294 -48115
rect 84240 -48233 84250 -48199
rect 84284 -48233 84294 -48199
rect 84240 -48245 84294 -48233
rect 84324 -48131 84378 -48115
rect 84324 -48165 84334 -48131
rect 84368 -48165 84378 -48131
rect 84324 -48199 84378 -48165
rect 84324 -48233 84334 -48199
rect 84368 -48233 84378 -48199
rect 84324 -48245 84378 -48233
rect 84408 -48199 84462 -48115
rect 84408 -48233 84418 -48199
rect 84452 -48233 84462 -48199
rect 84408 -48245 84462 -48233
rect 84492 -48131 84546 -48115
rect 84492 -48165 84502 -48131
rect 84536 -48165 84546 -48131
rect 84492 -48199 84546 -48165
rect 84492 -48233 84502 -48199
rect 84536 -48233 84546 -48199
rect 84492 -48245 84546 -48233
rect 84576 -48199 84630 -48115
rect 84576 -48233 84586 -48199
rect 84620 -48233 84630 -48199
rect 84576 -48245 84630 -48233
rect 84660 -48131 84714 -48115
rect 84660 -48165 84670 -48131
rect 84704 -48165 84714 -48131
rect 84660 -48199 84714 -48165
rect 84660 -48233 84670 -48199
rect 84704 -48233 84714 -48199
rect 84660 -48245 84714 -48233
rect 84744 -48199 84798 -48115
rect 84744 -48233 84754 -48199
rect 84788 -48233 84798 -48199
rect 84744 -48245 84798 -48233
rect 84828 -48131 84882 -48115
rect 84828 -48165 84838 -48131
rect 84872 -48165 84882 -48131
rect 84828 -48199 84882 -48165
rect 84828 -48233 84838 -48199
rect 84872 -48233 84882 -48199
rect 84828 -48245 84882 -48233
rect 84912 -48199 84966 -48115
rect 84912 -48233 84922 -48199
rect 84956 -48233 84966 -48199
rect 84912 -48245 84966 -48233
rect 84996 -48131 85050 -48115
rect 84996 -48165 85006 -48131
rect 85040 -48165 85050 -48131
rect 84996 -48199 85050 -48165
rect 84996 -48233 85006 -48199
rect 85040 -48233 85050 -48199
rect 84996 -48245 85050 -48233
rect 85080 -48199 85134 -48115
rect 85080 -48233 85090 -48199
rect 85124 -48233 85134 -48199
rect 85080 -48245 85134 -48233
rect 85164 -48131 85218 -48115
rect 85164 -48165 85174 -48131
rect 85208 -48165 85218 -48131
rect 85164 -48199 85218 -48165
rect 85164 -48233 85174 -48199
rect 85208 -48233 85218 -48199
rect 85164 -48245 85218 -48233
rect 85248 -48199 85302 -48115
rect 85248 -48233 85258 -48199
rect 85292 -48233 85302 -48199
rect 85248 -48245 85302 -48233
rect 85332 -48131 85386 -48115
rect 85332 -48165 85342 -48131
rect 85376 -48165 85386 -48131
rect 85332 -48199 85386 -48165
rect 85332 -48233 85342 -48199
rect 85376 -48233 85386 -48199
rect 85332 -48245 85386 -48233
rect 85416 -48131 85468 -48115
rect 85416 -48165 85426 -48131
rect 85460 -48165 85468 -48131
rect 85416 -48199 85468 -48165
rect 85416 -48233 85426 -48199
rect 85460 -48233 85468 -48199
rect 85416 -48245 85468 -48233
rect 85546 -48131 85598 -48115
rect 85546 -48165 85554 -48131
rect 85588 -48165 85598 -48131
rect 85546 -48199 85598 -48165
rect 85546 -48233 85554 -48199
rect 85588 -48233 85598 -48199
rect 85546 -48245 85598 -48233
rect 85628 -48131 85682 -48115
rect 85628 -48165 85638 -48131
rect 85672 -48165 85682 -48131
rect 85628 -48199 85682 -48165
rect 85628 -48233 85638 -48199
rect 85672 -48233 85682 -48199
rect 85628 -48245 85682 -48233
rect 85712 -48199 85766 -48115
rect 85712 -48233 85722 -48199
rect 85756 -48233 85766 -48199
rect 85712 -48245 85766 -48233
rect 85796 -48131 85850 -48115
rect 85796 -48165 85806 -48131
rect 85840 -48165 85850 -48131
rect 85796 -48199 85850 -48165
rect 85796 -48233 85806 -48199
rect 85840 -48233 85850 -48199
rect 85796 -48245 85850 -48233
rect 85880 -48199 85934 -48115
rect 85880 -48233 85890 -48199
rect 85924 -48233 85934 -48199
rect 85880 -48245 85934 -48233
rect 85964 -48131 86018 -48115
rect 85964 -48165 85974 -48131
rect 86008 -48165 86018 -48131
rect 85964 -48199 86018 -48165
rect 85964 -48233 85974 -48199
rect 86008 -48233 86018 -48199
rect 85964 -48245 86018 -48233
rect 86048 -48199 86102 -48115
rect 86048 -48233 86058 -48199
rect 86092 -48233 86102 -48199
rect 86048 -48245 86102 -48233
rect 86132 -48131 86186 -48115
rect 86132 -48165 86142 -48131
rect 86176 -48165 86186 -48131
rect 86132 -48199 86186 -48165
rect 86132 -48233 86142 -48199
rect 86176 -48233 86186 -48199
rect 86132 -48245 86186 -48233
rect 86216 -48199 86270 -48115
rect 86216 -48233 86226 -48199
rect 86260 -48233 86270 -48199
rect 86216 -48245 86270 -48233
rect 86300 -48131 86354 -48115
rect 86300 -48165 86310 -48131
rect 86344 -48165 86354 -48131
rect 86300 -48199 86354 -48165
rect 86300 -48233 86310 -48199
rect 86344 -48233 86354 -48199
rect 86300 -48245 86354 -48233
rect 86384 -48199 86438 -48115
rect 86384 -48233 86394 -48199
rect 86428 -48233 86438 -48199
rect 86384 -48245 86438 -48233
rect 86468 -48131 86522 -48115
rect 86468 -48165 86478 -48131
rect 86512 -48165 86522 -48131
rect 86468 -48199 86522 -48165
rect 86468 -48233 86478 -48199
rect 86512 -48233 86522 -48199
rect 86468 -48245 86522 -48233
rect 86552 -48199 86606 -48115
rect 86552 -48233 86562 -48199
rect 86596 -48233 86606 -48199
rect 86552 -48245 86606 -48233
rect 86636 -48131 86690 -48115
rect 86636 -48165 86646 -48131
rect 86680 -48165 86690 -48131
rect 86636 -48199 86690 -48165
rect 86636 -48233 86646 -48199
rect 86680 -48233 86690 -48199
rect 86636 -48245 86690 -48233
rect 86720 -48199 86774 -48115
rect 86720 -48233 86730 -48199
rect 86764 -48233 86774 -48199
rect 86720 -48245 86774 -48233
rect 86804 -48131 86858 -48115
rect 86804 -48165 86814 -48131
rect 86848 -48165 86858 -48131
rect 86804 -48199 86858 -48165
rect 86804 -48233 86814 -48199
rect 86848 -48233 86858 -48199
rect 86804 -48245 86858 -48233
rect 86888 -48131 86940 -48115
rect 86888 -48165 86898 -48131
rect 86932 -48165 86940 -48131
rect 86888 -48199 86940 -48165
rect 86888 -48233 86898 -48199
rect 86932 -48233 86940 -48199
rect 86888 -48245 86940 -48233
rect 87018 -48131 87070 -48115
rect 87018 -48165 87026 -48131
rect 87060 -48165 87070 -48131
rect 87018 -48199 87070 -48165
rect 87018 -48233 87026 -48199
rect 87060 -48233 87070 -48199
rect 87018 -48245 87070 -48233
rect 87100 -48131 87154 -48115
rect 87100 -48165 87110 -48131
rect 87144 -48165 87154 -48131
rect 87100 -48199 87154 -48165
rect 87100 -48233 87110 -48199
rect 87144 -48233 87154 -48199
rect 87100 -48245 87154 -48233
rect 87184 -48199 87238 -48115
rect 87184 -48233 87194 -48199
rect 87228 -48233 87238 -48199
rect 87184 -48245 87238 -48233
rect 87268 -48131 87322 -48115
rect 87268 -48165 87278 -48131
rect 87312 -48165 87322 -48131
rect 87268 -48199 87322 -48165
rect 87268 -48233 87278 -48199
rect 87312 -48233 87322 -48199
rect 87268 -48245 87322 -48233
rect 87352 -48199 87406 -48115
rect 87352 -48233 87362 -48199
rect 87396 -48233 87406 -48199
rect 87352 -48245 87406 -48233
rect 87436 -48131 87490 -48115
rect 87436 -48165 87446 -48131
rect 87480 -48165 87490 -48131
rect 87436 -48199 87490 -48165
rect 87436 -48233 87446 -48199
rect 87480 -48233 87490 -48199
rect 87436 -48245 87490 -48233
rect 87520 -48199 87574 -48115
rect 87520 -48233 87530 -48199
rect 87564 -48233 87574 -48199
rect 87520 -48245 87574 -48233
rect 87604 -48131 87658 -48115
rect 87604 -48165 87614 -48131
rect 87648 -48165 87658 -48131
rect 87604 -48199 87658 -48165
rect 87604 -48233 87614 -48199
rect 87648 -48233 87658 -48199
rect 87604 -48245 87658 -48233
rect 87688 -48199 87742 -48115
rect 87688 -48233 87698 -48199
rect 87732 -48233 87742 -48199
rect 87688 -48245 87742 -48233
rect 87772 -48131 87826 -48115
rect 87772 -48165 87782 -48131
rect 87816 -48165 87826 -48131
rect 87772 -48199 87826 -48165
rect 87772 -48233 87782 -48199
rect 87816 -48233 87826 -48199
rect 87772 -48245 87826 -48233
rect 87856 -48199 87910 -48115
rect 87856 -48233 87866 -48199
rect 87900 -48233 87910 -48199
rect 87856 -48245 87910 -48233
rect 87940 -48131 87994 -48115
rect 87940 -48165 87950 -48131
rect 87984 -48165 87994 -48131
rect 87940 -48199 87994 -48165
rect 87940 -48233 87950 -48199
rect 87984 -48233 87994 -48199
rect 87940 -48245 87994 -48233
rect 88024 -48199 88078 -48115
rect 88024 -48233 88034 -48199
rect 88068 -48233 88078 -48199
rect 88024 -48245 88078 -48233
rect 88108 -48131 88162 -48115
rect 88108 -48165 88118 -48131
rect 88152 -48165 88162 -48131
rect 88108 -48199 88162 -48165
rect 88108 -48233 88118 -48199
rect 88152 -48233 88162 -48199
rect 88108 -48245 88162 -48233
rect 88192 -48199 88246 -48115
rect 88192 -48233 88202 -48199
rect 88236 -48233 88246 -48199
rect 88192 -48245 88246 -48233
rect 88276 -48131 88330 -48115
rect 88276 -48165 88286 -48131
rect 88320 -48165 88330 -48131
rect 88276 -48199 88330 -48165
rect 88276 -48233 88286 -48199
rect 88320 -48233 88330 -48199
rect 88276 -48245 88330 -48233
rect 88360 -48131 88412 -48115
rect 88360 -48165 88370 -48131
rect 88404 -48165 88412 -48131
rect 88360 -48199 88412 -48165
rect 88360 -48233 88370 -48199
rect 88404 -48233 88412 -48199
rect 88360 -48245 88412 -48233
rect 88490 -48131 88542 -48115
rect 88490 -48165 88498 -48131
rect 88532 -48165 88542 -48131
rect 88490 -48199 88542 -48165
rect 88490 -48233 88498 -48199
rect 88532 -48233 88542 -48199
rect 88490 -48245 88542 -48233
rect 88572 -48131 88626 -48115
rect 88572 -48165 88582 -48131
rect 88616 -48165 88626 -48131
rect 88572 -48199 88626 -48165
rect 88572 -48233 88582 -48199
rect 88616 -48233 88626 -48199
rect 88572 -48245 88626 -48233
rect 88656 -48199 88710 -48115
rect 88656 -48233 88666 -48199
rect 88700 -48233 88710 -48199
rect 88656 -48245 88710 -48233
rect 88740 -48131 88794 -48115
rect 88740 -48165 88750 -48131
rect 88784 -48165 88794 -48131
rect 88740 -48199 88794 -48165
rect 88740 -48233 88750 -48199
rect 88784 -48233 88794 -48199
rect 88740 -48245 88794 -48233
rect 88824 -48199 88878 -48115
rect 88824 -48233 88834 -48199
rect 88868 -48233 88878 -48199
rect 88824 -48245 88878 -48233
rect 88908 -48131 88962 -48115
rect 88908 -48165 88918 -48131
rect 88952 -48165 88962 -48131
rect 88908 -48199 88962 -48165
rect 88908 -48233 88918 -48199
rect 88952 -48233 88962 -48199
rect 88908 -48245 88962 -48233
rect 88992 -48199 89046 -48115
rect 88992 -48233 89002 -48199
rect 89036 -48233 89046 -48199
rect 88992 -48245 89046 -48233
rect 89076 -48131 89130 -48115
rect 89076 -48165 89086 -48131
rect 89120 -48165 89130 -48131
rect 89076 -48199 89130 -48165
rect 89076 -48233 89086 -48199
rect 89120 -48233 89130 -48199
rect 89076 -48245 89130 -48233
rect 89160 -48199 89214 -48115
rect 89160 -48233 89170 -48199
rect 89204 -48233 89214 -48199
rect 89160 -48245 89214 -48233
rect 89244 -48131 89298 -48115
rect 89244 -48165 89254 -48131
rect 89288 -48165 89298 -48131
rect 89244 -48199 89298 -48165
rect 89244 -48233 89254 -48199
rect 89288 -48233 89298 -48199
rect 89244 -48245 89298 -48233
rect 89328 -48199 89382 -48115
rect 89328 -48233 89338 -48199
rect 89372 -48233 89382 -48199
rect 89328 -48245 89382 -48233
rect 89412 -48131 89466 -48115
rect 89412 -48165 89422 -48131
rect 89456 -48165 89466 -48131
rect 89412 -48199 89466 -48165
rect 89412 -48233 89422 -48199
rect 89456 -48233 89466 -48199
rect 89412 -48245 89466 -48233
rect 89496 -48199 89550 -48115
rect 89496 -48233 89506 -48199
rect 89540 -48233 89550 -48199
rect 89496 -48245 89550 -48233
rect 89580 -48131 89634 -48115
rect 89580 -48165 89590 -48131
rect 89624 -48165 89634 -48131
rect 89580 -48199 89634 -48165
rect 89580 -48233 89590 -48199
rect 89624 -48233 89634 -48199
rect 89580 -48245 89634 -48233
rect 89664 -48199 89718 -48115
rect 89664 -48233 89674 -48199
rect 89708 -48233 89718 -48199
rect 89664 -48245 89718 -48233
rect 89748 -48131 89802 -48115
rect 89748 -48165 89758 -48131
rect 89792 -48165 89802 -48131
rect 89748 -48199 89802 -48165
rect 89748 -48233 89758 -48199
rect 89792 -48233 89802 -48199
rect 89748 -48245 89802 -48233
rect 89832 -48131 89884 -48115
rect 89832 -48165 89842 -48131
rect 89876 -48165 89884 -48131
rect 89832 -48199 89884 -48165
rect 89832 -48233 89842 -48199
rect 89876 -48233 89884 -48199
rect 89832 -48245 89884 -48233
rect 89962 -48131 90014 -48115
rect 89962 -48165 89970 -48131
rect 90004 -48165 90014 -48131
rect 89962 -48199 90014 -48165
rect 89962 -48233 89970 -48199
rect 90004 -48233 90014 -48199
rect 89962 -48245 90014 -48233
rect 90044 -48131 90098 -48115
rect 90044 -48165 90054 -48131
rect 90088 -48165 90098 -48131
rect 90044 -48199 90098 -48165
rect 90044 -48233 90054 -48199
rect 90088 -48233 90098 -48199
rect 90044 -48245 90098 -48233
rect 90128 -48199 90182 -48115
rect 90128 -48233 90138 -48199
rect 90172 -48233 90182 -48199
rect 90128 -48245 90182 -48233
rect 90212 -48131 90266 -48115
rect 90212 -48165 90222 -48131
rect 90256 -48165 90266 -48131
rect 90212 -48199 90266 -48165
rect 90212 -48233 90222 -48199
rect 90256 -48233 90266 -48199
rect 90212 -48245 90266 -48233
rect 90296 -48199 90350 -48115
rect 90296 -48233 90306 -48199
rect 90340 -48233 90350 -48199
rect 90296 -48245 90350 -48233
rect 90380 -48131 90434 -48115
rect 90380 -48165 90390 -48131
rect 90424 -48165 90434 -48131
rect 90380 -48199 90434 -48165
rect 90380 -48233 90390 -48199
rect 90424 -48233 90434 -48199
rect 90380 -48245 90434 -48233
rect 90464 -48199 90518 -48115
rect 90464 -48233 90474 -48199
rect 90508 -48233 90518 -48199
rect 90464 -48245 90518 -48233
rect 90548 -48131 90602 -48115
rect 90548 -48165 90558 -48131
rect 90592 -48165 90602 -48131
rect 90548 -48199 90602 -48165
rect 90548 -48233 90558 -48199
rect 90592 -48233 90602 -48199
rect 90548 -48245 90602 -48233
rect 90632 -48199 90686 -48115
rect 90632 -48233 90642 -48199
rect 90676 -48233 90686 -48199
rect 90632 -48245 90686 -48233
rect 90716 -48131 90770 -48115
rect 90716 -48165 90726 -48131
rect 90760 -48165 90770 -48131
rect 90716 -48199 90770 -48165
rect 90716 -48233 90726 -48199
rect 90760 -48233 90770 -48199
rect 90716 -48245 90770 -48233
rect 90800 -48199 90854 -48115
rect 90800 -48233 90810 -48199
rect 90844 -48233 90854 -48199
rect 90800 -48245 90854 -48233
rect 90884 -48131 90938 -48115
rect 90884 -48165 90894 -48131
rect 90928 -48165 90938 -48131
rect 90884 -48199 90938 -48165
rect 90884 -48233 90894 -48199
rect 90928 -48233 90938 -48199
rect 90884 -48245 90938 -48233
rect 90968 -48199 91022 -48115
rect 90968 -48233 90978 -48199
rect 91012 -48233 91022 -48199
rect 90968 -48245 91022 -48233
rect 91052 -48131 91106 -48115
rect 91052 -48165 91062 -48131
rect 91096 -48165 91106 -48131
rect 91052 -48199 91106 -48165
rect 91052 -48233 91062 -48199
rect 91096 -48233 91106 -48199
rect 91052 -48245 91106 -48233
rect 91136 -48199 91190 -48115
rect 91136 -48233 91146 -48199
rect 91180 -48233 91190 -48199
rect 91136 -48245 91190 -48233
rect 91220 -48131 91274 -48115
rect 91220 -48165 91230 -48131
rect 91264 -48165 91274 -48131
rect 91220 -48199 91274 -48165
rect 91220 -48233 91230 -48199
rect 91264 -48233 91274 -48199
rect 91220 -48245 91274 -48233
rect 91304 -48131 91356 -48115
rect 91304 -48165 91314 -48131
rect 91348 -48165 91356 -48131
rect 91304 -48199 91356 -48165
rect 91304 -48233 91314 -48199
rect 91348 -48233 91356 -48199
rect 91304 -48245 91356 -48233
rect 77833 -48733 77885 -48715
rect 77637 -48771 77693 -48733
rect 77637 -48805 77649 -48771
rect 77683 -48805 77693 -48771
rect 77637 -48817 77693 -48805
rect 77723 -48817 77777 -48733
rect 77807 -48799 77885 -48733
rect 77807 -48817 77841 -48799
rect 77833 -48833 77841 -48817
rect 77875 -48833 77885 -48799
rect 77833 -48845 77885 -48833
rect 77915 -48799 77971 -48715
rect 77915 -48833 77925 -48799
rect 77959 -48833 77971 -48799
rect 77915 -48845 77971 -48833
rect 77833 -49027 77885 -49015
rect 77833 -49043 77841 -49027
rect 77637 -49055 77693 -49043
rect 77637 -49089 77649 -49055
rect 77683 -49089 77693 -49055
rect 77637 -49127 77693 -49089
rect 77723 -49127 77777 -49043
rect 77807 -49061 77841 -49043
rect 77875 -49061 77885 -49027
rect 77807 -49127 77885 -49061
rect 77833 -49145 77885 -49127
rect 77915 -49027 77971 -49015
rect 78426 -49021 78479 -49015
rect 77915 -49061 77925 -49027
rect 77959 -49061 77971 -49027
rect 77915 -49145 77971 -49061
rect 78065 -49051 78117 -49021
rect 78065 -49085 78073 -49051
rect 78107 -49085 78117 -49051
rect 78065 -49105 78117 -49085
rect 78147 -49045 78213 -49021
rect 78147 -49079 78163 -49045
rect 78197 -49079 78213 -49045
rect 78147 -49105 78213 -49079
rect 78243 -49031 78297 -49021
rect 78243 -49065 78253 -49031
rect 78287 -49065 78297 -49031
rect 78243 -49105 78297 -49065
rect 78327 -49045 78381 -49021
rect 78327 -49079 78337 -49045
rect 78371 -49079 78381 -49045
rect 78327 -49105 78381 -49079
rect 78411 -49031 78479 -49021
rect 78411 -49065 78431 -49031
rect 78465 -49065 78479 -49031
rect 78411 -49105 78479 -49065
rect 78426 -49145 78479 -49105
rect 78509 -49069 78563 -49015
rect 78509 -49103 78519 -49069
rect 78553 -49103 78563 -49069
rect 78509 -49145 78563 -49103
rect 77833 -49973 77885 -49955
rect 77637 -50011 77693 -49973
rect 77637 -50045 77649 -50011
rect 77683 -50045 77693 -50011
rect 77637 -50057 77693 -50045
rect 77723 -50057 77777 -49973
rect 77807 -50039 77885 -49973
rect 77807 -50057 77841 -50039
rect 77833 -50073 77841 -50057
rect 77875 -50073 77885 -50039
rect 77833 -50085 77885 -50073
rect 77915 -50039 77971 -49955
rect 77915 -50073 77925 -50039
rect 77959 -50073 77971 -50039
rect 77915 -50085 77971 -50073
rect 77835 -50281 77887 -50269
rect 77835 -50297 77843 -50281
rect 77639 -50309 77695 -50297
rect 77639 -50343 77651 -50309
rect 77685 -50343 77695 -50309
rect 77639 -50381 77695 -50343
rect 77725 -50381 77779 -50297
rect 77809 -50315 77843 -50297
rect 77877 -50315 77887 -50281
rect 77809 -50381 77887 -50315
rect 53452 -50790 53510 -50778
rect 53452 -51566 53464 -50790
rect 53498 -51566 53510 -50790
rect 53452 -51578 53510 -51566
rect 53630 -50790 53688 -50778
rect 53630 -51566 53642 -50790
rect 53676 -51566 53688 -50790
rect 53630 -51578 53688 -51566
rect 55278 -50852 55336 -50840
rect 55278 -51028 55290 -50852
rect 55324 -51028 55336 -50852
rect 55278 -51040 55336 -51028
rect 55366 -50852 55424 -50840
rect 55366 -51028 55378 -50852
rect 55412 -51028 55424 -50852
rect 55366 -51040 55424 -51028
rect 53930 -51378 54730 -51366
rect 53930 -51412 53942 -51378
rect 54718 -51412 54730 -51378
rect 53930 -51424 54730 -51412
rect 53930 -51556 54730 -51544
rect 53930 -51590 53942 -51556
rect 54718 -51590 54730 -51556
rect 53930 -51602 54730 -51590
rect 55808 -50740 55866 -50728
rect 55808 -51516 55820 -50740
rect 55854 -51516 55866 -50740
rect 55808 -51528 55866 -51516
rect 55986 -50740 56044 -50728
rect 55986 -51516 55998 -50740
rect 56032 -51516 56044 -50740
rect 55986 -51528 56044 -51516
rect 77835 -50399 77887 -50381
rect 77917 -50281 77973 -50269
rect 77917 -50315 77927 -50281
rect 77961 -50315 77973 -50281
rect 77917 -50399 77973 -50315
rect 57123 -51100 57175 -51055
rect 53452 -51808 53510 -51796
rect 53452 -52584 53464 -51808
rect 53498 -52584 53510 -51808
rect 53452 -52596 53510 -52584
rect 53630 -51808 53688 -51796
rect 53630 -52584 53642 -51808
rect 53676 -52584 53688 -51808
rect 53630 -52596 53688 -52584
rect 53930 -51784 54730 -51772
rect 53930 -51818 53942 -51784
rect 54718 -51818 54730 -51784
rect 53930 -51830 54730 -51818
rect 53930 -51962 54730 -51950
rect 53930 -51996 53942 -51962
rect 54718 -51996 54730 -51962
rect 53930 -52008 54730 -51996
rect 55268 -52348 55326 -52336
rect 55268 -52524 55280 -52348
rect 55314 -52524 55326 -52348
rect 55268 -52536 55326 -52524
rect 55356 -52348 55414 -52336
rect 55356 -52524 55368 -52348
rect 55402 -52524 55414 -52348
rect 55356 -52536 55414 -52524
rect 55808 -51854 55866 -51842
rect 55808 -52630 55820 -51854
rect 55854 -52630 55866 -51854
rect 55808 -52642 55866 -52630
rect 55986 -51854 56044 -51842
rect 55986 -52630 55998 -51854
rect 56032 -52630 56044 -51854
rect 55986 -52642 56044 -52630
rect 57123 -51134 57131 -51100
rect 57165 -51134 57175 -51100
rect 57123 -51159 57175 -51134
rect 57205 -51113 57263 -51055
rect 57205 -51147 57217 -51113
rect 57251 -51147 57263 -51113
rect 57205 -51159 57263 -51147
rect 57293 -51083 57345 -51055
rect 57293 -51117 57303 -51083
rect 57337 -51117 57345 -51083
rect 57293 -51159 57345 -51117
rect 59946 -50974 60346 -50962
rect 59946 -51008 59958 -50974
rect 60334 -51008 60346 -50974
rect 59946 -51020 60346 -51008
rect 59946 -51082 60346 -51070
rect 59946 -51116 59958 -51082
rect 60334 -51116 60346 -51082
rect 59946 -51128 60346 -51116
rect 59490 -51382 59548 -51370
rect 59490 -51450 59502 -51382
rect 59476 -51520 59502 -51450
rect 59490 -51558 59502 -51520
rect 59536 -51558 59548 -51382
rect 59490 -51570 59548 -51558
rect 59578 -51382 59636 -51370
rect 59578 -51558 59590 -51382
rect 59624 -51558 59636 -51382
rect 59578 -51570 59636 -51558
rect 59806 -51382 59864 -51370
rect 59806 -51558 59818 -51382
rect 59852 -51558 59864 -51382
rect 59806 -51570 59864 -51558
rect 59894 -51382 59952 -51370
rect 59894 -51558 59906 -51382
rect 59940 -51558 59952 -51382
rect 59894 -51570 59952 -51558
rect 78020 -51221 78113 -51205
rect 78020 -51251 78054 -51221
rect 77605 -51281 77657 -51251
rect 77605 -51315 77613 -51281
rect 77647 -51315 77657 -51281
rect 77605 -51335 77657 -51315
rect 77687 -51335 77745 -51251
rect 77775 -51335 77851 -51251
rect 77881 -51335 77947 -51251
rect 77977 -51255 78054 -51251
rect 78088 -51255 78113 -51221
rect 77977 -51289 78113 -51255
rect 77977 -51323 78054 -51289
rect 78088 -51323 78113 -51289
rect 77977 -51335 78113 -51323
rect 78143 -51221 78195 -51205
rect 78143 -51255 78153 -51221
rect 78187 -51255 78195 -51221
rect 78710 -51245 78763 -51205
rect 78143 -51289 78195 -51255
rect 78143 -51323 78153 -51289
rect 78187 -51323 78195 -51289
rect 78143 -51335 78195 -51323
rect 78349 -51265 78401 -51245
rect 78349 -51299 78357 -51265
rect 78391 -51299 78401 -51265
rect 78349 -51329 78401 -51299
rect 78431 -51271 78497 -51245
rect 78431 -51305 78447 -51271
rect 78481 -51305 78497 -51271
rect 78431 -51329 78497 -51305
rect 78527 -51285 78581 -51245
rect 78527 -51319 78537 -51285
rect 78571 -51319 78581 -51285
rect 78527 -51329 78581 -51319
rect 78611 -51271 78665 -51245
rect 78611 -51305 78621 -51271
rect 78655 -51305 78665 -51271
rect 78611 -51329 78665 -51305
rect 78695 -51285 78763 -51245
rect 78695 -51319 78715 -51285
rect 78749 -51319 78763 -51285
rect 78695 -51329 78763 -51319
rect 78710 -51335 78763 -51329
rect 78793 -51247 78847 -51205
rect 78793 -51281 78803 -51247
rect 78837 -51281 78847 -51247
rect 78793 -51335 78847 -51281
rect 77605 -51521 77657 -51501
rect 77605 -51555 77613 -51521
rect 77647 -51555 77657 -51521
rect 60191 -51573 60321 -51565
rect 60191 -51607 60203 -51573
rect 60237 -51607 60321 -51573
rect 60191 -51617 60321 -51607
rect 61131 -51573 61261 -51565
rect 61131 -51607 61215 -51573
rect 61249 -51607 61261 -51573
rect 77605 -51585 77657 -51555
rect 77687 -51585 77745 -51501
rect 77775 -51585 77851 -51501
rect 77881 -51585 77947 -51501
rect 77977 -51513 78113 -51501
rect 77977 -51547 78054 -51513
rect 78088 -51547 78113 -51513
rect 77977 -51581 78113 -51547
rect 77977 -51585 78054 -51581
rect 61131 -51617 61261 -51607
rect 60191 -51657 60321 -51647
rect 60191 -51691 60211 -51657
rect 60245 -51691 60321 -51657
rect 60191 -51701 60321 -51691
rect 61131 -51657 61261 -51647
rect 61131 -51691 61207 -51657
rect 61241 -51691 61261 -51657
rect 61131 -51701 61261 -51691
rect 57123 -52254 57175 -52229
rect 57123 -52288 57131 -52254
rect 57165 -52288 57175 -52254
rect 57123 -52333 57175 -52288
rect 57205 -52241 57263 -52229
rect 57205 -52275 57217 -52241
rect 57251 -52275 57263 -52241
rect 57205 -52333 57263 -52275
rect 57293 -52271 57345 -52229
rect 57293 -52305 57303 -52271
rect 57337 -52305 57345 -52271
rect 57293 -52333 57345 -52305
rect 78020 -51615 78054 -51585
rect 78088 -51615 78113 -51581
rect 78020 -51631 78113 -51615
rect 78143 -51513 78195 -51501
rect 78143 -51547 78153 -51513
rect 78187 -51547 78195 -51513
rect 78143 -51581 78195 -51547
rect 78143 -51615 78153 -51581
rect 78187 -51615 78195 -51581
rect 78143 -51631 78195 -51615
rect 60191 -51741 60321 -51731
rect 59489 -51895 59547 -51883
rect 59489 -52071 59501 -51895
rect 59535 -52071 59547 -51895
rect 59489 -52083 59547 -52071
rect 59577 -51895 59635 -51883
rect 59577 -52071 59589 -51895
rect 59623 -52071 59635 -51895
rect 59577 -52083 59635 -52071
rect 60191 -51775 60203 -51741
rect 60237 -51775 60321 -51741
rect 60191 -51785 60321 -51775
rect 61131 -51741 61261 -51731
rect 61131 -51775 61215 -51741
rect 61249 -51775 61261 -51741
rect 61131 -51785 61261 -51775
rect 59805 -51895 59863 -51883
rect 59805 -52071 59817 -51895
rect 59851 -52071 59863 -51895
rect 59805 -52083 59863 -52071
rect 59893 -51895 59951 -51883
rect 59893 -52071 59905 -51895
rect 59939 -52071 59951 -51895
rect 59893 -52083 59951 -52071
rect 60191 -51825 60321 -51815
rect 60191 -51859 60211 -51825
rect 60245 -51859 60321 -51825
rect 60191 -51869 60321 -51859
rect 61131 -51825 61261 -51815
rect 61131 -51859 61207 -51825
rect 61241 -51859 61261 -51825
rect 61131 -51869 61261 -51859
rect 60191 -51909 60321 -51899
rect 60191 -51943 60204 -51909
rect 60238 -51943 60321 -51909
rect 60191 -51951 60321 -51943
rect 61131 -51909 61261 -51899
rect 61131 -51943 61214 -51909
rect 61248 -51943 61261 -51909
rect 61131 -51951 61261 -51943
rect 83075 -51811 83127 -51765
rect 82894 -51839 82946 -51811
rect 82894 -51873 82902 -51839
rect 82936 -51873 82946 -51839
rect 82894 -51895 82946 -51873
rect 82976 -51839 83030 -51811
rect 82976 -51873 82986 -51839
rect 83020 -51873 83030 -51839
rect 82976 -51895 83030 -51873
rect 83060 -51839 83127 -51811
rect 83060 -51873 83082 -51839
rect 83116 -51873 83127 -51839
rect 83060 -51895 83127 -51873
rect 83157 -51779 83209 -51765
rect 83157 -51813 83167 -51779
rect 83201 -51813 83209 -51779
rect 83157 -51847 83209 -51813
rect 83157 -51881 83167 -51847
rect 83201 -51881 83209 -51847
rect 83157 -51895 83209 -51881
rect 83366 -51777 83418 -51765
rect 83366 -51811 83374 -51777
rect 83408 -51811 83418 -51777
rect 83366 -51845 83418 -51811
rect 83366 -51879 83374 -51845
rect 83408 -51879 83418 -51845
rect 83366 -51895 83418 -51879
rect 83448 -51777 83500 -51765
rect 83448 -51811 83458 -51777
rect 83492 -51811 83500 -51777
rect 83448 -51845 83500 -51811
rect 83448 -51879 83458 -51845
rect 83492 -51879 83500 -51845
rect 83448 -51895 83500 -51879
rect 83611 -51849 83663 -51765
rect 83611 -51883 83619 -51849
rect 83653 -51883 83663 -51849
rect 83611 -51895 83663 -51883
rect 83693 -51841 83747 -51765
rect 83693 -51875 83703 -51841
rect 83737 -51875 83747 -51841
rect 83693 -51895 83747 -51875
rect 83777 -51849 83831 -51765
rect 83777 -51883 83787 -51849
rect 83821 -51883 83831 -51849
rect 83777 -51895 83831 -51883
rect 83861 -51841 83915 -51765
rect 83861 -51875 83871 -51841
rect 83905 -51875 83915 -51841
rect 83861 -51895 83915 -51875
rect 83945 -51848 83997 -51765
rect 83945 -51882 83955 -51848
rect 83989 -51882 83997 -51848
rect 83945 -51895 83997 -51882
rect 84074 -51781 84126 -51765
rect 84074 -51815 84082 -51781
rect 84116 -51815 84126 -51781
rect 84074 -51849 84126 -51815
rect 84074 -51883 84082 -51849
rect 84116 -51883 84126 -51849
rect 84074 -51895 84126 -51883
rect 84156 -51781 84210 -51765
rect 84156 -51815 84166 -51781
rect 84200 -51815 84210 -51781
rect 84156 -51849 84210 -51815
rect 84156 -51883 84166 -51849
rect 84200 -51883 84210 -51849
rect 84156 -51895 84210 -51883
rect 84240 -51849 84294 -51765
rect 84240 -51883 84250 -51849
rect 84284 -51883 84294 -51849
rect 84240 -51895 84294 -51883
rect 84324 -51781 84378 -51765
rect 84324 -51815 84334 -51781
rect 84368 -51815 84378 -51781
rect 84324 -51849 84378 -51815
rect 84324 -51883 84334 -51849
rect 84368 -51883 84378 -51849
rect 84324 -51895 84378 -51883
rect 84408 -51849 84462 -51765
rect 84408 -51883 84418 -51849
rect 84452 -51883 84462 -51849
rect 84408 -51895 84462 -51883
rect 84492 -51781 84546 -51765
rect 84492 -51815 84502 -51781
rect 84536 -51815 84546 -51781
rect 84492 -51849 84546 -51815
rect 84492 -51883 84502 -51849
rect 84536 -51883 84546 -51849
rect 84492 -51895 84546 -51883
rect 84576 -51849 84630 -51765
rect 84576 -51883 84586 -51849
rect 84620 -51883 84630 -51849
rect 84576 -51895 84630 -51883
rect 84660 -51781 84714 -51765
rect 84660 -51815 84670 -51781
rect 84704 -51815 84714 -51781
rect 84660 -51849 84714 -51815
rect 84660 -51883 84670 -51849
rect 84704 -51883 84714 -51849
rect 84660 -51895 84714 -51883
rect 84744 -51849 84798 -51765
rect 84744 -51883 84754 -51849
rect 84788 -51883 84798 -51849
rect 84744 -51895 84798 -51883
rect 84828 -51781 84882 -51765
rect 84828 -51815 84838 -51781
rect 84872 -51815 84882 -51781
rect 84828 -51849 84882 -51815
rect 84828 -51883 84838 -51849
rect 84872 -51883 84882 -51849
rect 84828 -51895 84882 -51883
rect 84912 -51849 84966 -51765
rect 84912 -51883 84922 -51849
rect 84956 -51883 84966 -51849
rect 84912 -51895 84966 -51883
rect 84996 -51781 85050 -51765
rect 84996 -51815 85006 -51781
rect 85040 -51815 85050 -51781
rect 84996 -51849 85050 -51815
rect 84996 -51883 85006 -51849
rect 85040 -51883 85050 -51849
rect 84996 -51895 85050 -51883
rect 85080 -51849 85134 -51765
rect 85080 -51883 85090 -51849
rect 85124 -51883 85134 -51849
rect 85080 -51895 85134 -51883
rect 85164 -51781 85218 -51765
rect 85164 -51815 85174 -51781
rect 85208 -51815 85218 -51781
rect 85164 -51849 85218 -51815
rect 85164 -51883 85174 -51849
rect 85208 -51883 85218 -51849
rect 85164 -51895 85218 -51883
rect 85248 -51849 85302 -51765
rect 85248 -51883 85258 -51849
rect 85292 -51883 85302 -51849
rect 85248 -51895 85302 -51883
rect 85332 -51781 85386 -51765
rect 85332 -51815 85342 -51781
rect 85376 -51815 85386 -51781
rect 85332 -51849 85386 -51815
rect 85332 -51883 85342 -51849
rect 85376 -51883 85386 -51849
rect 85332 -51895 85386 -51883
rect 85416 -51781 85468 -51765
rect 85416 -51815 85426 -51781
rect 85460 -51815 85468 -51781
rect 85416 -51849 85468 -51815
rect 85416 -51883 85426 -51849
rect 85460 -51883 85468 -51849
rect 85416 -51895 85468 -51883
rect 85546 -51781 85598 -51765
rect 85546 -51815 85554 -51781
rect 85588 -51815 85598 -51781
rect 85546 -51849 85598 -51815
rect 85546 -51883 85554 -51849
rect 85588 -51883 85598 -51849
rect 85546 -51895 85598 -51883
rect 85628 -51781 85682 -51765
rect 85628 -51815 85638 -51781
rect 85672 -51815 85682 -51781
rect 85628 -51849 85682 -51815
rect 85628 -51883 85638 -51849
rect 85672 -51883 85682 -51849
rect 85628 -51895 85682 -51883
rect 85712 -51849 85766 -51765
rect 85712 -51883 85722 -51849
rect 85756 -51883 85766 -51849
rect 85712 -51895 85766 -51883
rect 85796 -51781 85850 -51765
rect 85796 -51815 85806 -51781
rect 85840 -51815 85850 -51781
rect 85796 -51849 85850 -51815
rect 85796 -51883 85806 -51849
rect 85840 -51883 85850 -51849
rect 85796 -51895 85850 -51883
rect 85880 -51849 85934 -51765
rect 85880 -51883 85890 -51849
rect 85924 -51883 85934 -51849
rect 85880 -51895 85934 -51883
rect 85964 -51781 86018 -51765
rect 85964 -51815 85974 -51781
rect 86008 -51815 86018 -51781
rect 85964 -51849 86018 -51815
rect 85964 -51883 85974 -51849
rect 86008 -51883 86018 -51849
rect 85964 -51895 86018 -51883
rect 86048 -51849 86102 -51765
rect 86048 -51883 86058 -51849
rect 86092 -51883 86102 -51849
rect 86048 -51895 86102 -51883
rect 86132 -51781 86186 -51765
rect 86132 -51815 86142 -51781
rect 86176 -51815 86186 -51781
rect 86132 -51849 86186 -51815
rect 86132 -51883 86142 -51849
rect 86176 -51883 86186 -51849
rect 86132 -51895 86186 -51883
rect 86216 -51849 86270 -51765
rect 86216 -51883 86226 -51849
rect 86260 -51883 86270 -51849
rect 86216 -51895 86270 -51883
rect 86300 -51781 86354 -51765
rect 86300 -51815 86310 -51781
rect 86344 -51815 86354 -51781
rect 86300 -51849 86354 -51815
rect 86300 -51883 86310 -51849
rect 86344 -51883 86354 -51849
rect 86300 -51895 86354 -51883
rect 86384 -51849 86438 -51765
rect 86384 -51883 86394 -51849
rect 86428 -51883 86438 -51849
rect 86384 -51895 86438 -51883
rect 86468 -51781 86522 -51765
rect 86468 -51815 86478 -51781
rect 86512 -51815 86522 -51781
rect 86468 -51849 86522 -51815
rect 86468 -51883 86478 -51849
rect 86512 -51883 86522 -51849
rect 86468 -51895 86522 -51883
rect 86552 -51849 86606 -51765
rect 86552 -51883 86562 -51849
rect 86596 -51883 86606 -51849
rect 86552 -51895 86606 -51883
rect 86636 -51781 86690 -51765
rect 86636 -51815 86646 -51781
rect 86680 -51815 86690 -51781
rect 86636 -51849 86690 -51815
rect 86636 -51883 86646 -51849
rect 86680 -51883 86690 -51849
rect 86636 -51895 86690 -51883
rect 86720 -51849 86774 -51765
rect 86720 -51883 86730 -51849
rect 86764 -51883 86774 -51849
rect 86720 -51895 86774 -51883
rect 86804 -51781 86858 -51765
rect 86804 -51815 86814 -51781
rect 86848 -51815 86858 -51781
rect 86804 -51849 86858 -51815
rect 86804 -51883 86814 -51849
rect 86848 -51883 86858 -51849
rect 86804 -51895 86858 -51883
rect 86888 -51781 86940 -51765
rect 86888 -51815 86898 -51781
rect 86932 -51815 86940 -51781
rect 86888 -51849 86940 -51815
rect 86888 -51883 86898 -51849
rect 86932 -51883 86940 -51849
rect 86888 -51895 86940 -51883
rect 87018 -51781 87070 -51765
rect 87018 -51815 87026 -51781
rect 87060 -51815 87070 -51781
rect 87018 -51849 87070 -51815
rect 87018 -51883 87026 -51849
rect 87060 -51883 87070 -51849
rect 87018 -51895 87070 -51883
rect 87100 -51781 87154 -51765
rect 87100 -51815 87110 -51781
rect 87144 -51815 87154 -51781
rect 87100 -51849 87154 -51815
rect 87100 -51883 87110 -51849
rect 87144 -51883 87154 -51849
rect 87100 -51895 87154 -51883
rect 87184 -51849 87238 -51765
rect 87184 -51883 87194 -51849
rect 87228 -51883 87238 -51849
rect 87184 -51895 87238 -51883
rect 87268 -51781 87322 -51765
rect 87268 -51815 87278 -51781
rect 87312 -51815 87322 -51781
rect 87268 -51849 87322 -51815
rect 87268 -51883 87278 -51849
rect 87312 -51883 87322 -51849
rect 87268 -51895 87322 -51883
rect 87352 -51849 87406 -51765
rect 87352 -51883 87362 -51849
rect 87396 -51883 87406 -51849
rect 87352 -51895 87406 -51883
rect 87436 -51781 87490 -51765
rect 87436 -51815 87446 -51781
rect 87480 -51815 87490 -51781
rect 87436 -51849 87490 -51815
rect 87436 -51883 87446 -51849
rect 87480 -51883 87490 -51849
rect 87436 -51895 87490 -51883
rect 87520 -51849 87574 -51765
rect 87520 -51883 87530 -51849
rect 87564 -51883 87574 -51849
rect 87520 -51895 87574 -51883
rect 87604 -51781 87658 -51765
rect 87604 -51815 87614 -51781
rect 87648 -51815 87658 -51781
rect 87604 -51849 87658 -51815
rect 87604 -51883 87614 -51849
rect 87648 -51883 87658 -51849
rect 87604 -51895 87658 -51883
rect 87688 -51849 87742 -51765
rect 87688 -51883 87698 -51849
rect 87732 -51883 87742 -51849
rect 87688 -51895 87742 -51883
rect 87772 -51781 87826 -51765
rect 87772 -51815 87782 -51781
rect 87816 -51815 87826 -51781
rect 87772 -51849 87826 -51815
rect 87772 -51883 87782 -51849
rect 87816 -51883 87826 -51849
rect 87772 -51895 87826 -51883
rect 87856 -51849 87910 -51765
rect 87856 -51883 87866 -51849
rect 87900 -51883 87910 -51849
rect 87856 -51895 87910 -51883
rect 87940 -51781 87994 -51765
rect 87940 -51815 87950 -51781
rect 87984 -51815 87994 -51781
rect 87940 -51849 87994 -51815
rect 87940 -51883 87950 -51849
rect 87984 -51883 87994 -51849
rect 87940 -51895 87994 -51883
rect 88024 -51849 88078 -51765
rect 88024 -51883 88034 -51849
rect 88068 -51883 88078 -51849
rect 88024 -51895 88078 -51883
rect 88108 -51781 88162 -51765
rect 88108 -51815 88118 -51781
rect 88152 -51815 88162 -51781
rect 88108 -51849 88162 -51815
rect 88108 -51883 88118 -51849
rect 88152 -51883 88162 -51849
rect 88108 -51895 88162 -51883
rect 88192 -51849 88246 -51765
rect 88192 -51883 88202 -51849
rect 88236 -51883 88246 -51849
rect 88192 -51895 88246 -51883
rect 88276 -51781 88330 -51765
rect 88276 -51815 88286 -51781
rect 88320 -51815 88330 -51781
rect 88276 -51849 88330 -51815
rect 88276 -51883 88286 -51849
rect 88320 -51883 88330 -51849
rect 88276 -51895 88330 -51883
rect 88360 -51781 88412 -51765
rect 88360 -51815 88370 -51781
rect 88404 -51815 88412 -51781
rect 88360 -51849 88412 -51815
rect 88360 -51883 88370 -51849
rect 88404 -51883 88412 -51849
rect 88360 -51895 88412 -51883
rect 88490 -51781 88542 -51765
rect 88490 -51815 88498 -51781
rect 88532 -51815 88542 -51781
rect 88490 -51849 88542 -51815
rect 88490 -51883 88498 -51849
rect 88532 -51883 88542 -51849
rect 88490 -51895 88542 -51883
rect 88572 -51781 88626 -51765
rect 88572 -51815 88582 -51781
rect 88616 -51815 88626 -51781
rect 88572 -51849 88626 -51815
rect 88572 -51883 88582 -51849
rect 88616 -51883 88626 -51849
rect 88572 -51895 88626 -51883
rect 88656 -51849 88710 -51765
rect 88656 -51883 88666 -51849
rect 88700 -51883 88710 -51849
rect 88656 -51895 88710 -51883
rect 88740 -51781 88794 -51765
rect 88740 -51815 88750 -51781
rect 88784 -51815 88794 -51781
rect 88740 -51849 88794 -51815
rect 88740 -51883 88750 -51849
rect 88784 -51883 88794 -51849
rect 88740 -51895 88794 -51883
rect 88824 -51849 88878 -51765
rect 88824 -51883 88834 -51849
rect 88868 -51883 88878 -51849
rect 88824 -51895 88878 -51883
rect 88908 -51781 88962 -51765
rect 88908 -51815 88918 -51781
rect 88952 -51815 88962 -51781
rect 88908 -51849 88962 -51815
rect 88908 -51883 88918 -51849
rect 88952 -51883 88962 -51849
rect 88908 -51895 88962 -51883
rect 88992 -51849 89046 -51765
rect 88992 -51883 89002 -51849
rect 89036 -51883 89046 -51849
rect 88992 -51895 89046 -51883
rect 89076 -51781 89130 -51765
rect 89076 -51815 89086 -51781
rect 89120 -51815 89130 -51781
rect 89076 -51849 89130 -51815
rect 89076 -51883 89086 -51849
rect 89120 -51883 89130 -51849
rect 89076 -51895 89130 -51883
rect 89160 -51849 89214 -51765
rect 89160 -51883 89170 -51849
rect 89204 -51883 89214 -51849
rect 89160 -51895 89214 -51883
rect 89244 -51781 89298 -51765
rect 89244 -51815 89254 -51781
rect 89288 -51815 89298 -51781
rect 89244 -51849 89298 -51815
rect 89244 -51883 89254 -51849
rect 89288 -51883 89298 -51849
rect 89244 -51895 89298 -51883
rect 89328 -51849 89382 -51765
rect 89328 -51883 89338 -51849
rect 89372 -51883 89382 -51849
rect 89328 -51895 89382 -51883
rect 89412 -51781 89466 -51765
rect 89412 -51815 89422 -51781
rect 89456 -51815 89466 -51781
rect 89412 -51849 89466 -51815
rect 89412 -51883 89422 -51849
rect 89456 -51883 89466 -51849
rect 89412 -51895 89466 -51883
rect 89496 -51849 89550 -51765
rect 89496 -51883 89506 -51849
rect 89540 -51883 89550 -51849
rect 89496 -51895 89550 -51883
rect 89580 -51781 89634 -51765
rect 89580 -51815 89590 -51781
rect 89624 -51815 89634 -51781
rect 89580 -51849 89634 -51815
rect 89580 -51883 89590 -51849
rect 89624 -51883 89634 -51849
rect 89580 -51895 89634 -51883
rect 89664 -51849 89718 -51765
rect 89664 -51883 89674 -51849
rect 89708 -51883 89718 -51849
rect 89664 -51895 89718 -51883
rect 89748 -51781 89802 -51765
rect 89748 -51815 89758 -51781
rect 89792 -51815 89802 -51781
rect 89748 -51849 89802 -51815
rect 89748 -51883 89758 -51849
rect 89792 -51883 89802 -51849
rect 89748 -51895 89802 -51883
rect 89832 -51781 89884 -51765
rect 89832 -51815 89842 -51781
rect 89876 -51815 89884 -51781
rect 89832 -51849 89884 -51815
rect 89832 -51883 89842 -51849
rect 89876 -51883 89884 -51849
rect 89832 -51895 89884 -51883
rect 89962 -51781 90014 -51765
rect 89962 -51815 89970 -51781
rect 90004 -51815 90014 -51781
rect 89962 -51849 90014 -51815
rect 89962 -51883 89970 -51849
rect 90004 -51883 90014 -51849
rect 89962 -51895 90014 -51883
rect 90044 -51781 90098 -51765
rect 90044 -51815 90054 -51781
rect 90088 -51815 90098 -51781
rect 90044 -51849 90098 -51815
rect 90044 -51883 90054 -51849
rect 90088 -51883 90098 -51849
rect 90044 -51895 90098 -51883
rect 90128 -51849 90182 -51765
rect 90128 -51883 90138 -51849
rect 90172 -51883 90182 -51849
rect 90128 -51895 90182 -51883
rect 90212 -51781 90266 -51765
rect 90212 -51815 90222 -51781
rect 90256 -51815 90266 -51781
rect 90212 -51849 90266 -51815
rect 90212 -51883 90222 -51849
rect 90256 -51883 90266 -51849
rect 90212 -51895 90266 -51883
rect 90296 -51849 90350 -51765
rect 90296 -51883 90306 -51849
rect 90340 -51883 90350 -51849
rect 90296 -51895 90350 -51883
rect 90380 -51781 90434 -51765
rect 90380 -51815 90390 -51781
rect 90424 -51815 90434 -51781
rect 90380 -51849 90434 -51815
rect 90380 -51883 90390 -51849
rect 90424 -51883 90434 -51849
rect 90380 -51895 90434 -51883
rect 90464 -51849 90518 -51765
rect 90464 -51883 90474 -51849
rect 90508 -51883 90518 -51849
rect 90464 -51895 90518 -51883
rect 90548 -51781 90602 -51765
rect 90548 -51815 90558 -51781
rect 90592 -51815 90602 -51781
rect 90548 -51849 90602 -51815
rect 90548 -51883 90558 -51849
rect 90592 -51883 90602 -51849
rect 90548 -51895 90602 -51883
rect 90632 -51849 90686 -51765
rect 90632 -51883 90642 -51849
rect 90676 -51883 90686 -51849
rect 90632 -51895 90686 -51883
rect 90716 -51781 90770 -51765
rect 90716 -51815 90726 -51781
rect 90760 -51815 90770 -51781
rect 90716 -51849 90770 -51815
rect 90716 -51883 90726 -51849
rect 90760 -51883 90770 -51849
rect 90716 -51895 90770 -51883
rect 90800 -51849 90854 -51765
rect 90800 -51883 90810 -51849
rect 90844 -51883 90854 -51849
rect 90800 -51895 90854 -51883
rect 90884 -51781 90938 -51765
rect 90884 -51815 90894 -51781
rect 90928 -51815 90938 -51781
rect 90884 -51849 90938 -51815
rect 90884 -51883 90894 -51849
rect 90928 -51883 90938 -51849
rect 90884 -51895 90938 -51883
rect 90968 -51849 91022 -51765
rect 90968 -51883 90978 -51849
rect 91012 -51883 91022 -51849
rect 90968 -51895 91022 -51883
rect 91052 -51781 91106 -51765
rect 91052 -51815 91062 -51781
rect 91096 -51815 91106 -51781
rect 91052 -51849 91106 -51815
rect 91052 -51883 91062 -51849
rect 91096 -51883 91106 -51849
rect 91052 -51895 91106 -51883
rect 91136 -51849 91190 -51765
rect 91136 -51883 91146 -51849
rect 91180 -51883 91190 -51849
rect 91136 -51895 91190 -51883
rect 91220 -51781 91274 -51765
rect 91220 -51815 91230 -51781
rect 91264 -51815 91274 -51781
rect 91220 -51849 91274 -51815
rect 91220 -51883 91230 -51849
rect 91264 -51883 91274 -51849
rect 91220 -51895 91274 -51883
rect 91304 -51781 91356 -51765
rect 91304 -51815 91314 -51781
rect 91348 -51815 91356 -51781
rect 91304 -51849 91356 -51815
rect 91304 -51883 91314 -51849
rect 91348 -51883 91356 -51849
rect 91304 -51895 91356 -51883
rect 59946 -52340 60346 -52328
rect 59946 -52374 59958 -52340
rect 60334 -52374 60346 -52340
rect 59946 -52386 60346 -52374
rect 59946 -52448 60346 -52436
rect 59946 -52482 59958 -52448
rect 60334 -52482 60346 -52448
rect 59946 -52494 60346 -52482
rect 78020 -52453 78113 -52437
rect 78020 -52483 78054 -52453
rect 77605 -52513 77657 -52483
rect 77605 -52547 77613 -52513
rect 77647 -52547 77657 -52513
rect 77605 -52567 77657 -52547
rect 77687 -52567 77745 -52483
rect 77775 -52567 77851 -52483
rect 77881 -52567 77947 -52483
rect 77977 -52487 78054 -52483
rect 78088 -52487 78113 -52453
rect 77977 -52521 78113 -52487
rect 77977 -52555 78054 -52521
rect 78088 -52555 78113 -52521
rect 77977 -52567 78113 -52555
rect 78143 -52453 78195 -52437
rect 78143 -52487 78153 -52453
rect 78187 -52487 78195 -52453
rect 78143 -52521 78195 -52487
rect 78143 -52555 78153 -52521
rect 78187 -52555 78195 -52521
rect 78143 -52567 78195 -52555
rect 77605 -52755 77657 -52735
rect 77605 -52789 77613 -52755
rect 77647 -52789 77657 -52755
rect 77605 -52819 77657 -52789
rect 77687 -52819 77745 -52735
rect 77775 -52819 77851 -52735
rect 77881 -52819 77947 -52735
rect 77977 -52747 78113 -52735
rect 77977 -52781 78054 -52747
rect 78088 -52781 78113 -52747
rect 77977 -52815 78113 -52781
rect 77977 -52819 78054 -52815
rect 78020 -52849 78054 -52819
rect 78088 -52849 78113 -52815
rect 78020 -52865 78113 -52849
rect 78143 -52747 78195 -52735
rect 78143 -52781 78153 -52747
rect 78187 -52781 78195 -52747
rect 78143 -52815 78195 -52781
rect 78143 -52849 78153 -52815
rect 78187 -52849 78195 -52815
rect 78143 -52865 78195 -52849
rect 55288 -53158 55488 -53146
rect 55288 -53192 55300 -53158
rect 55476 -53192 55488 -53158
rect 55288 -53204 55488 -53192
rect 55288 -53246 55488 -53234
rect 55288 -53280 55300 -53246
rect 55476 -53280 55488 -53246
rect 55288 -53292 55488 -53280
rect 77879 -53721 77929 -53675
rect 77605 -53759 77657 -53721
rect 77605 -53793 77613 -53759
rect 77647 -53793 77657 -53759
rect 77605 -53805 77657 -53793
rect 77687 -53805 77729 -53721
rect 77759 -53805 77801 -53721
rect 77831 -53743 77929 -53721
rect 77831 -53777 77885 -53743
rect 77919 -53777 77929 -53743
rect 77831 -53805 77929 -53777
rect 77959 -53733 78011 -53675
rect 78293 -53693 78345 -53675
rect 77959 -53767 77969 -53733
rect 78003 -53767 78011 -53733
rect 77959 -53805 78011 -53767
rect 78097 -53731 78153 -53693
rect 78097 -53765 78109 -53731
rect 78143 -53765 78153 -53731
rect 78097 -53777 78153 -53765
rect 78183 -53777 78237 -53693
rect 78267 -53759 78345 -53693
rect 78267 -53777 78301 -53759
rect 78293 -53793 78301 -53777
rect 78335 -53793 78345 -53759
rect 78293 -53805 78345 -53793
rect 78375 -53759 78431 -53675
rect 78886 -53715 78939 -53675
rect 78375 -53793 78385 -53759
rect 78419 -53793 78431 -53759
rect 78375 -53805 78431 -53793
rect 78525 -53735 78577 -53715
rect 78525 -53769 78533 -53735
rect 78567 -53769 78577 -53735
rect 78525 -53799 78577 -53769
rect 78607 -53741 78673 -53715
rect 78607 -53775 78623 -53741
rect 78657 -53775 78673 -53741
rect 78607 -53799 78673 -53775
rect 78703 -53755 78757 -53715
rect 78703 -53789 78713 -53755
rect 78747 -53789 78757 -53755
rect 78703 -53799 78757 -53789
rect 78787 -53741 78841 -53715
rect 78787 -53775 78797 -53741
rect 78831 -53775 78841 -53741
rect 78787 -53799 78841 -53775
rect 78871 -53755 78939 -53715
rect 78871 -53789 78891 -53755
rect 78925 -53789 78939 -53755
rect 78871 -53799 78939 -53789
rect 78886 -53805 78939 -53799
rect 78969 -53717 79023 -53675
rect 78969 -53751 78979 -53717
rect 79013 -53751 79023 -53717
rect 78969 -53805 79023 -53751
rect 53452 -56190 53510 -56178
rect 53452 -56966 53464 -56190
rect 53498 -56966 53510 -56190
rect 53452 -56978 53510 -56966
rect 53630 -56190 53688 -56178
rect 53630 -56966 53642 -56190
rect 53676 -56966 53688 -56190
rect 53630 -56978 53688 -56966
rect 55278 -56252 55336 -56240
rect 55278 -56428 55290 -56252
rect 55324 -56428 55336 -56252
rect 55278 -56440 55336 -56428
rect 55366 -56252 55424 -56240
rect 55366 -56428 55378 -56252
rect 55412 -56428 55424 -56252
rect 55366 -56440 55424 -56428
rect 53930 -56778 54730 -56766
rect 53930 -56812 53942 -56778
rect 54718 -56812 54730 -56778
rect 53930 -56824 54730 -56812
rect 53930 -56956 54730 -56944
rect 53930 -56990 53942 -56956
rect 54718 -56990 54730 -56956
rect 53930 -57002 54730 -56990
rect 55808 -56140 55866 -56128
rect 55808 -56916 55820 -56140
rect 55854 -56916 55866 -56140
rect 55808 -56928 55866 -56916
rect 55986 -56140 56044 -56128
rect 55986 -56916 55998 -56140
rect 56032 -56916 56044 -56140
rect 55986 -56928 56044 -56916
rect 57123 -56500 57175 -56455
rect 53452 -57208 53510 -57196
rect 53452 -57984 53464 -57208
rect 53498 -57984 53510 -57208
rect 53452 -57996 53510 -57984
rect 53630 -57208 53688 -57196
rect 53630 -57984 53642 -57208
rect 53676 -57984 53688 -57208
rect 53630 -57996 53688 -57984
rect 53930 -57184 54730 -57172
rect 53930 -57218 53942 -57184
rect 54718 -57218 54730 -57184
rect 53930 -57230 54730 -57218
rect 53930 -57362 54730 -57350
rect 53930 -57396 53942 -57362
rect 54718 -57396 54730 -57362
rect 53930 -57408 54730 -57396
rect 55268 -57748 55326 -57736
rect 55268 -57924 55280 -57748
rect 55314 -57924 55326 -57748
rect 55268 -57936 55326 -57924
rect 55356 -57748 55414 -57736
rect 55356 -57924 55368 -57748
rect 55402 -57924 55414 -57748
rect 55356 -57936 55414 -57924
rect 55808 -57254 55866 -57242
rect 55808 -58030 55820 -57254
rect 55854 -58030 55866 -57254
rect 55808 -58042 55866 -58030
rect 55986 -57254 56044 -57242
rect 55986 -58030 55998 -57254
rect 56032 -58030 56044 -57254
rect 55986 -58042 56044 -58030
rect 57123 -56534 57131 -56500
rect 57165 -56534 57175 -56500
rect 57123 -56559 57175 -56534
rect 57205 -56513 57263 -56455
rect 57205 -56547 57217 -56513
rect 57251 -56547 57263 -56513
rect 57205 -56559 57263 -56547
rect 57293 -56483 57345 -56455
rect 57293 -56517 57303 -56483
rect 57337 -56517 57345 -56483
rect 57293 -56559 57345 -56517
rect 59946 -56374 60346 -56362
rect 59946 -56408 59958 -56374
rect 60334 -56408 60346 -56374
rect 59946 -56420 60346 -56408
rect 59946 -56482 60346 -56470
rect 59946 -56516 59958 -56482
rect 60334 -56516 60346 -56482
rect 59946 -56528 60346 -56516
rect 59490 -56782 59548 -56770
rect 59490 -56850 59502 -56782
rect 59476 -56920 59502 -56850
rect 59490 -56958 59502 -56920
rect 59536 -56958 59548 -56782
rect 59490 -56970 59548 -56958
rect 59578 -56782 59636 -56770
rect 59578 -56958 59590 -56782
rect 59624 -56958 59636 -56782
rect 59578 -56970 59636 -56958
rect 59806 -56782 59864 -56770
rect 59806 -56958 59818 -56782
rect 59852 -56958 59864 -56782
rect 59806 -56970 59864 -56958
rect 59894 -56782 59952 -56770
rect 59894 -56958 59906 -56782
rect 59940 -56958 59952 -56782
rect 59894 -56970 59952 -56958
rect 60191 -56973 60321 -56965
rect 60191 -57007 60203 -56973
rect 60237 -57007 60321 -56973
rect 60191 -57017 60321 -57007
rect 61131 -56973 61261 -56965
rect 61131 -57007 61215 -56973
rect 61249 -57007 61261 -56973
rect 61131 -57017 61261 -57007
rect 60191 -57057 60321 -57047
rect 60191 -57091 60211 -57057
rect 60245 -57091 60321 -57057
rect 60191 -57101 60321 -57091
rect 61131 -57057 61261 -57047
rect 61131 -57091 61207 -57057
rect 61241 -57091 61261 -57057
rect 61131 -57101 61261 -57091
rect 57123 -57654 57175 -57629
rect 57123 -57688 57131 -57654
rect 57165 -57688 57175 -57654
rect 57123 -57733 57175 -57688
rect 57205 -57641 57263 -57629
rect 57205 -57675 57217 -57641
rect 57251 -57675 57263 -57641
rect 57205 -57733 57263 -57675
rect 57293 -57671 57345 -57629
rect 57293 -57705 57303 -57671
rect 57337 -57705 57345 -57671
rect 57293 -57733 57345 -57705
rect 60191 -57141 60321 -57131
rect 59489 -57295 59547 -57283
rect 59489 -57471 59501 -57295
rect 59535 -57471 59547 -57295
rect 59489 -57483 59547 -57471
rect 59577 -57295 59635 -57283
rect 59577 -57471 59589 -57295
rect 59623 -57471 59635 -57295
rect 59577 -57483 59635 -57471
rect 60191 -57175 60203 -57141
rect 60237 -57175 60321 -57141
rect 60191 -57185 60321 -57175
rect 61131 -57141 61261 -57131
rect 61131 -57175 61215 -57141
rect 61249 -57175 61261 -57141
rect 61131 -57185 61261 -57175
rect 59805 -57295 59863 -57283
rect 59805 -57471 59817 -57295
rect 59851 -57471 59863 -57295
rect 59805 -57483 59863 -57471
rect 59893 -57295 59951 -57283
rect 59893 -57471 59905 -57295
rect 59939 -57471 59951 -57295
rect 59893 -57483 59951 -57471
rect 60191 -57225 60321 -57215
rect 60191 -57259 60211 -57225
rect 60245 -57259 60321 -57225
rect 60191 -57269 60321 -57259
rect 61131 -57225 61261 -57215
rect 61131 -57259 61207 -57225
rect 61241 -57259 61261 -57225
rect 61131 -57269 61261 -57259
rect 60191 -57309 60321 -57299
rect 60191 -57343 60204 -57309
rect 60238 -57343 60321 -57309
rect 60191 -57351 60321 -57343
rect 61131 -57309 61261 -57299
rect 61131 -57343 61214 -57309
rect 61248 -57343 61261 -57309
rect 61131 -57351 61261 -57343
rect 59946 -57740 60346 -57728
rect 59946 -57774 59958 -57740
rect 60334 -57774 60346 -57740
rect 59946 -57786 60346 -57774
rect 59946 -57848 60346 -57836
rect 59946 -57882 59958 -57848
rect 60334 -57882 60346 -57848
rect 59946 -57894 60346 -57882
rect 55288 -58558 55488 -58546
rect 55288 -58592 55300 -58558
rect 55476 -58592 55488 -58558
rect 55288 -58604 55488 -58592
rect 55288 -58646 55488 -58634
rect 55288 -58680 55300 -58646
rect 55476 -58680 55488 -58646
rect 55288 -58692 55488 -58680
rect 53452 -61590 53510 -61578
rect 53452 -62366 53464 -61590
rect 53498 -62366 53510 -61590
rect 53452 -62378 53510 -62366
rect 53630 -61590 53688 -61578
rect 53630 -62366 53642 -61590
rect 53676 -62366 53688 -61590
rect 53630 -62378 53688 -62366
rect 55278 -61652 55336 -61640
rect 55278 -61828 55290 -61652
rect 55324 -61828 55336 -61652
rect 55278 -61840 55336 -61828
rect 55366 -61652 55424 -61640
rect 55366 -61828 55378 -61652
rect 55412 -61828 55424 -61652
rect 55366 -61840 55424 -61828
rect 53930 -62178 54730 -62166
rect 53930 -62212 53942 -62178
rect 54718 -62212 54730 -62178
rect 53930 -62224 54730 -62212
rect 53930 -62356 54730 -62344
rect 53930 -62390 53942 -62356
rect 54718 -62390 54730 -62356
rect 53930 -62402 54730 -62390
rect 55808 -61540 55866 -61528
rect 55808 -62316 55820 -61540
rect 55854 -62316 55866 -61540
rect 55808 -62328 55866 -62316
rect 55986 -61540 56044 -61528
rect 55986 -62316 55998 -61540
rect 56032 -62316 56044 -61540
rect 55986 -62328 56044 -62316
rect 57123 -61900 57175 -61855
rect 53452 -62608 53510 -62596
rect 53452 -63384 53464 -62608
rect 53498 -63384 53510 -62608
rect 53452 -63396 53510 -63384
rect 53630 -62608 53688 -62596
rect 53630 -63384 53642 -62608
rect 53676 -63384 53688 -62608
rect 53630 -63396 53688 -63384
rect 53930 -62584 54730 -62572
rect 53930 -62618 53942 -62584
rect 54718 -62618 54730 -62584
rect 53930 -62630 54730 -62618
rect 53930 -62762 54730 -62750
rect 53930 -62796 53942 -62762
rect 54718 -62796 54730 -62762
rect 53930 -62808 54730 -62796
rect 55268 -63148 55326 -63136
rect 55268 -63324 55280 -63148
rect 55314 -63324 55326 -63148
rect 55268 -63336 55326 -63324
rect 55356 -63148 55414 -63136
rect 55356 -63324 55368 -63148
rect 55402 -63324 55414 -63148
rect 55356 -63336 55414 -63324
rect 55808 -62654 55866 -62642
rect 55808 -63430 55820 -62654
rect 55854 -63430 55866 -62654
rect 55808 -63442 55866 -63430
rect 55986 -62654 56044 -62642
rect 55986 -63430 55998 -62654
rect 56032 -63430 56044 -62654
rect 55986 -63442 56044 -63430
rect 57123 -61934 57131 -61900
rect 57165 -61934 57175 -61900
rect 57123 -61959 57175 -61934
rect 57205 -61913 57263 -61855
rect 57205 -61947 57217 -61913
rect 57251 -61947 57263 -61913
rect 57205 -61959 57263 -61947
rect 57293 -61883 57345 -61855
rect 57293 -61917 57303 -61883
rect 57337 -61917 57345 -61883
rect 57293 -61959 57345 -61917
rect 59946 -61774 60346 -61762
rect 59946 -61808 59958 -61774
rect 60334 -61808 60346 -61774
rect 59946 -61820 60346 -61808
rect 59946 -61882 60346 -61870
rect 59946 -61916 59958 -61882
rect 60334 -61916 60346 -61882
rect 59946 -61928 60346 -61916
rect 59490 -62182 59548 -62170
rect 59490 -62250 59502 -62182
rect 59476 -62320 59502 -62250
rect 59490 -62358 59502 -62320
rect 59536 -62358 59548 -62182
rect 59490 -62370 59548 -62358
rect 59578 -62182 59636 -62170
rect 59578 -62358 59590 -62182
rect 59624 -62358 59636 -62182
rect 59578 -62370 59636 -62358
rect 59806 -62182 59864 -62170
rect 59806 -62358 59818 -62182
rect 59852 -62358 59864 -62182
rect 59806 -62370 59864 -62358
rect 59894 -62182 59952 -62170
rect 59894 -62358 59906 -62182
rect 59940 -62358 59952 -62182
rect 59894 -62370 59952 -62358
rect 60191 -62373 60321 -62365
rect 60191 -62407 60203 -62373
rect 60237 -62407 60321 -62373
rect 60191 -62417 60321 -62407
rect 61131 -62373 61261 -62365
rect 61131 -62407 61215 -62373
rect 61249 -62407 61261 -62373
rect 61131 -62417 61261 -62407
rect 60191 -62457 60321 -62447
rect 60191 -62491 60211 -62457
rect 60245 -62491 60321 -62457
rect 60191 -62501 60321 -62491
rect 61131 -62457 61261 -62447
rect 61131 -62491 61207 -62457
rect 61241 -62491 61261 -62457
rect 61131 -62501 61261 -62491
rect 57123 -63054 57175 -63029
rect 57123 -63088 57131 -63054
rect 57165 -63088 57175 -63054
rect 57123 -63133 57175 -63088
rect 57205 -63041 57263 -63029
rect 57205 -63075 57217 -63041
rect 57251 -63075 57263 -63041
rect 57205 -63133 57263 -63075
rect 57293 -63071 57345 -63029
rect 57293 -63105 57303 -63071
rect 57337 -63105 57345 -63071
rect 57293 -63133 57345 -63105
rect 60191 -62541 60321 -62531
rect 59489 -62695 59547 -62683
rect 59489 -62871 59501 -62695
rect 59535 -62871 59547 -62695
rect 59489 -62883 59547 -62871
rect 59577 -62695 59635 -62683
rect 59577 -62871 59589 -62695
rect 59623 -62871 59635 -62695
rect 59577 -62883 59635 -62871
rect 60191 -62575 60203 -62541
rect 60237 -62575 60321 -62541
rect 60191 -62585 60321 -62575
rect 61131 -62541 61261 -62531
rect 61131 -62575 61215 -62541
rect 61249 -62575 61261 -62541
rect 61131 -62585 61261 -62575
rect 59805 -62695 59863 -62683
rect 59805 -62871 59817 -62695
rect 59851 -62871 59863 -62695
rect 59805 -62883 59863 -62871
rect 59893 -62695 59951 -62683
rect 59893 -62871 59905 -62695
rect 59939 -62871 59951 -62695
rect 59893 -62883 59951 -62871
rect 60191 -62625 60321 -62615
rect 60191 -62659 60211 -62625
rect 60245 -62659 60321 -62625
rect 60191 -62669 60321 -62659
rect 61131 -62625 61261 -62615
rect 61131 -62659 61207 -62625
rect 61241 -62659 61261 -62625
rect 61131 -62669 61261 -62659
rect 60191 -62709 60321 -62699
rect 60191 -62743 60204 -62709
rect 60238 -62743 60321 -62709
rect 60191 -62751 60321 -62743
rect 61131 -62709 61261 -62699
rect 61131 -62743 61214 -62709
rect 61248 -62743 61261 -62709
rect 61131 -62751 61261 -62743
rect 59946 -63140 60346 -63128
rect 59946 -63174 59958 -63140
rect 60334 -63174 60346 -63140
rect 59946 -63186 60346 -63174
rect 59946 -63248 60346 -63236
rect 59946 -63282 59958 -63248
rect 60334 -63282 60346 -63248
rect 59946 -63294 60346 -63282
rect 55288 -63958 55488 -63946
rect 55288 -63992 55300 -63958
rect 55476 -63992 55488 -63958
rect 55288 -64004 55488 -63992
rect 55288 -64046 55488 -64034
rect 55288 -64080 55300 -64046
rect 55476 -64080 55488 -64046
rect 55288 -64092 55488 -64080
rect 53452 -66990 53510 -66978
rect 53452 -67766 53464 -66990
rect 53498 -67766 53510 -66990
rect 53452 -67778 53510 -67766
rect 53630 -66990 53688 -66978
rect 53630 -67766 53642 -66990
rect 53676 -67766 53688 -66990
rect 53630 -67778 53688 -67766
rect 55278 -67052 55336 -67040
rect 55278 -67228 55290 -67052
rect 55324 -67228 55336 -67052
rect 55278 -67240 55336 -67228
rect 55366 -67052 55424 -67040
rect 55366 -67228 55378 -67052
rect 55412 -67228 55424 -67052
rect 55366 -67240 55424 -67228
rect 53930 -67578 54730 -67566
rect 53930 -67612 53942 -67578
rect 54718 -67612 54730 -67578
rect 53930 -67624 54730 -67612
rect 53930 -67756 54730 -67744
rect 53930 -67790 53942 -67756
rect 54718 -67790 54730 -67756
rect 53930 -67802 54730 -67790
rect 55808 -66940 55866 -66928
rect 55808 -67716 55820 -66940
rect 55854 -67716 55866 -66940
rect 55808 -67728 55866 -67716
rect 55986 -66940 56044 -66928
rect 55986 -67716 55998 -66940
rect 56032 -67716 56044 -66940
rect 55986 -67728 56044 -67716
rect 57123 -67300 57175 -67255
rect 53452 -68008 53510 -67996
rect 53452 -68784 53464 -68008
rect 53498 -68784 53510 -68008
rect 53452 -68796 53510 -68784
rect 53630 -68008 53688 -67996
rect 53630 -68784 53642 -68008
rect 53676 -68784 53688 -68008
rect 53630 -68796 53688 -68784
rect 53930 -67984 54730 -67972
rect 53930 -68018 53942 -67984
rect 54718 -68018 54730 -67984
rect 53930 -68030 54730 -68018
rect 53930 -68162 54730 -68150
rect 53930 -68196 53942 -68162
rect 54718 -68196 54730 -68162
rect 53930 -68208 54730 -68196
rect 55268 -68548 55326 -68536
rect 55268 -68724 55280 -68548
rect 55314 -68724 55326 -68548
rect 55268 -68736 55326 -68724
rect 55356 -68548 55414 -68536
rect 55356 -68724 55368 -68548
rect 55402 -68724 55414 -68548
rect 55356 -68736 55414 -68724
rect 55808 -68054 55866 -68042
rect 55808 -68830 55820 -68054
rect 55854 -68830 55866 -68054
rect 55808 -68842 55866 -68830
rect 55986 -68054 56044 -68042
rect 55986 -68830 55998 -68054
rect 56032 -68830 56044 -68054
rect 55986 -68842 56044 -68830
rect 57123 -67334 57131 -67300
rect 57165 -67334 57175 -67300
rect 57123 -67359 57175 -67334
rect 57205 -67313 57263 -67255
rect 57205 -67347 57217 -67313
rect 57251 -67347 57263 -67313
rect 57205 -67359 57263 -67347
rect 57293 -67283 57345 -67255
rect 57293 -67317 57303 -67283
rect 57337 -67317 57345 -67283
rect 57293 -67359 57345 -67317
rect 59946 -67174 60346 -67162
rect 59946 -67208 59958 -67174
rect 60334 -67208 60346 -67174
rect 59946 -67220 60346 -67208
rect 59946 -67282 60346 -67270
rect 59946 -67316 59958 -67282
rect 60334 -67316 60346 -67282
rect 59946 -67328 60346 -67316
rect 59490 -67582 59548 -67570
rect 59490 -67650 59502 -67582
rect 59476 -67720 59502 -67650
rect 59490 -67758 59502 -67720
rect 59536 -67758 59548 -67582
rect 59490 -67770 59548 -67758
rect 59578 -67582 59636 -67570
rect 59578 -67758 59590 -67582
rect 59624 -67758 59636 -67582
rect 59578 -67770 59636 -67758
rect 59806 -67582 59864 -67570
rect 59806 -67758 59818 -67582
rect 59852 -67758 59864 -67582
rect 59806 -67770 59864 -67758
rect 59894 -67582 59952 -67570
rect 59894 -67758 59906 -67582
rect 59940 -67758 59952 -67582
rect 59894 -67770 59952 -67758
rect 60191 -67773 60321 -67765
rect 60191 -67807 60203 -67773
rect 60237 -67807 60321 -67773
rect 60191 -67817 60321 -67807
rect 61131 -67773 61261 -67765
rect 61131 -67807 61215 -67773
rect 61249 -67807 61261 -67773
rect 61131 -67817 61261 -67807
rect 60191 -67857 60321 -67847
rect 60191 -67891 60211 -67857
rect 60245 -67891 60321 -67857
rect 60191 -67901 60321 -67891
rect 61131 -67857 61261 -67847
rect 61131 -67891 61207 -67857
rect 61241 -67891 61261 -67857
rect 61131 -67901 61261 -67891
rect 57123 -68454 57175 -68429
rect 57123 -68488 57131 -68454
rect 57165 -68488 57175 -68454
rect 57123 -68533 57175 -68488
rect 57205 -68441 57263 -68429
rect 57205 -68475 57217 -68441
rect 57251 -68475 57263 -68441
rect 57205 -68533 57263 -68475
rect 57293 -68471 57345 -68429
rect 57293 -68505 57303 -68471
rect 57337 -68505 57345 -68471
rect 57293 -68533 57345 -68505
rect 60191 -67941 60321 -67931
rect 59489 -68095 59547 -68083
rect 59489 -68271 59501 -68095
rect 59535 -68271 59547 -68095
rect 59489 -68283 59547 -68271
rect 59577 -68095 59635 -68083
rect 59577 -68271 59589 -68095
rect 59623 -68271 59635 -68095
rect 59577 -68283 59635 -68271
rect 60191 -67975 60203 -67941
rect 60237 -67975 60321 -67941
rect 60191 -67985 60321 -67975
rect 61131 -67941 61261 -67931
rect 61131 -67975 61215 -67941
rect 61249 -67975 61261 -67941
rect 61131 -67985 61261 -67975
rect 59805 -68095 59863 -68083
rect 59805 -68271 59817 -68095
rect 59851 -68271 59863 -68095
rect 59805 -68283 59863 -68271
rect 59893 -68095 59951 -68083
rect 59893 -68271 59905 -68095
rect 59939 -68271 59951 -68095
rect 59893 -68283 59951 -68271
rect 60191 -68025 60321 -68015
rect 60191 -68059 60211 -68025
rect 60245 -68059 60321 -68025
rect 60191 -68069 60321 -68059
rect 61131 -68025 61261 -68015
rect 61131 -68059 61207 -68025
rect 61241 -68059 61261 -68025
rect 61131 -68069 61261 -68059
rect 60191 -68109 60321 -68099
rect 60191 -68143 60204 -68109
rect 60238 -68143 60321 -68109
rect 60191 -68151 60321 -68143
rect 61131 -68109 61261 -68099
rect 61131 -68143 61214 -68109
rect 61248 -68143 61261 -68109
rect 61131 -68151 61261 -68143
rect 59946 -68540 60346 -68528
rect 59946 -68574 59958 -68540
rect 60334 -68574 60346 -68540
rect 59946 -68586 60346 -68574
rect 59946 -68648 60346 -68636
rect 59946 -68682 59958 -68648
rect 60334 -68682 60346 -68648
rect 59946 -68694 60346 -68682
rect 55288 -69358 55488 -69346
rect 55288 -69392 55300 -69358
rect 55476 -69392 55488 -69358
rect 55288 -69404 55488 -69392
rect 55288 -69446 55488 -69434
rect 55288 -69480 55300 -69446
rect 55476 -69480 55488 -69446
rect 55288 -69492 55488 -69480
rect 53452 -72390 53510 -72378
rect 53452 -73166 53464 -72390
rect 53498 -73166 53510 -72390
rect 53452 -73178 53510 -73166
rect 53630 -72390 53688 -72378
rect 53630 -73166 53642 -72390
rect 53676 -73166 53688 -72390
rect 53630 -73178 53688 -73166
rect 55278 -72452 55336 -72440
rect 55278 -72628 55290 -72452
rect 55324 -72628 55336 -72452
rect 55278 -72640 55336 -72628
rect 55366 -72452 55424 -72440
rect 55366 -72628 55378 -72452
rect 55412 -72628 55424 -72452
rect 55366 -72640 55424 -72628
rect 53930 -72978 54730 -72966
rect 53930 -73012 53942 -72978
rect 54718 -73012 54730 -72978
rect 53930 -73024 54730 -73012
rect 53930 -73156 54730 -73144
rect 53930 -73190 53942 -73156
rect 54718 -73190 54730 -73156
rect 53930 -73202 54730 -73190
rect 55808 -72340 55866 -72328
rect 55808 -73116 55820 -72340
rect 55854 -73116 55866 -72340
rect 55808 -73128 55866 -73116
rect 55986 -72340 56044 -72328
rect 55986 -73116 55998 -72340
rect 56032 -73116 56044 -72340
rect 55986 -73128 56044 -73116
rect 57123 -72700 57175 -72655
rect 53452 -73408 53510 -73396
rect 53452 -74184 53464 -73408
rect 53498 -74184 53510 -73408
rect 53452 -74196 53510 -74184
rect 53630 -73408 53688 -73396
rect 53630 -74184 53642 -73408
rect 53676 -74184 53688 -73408
rect 53630 -74196 53688 -74184
rect 53930 -73384 54730 -73372
rect 53930 -73418 53942 -73384
rect 54718 -73418 54730 -73384
rect 53930 -73430 54730 -73418
rect 53930 -73562 54730 -73550
rect 53930 -73596 53942 -73562
rect 54718 -73596 54730 -73562
rect 53930 -73608 54730 -73596
rect 55268 -73948 55326 -73936
rect 55268 -74124 55280 -73948
rect 55314 -74124 55326 -73948
rect 55268 -74136 55326 -74124
rect 55356 -73948 55414 -73936
rect 55356 -74124 55368 -73948
rect 55402 -74124 55414 -73948
rect 55356 -74136 55414 -74124
rect 55808 -73454 55866 -73442
rect 55808 -74230 55820 -73454
rect 55854 -74230 55866 -73454
rect 55808 -74242 55866 -74230
rect 55986 -73454 56044 -73442
rect 55986 -74230 55998 -73454
rect 56032 -74230 56044 -73454
rect 55986 -74242 56044 -74230
rect 57123 -72734 57131 -72700
rect 57165 -72734 57175 -72700
rect 57123 -72759 57175 -72734
rect 57205 -72713 57263 -72655
rect 57205 -72747 57217 -72713
rect 57251 -72747 57263 -72713
rect 57205 -72759 57263 -72747
rect 57293 -72683 57345 -72655
rect 57293 -72717 57303 -72683
rect 57337 -72717 57345 -72683
rect 57293 -72759 57345 -72717
rect 59946 -72574 60346 -72562
rect 59946 -72608 59958 -72574
rect 60334 -72608 60346 -72574
rect 59946 -72620 60346 -72608
rect 59946 -72682 60346 -72670
rect 59946 -72716 59958 -72682
rect 60334 -72716 60346 -72682
rect 59946 -72728 60346 -72716
rect 59490 -72982 59548 -72970
rect 59490 -73050 59502 -72982
rect 59476 -73120 59502 -73050
rect 59490 -73158 59502 -73120
rect 59536 -73158 59548 -72982
rect 59490 -73170 59548 -73158
rect 59578 -72982 59636 -72970
rect 59578 -73158 59590 -72982
rect 59624 -73158 59636 -72982
rect 59578 -73170 59636 -73158
rect 59806 -72982 59864 -72970
rect 59806 -73158 59818 -72982
rect 59852 -73158 59864 -72982
rect 59806 -73170 59864 -73158
rect 59894 -72982 59952 -72970
rect 59894 -73158 59906 -72982
rect 59940 -73158 59952 -72982
rect 59894 -73170 59952 -73158
rect 60191 -73173 60321 -73165
rect 60191 -73207 60203 -73173
rect 60237 -73207 60321 -73173
rect 60191 -73217 60321 -73207
rect 61131 -73173 61261 -73165
rect 61131 -73207 61215 -73173
rect 61249 -73207 61261 -73173
rect 61131 -73217 61261 -73207
rect 60191 -73257 60321 -73247
rect 60191 -73291 60211 -73257
rect 60245 -73291 60321 -73257
rect 60191 -73301 60321 -73291
rect 61131 -73257 61261 -73247
rect 61131 -73291 61207 -73257
rect 61241 -73291 61261 -73257
rect 61131 -73301 61261 -73291
rect 57123 -73854 57175 -73829
rect 57123 -73888 57131 -73854
rect 57165 -73888 57175 -73854
rect 57123 -73933 57175 -73888
rect 57205 -73841 57263 -73829
rect 57205 -73875 57217 -73841
rect 57251 -73875 57263 -73841
rect 57205 -73933 57263 -73875
rect 57293 -73871 57345 -73829
rect 57293 -73905 57303 -73871
rect 57337 -73905 57345 -73871
rect 57293 -73933 57345 -73905
rect 60191 -73341 60321 -73331
rect 59489 -73495 59547 -73483
rect 59489 -73671 59501 -73495
rect 59535 -73671 59547 -73495
rect 59489 -73683 59547 -73671
rect 59577 -73495 59635 -73483
rect 59577 -73671 59589 -73495
rect 59623 -73671 59635 -73495
rect 59577 -73683 59635 -73671
rect 60191 -73375 60203 -73341
rect 60237 -73375 60321 -73341
rect 60191 -73385 60321 -73375
rect 61131 -73341 61261 -73331
rect 61131 -73375 61215 -73341
rect 61249 -73375 61261 -73341
rect 61131 -73385 61261 -73375
rect 59805 -73495 59863 -73483
rect 59805 -73671 59817 -73495
rect 59851 -73671 59863 -73495
rect 59805 -73683 59863 -73671
rect 59893 -73495 59951 -73483
rect 59893 -73671 59905 -73495
rect 59939 -73671 59951 -73495
rect 59893 -73683 59951 -73671
rect 60191 -73425 60321 -73415
rect 60191 -73459 60211 -73425
rect 60245 -73459 60321 -73425
rect 60191 -73469 60321 -73459
rect 61131 -73425 61261 -73415
rect 61131 -73459 61207 -73425
rect 61241 -73459 61261 -73425
rect 61131 -73469 61261 -73459
rect 60191 -73509 60321 -73499
rect 60191 -73543 60204 -73509
rect 60238 -73543 60321 -73509
rect 60191 -73551 60321 -73543
rect 61131 -73509 61261 -73499
rect 61131 -73543 61214 -73509
rect 61248 -73543 61261 -73509
rect 61131 -73551 61261 -73543
rect 59946 -73940 60346 -73928
rect 59946 -73974 59958 -73940
rect 60334 -73974 60346 -73940
rect 59946 -73986 60346 -73974
rect 59946 -74048 60346 -74036
rect 59946 -74082 59958 -74048
rect 60334 -74082 60346 -74048
rect 59946 -74094 60346 -74082
rect 55288 -74758 55488 -74746
rect 55288 -74792 55300 -74758
rect 55476 -74792 55488 -74758
rect 55288 -74804 55488 -74792
rect 55288 -74846 55488 -74834
rect 55288 -74880 55300 -74846
rect 55476 -74880 55488 -74846
rect 55288 -74892 55488 -74880
rect 53452 -77790 53510 -77778
rect 53452 -78566 53464 -77790
rect 53498 -78566 53510 -77790
rect 53452 -78578 53510 -78566
rect 53630 -77790 53688 -77778
rect 53630 -78566 53642 -77790
rect 53676 -78566 53688 -77790
rect 53630 -78578 53688 -78566
rect 55278 -77852 55336 -77840
rect 55278 -78028 55290 -77852
rect 55324 -78028 55336 -77852
rect 55278 -78040 55336 -78028
rect 55366 -77852 55424 -77840
rect 55366 -78028 55378 -77852
rect 55412 -78028 55424 -77852
rect 55366 -78040 55424 -78028
rect 53930 -78378 54730 -78366
rect 53930 -78412 53942 -78378
rect 54718 -78412 54730 -78378
rect 53930 -78424 54730 -78412
rect 53930 -78556 54730 -78544
rect 53930 -78590 53942 -78556
rect 54718 -78590 54730 -78556
rect 53930 -78602 54730 -78590
rect 55808 -77740 55866 -77728
rect 55808 -78516 55820 -77740
rect 55854 -78516 55866 -77740
rect 55808 -78528 55866 -78516
rect 55986 -77740 56044 -77728
rect 55986 -78516 55998 -77740
rect 56032 -78516 56044 -77740
rect 55986 -78528 56044 -78516
rect 57123 -78100 57175 -78055
rect 53452 -78808 53510 -78796
rect 53452 -79584 53464 -78808
rect 53498 -79584 53510 -78808
rect 53452 -79596 53510 -79584
rect 53630 -78808 53688 -78796
rect 53630 -79584 53642 -78808
rect 53676 -79584 53688 -78808
rect 53630 -79596 53688 -79584
rect 53930 -78784 54730 -78772
rect 53930 -78818 53942 -78784
rect 54718 -78818 54730 -78784
rect 53930 -78830 54730 -78818
rect 53930 -78962 54730 -78950
rect 53930 -78996 53942 -78962
rect 54718 -78996 54730 -78962
rect 53930 -79008 54730 -78996
rect 55268 -79348 55326 -79336
rect 55268 -79524 55280 -79348
rect 55314 -79524 55326 -79348
rect 55268 -79536 55326 -79524
rect 55356 -79348 55414 -79336
rect 55356 -79524 55368 -79348
rect 55402 -79524 55414 -79348
rect 55356 -79536 55414 -79524
rect 55808 -78854 55866 -78842
rect 55808 -79630 55820 -78854
rect 55854 -79630 55866 -78854
rect 55808 -79642 55866 -79630
rect 55986 -78854 56044 -78842
rect 55986 -79630 55998 -78854
rect 56032 -79630 56044 -78854
rect 55986 -79642 56044 -79630
rect 57123 -78134 57131 -78100
rect 57165 -78134 57175 -78100
rect 57123 -78159 57175 -78134
rect 57205 -78113 57263 -78055
rect 57205 -78147 57217 -78113
rect 57251 -78147 57263 -78113
rect 57205 -78159 57263 -78147
rect 57293 -78083 57345 -78055
rect 57293 -78117 57303 -78083
rect 57337 -78117 57345 -78083
rect 57293 -78159 57345 -78117
rect 59946 -77974 60346 -77962
rect 59946 -78008 59958 -77974
rect 60334 -78008 60346 -77974
rect 59946 -78020 60346 -78008
rect 59946 -78082 60346 -78070
rect 59946 -78116 59958 -78082
rect 60334 -78116 60346 -78082
rect 59946 -78128 60346 -78116
rect 59490 -78382 59548 -78370
rect 59490 -78450 59502 -78382
rect 59476 -78520 59502 -78450
rect 59490 -78558 59502 -78520
rect 59536 -78558 59548 -78382
rect 59490 -78570 59548 -78558
rect 59578 -78382 59636 -78370
rect 59578 -78558 59590 -78382
rect 59624 -78558 59636 -78382
rect 59578 -78570 59636 -78558
rect 59806 -78382 59864 -78370
rect 59806 -78558 59818 -78382
rect 59852 -78558 59864 -78382
rect 59806 -78570 59864 -78558
rect 59894 -78382 59952 -78370
rect 59894 -78558 59906 -78382
rect 59940 -78558 59952 -78382
rect 59894 -78570 59952 -78558
rect 60191 -78573 60321 -78565
rect 60191 -78607 60203 -78573
rect 60237 -78607 60321 -78573
rect 60191 -78617 60321 -78607
rect 61131 -78573 61261 -78565
rect 61131 -78607 61215 -78573
rect 61249 -78607 61261 -78573
rect 61131 -78617 61261 -78607
rect 60191 -78657 60321 -78647
rect 60191 -78691 60211 -78657
rect 60245 -78691 60321 -78657
rect 60191 -78701 60321 -78691
rect 61131 -78657 61261 -78647
rect 61131 -78691 61207 -78657
rect 61241 -78691 61261 -78657
rect 61131 -78701 61261 -78691
rect 57123 -79254 57175 -79229
rect 57123 -79288 57131 -79254
rect 57165 -79288 57175 -79254
rect 57123 -79333 57175 -79288
rect 57205 -79241 57263 -79229
rect 57205 -79275 57217 -79241
rect 57251 -79275 57263 -79241
rect 57205 -79333 57263 -79275
rect 57293 -79271 57345 -79229
rect 57293 -79305 57303 -79271
rect 57337 -79305 57345 -79271
rect 57293 -79333 57345 -79305
rect 60191 -78741 60321 -78731
rect 59489 -78895 59547 -78883
rect 59489 -79071 59501 -78895
rect 59535 -79071 59547 -78895
rect 59489 -79083 59547 -79071
rect 59577 -78895 59635 -78883
rect 59577 -79071 59589 -78895
rect 59623 -79071 59635 -78895
rect 59577 -79083 59635 -79071
rect 60191 -78775 60203 -78741
rect 60237 -78775 60321 -78741
rect 60191 -78785 60321 -78775
rect 61131 -78741 61261 -78731
rect 61131 -78775 61215 -78741
rect 61249 -78775 61261 -78741
rect 61131 -78785 61261 -78775
rect 59805 -78895 59863 -78883
rect 59805 -79071 59817 -78895
rect 59851 -79071 59863 -78895
rect 59805 -79083 59863 -79071
rect 59893 -78895 59951 -78883
rect 59893 -79071 59905 -78895
rect 59939 -79071 59951 -78895
rect 59893 -79083 59951 -79071
rect 60191 -78825 60321 -78815
rect 60191 -78859 60211 -78825
rect 60245 -78859 60321 -78825
rect 60191 -78869 60321 -78859
rect 61131 -78825 61261 -78815
rect 61131 -78859 61207 -78825
rect 61241 -78859 61261 -78825
rect 61131 -78869 61261 -78859
rect 60191 -78909 60321 -78899
rect 60191 -78943 60204 -78909
rect 60238 -78943 60321 -78909
rect 60191 -78951 60321 -78943
rect 61131 -78909 61261 -78899
rect 61131 -78943 61214 -78909
rect 61248 -78943 61261 -78909
rect 61131 -78951 61261 -78943
rect 59946 -79340 60346 -79328
rect 59946 -79374 59958 -79340
rect 60334 -79374 60346 -79340
rect 59946 -79386 60346 -79374
rect 59946 -79448 60346 -79436
rect 59946 -79482 59958 -79448
rect 60334 -79482 60346 -79448
rect 59946 -79494 60346 -79482
rect 55288 -80158 55488 -80146
rect 55288 -80192 55300 -80158
rect 55476 -80192 55488 -80158
rect 55288 -80204 55488 -80192
rect 55288 -80246 55488 -80234
rect 55288 -80280 55300 -80246
rect 55476 -80280 55488 -80246
rect 55288 -80292 55488 -80280
rect 53452 -83190 53510 -83178
rect 53452 -83966 53464 -83190
rect 53498 -83966 53510 -83190
rect 53452 -83978 53510 -83966
rect 53630 -83190 53688 -83178
rect 53630 -83966 53642 -83190
rect 53676 -83966 53688 -83190
rect 53630 -83978 53688 -83966
rect 55278 -83252 55336 -83240
rect 55278 -83428 55290 -83252
rect 55324 -83428 55336 -83252
rect 55278 -83440 55336 -83428
rect 55366 -83252 55424 -83240
rect 55366 -83428 55378 -83252
rect 55412 -83428 55424 -83252
rect 55366 -83440 55424 -83428
rect 53930 -83778 54730 -83766
rect 53930 -83812 53942 -83778
rect 54718 -83812 54730 -83778
rect 53930 -83824 54730 -83812
rect 53930 -83956 54730 -83944
rect 53930 -83990 53942 -83956
rect 54718 -83990 54730 -83956
rect 53930 -84002 54730 -83990
rect 55808 -83140 55866 -83128
rect 55808 -83916 55820 -83140
rect 55854 -83916 55866 -83140
rect 55808 -83928 55866 -83916
rect 55986 -83140 56044 -83128
rect 55986 -83916 55998 -83140
rect 56032 -83916 56044 -83140
rect 55986 -83928 56044 -83916
rect 57123 -83500 57175 -83455
rect 53452 -84208 53510 -84196
rect 53452 -84984 53464 -84208
rect 53498 -84984 53510 -84208
rect 53452 -84996 53510 -84984
rect 53630 -84208 53688 -84196
rect 53630 -84984 53642 -84208
rect 53676 -84984 53688 -84208
rect 53630 -84996 53688 -84984
rect 53930 -84184 54730 -84172
rect 53930 -84218 53942 -84184
rect 54718 -84218 54730 -84184
rect 53930 -84230 54730 -84218
rect 53930 -84362 54730 -84350
rect 53930 -84396 53942 -84362
rect 54718 -84396 54730 -84362
rect 53930 -84408 54730 -84396
rect 55268 -84748 55326 -84736
rect 55268 -84924 55280 -84748
rect 55314 -84924 55326 -84748
rect 55268 -84936 55326 -84924
rect 55356 -84748 55414 -84736
rect 55356 -84924 55368 -84748
rect 55402 -84924 55414 -84748
rect 55356 -84936 55414 -84924
rect 55808 -84254 55866 -84242
rect 55808 -85030 55820 -84254
rect 55854 -85030 55866 -84254
rect 55808 -85042 55866 -85030
rect 55986 -84254 56044 -84242
rect 55986 -85030 55998 -84254
rect 56032 -85030 56044 -84254
rect 55986 -85042 56044 -85030
rect 57123 -83534 57131 -83500
rect 57165 -83534 57175 -83500
rect 57123 -83559 57175 -83534
rect 57205 -83513 57263 -83455
rect 57205 -83547 57217 -83513
rect 57251 -83547 57263 -83513
rect 57205 -83559 57263 -83547
rect 57293 -83483 57345 -83455
rect 57293 -83517 57303 -83483
rect 57337 -83517 57345 -83483
rect 57293 -83559 57345 -83517
rect 59946 -83374 60346 -83362
rect 59946 -83408 59958 -83374
rect 60334 -83408 60346 -83374
rect 59946 -83420 60346 -83408
rect 59946 -83482 60346 -83470
rect 59946 -83516 59958 -83482
rect 60334 -83516 60346 -83482
rect 59946 -83528 60346 -83516
rect 59490 -83782 59548 -83770
rect 59490 -83850 59502 -83782
rect 59476 -83920 59502 -83850
rect 59490 -83958 59502 -83920
rect 59536 -83958 59548 -83782
rect 59490 -83970 59548 -83958
rect 59578 -83782 59636 -83770
rect 59578 -83958 59590 -83782
rect 59624 -83958 59636 -83782
rect 59578 -83970 59636 -83958
rect 59806 -83782 59864 -83770
rect 59806 -83958 59818 -83782
rect 59852 -83958 59864 -83782
rect 59806 -83970 59864 -83958
rect 59894 -83782 59952 -83770
rect 59894 -83958 59906 -83782
rect 59940 -83958 59952 -83782
rect 59894 -83970 59952 -83958
rect 60191 -83973 60321 -83965
rect 60191 -84007 60203 -83973
rect 60237 -84007 60321 -83973
rect 60191 -84017 60321 -84007
rect 61131 -83973 61261 -83965
rect 61131 -84007 61215 -83973
rect 61249 -84007 61261 -83973
rect 61131 -84017 61261 -84007
rect 60191 -84057 60321 -84047
rect 60191 -84091 60211 -84057
rect 60245 -84091 60321 -84057
rect 60191 -84101 60321 -84091
rect 61131 -84057 61261 -84047
rect 61131 -84091 61207 -84057
rect 61241 -84091 61261 -84057
rect 61131 -84101 61261 -84091
rect 57123 -84654 57175 -84629
rect 57123 -84688 57131 -84654
rect 57165 -84688 57175 -84654
rect 57123 -84733 57175 -84688
rect 57205 -84641 57263 -84629
rect 57205 -84675 57217 -84641
rect 57251 -84675 57263 -84641
rect 57205 -84733 57263 -84675
rect 57293 -84671 57345 -84629
rect 57293 -84705 57303 -84671
rect 57337 -84705 57345 -84671
rect 57293 -84733 57345 -84705
rect 60191 -84141 60321 -84131
rect 59489 -84295 59547 -84283
rect 59489 -84471 59501 -84295
rect 59535 -84471 59547 -84295
rect 59489 -84483 59547 -84471
rect 59577 -84295 59635 -84283
rect 59577 -84471 59589 -84295
rect 59623 -84471 59635 -84295
rect 59577 -84483 59635 -84471
rect 60191 -84175 60203 -84141
rect 60237 -84175 60321 -84141
rect 60191 -84185 60321 -84175
rect 61131 -84141 61261 -84131
rect 61131 -84175 61215 -84141
rect 61249 -84175 61261 -84141
rect 61131 -84185 61261 -84175
rect 59805 -84295 59863 -84283
rect 59805 -84471 59817 -84295
rect 59851 -84471 59863 -84295
rect 59805 -84483 59863 -84471
rect 59893 -84295 59951 -84283
rect 59893 -84471 59905 -84295
rect 59939 -84471 59951 -84295
rect 59893 -84483 59951 -84471
rect 60191 -84225 60321 -84215
rect 60191 -84259 60211 -84225
rect 60245 -84259 60321 -84225
rect 60191 -84269 60321 -84259
rect 61131 -84225 61261 -84215
rect 61131 -84259 61207 -84225
rect 61241 -84259 61261 -84225
rect 61131 -84269 61261 -84259
rect 60191 -84309 60321 -84299
rect 60191 -84343 60204 -84309
rect 60238 -84343 60321 -84309
rect 60191 -84351 60321 -84343
rect 61131 -84309 61261 -84299
rect 61131 -84343 61214 -84309
rect 61248 -84343 61261 -84309
rect 61131 -84351 61261 -84343
rect 59946 -84740 60346 -84728
rect 59946 -84774 59958 -84740
rect 60334 -84774 60346 -84740
rect 59946 -84786 60346 -84774
rect 59946 -84848 60346 -84836
rect 59946 -84882 59958 -84848
rect 60334 -84882 60346 -84848
rect 59946 -84894 60346 -84882
rect 55288 -85558 55488 -85546
rect 55288 -85592 55300 -85558
rect 55476 -85592 55488 -85558
rect 55288 -85604 55488 -85592
rect 55288 -85646 55488 -85634
rect 55288 -85680 55300 -85646
rect 55476 -85680 55488 -85646
rect 55288 -85692 55488 -85680
<< pdiff >>
rect 54079 -1672 54879 -1660
rect 54079 -1706 54091 -1672
rect 54867 -1706 54879 -1672
rect 54079 -1718 54879 -1706
rect 54079 -1800 54879 -1788
rect 54079 -1834 54091 -1800
rect 54867 -1834 54879 -1800
rect 54079 -1846 54879 -1834
rect 54079 -2028 54879 -2016
rect 54079 -2062 54091 -2028
rect 54867 -2062 54879 -2028
rect 54079 -2074 54879 -2062
rect 54079 -2156 54879 -2144
rect 54079 -2190 54091 -2156
rect 54867 -2190 54879 -2156
rect 54079 -2202 54879 -2190
rect 57123 -2129 57175 -2109
rect 57123 -2163 57131 -2129
rect 57165 -2163 57175 -2129
rect 57123 -2197 57175 -2163
rect 57123 -2231 57131 -2197
rect 57165 -2231 57175 -2197
rect 57123 -2267 57175 -2231
rect 57205 -2129 57263 -2109
rect 57205 -2163 57217 -2129
rect 57251 -2163 57263 -2129
rect 57205 -2197 57263 -2163
rect 57205 -2231 57217 -2197
rect 57251 -2231 57263 -2197
rect 57205 -2267 57263 -2231
rect 57293 -2129 57345 -2109
rect 57293 -2163 57303 -2129
rect 57337 -2163 57345 -2129
rect 57293 -2210 57345 -2163
rect 57293 -2244 57303 -2210
rect 57337 -2244 57345 -2210
rect 57293 -2267 57345 -2244
rect 59113 -2047 59513 -2035
rect 59113 -2081 59125 -2047
rect 59501 -2081 59513 -2047
rect 59113 -2093 59513 -2081
rect 59113 -2155 59513 -2143
rect 59113 -2189 59125 -2155
rect 59501 -2189 59513 -2155
rect 59113 -2201 59513 -2189
rect 59113 -2263 59513 -2251
rect 59113 -2297 59125 -2263
rect 59501 -2297 59513 -2263
rect 59113 -2309 59513 -2297
rect 54069 -3988 54869 -3976
rect 54069 -4022 54081 -3988
rect 54857 -4022 54869 -3988
rect 54069 -4034 54869 -4022
rect 54069 -4116 54869 -4104
rect 54069 -4150 54081 -4116
rect 54857 -4150 54869 -4116
rect 54069 -4162 54869 -4150
rect 56418 -2699 56476 -2687
rect 56418 -3475 56430 -2699
rect 56464 -3475 56476 -2699
rect 56418 -3487 56476 -3475
rect 56546 -2699 56604 -2687
rect 56546 -3475 56558 -2699
rect 56592 -3475 56604 -2699
rect 56546 -3487 56604 -3475
rect 59032 -2571 59090 -2559
rect 59032 -2947 59044 -2571
rect 59078 -2947 59090 -2571
rect 59032 -2959 59090 -2947
rect 59150 -2571 59208 -2559
rect 59150 -2947 59162 -2571
rect 59196 -2947 59208 -2571
rect 59150 -2959 59208 -2947
rect 60441 -2973 60641 -2965
rect 60441 -3007 60459 -2973
rect 60493 -3007 60527 -2973
rect 60561 -3007 60595 -2973
rect 60629 -3007 60641 -2973
rect 60441 -3017 60641 -3007
rect 60811 -2973 61011 -2965
rect 60811 -3007 60823 -2973
rect 60857 -3007 60891 -2973
rect 60925 -3007 60959 -2973
rect 60993 -3007 61011 -2973
rect 60811 -3017 61011 -3007
rect 60441 -3057 60641 -3047
rect 60441 -3091 60459 -3057
rect 60493 -3091 60527 -3057
rect 60561 -3091 60595 -3057
rect 60629 -3091 60641 -3057
rect 60441 -3101 60641 -3091
rect 60811 -3057 61011 -3047
rect 60811 -3091 60823 -3057
rect 60857 -3091 60891 -3057
rect 60925 -3091 60959 -3057
rect 60993 -3091 61011 -3057
rect 60811 -3101 61011 -3091
rect 59032 -3301 59090 -3289
rect 59032 -3677 59044 -3301
rect 59078 -3677 59090 -3301
rect 59032 -3689 59090 -3677
rect 59150 -3301 59208 -3289
rect 59150 -3677 59162 -3301
rect 59196 -3677 59208 -3301
rect 59150 -3689 59208 -3677
rect 60441 -3141 60641 -3131
rect 60441 -3175 60527 -3141
rect 60561 -3175 60595 -3141
rect 60629 -3175 60641 -3141
rect 60441 -3185 60641 -3175
rect 60811 -3141 61011 -3131
rect 60811 -3175 60823 -3141
rect 60857 -3175 60891 -3141
rect 60925 -3175 61011 -3141
rect 60811 -3185 61011 -3175
rect 60441 -3225 60641 -3215
rect 60441 -3259 60459 -3225
rect 60493 -3259 60527 -3225
rect 60561 -3259 60595 -3225
rect 60629 -3259 60641 -3225
rect 60441 -3269 60641 -3259
rect 60811 -3225 61011 -3215
rect 60811 -3259 60823 -3225
rect 60857 -3259 60891 -3225
rect 60925 -3259 60959 -3225
rect 60993 -3259 61011 -3225
rect 60811 -3269 61011 -3259
rect 60441 -3309 60641 -3299
rect 60441 -3343 60595 -3309
rect 60629 -3343 60641 -3309
rect 60441 -3351 60641 -3343
rect 60811 -3309 61011 -3299
rect 60811 -3343 60823 -3309
rect 60857 -3343 61011 -3309
rect 60811 -3351 61011 -3343
rect 57123 -3957 57175 -3921
rect 57123 -3991 57131 -3957
rect 57165 -3991 57175 -3957
rect 57123 -4025 57175 -3991
rect 57123 -4059 57131 -4025
rect 57165 -4059 57175 -4025
rect 57123 -4079 57175 -4059
rect 57205 -3957 57263 -3921
rect 57205 -3991 57217 -3957
rect 57251 -3991 57263 -3957
rect 57205 -4025 57263 -3991
rect 57205 -4059 57217 -4025
rect 57251 -4059 57263 -4025
rect 57205 -4079 57263 -4059
rect 57293 -3944 57345 -3921
rect 57293 -3978 57303 -3944
rect 57337 -3978 57345 -3944
rect 57293 -4025 57345 -3978
rect 57293 -4059 57303 -4025
rect 57337 -4059 57345 -4025
rect 57293 -4079 57345 -4059
rect 59113 -3954 59513 -3942
rect 59113 -3988 59125 -3954
rect 59501 -3988 59513 -3954
rect 59113 -4000 59513 -3988
rect 59113 -4062 59513 -4050
rect 59113 -4096 59125 -4062
rect 59501 -4096 59513 -4062
rect 59113 -4108 59513 -4096
rect 59113 -4170 59513 -4158
rect 59113 -4204 59125 -4170
rect 59501 -4204 59513 -4170
rect 59113 -4216 59513 -4204
rect 54069 -4344 54869 -4332
rect 54069 -4378 54081 -4344
rect 54857 -4378 54869 -4344
rect 54069 -4390 54869 -4378
rect 54069 -4472 54869 -4460
rect 54069 -4506 54081 -4472
rect 54857 -4506 54869 -4472
rect 54069 -4518 54869 -4506
rect 54079 -7072 54879 -7060
rect 54079 -7106 54091 -7072
rect 54867 -7106 54879 -7072
rect 54079 -7118 54879 -7106
rect 54079 -7200 54879 -7188
rect 54079 -7234 54091 -7200
rect 54867 -7234 54879 -7200
rect 54079 -7246 54879 -7234
rect 20834 -7868 20892 -7856
rect 20834 -11644 20846 -7868
rect 20880 -11644 20892 -7868
rect 20834 -11656 20892 -11644
rect 21092 -7868 21150 -7856
rect 21092 -11644 21104 -7868
rect 21138 -11644 21150 -7868
rect 21092 -11656 21150 -11644
rect 21320 -7868 21378 -7856
rect 21320 -11644 21332 -7868
rect 21366 -11644 21378 -7868
rect 21320 -11656 21378 -11644
rect 21578 -7868 21636 -7856
rect 21578 -11644 21590 -7868
rect 21624 -11644 21636 -7868
rect 21578 -11656 21636 -11644
rect 21806 -7868 21864 -7856
rect 21806 -11644 21818 -7868
rect 21852 -11644 21864 -7868
rect 21806 -11656 21864 -11644
rect 22064 -7868 22122 -7856
rect 22064 -11644 22076 -7868
rect 22110 -11644 22122 -7868
rect 22064 -11656 22122 -11644
rect 54079 -7428 54879 -7416
rect 54079 -7462 54091 -7428
rect 54867 -7462 54879 -7428
rect 54079 -7474 54879 -7462
rect 54079 -7556 54879 -7544
rect 54079 -7590 54091 -7556
rect 54867 -7590 54879 -7556
rect 54079 -7602 54879 -7590
rect 57123 -7529 57175 -7509
rect 57123 -7563 57131 -7529
rect 57165 -7563 57175 -7529
rect 57123 -7597 57175 -7563
rect 57123 -7631 57131 -7597
rect 57165 -7631 57175 -7597
rect 57123 -7667 57175 -7631
rect 57205 -7529 57263 -7509
rect 57205 -7563 57217 -7529
rect 57251 -7563 57263 -7529
rect 57205 -7597 57263 -7563
rect 57205 -7631 57217 -7597
rect 57251 -7631 57263 -7597
rect 57205 -7667 57263 -7631
rect 57293 -7529 57345 -7509
rect 57293 -7563 57303 -7529
rect 57337 -7563 57345 -7529
rect 57293 -7610 57345 -7563
rect 57293 -7644 57303 -7610
rect 57337 -7644 57345 -7610
rect 57293 -7667 57345 -7644
rect 59113 -7447 59513 -7435
rect 59113 -7481 59125 -7447
rect 59501 -7481 59513 -7447
rect 59113 -7493 59513 -7481
rect 59113 -7555 59513 -7543
rect 59113 -7589 59125 -7555
rect 59501 -7589 59513 -7555
rect 59113 -7601 59513 -7589
rect 59113 -7663 59513 -7651
rect 59113 -7697 59125 -7663
rect 59501 -7697 59513 -7663
rect 59113 -7709 59513 -7697
rect 54069 -9388 54869 -9376
rect 54069 -9422 54081 -9388
rect 54857 -9422 54869 -9388
rect 54069 -9434 54869 -9422
rect 54069 -9516 54869 -9504
rect 54069 -9550 54081 -9516
rect 54857 -9550 54869 -9516
rect 54069 -9562 54869 -9550
rect 56418 -8099 56476 -8087
rect 56418 -8875 56430 -8099
rect 56464 -8875 56476 -8099
rect 56418 -8887 56476 -8875
rect 56546 -8099 56604 -8087
rect 56546 -8875 56558 -8099
rect 56592 -8875 56604 -8099
rect 56546 -8887 56604 -8875
rect 59032 -7971 59090 -7959
rect 59032 -8347 59044 -7971
rect 59078 -8347 59090 -7971
rect 59032 -8359 59090 -8347
rect 59150 -7971 59208 -7959
rect 59150 -8347 59162 -7971
rect 59196 -8347 59208 -7971
rect 59150 -8359 59208 -8347
rect 60441 -8373 60641 -8365
rect 60441 -8407 60459 -8373
rect 60493 -8407 60527 -8373
rect 60561 -8407 60595 -8373
rect 60629 -8407 60641 -8373
rect 60441 -8417 60641 -8407
rect 60811 -8373 61011 -8365
rect 60811 -8407 60823 -8373
rect 60857 -8407 60891 -8373
rect 60925 -8407 60959 -8373
rect 60993 -8407 61011 -8373
rect 60811 -8417 61011 -8407
rect 60441 -8457 60641 -8447
rect 60441 -8491 60459 -8457
rect 60493 -8491 60527 -8457
rect 60561 -8491 60595 -8457
rect 60629 -8491 60641 -8457
rect 60441 -8501 60641 -8491
rect 60811 -8457 61011 -8447
rect 60811 -8491 60823 -8457
rect 60857 -8491 60891 -8457
rect 60925 -8491 60959 -8457
rect 60993 -8491 61011 -8457
rect 60811 -8501 61011 -8491
rect 59032 -8701 59090 -8689
rect 59032 -9077 59044 -8701
rect 59078 -9077 59090 -8701
rect 59032 -9089 59090 -9077
rect 59150 -8701 59208 -8689
rect 59150 -9077 59162 -8701
rect 59196 -9077 59208 -8701
rect 59150 -9089 59208 -9077
rect 60441 -8541 60641 -8531
rect 60441 -8575 60527 -8541
rect 60561 -8575 60595 -8541
rect 60629 -8575 60641 -8541
rect 60441 -8585 60641 -8575
rect 60811 -8541 61011 -8531
rect 60811 -8575 60823 -8541
rect 60857 -8575 60891 -8541
rect 60925 -8575 61011 -8541
rect 60811 -8585 61011 -8575
rect 60441 -8625 60641 -8615
rect 60441 -8659 60459 -8625
rect 60493 -8659 60527 -8625
rect 60561 -8659 60595 -8625
rect 60629 -8659 60641 -8625
rect 60441 -8669 60641 -8659
rect 60811 -8625 61011 -8615
rect 60811 -8659 60823 -8625
rect 60857 -8659 60891 -8625
rect 60925 -8659 60959 -8625
rect 60993 -8659 61011 -8625
rect 60811 -8669 61011 -8659
rect 60441 -8709 60641 -8699
rect 60441 -8743 60595 -8709
rect 60629 -8743 60641 -8709
rect 60441 -8751 60641 -8743
rect 60811 -8709 61011 -8699
rect 60811 -8743 60823 -8709
rect 60857 -8743 61011 -8709
rect 60811 -8751 61011 -8743
rect 57123 -9357 57175 -9321
rect 57123 -9391 57131 -9357
rect 57165 -9391 57175 -9357
rect 57123 -9425 57175 -9391
rect 57123 -9459 57131 -9425
rect 57165 -9459 57175 -9425
rect 57123 -9479 57175 -9459
rect 57205 -9357 57263 -9321
rect 57205 -9391 57217 -9357
rect 57251 -9391 57263 -9357
rect 57205 -9425 57263 -9391
rect 57205 -9459 57217 -9425
rect 57251 -9459 57263 -9425
rect 57205 -9479 57263 -9459
rect 57293 -9344 57345 -9321
rect 57293 -9378 57303 -9344
rect 57337 -9378 57345 -9344
rect 57293 -9425 57345 -9378
rect 57293 -9459 57303 -9425
rect 57337 -9459 57345 -9425
rect 57293 -9479 57345 -9459
rect 59113 -9354 59513 -9342
rect 59113 -9388 59125 -9354
rect 59501 -9388 59513 -9354
rect 59113 -9400 59513 -9388
rect 59113 -9462 59513 -9450
rect 59113 -9496 59125 -9462
rect 59501 -9496 59513 -9462
rect 59113 -9508 59513 -9496
rect 59113 -9570 59513 -9558
rect 59113 -9604 59125 -9570
rect 59501 -9604 59513 -9570
rect 59113 -9616 59513 -9604
rect 54069 -9744 54869 -9732
rect 54069 -9778 54081 -9744
rect 54857 -9778 54869 -9744
rect 54069 -9790 54869 -9778
rect 54069 -9872 54869 -9860
rect 54069 -9906 54081 -9872
rect 54857 -9906 54869 -9872
rect 54069 -9918 54869 -9906
rect 54079 -12472 54879 -12460
rect 54079 -12506 54091 -12472
rect 54867 -12506 54879 -12472
rect 54079 -12518 54879 -12506
rect 54079 -12600 54879 -12588
rect 54079 -12634 54091 -12600
rect 54867 -12634 54879 -12600
rect 54079 -12646 54879 -12634
rect 54079 -12828 54879 -12816
rect 54079 -12862 54091 -12828
rect 54867 -12862 54879 -12828
rect 54079 -12874 54879 -12862
rect 54079 -12956 54879 -12944
rect 54079 -12990 54091 -12956
rect 54867 -12990 54879 -12956
rect 54079 -13002 54879 -12990
rect 57123 -12929 57175 -12909
rect 57123 -12963 57131 -12929
rect 57165 -12963 57175 -12929
rect 57123 -12997 57175 -12963
rect 57123 -13031 57131 -12997
rect 57165 -13031 57175 -12997
rect 57123 -13067 57175 -13031
rect 57205 -12929 57263 -12909
rect 57205 -12963 57217 -12929
rect 57251 -12963 57263 -12929
rect 57205 -12997 57263 -12963
rect 57205 -13031 57217 -12997
rect 57251 -13031 57263 -12997
rect 57205 -13067 57263 -13031
rect 57293 -12929 57345 -12909
rect 57293 -12963 57303 -12929
rect 57337 -12963 57345 -12929
rect 57293 -13010 57345 -12963
rect 57293 -13044 57303 -13010
rect 57337 -13044 57345 -13010
rect 57293 -13067 57345 -13044
rect 59113 -12847 59513 -12835
rect 59113 -12881 59125 -12847
rect 59501 -12881 59513 -12847
rect 59113 -12893 59513 -12881
rect 59113 -12955 59513 -12943
rect 59113 -12989 59125 -12955
rect 59501 -12989 59513 -12955
rect 59113 -13001 59513 -12989
rect 59113 -13063 59513 -13051
rect 59113 -13097 59125 -13063
rect 59501 -13097 59513 -13063
rect 59113 -13109 59513 -13097
rect 54069 -14788 54869 -14776
rect 54069 -14822 54081 -14788
rect 54857 -14822 54869 -14788
rect 54069 -14834 54869 -14822
rect 54069 -14916 54869 -14904
rect 54069 -14950 54081 -14916
rect 54857 -14950 54869 -14916
rect 54069 -14962 54869 -14950
rect 56418 -13499 56476 -13487
rect 56418 -14275 56430 -13499
rect 56464 -14275 56476 -13499
rect 56418 -14287 56476 -14275
rect 56546 -13499 56604 -13487
rect 56546 -14275 56558 -13499
rect 56592 -14275 56604 -13499
rect 56546 -14287 56604 -14275
rect 59032 -13371 59090 -13359
rect 59032 -13747 59044 -13371
rect 59078 -13747 59090 -13371
rect 59032 -13759 59090 -13747
rect 59150 -13371 59208 -13359
rect 59150 -13747 59162 -13371
rect 59196 -13747 59208 -13371
rect 59150 -13759 59208 -13747
rect 60441 -13773 60641 -13765
rect 60441 -13807 60459 -13773
rect 60493 -13807 60527 -13773
rect 60561 -13807 60595 -13773
rect 60629 -13807 60641 -13773
rect 60441 -13817 60641 -13807
rect 60811 -13773 61011 -13765
rect 60811 -13807 60823 -13773
rect 60857 -13807 60891 -13773
rect 60925 -13807 60959 -13773
rect 60993 -13807 61011 -13773
rect 60811 -13817 61011 -13807
rect 60441 -13857 60641 -13847
rect 60441 -13891 60459 -13857
rect 60493 -13891 60527 -13857
rect 60561 -13891 60595 -13857
rect 60629 -13891 60641 -13857
rect 60441 -13901 60641 -13891
rect 60811 -13857 61011 -13847
rect 60811 -13891 60823 -13857
rect 60857 -13891 60891 -13857
rect 60925 -13891 60959 -13857
rect 60993 -13891 61011 -13857
rect 60811 -13901 61011 -13891
rect 59032 -14101 59090 -14089
rect 59032 -14477 59044 -14101
rect 59078 -14477 59090 -14101
rect 59032 -14489 59090 -14477
rect 59150 -14101 59208 -14089
rect 59150 -14477 59162 -14101
rect 59196 -14477 59208 -14101
rect 59150 -14489 59208 -14477
rect 60441 -13941 60641 -13931
rect 60441 -13975 60527 -13941
rect 60561 -13975 60595 -13941
rect 60629 -13975 60641 -13941
rect 60441 -13985 60641 -13975
rect 60811 -13941 61011 -13931
rect 60811 -13975 60823 -13941
rect 60857 -13975 60891 -13941
rect 60925 -13975 61011 -13941
rect 60811 -13985 61011 -13975
rect 60441 -14025 60641 -14015
rect 60441 -14059 60459 -14025
rect 60493 -14059 60527 -14025
rect 60561 -14059 60595 -14025
rect 60629 -14059 60641 -14025
rect 60441 -14069 60641 -14059
rect 60811 -14025 61011 -14015
rect 60811 -14059 60823 -14025
rect 60857 -14059 60891 -14025
rect 60925 -14059 60959 -14025
rect 60993 -14059 61011 -14025
rect 60811 -14069 61011 -14059
rect 60441 -14109 60641 -14099
rect 60441 -14143 60595 -14109
rect 60629 -14143 60641 -14109
rect 60441 -14151 60641 -14143
rect 60811 -14109 61011 -14099
rect 60811 -14143 60823 -14109
rect 60857 -14143 61011 -14109
rect 60811 -14151 61011 -14143
rect 57123 -14757 57175 -14721
rect 57123 -14791 57131 -14757
rect 57165 -14791 57175 -14757
rect 57123 -14825 57175 -14791
rect 57123 -14859 57131 -14825
rect 57165 -14859 57175 -14825
rect 57123 -14879 57175 -14859
rect 57205 -14757 57263 -14721
rect 57205 -14791 57217 -14757
rect 57251 -14791 57263 -14757
rect 57205 -14825 57263 -14791
rect 57205 -14859 57217 -14825
rect 57251 -14859 57263 -14825
rect 57205 -14879 57263 -14859
rect 57293 -14744 57345 -14721
rect 57293 -14778 57303 -14744
rect 57337 -14778 57345 -14744
rect 57293 -14825 57345 -14778
rect 57293 -14859 57303 -14825
rect 57337 -14859 57345 -14825
rect 57293 -14879 57345 -14859
rect 59113 -14754 59513 -14742
rect 59113 -14788 59125 -14754
rect 59501 -14788 59513 -14754
rect 59113 -14800 59513 -14788
rect 59113 -14862 59513 -14850
rect 59113 -14896 59125 -14862
rect 59501 -14896 59513 -14862
rect 59113 -14908 59513 -14896
rect 59113 -14970 59513 -14958
rect 59113 -15004 59125 -14970
rect 59501 -15004 59513 -14970
rect 59113 -15016 59513 -15004
rect 54069 -15144 54869 -15132
rect 54069 -15178 54081 -15144
rect 54857 -15178 54869 -15144
rect 54069 -15190 54869 -15178
rect 54069 -15272 54869 -15260
rect 54069 -15306 54081 -15272
rect 54857 -15306 54869 -15272
rect 54069 -15318 54869 -15306
rect 54079 -17872 54879 -17860
rect 54079 -17906 54091 -17872
rect 54867 -17906 54879 -17872
rect 54079 -17918 54879 -17906
rect 54079 -18000 54879 -17988
rect 54079 -18034 54091 -18000
rect 54867 -18034 54879 -18000
rect 54079 -18046 54879 -18034
rect 54079 -18228 54879 -18216
rect 54079 -18262 54091 -18228
rect 54867 -18262 54879 -18228
rect 54079 -18274 54879 -18262
rect 54079 -18356 54879 -18344
rect 54079 -18390 54091 -18356
rect 54867 -18390 54879 -18356
rect 54079 -18402 54879 -18390
rect 57123 -18329 57175 -18309
rect 57123 -18363 57131 -18329
rect 57165 -18363 57175 -18329
rect 57123 -18397 57175 -18363
rect 57123 -18431 57131 -18397
rect 57165 -18431 57175 -18397
rect 57123 -18467 57175 -18431
rect 57205 -18329 57263 -18309
rect 57205 -18363 57217 -18329
rect 57251 -18363 57263 -18329
rect 57205 -18397 57263 -18363
rect 57205 -18431 57217 -18397
rect 57251 -18431 57263 -18397
rect 57205 -18467 57263 -18431
rect 57293 -18329 57345 -18309
rect 57293 -18363 57303 -18329
rect 57337 -18363 57345 -18329
rect 57293 -18410 57345 -18363
rect 57293 -18444 57303 -18410
rect 57337 -18444 57345 -18410
rect 57293 -18467 57345 -18444
rect 59113 -18247 59513 -18235
rect 59113 -18281 59125 -18247
rect 59501 -18281 59513 -18247
rect 59113 -18293 59513 -18281
rect 59113 -18355 59513 -18343
rect 59113 -18389 59125 -18355
rect 59501 -18389 59513 -18355
rect 59113 -18401 59513 -18389
rect 59113 -18463 59513 -18451
rect 59113 -18497 59125 -18463
rect 59501 -18497 59513 -18463
rect 59113 -18509 59513 -18497
rect 54069 -20188 54869 -20176
rect 54069 -20222 54081 -20188
rect 54857 -20222 54869 -20188
rect 54069 -20234 54869 -20222
rect 54069 -20316 54869 -20304
rect 54069 -20350 54081 -20316
rect 54857 -20350 54869 -20316
rect 54069 -20362 54869 -20350
rect 56418 -18899 56476 -18887
rect 56418 -19675 56430 -18899
rect 56464 -19675 56476 -18899
rect 56418 -19687 56476 -19675
rect 56546 -18899 56604 -18887
rect 56546 -19675 56558 -18899
rect 56592 -19675 56604 -18899
rect 56546 -19687 56604 -19675
rect 59032 -18771 59090 -18759
rect 59032 -19147 59044 -18771
rect 59078 -19147 59090 -18771
rect 59032 -19159 59090 -19147
rect 59150 -18771 59208 -18759
rect 59150 -19147 59162 -18771
rect 59196 -19147 59208 -18771
rect 59150 -19159 59208 -19147
rect 60441 -19173 60641 -19165
rect 60441 -19207 60459 -19173
rect 60493 -19207 60527 -19173
rect 60561 -19207 60595 -19173
rect 60629 -19207 60641 -19173
rect 60441 -19217 60641 -19207
rect 60811 -19173 61011 -19165
rect 60811 -19207 60823 -19173
rect 60857 -19207 60891 -19173
rect 60925 -19207 60959 -19173
rect 60993 -19207 61011 -19173
rect 60811 -19217 61011 -19207
rect 60441 -19257 60641 -19247
rect 60441 -19291 60459 -19257
rect 60493 -19291 60527 -19257
rect 60561 -19291 60595 -19257
rect 60629 -19291 60641 -19257
rect 60441 -19301 60641 -19291
rect 60811 -19257 61011 -19247
rect 60811 -19291 60823 -19257
rect 60857 -19291 60891 -19257
rect 60925 -19291 60959 -19257
rect 60993 -19291 61011 -19257
rect 60811 -19301 61011 -19291
rect 59032 -19501 59090 -19489
rect 59032 -19877 59044 -19501
rect 59078 -19877 59090 -19501
rect 59032 -19889 59090 -19877
rect 59150 -19501 59208 -19489
rect 59150 -19877 59162 -19501
rect 59196 -19877 59208 -19501
rect 59150 -19889 59208 -19877
rect 60441 -19341 60641 -19331
rect 60441 -19375 60527 -19341
rect 60561 -19375 60595 -19341
rect 60629 -19375 60641 -19341
rect 60441 -19385 60641 -19375
rect 60811 -19341 61011 -19331
rect 60811 -19375 60823 -19341
rect 60857 -19375 60891 -19341
rect 60925 -19375 61011 -19341
rect 60811 -19385 61011 -19375
rect 60441 -19425 60641 -19415
rect 60441 -19459 60459 -19425
rect 60493 -19459 60527 -19425
rect 60561 -19459 60595 -19425
rect 60629 -19459 60641 -19425
rect 60441 -19469 60641 -19459
rect 60811 -19425 61011 -19415
rect 60811 -19459 60823 -19425
rect 60857 -19459 60891 -19425
rect 60925 -19459 60959 -19425
rect 60993 -19459 61011 -19425
rect 60811 -19469 61011 -19459
rect 60441 -19509 60641 -19499
rect 60441 -19543 60595 -19509
rect 60629 -19543 60641 -19509
rect 60441 -19551 60641 -19543
rect 60811 -19509 61011 -19499
rect 60811 -19543 60823 -19509
rect 60857 -19543 61011 -19509
rect 60811 -19551 61011 -19543
rect 57123 -20157 57175 -20121
rect 57123 -20191 57131 -20157
rect 57165 -20191 57175 -20157
rect 57123 -20225 57175 -20191
rect 57123 -20259 57131 -20225
rect 57165 -20259 57175 -20225
rect 57123 -20279 57175 -20259
rect 57205 -20157 57263 -20121
rect 57205 -20191 57217 -20157
rect 57251 -20191 57263 -20157
rect 57205 -20225 57263 -20191
rect 57205 -20259 57217 -20225
rect 57251 -20259 57263 -20225
rect 57205 -20279 57263 -20259
rect 57293 -20144 57345 -20121
rect 57293 -20178 57303 -20144
rect 57337 -20178 57345 -20144
rect 57293 -20225 57345 -20178
rect 57293 -20259 57303 -20225
rect 57337 -20259 57345 -20225
rect 57293 -20279 57345 -20259
rect 59113 -20154 59513 -20142
rect 59113 -20188 59125 -20154
rect 59501 -20188 59513 -20154
rect 59113 -20200 59513 -20188
rect 59113 -20262 59513 -20250
rect 59113 -20296 59125 -20262
rect 59501 -20296 59513 -20262
rect 59113 -20308 59513 -20296
rect 59113 -20370 59513 -20358
rect 59113 -20404 59125 -20370
rect 59501 -20404 59513 -20370
rect 59113 -20416 59513 -20404
rect 54069 -20544 54869 -20532
rect 54069 -20578 54081 -20544
rect 54857 -20578 54869 -20544
rect 54069 -20590 54869 -20578
rect 54069 -20672 54869 -20660
rect 54069 -20706 54081 -20672
rect 54857 -20706 54869 -20672
rect 54069 -20718 54869 -20706
rect 54079 -23272 54879 -23260
rect 54079 -23306 54091 -23272
rect 54867 -23306 54879 -23272
rect 54079 -23318 54879 -23306
rect 54079 -23400 54879 -23388
rect 54079 -23434 54091 -23400
rect 54867 -23434 54879 -23400
rect 54079 -23446 54879 -23434
rect 54079 -23628 54879 -23616
rect 54079 -23662 54091 -23628
rect 54867 -23662 54879 -23628
rect 54079 -23674 54879 -23662
rect 54079 -23756 54879 -23744
rect 54079 -23790 54091 -23756
rect 54867 -23790 54879 -23756
rect 54079 -23802 54879 -23790
rect 57123 -23729 57175 -23709
rect 57123 -23763 57131 -23729
rect 57165 -23763 57175 -23729
rect 57123 -23797 57175 -23763
rect 57123 -23831 57131 -23797
rect 57165 -23831 57175 -23797
rect 57123 -23867 57175 -23831
rect 57205 -23729 57263 -23709
rect 57205 -23763 57217 -23729
rect 57251 -23763 57263 -23729
rect 57205 -23797 57263 -23763
rect 57205 -23831 57217 -23797
rect 57251 -23831 57263 -23797
rect 57205 -23867 57263 -23831
rect 57293 -23729 57345 -23709
rect 57293 -23763 57303 -23729
rect 57337 -23763 57345 -23729
rect 57293 -23810 57345 -23763
rect 57293 -23844 57303 -23810
rect 57337 -23844 57345 -23810
rect 57293 -23867 57345 -23844
rect 59113 -23647 59513 -23635
rect 59113 -23681 59125 -23647
rect 59501 -23681 59513 -23647
rect 59113 -23693 59513 -23681
rect 59113 -23755 59513 -23743
rect 59113 -23789 59125 -23755
rect 59501 -23789 59513 -23755
rect 59113 -23801 59513 -23789
rect 59113 -23863 59513 -23851
rect 59113 -23897 59125 -23863
rect 59501 -23897 59513 -23863
rect 59113 -23909 59513 -23897
rect 54069 -25588 54869 -25576
rect 54069 -25622 54081 -25588
rect 54857 -25622 54869 -25588
rect 54069 -25634 54869 -25622
rect 54069 -25716 54869 -25704
rect 54069 -25750 54081 -25716
rect 54857 -25750 54869 -25716
rect 54069 -25762 54869 -25750
rect 56418 -24299 56476 -24287
rect 56418 -25075 56430 -24299
rect 56464 -25075 56476 -24299
rect 56418 -25087 56476 -25075
rect 56546 -24299 56604 -24287
rect 56546 -25075 56558 -24299
rect 56592 -25075 56604 -24299
rect 56546 -25087 56604 -25075
rect 59032 -24171 59090 -24159
rect 59032 -24547 59044 -24171
rect 59078 -24547 59090 -24171
rect 59032 -24559 59090 -24547
rect 59150 -24171 59208 -24159
rect 59150 -24547 59162 -24171
rect 59196 -24547 59208 -24171
rect 59150 -24559 59208 -24547
rect 60441 -24573 60641 -24565
rect 60441 -24607 60459 -24573
rect 60493 -24607 60527 -24573
rect 60561 -24607 60595 -24573
rect 60629 -24607 60641 -24573
rect 60441 -24617 60641 -24607
rect 60811 -24573 61011 -24565
rect 60811 -24607 60823 -24573
rect 60857 -24607 60891 -24573
rect 60925 -24607 60959 -24573
rect 60993 -24607 61011 -24573
rect 60811 -24617 61011 -24607
rect 60441 -24657 60641 -24647
rect 60441 -24691 60459 -24657
rect 60493 -24691 60527 -24657
rect 60561 -24691 60595 -24657
rect 60629 -24691 60641 -24657
rect 60441 -24701 60641 -24691
rect 60811 -24657 61011 -24647
rect 60811 -24691 60823 -24657
rect 60857 -24691 60891 -24657
rect 60925 -24691 60959 -24657
rect 60993 -24691 61011 -24657
rect 60811 -24701 61011 -24691
rect 59032 -24901 59090 -24889
rect 59032 -25277 59044 -24901
rect 59078 -25277 59090 -24901
rect 59032 -25289 59090 -25277
rect 59150 -24901 59208 -24889
rect 59150 -25277 59162 -24901
rect 59196 -25277 59208 -24901
rect 59150 -25289 59208 -25277
rect 60441 -24741 60641 -24731
rect 60441 -24775 60527 -24741
rect 60561 -24775 60595 -24741
rect 60629 -24775 60641 -24741
rect 60441 -24785 60641 -24775
rect 60811 -24741 61011 -24731
rect 60811 -24775 60823 -24741
rect 60857 -24775 60891 -24741
rect 60925 -24775 61011 -24741
rect 60811 -24785 61011 -24775
rect 60441 -24825 60641 -24815
rect 60441 -24859 60459 -24825
rect 60493 -24859 60527 -24825
rect 60561 -24859 60595 -24825
rect 60629 -24859 60641 -24825
rect 60441 -24869 60641 -24859
rect 60811 -24825 61011 -24815
rect 60811 -24859 60823 -24825
rect 60857 -24859 60891 -24825
rect 60925 -24859 60959 -24825
rect 60993 -24859 61011 -24825
rect 60811 -24869 61011 -24859
rect 60441 -24909 60641 -24899
rect 60441 -24943 60595 -24909
rect 60629 -24943 60641 -24909
rect 60441 -24951 60641 -24943
rect 60811 -24909 61011 -24899
rect 60811 -24943 60823 -24909
rect 60857 -24943 61011 -24909
rect 60811 -24951 61011 -24943
rect 57123 -25557 57175 -25521
rect 57123 -25591 57131 -25557
rect 57165 -25591 57175 -25557
rect 57123 -25625 57175 -25591
rect 57123 -25659 57131 -25625
rect 57165 -25659 57175 -25625
rect 57123 -25679 57175 -25659
rect 57205 -25557 57263 -25521
rect 57205 -25591 57217 -25557
rect 57251 -25591 57263 -25557
rect 57205 -25625 57263 -25591
rect 57205 -25659 57217 -25625
rect 57251 -25659 57263 -25625
rect 57205 -25679 57263 -25659
rect 57293 -25544 57345 -25521
rect 57293 -25578 57303 -25544
rect 57337 -25578 57345 -25544
rect 57293 -25625 57345 -25578
rect 57293 -25659 57303 -25625
rect 57337 -25659 57345 -25625
rect 57293 -25679 57345 -25659
rect 59113 -25554 59513 -25542
rect 59113 -25588 59125 -25554
rect 59501 -25588 59513 -25554
rect 59113 -25600 59513 -25588
rect 59113 -25662 59513 -25650
rect 59113 -25696 59125 -25662
rect 59501 -25696 59513 -25662
rect 59113 -25708 59513 -25696
rect 59113 -25770 59513 -25758
rect 59113 -25804 59125 -25770
rect 59501 -25804 59513 -25770
rect 59113 -25816 59513 -25804
rect 54069 -25944 54869 -25932
rect 54069 -25978 54081 -25944
rect 54857 -25978 54869 -25944
rect 54069 -25990 54869 -25978
rect 54069 -26072 54869 -26060
rect 54069 -26106 54081 -26072
rect 54857 -26106 54869 -26072
rect 54069 -26118 54869 -26106
rect 54079 -28672 54879 -28660
rect 54079 -28706 54091 -28672
rect 54867 -28706 54879 -28672
rect 54079 -28718 54879 -28706
rect 54079 -28800 54879 -28788
rect 54079 -28834 54091 -28800
rect 54867 -28834 54879 -28800
rect 54079 -28846 54879 -28834
rect 54079 -29028 54879 -29016
rect 54079 -29062 54091 -29028
rect 54867 -29062 54879 -29028
rect 54079 -29074 54879 -29062
rect 54079 -29156 54879 -29144
rect 54079 -29190 54091 -29156
rect 54867 -29190 54879 -29156
rect 54079 -29202 54879 -29190
rect 57123 -29129 57175 -29109
rect 57123 -29163 57131 -29129
rect 57165 -29163 57175 -29129
rect 57123 -29197 57175 -29163
rect 57123 -29231 57131 -29197
rect 57165 -29231 57175 -29197
rect 57123 -29267 57175 -29231
rect 57205 -29129 57263 -29109
rect 57205 -29163 57217 -29129
rect 57251 -29163 57263 -29129
rect 57205 -29197 57263 -29163
rect 57205 -29231 57217 -29197
rect 57251 -29231 57263 -29197
rect 57205 -29267 57263 -29231
rect 57293 -29129 57345 -29109
rect 57293 -29163 57303 -29129
rect 57337 -29163 57345 -29129
rect 57293 -29210 57345 -29163
rect 57293 -29244 57303 -29210
rect 57337 -29244 57345 -29210
rect 57293 -29267 57345 -29244
rect 59113 -29047 59513 -29035
rect 59113 -29081 59125 -29047
rect 59501 -29081 59513 -29047
rect 59113 -29093 59513 -29081
rect 59113 -29155 59513 -29143
rect 59113 -29189 59125 -29155
rect 59501 -29189 59513 -29155
rect 59113 -29201 59513 -29189
rect 59113 -29263 59513 -29251
rect 59113 -29297 59125 -29263
rect 59501 -29297 59513 -29263
rect 59113 -29309 59513 -29297
rect 54069 -30988 54869 -30976
rect 54069 -31022 54081 -30988
rect 54857 -31022 54869 -30988
rect 54069 -31034 54869 -31022
rect 54069 -31116 54869 -31104
rect 54069 -31150 54081 -31116
rect 54857 -31150 54869 -31116
rect 54069 -31162 54869 -31150
rect 56418 -29699 56476 -29687
rect 56418 -30475 56430 -29699
rect 56464 -30475 56476 -29699
rect 56418 -30487 56476 -30475
rect 56546 -29699 56604 -29687
rect 56546 -30475 56558 -29699
rect 56592 -30475 56604 -29699
rect 56546 -30487 56604 -30475
rect 59032 -29571 59090 -29559
rect 59032 -29947 59044 -29571
rect 59078 -29947 59090 -29571
rect 59032 -29959 59090 -29947
rect 59150 -29571 59208 -29559
rect 59150 -29947 59162 -29571
rect 59196 -29947 59208 -29571
rect 59150 -29959 59208 -29947
rect 60441 -29973 60641 -29965
rect 60441 -30007 60459 -29973
rect 60493 -30007 60527 -29973
rect 60561 -30007 60595 -29973
rect 60629 -30007 60641 -29973
rect 60441 -30017 60641 -30007
rect 60811 -29973 61011 -29965
rect 60811 -30007 60823 -29973
rect 60857 -30007 60891 -29973
rect 60925 -30007 60959 -29973
rect 60993 -30007 61011 -29973
rect 60811 -30017 61011 -30007
rect 60441 -30057 60641 -30047
rect 60441 -30091 60459 -30057
rect 60493 -30091 60527 -30057
rect 60561 -30091 60595 -30057
rect 60629 -30091 60641 -30057
rect 60441 -30101 60641 -30091
rect 60811 -30057 61011 -30047
rect 60811 -30091 60823 -30057
rect 60857 -30091 60891 -30057
rect 60925 -30091 60959 -30057
rect 60993 -30091 61011 -30057
rect 60811 -30101 61011 -30091
rect 59032 -30301 59090 -30289
rect 59032 -30677 59044 -30301
rect 59078 -30677 59090 -30301
rect 59032 -30689 59090 -30677
rect 59150 -30301 59208 -30289
rect 59150 -30677 59162 -30301
rect 59196 -30677 59208 -30301
rect 59150 -30689 59208 -30677
rect 60441 -30141 60641 -30131
rect 60441 -30175 60527 -30141
rect 60561 -30175 60595 -30141
rect 60629 -30175 60641 -30141
rect 60441 -30185 60641 -30175
rect 60811 -30141 61011 -30131
rect 60811 -30175 60823 -30141
rect 60857 -30175 60891 -30141
rect 60925 -30175 61011 -30141
rect 60811 -30185 61011 -30175
rect 60441 -30225 60641 -30215
rect 60441 -30259 60459 -30225
rect 60493 -30259 60527 -30225
rect 60561 -30259 60595 -30225
rect 60629 -30259 60641 -30225
rect 60441 -30269 60641 -30259
rect 60811 -30225 61011 -30215
rect 60811 -30259 60823 -30225
rect 60857 -30259 60891 -30225
rect 60925 -30259 60959 -30225
rect 60993 -30259 61011 -30225
rect 60811 -30269 61011 -30259
rect 60441 -30309 60641 -30299
rect 60441 -30343 60595 -30309
rect 60629 -30343 60641 -30309
rect 60441 -30351 60641 -30343
rect 60811 -30309 61011 -30299
rect 60811 -30343 60823 -30309
rect 60857 -30343 61011 -30309
rect 60811 -30351 61011 -30343
rect 57123 -30957 57175 -30921
rect 57123 -30991 57131 -30957
rect 57165 -30991 57175 -30957
rect 57123 -31025 57175 -30991
rect 57123 -31059 57131 -31025
rect 57165 -31059 57175 -31025
rect 57123 -31079 57175 -31059
rect 57205 -30957 57263 -30921
rect 57205 -30991 57217 -30957
rect 57251 -30991 57263 -30957
rect 57205 -31025 57263 -30991
rect 57205 -31059 57217 -31025
rect 57251 -31059 57263 -31025
rect 57205 -31079 57263 -31059
rect 57293 -30944 57345 -30921
rect 57293 -30978 57303 -30944
rect 57337 -30978 57345 -30944
rect 57293 -31025 57345 -30978
rect 57293 -31059 57303 -31025
rect 57337 -31059 57345 -31025
rect 57293 -31079 57345 -31059
rect 59113 -30954 59513 -30942
rect 59113 -30988 59125 -30954
rect 59501 -30988 59513 -30954
rect 59113 -31000 59513 -30988
rect 59113 -31062 59513 -31050
rect 59113 -31096 59125 -31062
rect 59501 -31096 59513 -31062
rect 59113 -31108 59513 -31096
rect 59113 -31170 59513 -31158
rect 59113 -31204 59125 -31170
rect 59501 -31204 59513 -31170
rect 59113 -31216 59513 -31204
rect 54069 -31344 54869 -31332
rect 54069 -31378 54081 -31344
rect 54857 -31378 54869 -31344
rect 54069 -31390 54869 -31378
rect 54069 -31472 54869 -31460
rect 54069 -31506 54081 -31472
rect 54857 -31506 54869 -31472
rect 54069 -31518 54869 -31506
rect 54079 -34072 54879 -34060
rect 54079 -34106 54091 -34072
rect 54867 -34106 54879 -34072
rect 54079 -34118 54879 -34106
rect 54079 -34200 54879 -34188
rect 54079 -34234 54091 -34200
rect 54867 -34234 54879 -34200
rect 54079 -34246 54879 -34234
rect 54079 -34428 54879 -34416
rect 54079 -34462 54091 -34428
rect 54867 -34462 54879 -34428
rect 54079 -34474 54879 -34462
rect 54079 -34556 54879 -34544
rect 54079 -34590 54091 -34556
rect 54867 -34590 54879 -34556
rect 54079 -34602 54879 -34590
rect 57123 -34529 57175 -34509
rect 57123 -34563 57131 -34529
rect 57165 -34563 57175 -34529
rect 57123 -34597 57175 -34563
rect 57123 -34631 57131 -34597
rect 57165 -34631 57175 -34597
rect 57123 -34667 57175 -34631
rect 57205 -34529 57263 -34509
rect 57205 -34563 57217 -34529
rect 57251 -34563 57263 -34529
rect 57205 -34597 57263 -34563
rect 57205 -34631 57217 -34597
rect 57251 -34631 57263 -34597
rect 57205 -34667 57263 -34631
rect 57293 -34529 57345 -34509
rect 57293 -34563 57303 -34529
rect 57337 -34563 57345 -34529
rect 57293 -34610 57345 -34563
rect 57293 -34644 57303 -34610
rect 57337 -34644 57345 -34610
rect 57293 -34667 57345 -34644
rect 59113 -34447 59513 -34435
rect 59113 -34481 59125 -34447
rect 59501 -34481 59513 -34447
rect 59113 -34493 59513 -34481
rect 59113 -34555 59513 -34543
rect 59113 -34589 59125 -34555
rect 59501 -34589 59513 -34555
rect 59113 -34601 59513 -34589
rect 59113 -34663 59513 -34651
rect 59113 -34697 59125 -34663
rect 59501 -34697 59513 -34663
rect 59113 -34709 59513 -34697
rect 54069 -36388 54869 -36376
rect 54069 -36422 54081 -36388
rect 54857 -36422 54869 -36388
rect 54069 -36434 54869 -36422
rect 54069 -36516 54869 -36504
rect 54069 -36550 54081 -36516
rect 54857 -36550 54869 -36516
rect 54069 -36562 54869 -36550
rect 56418 -35099 56476 -35087
rect 56418 -35875 56430 -35099
rect 56464 -35875 56476 -35099
rect 56418 -35887 56476 -35875
rect 56546 -35099 56604 -35087
rect 56546 -35875 56558 -35099
rect 56592 -35875 56604 -35099
rect 56546 -35887 56604 -35875
rect 59032 -34971 59090 -34959
rect 59032 -35347 59044 -34971
rect 59078 -35347 59090 -34971
rect 59032 -35359 59090 -35347
rect 59150 -34971 59208 -34959
rect 59150 -35347 59162 -34971
rect 59196 -35347 59208 -34971
rect 59150 -35359 59208 -35347
rect 60441 -35373 60641 -35365
rect 60441 -35407 60459 -35373
rect 60493 -35407 60527 -35373
rect 60561 -35407 60595 -35373
rect 60629 -35407 60641 -35373
rect 60441 -35417 60641 -35407
rect 60811 -35373 61011 -35365
rect 60811 -35407 60823 -35373
rect 60857 -35407 60891 -35373
rect 60925 -35407 60959 -35373
rect 60993 -35407 61011 -35373
rect 60811 -35417 61011 -35407
rect 60441 -35457 60641 -35447
rect 60441 -35491 60459 -35457
rect 60493 -35491 60527 -35457
rect 60561 -35491 60595 -35457
rect 60629 -35491 60641 -35457
rect 60441 -35501 60641 -35491
rect 60811 -35457 61011 -35447
rect 60811 -35491 60823 -35457
rect 60857 -35491 60891 -35457
rect 60925 -35491 60959 -35457
rect 60993 -35491 61011 -35457
rect 60811 -35501 61011 -35491
rect 59032 -35701 59090 -35689
rect 59032 -36077 59044 -35701
rect 59078 -36077 59090 -35701
rect 59032 -36089 59090 -36077
rect 59150 -35701 59208 -35689
rect 59150 -36077 59162 -35701
rect 59196 -36077 59208 -35701
rect 59150 -36089 59208 -36077
rect 60441 -35541 60641 -35531
rect 60441 -35575 60527 -35541
rect 60561 -35575 60595 -35541
rect 60629 -35575 60641 -35541
rect 60441 -35585 60641 -35575
rect 60811 -35541 61011 -35531
rect 60811 -35575 60823 -35541
rect 60857 -35575 60891 -35541
rect 60925 -35575 61011 -35541
rect 60811 -35585 61011 -35575
rect 60441 -35625 60641 -35615
rect 60441 -35659 60459 -35625
rect 60493 -35659 60527 -35625
rect 60561 -35659 60595 -35625
rect 60629 -35659 60641 -35625
rect 60441 -35669 60641 -35659
rect 60811 -35625 61011 -35615
rect 60811 -35659 60823 -35625
rect 60857 -35659 60891 -35625
rect 60925 -35659 60959 -35625
rect 60993 -35659 61011 -35625
rect 60811 -35669 61011 -35659
rect 60441 -35709 60641 -35699
rect 60441 -35743 60595 -35709
rect 60629 -35743 60641 -35709
rect 60441 -35751 60641 -35743
rect 60811 -35709 61011 -35699
rect 60811 -35743 60823 -35709
rect 60857 -35743 61011 -35709
rect 60811 -35751 61011 -35743
rect 57123 -36357 57175 -36321
rect 57123 -36391 57131 -36357
rect 57165 -36391 57175 -36357
rect 57123 -36425 57175 -36391
rect 57123 -36459 57131 -36425
rect 57165 -36459 57175 -36425
rect 57123 -36479 57175 -36459
rect 57205 -36357 57263 -36321
rect 57205 -36391 57217 -36357
rect 57251 -36391 57263 -36357
rect 57205 -36425 57263 -36391
rect 57205 -36459 57217 -36425
rect 57251 -36459 57263 -36425
rect 57205 -36479 57263 -36459
rect 57293 -36344 57345 -36321
rect 57293 -36378 57303 -36344
rect 57337 -36378 57345 -36344
rect 57293 -36425 57345 -36378
rect 57293 -36459 57303 -36425
rect 57337 -36459 57345 -36425
rect 57293 -36479 57345 -36459
rect 59113 -36354 59513 -36342
rect 59113 -36388 59125 -36354
rect 59501 -36388 59513 -36354
rect 59113 -36400 59513 -36388
rect 59113 -36462 59513 -36450
rect 59113 -36496 59125 -36462
rect 59501 -36496 59513 -36462
rect 59113 -36508 59513 -36496
rect 59113 -36570 59513 -36558
rect 59113 -36604 59125 -36570
rect 59501 -36604 59513 -36570
rect 59113 -36616 59513 -36604
rect 54069 -36744 54869 -36732
rect 54069 -36778 54081 -36744
rect 54857 -36778 54869 -36744
rect 54069 -36790 54869 -36778
rect 54069 -36872 54869 -36860
rect 54069 -36906 54081 -36872
rect 54857 -36906 54869 -36872
rect 54069 -36918 54869 -36906
rect 75574 -38703 75626 -38685
rect 75574 -38737 75582 -38703
rect 75616 -38737 75626 -38703
rect 75574 -38771 75626 -38737
rect 75574 -38805 75582 -38771
rect 75616 -38805 75626 -38771
rect 75574 -38839 75626 -38805
rect 75574 -38873 75582 -38839
rect 75616 -38873 75626 -38839
rect 75574 -38885 75626 -38873
rect 75656 -38703 75708 -38685
rect 75656 -38737 75666 -38703
rect 75700 -38737 75708 -38703
rect 75656 -38771 75708 -38737
rect 75656 -38805 75666 -38771
rect 75700 -38805 75708 -38771
rect 75656 -38839 75708 -38805
rect 75656 -38873 75666 -38839
rect 75700 -38873 75708 -38839
rect 75656 -38885 75708 -38873
rect 75850 -38703 75902 -38685
rect 75850 -38737 75858 -38703
rect 75892 -38737 75902 -38703
rect 75850 -38771 75902 -38737
rect 75850 -38805 75858 -38771
rect 75892 -38805 75902 -38771
rect 75850 -38839 75902 -38805
rect 75850 -38873 75858 -38839
rect 75892 -38873 75902 -38839
rect 75850 -38885 75902 -38873
rect 75932 -38703 75984 -38685
rect 75932 -38737 75942 -38703
rect 75976 -38737 75984 -38703
rect 75932 -38771 75984 -38737
rect 75932 -38805 75942 -38771
rect 75976 -38805 75984 -38771
rect 75932 -38839 75984 -38805
rect 75932 -38873 75942 -38839
rect 75976 -38873 75984 -38839
rect 75932 -38885 75984 -38873
rect 76124 -38703 76176 -38685
rect 76124 -38737 76132 -38703
rect 76166 -38737 76176 -38703
rect 76124 -38771 76176 -38737
rect 76124 -38805 76132 -38771
rect 76166 -38805 76176 -38771
rect 76124 -38839 76176 -38805
rect 76124 -38873 76132 -38839
rect 76166 -38873 76176 -38839
rect 76124 -38885 76176 -38873
rect 76206 -38703 76258 -38685
rect 76206 -38737 76216 -38703
rect 76250 -38737 76258 -38703
rect 76206 -38771 76258 -38737
rect 76206 -38805 76216 -38771
rect 76250 -38805 76258 -38771
rect 76206 -38839 76258 -38805
rect 76206 -38873 76216 -38839
rect 76250 -38873 76258 -38839
rect 76206 -38885 76258 -38873
rect 76400 -38703 76452 -38685
rect 76400 -38737 76408 -38703
rect 76442 -38737 76452 -38703
rect 76400 -38771 76452 -38737
rect 76400 -38805 76408 -38771
rect 76442 -38805 76452 -38771
rect 76400 -38839 76452 -38805
rect 76400 -38873 76408 -38839
rect 76442 -38873 76452 -38839
rect 76400 -38885 76452 -38873
rect 76482 -38703 76534 -38685
rect 76482 -38737 76492 -38703
rect 76526 -38737 76534 -38703
rect 76482 -38771 76534 -38737
rect 76482 -38805 76492 -38771
rect 76526 -38805 76534 -38771
rect 76482 -38839 76534 -38805
rect 76482 -38873 76492 -38839
rect 76526 -38873 76534 -38839
rect 76482 -38885 76534 -38873
rect 76676 -38703 76728 -38685
rect 76676 -38737 76684 -38703
rect 76718 -38737 76728 -38703
rect 76676 -38771 76728 -38737
rect 76676 -38805 76684 -38771
rect 76718 -38805 76728 -38771
rect 76676 -38839 76728 -38805
rect 76676 -38873 76684 -38839
rect 76718 -38873 76728 -38839
rect 76676 -38885 76728 -38873
rect 76758 -38703 76810 -38685
rect 76758 -38737 76768 -38703
rect 76802 -38737 76810 -38703
rect 76758 -38771 76810 -38737
rect 76758 -38805 76768 -38771
rect 76802 -38805 76810 -38771
rect 76758 -38839 76810 -38805
rect 76758 -38873 76768 -38839
rect 76802 -38873 76810 -38839
rect 76758 -38885 76810 -38873
rect 77966 -39117 78019 -39105
rect 77966 -39151 77974 -39117
rect 78008 -39151 78019 -39117
rect 77966 -39185 78019 -39151
rect 77966 -39219 77974 -39185
rect 78008 -39219 78019 -39185
rect 77966 -39221 78019 -39219
rect 77605 -39248 77657 -39221
rect 77605 -39282 77613 -39248
rect 77647 -39282 77657 -39248
rect 77605 -39305 77657 -39282
rect 77687 -39305 77753 -39221
rect 77783 -39305 77825 -39221
rect 77855 -39305 77921 -39221
rect 77951 -39305 78019 -39221
rect 78049 -39148 78103 -39105
rect 78424 -39117 78477 -39105
rect 78049 -39182 78059 -39148
rect 78093 -39182 78103 -39148
rect 78424 -39151 78432 -39117
rect 78466 -39151 78477 -39117
rect 78049 -39216 78103 -39182
rect 78049 -39250 78059 -39216
rect 78093 -39250 78103 -39216
rect 78424 -39185 78477 -39151
rect 78424 -39219 78432 -39185
rect 78466 -39219 78477 -39185
rect 78424 -39221 78477 -39219
rect 78049 -39305 78103 -39250
rect 78159 -39248 78211 -39221
rect 78159 -39282 78167 -39248
rect 78201 -39282 78211 -39248
rect 78159 -39305 78211 -39282
rect 78241 -39305 78283 -39221
rect 78313 -39305 78379 -39221
rect 78409 -39305 78477 -39221
rect 78507 -39148 78563 -39105
rect 78845 -39117 78897 -39105
rect 78845 -39147 78853 -39117
rect 78507 -39182 78517 -39148
rect 78551 -39182 78563 -39148
rect 78507 -39216 78563 -39182
rect 78507 -39250 78517 -39216
rect 78551 -39250 78563 -39216
rect 78649 -39159 78705 -39147
rect 78649 -39193 78661 -39159
rect 78695 -39193 78705 -39159
rect 78649 -39231 78705 -39193
rect 78735 -39159 78789 -39147
rect 78735 -39193 78745 -39159
rect 78779 -39193 78789 -39159
rect 78735 -39231 78789 -39193
rect 78819 -39151 78853 -39147
rect 78887 -39151 78897 -39117
rect 78819 -39185 78897 -39151
rect 78819 -39219 78853 -39185
rect 78887 -39219 78897 -39185
rect 78819 -39231 78897 -39219
rect 78507 -39305 78563 -39250
rect 54079 -39472 54879 -39460
rect 54079 -39506 54091 -39472
rect 54867 -39506 54879 -39472
rect 54079 -39518 54879 -39506
rect 54079 -39600 54879 -39588
rect 54079 -39634 54091 -39600
rect 54867 -39634 54879 -39600
rect 54079 -39646 54879 -39634
rect 78835 -39305 78897 -39231
rect 78927 -39117 79022 -39105
rect 78927 -39151 78957 -39117
rect 78991 -39151 79022 -39117
rect 78927 -39185 79022 -39151
rect 78927 -39219 78957 -39185
rect 78991 -39219 79022 -39185
rect 78927 -39305 79022 -39219
rect 80806 -39167 80858 -39155
rect 80806 -39201 80814 -39167
rect 80848 -39201 80858 -39167
rect 80806 -39235 80858 -39201
rect 80806 -39269 80814 -39235
rect 80848 -39269 80858 -39235
rect 80806 -39303 80858 -39269
rect 80806 -39337 80814 -39303
rect 80848 -39337 80858 -39303
rect 80806 -39355 80858 -39337
rect 80888 -39167 80940 -39155
rect 80888 -39201 80898 -39167
rect 80932 -39201 80940 -39167
rect 80888 -39235 80940 -39201
rect 80888 -39269 80898 -39235
rect 80932 -39269 80940 -39235
rect 80888 -39303 80940 -39269
rect 80888 -39337 80898 -39303
rect 80932 -39337 80940 -39303
rect 80888 -39355 80940 -39337
rect 81051 -39167 81103 -39155
rect 81051 -39201 81059 -39167
rect 81093 -39201 81103 -39167
rect 81051 -39235 81103 -39201
rect 81051 -39269 81059 -39235
rect 81093 -39269 81103 -39235
rect 81051 -39303 81103 -39269
rect 81051 -39337 81059 -39303
rect 81093 -39337 81103 -39303
rect 81051 -39355 81103 -39337
rect 81133 -39167 81187 -39155
rect 81133 -39201 81143 -39167
rect 81177 -39201 81187 -39167
rect 81133 -39235 81187 -39201
rect 81133 -39269 81143 -39235
rect 81177 -39269 81187 -39235
rect 81133 -39303 81187 -39269
rect 81133 -39337 81143 -39303
rect 81177 -39337 81187 -39303
rect 81133 -39355 81187 -39337
rect 81217 -39167 81271 -39155
rect 81217 -39201 81227 -39167
rect 81261 -39201 81271 -39167
rect 81217 -39235 81271 -39201
rect 81217 -39269 81227 -39235
rect 81261 -39269 81271 -39235
rect 81217 -39355 81271 -39269
rect 81301 -39167 81355 -39155
rect 81301 -39201 81311 -39167
rect 81345 -39201 81355 -39167
rect 81301 -39235 81355 -39201
rect 81301 -39269 81311 -39235
rect 81345 -39269 81355 -39235
rect 81301 -39303 81355 -39269
rect 81301 -39337 81311 -39303
rect 81345 -39337 81355 -39303
rect 81301 -39355 81355 -39337
rect 81385 -39167 81437 -39155
rect 81385 -39201 81395 -39167
rect 81429 -39201 81437 -39167
rect 81385 -39355 81437 -39201
rect 81514 -39167 81566 -39155
rect 81514 -39201 81522 -39167
rect 81556 -39201 81566 -39167
rect 81514 -39235 81566 -39201
rect 81514 -39269 81522 -39235
rect 81556 -39269 81566 -39235
rect 81514 -39305 81566 -39269
rect 81514 -39339 81522 -39305
rect 81556 -39339 81566 -39305
rect 81514 -39355 81566 -39339
rect 81596 -39167 81650 -39155
rect 81596 -39201 81606 -39167
rect 81640 -39201 81650 -39167
rect 81596 -39235 81650 -39201
rect 81596 -39269 81606 -39235
rect 81640 -39269 81650 -39235
rect 81596 -39305 81650 -39269
rect 81596 -39339 81606 -39305
rect 81640 -39339 81650 -39305
rect 81596 -39355 81650 -39339
rect 81680 -39167 81734 -39155
rect 81680 -39201 81690 -39167
rect 81724 -39201 81734 -39167
rect 81680 -39235 81734 -39201
rect 81680 -39269 81690 -39235
rect 81724 -39269 81734 -39235
rect 81680 -39355 81734 -39269
rect 81764 -39167 81818 -39155
rect 81764 -39201 81774 -39167
rect 81808 -39201 81818 -39167
rect 81764 -39235 81818 -39201
rect 81764 -39269 81774 -39235
rect 81808 -39269 81818 -39235
rect 81764 -39305 81818 -39269
rect 81764 -39339 81774 -39305
rect 81808 -39339 81818 -39305
rect 81764 -39355 81818 -39339
rect 81848 -39167 81902 -39155
rect 81848 -39201 81858 -39167
rect 81892 -39201 81902 -39167
rect 81848 -39235 81902 -39201
rect 81848 -39269 81858 -39235
rect 81892 -39269 81902 -39235
rect 81848 -39355 81902 -39269
rect 81932 -39167 81986 -39155
rect 81932 -39201 81942 -39167
rect 81976 -39201 81986 -39167
rect 81932 -39235 81986 -39201
rect 81932 -39269 81942 -39235
rect 81976 -39269 81986 -39235
rect 81932 -39305 81986 -39269
rect 81932 -39339 81942 -39305
rect 81976 -39339 81986 -39305
rect 81932 -39355 81986 -39339
rect 82016 -39167 82070 -39155
rect 82016 -39201 82026 -39167
rect 82060 -39201 82070 -39167
rect 82016 -39235 82070 -39201
rect 82016 -39269 82026 -39235
rect 82060 -39269 82070 -39235
rect 82016 -39355 82070 -39269
rect 82100 -39167 82154 -39155
rect 82100 -39201 82110 -39167
rect 82144 -39201 82154 -39167
rect 82100 -39235 82154 -39201
rect 82100 -39269 82110 -39235
rect 82144 -39269 82154 -39235
rect 82100 -39305 82154 -39269
rect 82100 -39339 82110 -39305
rect 82144 -39339 82154 -39305
rect 82100 -39355 82154 -39339
rect 82184 -39167 82238 -39155
rect 82184 -39201 82194 -39167
rect 82228 -39201 82238 -39167
rect 82184 -39235 82238 -39201
rect 82184 -39269 82194 -39235
rect 82228 -39269 82238 -39235
rect 82184 -39355 82238 -39269
rect 82268 -39167 82322 -39155
rect 82268 -39201 82278 -39167
rect 82312 -39201 82322 -39167
rect 82268 -39235 82322 -39201
rect 82268 -39269 82278 -39235
rect 82312 -39269 82322 -39235
rect 82268 -39305 82322 -39269
rect 82268 -39339 82278 -39305
rect 82312 -39339 82322 -39305
rect 82268 -39355 82322 -39339
rect 82352 -39167 82406 -39155
rect 82352 -39201 82362 -39167
rect 82396 -39201 82406 -39167
rect 82352 -39235 82406 -39201
rect 82352 -39269 82362 -39235
rect 82396 -39269 82406 -39235
rect 82352 -39355 82406 -39269
rect 82436 -39167 82490 -39155
rect 82436 -39201 82446 -39167
rect 82480 -39201 82490 -39167
rect 82436 -39235 82490 -39201
rect 82436 -39269 82446 -39235
rect 82480 -39269 82490 -39235
rect 82436 -39305 82490 -39269
rect 82436 -39339 82446 -39305
rect 82480 -39339 82490 -39305
rect 82436 -39355 82490 -39339
rect 82520 -39167 82574 -39155
rect 82520 -39201 82530 -39167
rect 82564 -39201 82574 -39167
rect 82520 -39235 82574 -39201
rect 82520 -39269 82530 -39235
rect 82564 -39269 82574 -39235
rect 82520 -39355 82574 -39269
rect 82604 -39167 82658 -39155
rect 82604 -39201 82614 -39167
rect 82648 -39201 82658 -39167
rect 82604 -39235 82658 -39201
rect 82604 -39269 82614 -39235
rect 82648 -39269 82658 -39235
rect 82604 -39305 82658 -39269
rect 82604 -39339 82614 -39305
rect 82648 -39339 82658 -39305
rect 82604 -39355 82658 -39339
rect 82688 -39167 82742 -39155
rect 82688 -39201 82698 -39167
rect 82732 -39201 82742 -39167
rect 82688 -39235 82742 -39201
rect 82688 -39269 82698 -39235
rect 82732 -39269 82742 -39235
rect 82688 -39355 82742 -39269
rect 82772 -39167 82826 -39155
rect 82772 -39201 82782 -39167
rect 82816 -39201 82826 -39167
rect 82772 -39235 82826 -39201
rect 82772 -39269 82782 -39235
rect 82816 -39269 82826 -39235
rect 82772 -39305 82826 -39269
rect 82772 -39339 82782 -39305
rect 82816 -39339 82826 -39305
rect 82772 -39355 82826 -39339
rect 82856 -39167 82908 -39155
rect 82856 -39201 82866 -39167
rect 82900 -39201 82908 -39167
rect 82856 -39235 82908 -39201
rect 82856 -39269 82866 -39235
rect 82900 -39269 82908 -39235
rect 82856 -39355 82908 -39269
rect 82986 -39167 83038 -39155
rect 82986 -39201 82994 -39167
rect 83028 -39201 83038 -39167
rect 82986 -39235 83038 -39201
rect 82986 -39269 82994 -39235
rect 83028 -39269 83038 -39235
rect 82986 -39305 83038 -39269
rect 82986 -39339 82994 -39305
rect 83028 -39339 83038 -39305
rect 82986 -39355 83038 -39339
rect 83068 -39167 83122 -39155
rect 83068 -39201 83078 -39167
rect 83112 -39201 83122 -39167
rect 83068 -39235 83122 -39201
rect 83068 -39269 83078 -39235
rect 83112 -39269 83122 -39235
rect 83068 -39305 83122 -39269
rect 83068 -39339 83078 -39305
rect 83112 -39339 83122 -39305
rect 83068 -39355 83122 -39339
rect 83152 -39167 83206 -39155
rect 83152 -39201 83162 -39167
rect 83196 -39201 83206 -39167
rect 83152 -39235 83206 -39201
rect 83152 -39269 83162 -39235
rect 83196 -39269 83206 -39235
rect 83152 -39355 83206 -39269
rect 83236 -39167 83290 -39155
rect 83236 -39201 83246 -39167
rect 83280 -39201 83290 -39167
rect 83236 -39235 83290 -39201
rect 83236 -39269 83246 -39235
rect 83280 -39269 83290 -39235
rect 83236 -39305 83290 -39269
rect 83236 -39339 83246 -39305
rect 83280 -39339 83290 -39305
rect 83236 -39355 83290 -39339
rect 83320 -39167 83374 -39155
rect 83320 -39201 83330 -39167
rect 83364 -39201 83374 -39167
rect 83320 -39235 83374 -39201
rect 83320 -39269 83330 -39235
rect 83364 -39269 83374 -39235
rect 83320 -39355 83374 -39269
rect 83404 -39167 83458 -39155
rect 83404 -39201 83414 -39167
rect 83448 -39201 83458 -39167
rect 83404 -39235 83458 -39201
rect 83404 -39269 83414 -39235
rect 83448 -39269 83458 -39235
rect 83404 -39305 83458 -39269
rect 83404 -39339 83414 -39305
rect 83448 -39339 83458 -39305
rect 83404 -39355 83458 -39339
rect 83488 -39167 83542 -39155
rect 83488 -39201 83498 -39167
rect 83532 -39201 83542 -39167
rect 83488 -39235 83542 -39201
rect 83488 -39269 83498 -39235
rect 83532 -39269 83542 -39235
rect 83488 -39355 83542 -39269
rect 83572 -39167 83626 -39155
rect 83572 -39201 83582 -39167
rect 83616 -39201 83626 -39167
rect 83572 -39235 83626 -39201
rect 83572 -39269 83582 -39235
rect 83616 -39269 83626 -39235
rect 83572 -39305 83626 -39269
rect 83572 -39339 83582 -39305
rect 83616 -39339 83626 -39305
rect 83572 -39355 83626 -39339
rect 83656 -39167 83710 -39155
rect 83656 -39201 83666 -39167
rect 83700 -39201 83710 -39167
rect 83656 -39235 83710 -39201
rect 83656 -39269 83666 -39235
rect 83700 -39269 83710 -39235
rect 83656 -39355 83710 -39269
rect 83740 -39167 83794 -39155
rect 83740 -39201 83750 -39167
rect 83784 -39201 83794 -39167
rect 83740 -39235 83794 -39201
rect 83740 -39269 83750 -39235
rect 83784 -39269 83794 -39235
rect 83740 -39305 83794 -39269
rect 83740 -39339 83750 -39305
rect 83784 -39339 83794 -39305
rect 83740 -39355 83794 -39339
rect 83824 -39167 83878 -39155
rect 83824 -39201 83834 -39167
rect 83868 -39201 83878 -39167
rect 83824 -39235 83878 -39201
rect 83824 -39269 83834 -39235
rect 83868 -39269 83878 -39235
rect 83824 -39355 83878 -39269
rect 83908 -39167 83962 -39155
rect 83908 -39201 83918 -39167
rect 83952 -39201 83962 -39167
rect 83908 -39235 83962 -39201
rect 83908 -39269 83918 -39235
rect 83952 -39269 83962 -39235
rect 83908 -39305 83962 -39269
rect 83908 -39339 83918 -39305
rect 83952 -39339 83962 -39305
rect 83908 -39355 83962 -39339
rect 83992 -39167 84046 -39155
rect 83992 -39201 84002 -39167
rect 84036 -39201 84046 -39167
rect 83992 -39235 84046 -39201
rect 83992 -39269 84002 -39235
rect 84036 -39269 84046 -39235
rect 83992 -39355 84046 -39269
rect 84076 -39167 84130 -39155
rect 84076 -39201 84086 -39167
rect 84120 -39201 84130 -39167
rect 84076 -39235 84130 -39201
rect 84076 -39269 84086 -39235
rect 84120 -39269 84130 -39235
rect 84076 -39305 84130 -39269
rect 84076 -39339 84086 -39305
rect 84120 -39339 84130 -39305
rect 84076 -39355 84130 -39339
rect 84160 -39167 84214 -39155
rect 84160 -39201 84170 -39167
rect 84204 -39201 84214 -39167
rect 84160 -39235 84214 -39201
rect 84160 -39269 84170 -39235
rect 84204 -39269 84214 -39235
rect 84160 -39355 84214 -39269
rect 84244 -39167 84298 -39155
rect 84244 -39201 84254 -39167
rect 84288 -39201 84298 -39167
rect 84244 -39235 84298 -39201
rect 84244 -39269 84254 -39235
rect 84288 -39269 84298 -39235
rect 84244 -39305 84298 -39269
rect 84244 -39339 84254 -39305
rect 84288 -39339 84298 -39305
rect 84244 -39355 84298 -39339
rect 84328 -39167 84380 -39155
rect 84328 -39201 84338 -39167
rect 84372 -39201 84380 -39167
rect 84328 -39235 84380 -39201
rect 84328 -39269 84338 -39235
rect 84372 -39269 84380 -39235
rect 84328 -39355 84380 -39269
rect 84458 -39167 84510 -39155
rect 84458 -39201 84466 -39167
rect 84500 -39201 84510 -39167
rect 84458 -39235 84510 -39201
rect 84458 -39269 84466 -39235
rect 84500 -39269 84510 -39235
rect 84458 -39305 84510 -39269
rect 84458 -39339 84466 -39305
rect 84500 -39339 84510 -39305
rect 84458 -39355 84510 -39339
rect 84540 -39167 84594 -39155
rect 84540 -39201 84550 -39167
rect 84584 -39201 84594 -39167
rect 84540 -39235 84594 -39201
rect 84540 -39269 84550 -39235
rect 84584 -39269 84594 -39235
rect 84540 -39305 84594 -39269
rect 84540 -39339 84550 -39305
rect 84584 -39339 84594 -39305
rect 84540 -39355 84594 -39339
rect 84624 -39167 84678 -39155
rect 84624 -39201 84634 -39167
rect 84668 -39201 84678 -39167
rect 84624 -39235 84678 -39201
rect 84624 -39269 84634 -39235
rect 84668 -39269 84678 -39235
rect 84624 -39355 84678 -39269
rect 84708 -39167 84762 -39155
rect 84708 -39201 84718 -39167
rect 84752 -39201 84762 -39167
rect 84708 -39235 84762 -39201
rect 84708 -39269 84718 -39235
rect 84752 -39269 84762 -39235
rect 84708 -39305 84762 -39269
rect 84708 -39339 84718 -39305
rect 84752 -39339 84762 -39305
rect 84708 -39355 84762 -39339
rect 84792 -39167 84846 -39155
rect 84792 -39201 84802 -39167
rect 84836 -39201 84846 -39167
rect 84792 -39235 84846 -39201
rect 84792 -39269 84802 -39235
rect 84836 -39269 84846 -39235
rect 84792 -39355 84846 -39269
rect 84876 -39167 84930 -39155
rect 84876 -39201 84886 -39167
rect 84920 -39201 84930 -39167
rect 84876 -39235 84930 -39201
rect 84876 -39269 84886 -39235
rect 84920 -39269 84930 -39235
rect 84876 -39305 84930 -39269
rect 84876 -39339 84886 -39305
rect 84920 -39339 84930 -39305
rect 84876 -39355 84930 -39339
rect 84960 -39167 85014 -39155
rect 84960 -39201 84970 -39167
rect 85004 -39201 85014 -39167
rect 84960 -39235 85014 -39201
rect 84960 -39269 84970 -39235
rect 85004 -39269 85014 -39235
rect 84960 -39355 85014 -39269
rect 85044 -39167 85098 -39155
rect 85044 -39201 85054 -39167
rect 85088 -39201 85098 -39167
rect 85044 -39235 85098 -39201
rect 85044 -39269 85054 -39235
rect 85088 -39269 85098 -39235
rect 85044 -39305 85098 -39269
rect 85044 -39339 85054 -39305
rect 85088 -39339 85098 -39305
rect 85044 -39355 85098 -39339
rect 85128 -39167 85182 -39155
rect 85128 -39201 85138 -39167
rect 85172 -39201 85182 -39167
rect 85128 -39235 85182 -39201
rect 85128 -39269 85138 -39235
rect 85172 -39269 85182 -39235
rect 85128 -39355 85182 -39269
rect 85212 -39167 85266 -39155
rect 85212 -39201 85222 -39167
rect 85256 -39201 85266 -39167
rect 85212 -39235 85266 -39201
rect 85212 -39269 85222 -39235
rect 85256 -39269 85266 -39235
rect 85212 -39305 85266 -39269
rect 85212 -39339 85222 -39305
rect 85256 -39339 85266 -39305
rect 85212 -39355 85266 -39339
rect 85296 -39167 85350 -39155
rect 85296 -39201 85306 -39167
rect 85340 -39201 85350 -39167
rect 85296 -39235 85350 -39201
rect 85296 -39269 85306 -39235
rect 85340 -39269 85350 -39235
rect 85296 -39355 85350 -39269
rect 85380 -39167 85434 -39155
rect 85380 -39201 85390 -39167
rect 85424 -39201 85434 -39167
rect 85380 -39235 85434 -39201
rect 85380 -39269 85390 -39235
rect 85424 -39269 85434 -39235
rect 85380 -39305 85434 -39269
rect 85380 -39339 85390 -39305
rect 85424 -39339 85434 -39305
rect 85380 -39355 85434 -39339
rect 85464 -39167 85518 -39155
rect 85464 -39201 85474 -39167
rect 85508 -39201 85518 -39167
rect 85464 -39235 85518 -39201
rect 85464 -39269 85474 -39235
rect 85508 -39269 85518 -39235
rect 85464 -39355 85518 -39269
rect 85548 -39167 85602 -39155
rect 85548 -39201 85558 -39167
rect 85592 -39201 85602 -39167
rect 85548 -39235 85602 -39201
rect 85548 -39269 85558 -39235
rect 85592 -39269 85602 -39235
rect 85548 -39305 85602 -39269
rect 85548 -39339 85558 -39305
rect 85592 -39339 85602 -39305
rect 85548 -39355 85602 -39339
rect 85632 -39167 85686 -39155
rect 85632 -39201 85642 -39167
rect 85676 -39201 85686 -39167
rect 85632 -39235 85686 -39201
rect 85632 -39269 85642 -39235
rect 85676 -39269 85686 -39235
rect 85632 -39355 85686 -39269
rect 85716 -39167 85770 -39155
rect 85716 -39201 85726 -39167
rect 85760 -39201 85770 -39167
rect 85716 -39235 85770 -39201
rect 85716 -39269 85726 -39235
rect 85760 -39269 85770 -39235
rect 85716 -39305 85770 -39269
rect 85716 -39339 85726 -39305
rect 85760 -39339 85770 -39305
rect 85716 -39355 85770 -39339
rect 85800 -39167 85852 -39155
rect 85800 -39201 85810 -39167
rect 85844 -39201 85852 -39167
rect 85800 -39235 85852 -39201
rect 85800 -39269 85810 -39235
rect 85844 -39269 85852 -39235
rect 85800 -39355 85852 -39269
rect 85930 -39167 85982 -39155
rect 85930 -39201 85938 -39167
rect 85972 -39201 85982 -39167
rect 85930 -39235 85982 -39201
rect 85930 -39269 85938 -39235
rect 85972 -39269 85982 -39235
rect 85930 -39305 85982 -39269
rect 85930 -39339 85938 -39305
rect 85972 -39339 85982 -39305
rect 85930 -39355 85982 -39339
rect 86012 -39167 86066 -39155
rect 86012 -39201 86022 -39167
rect 86056 -39201 86066 -39167
rect 86012 -39235 86066 -39201
rect 86012 -39269 86022 -39235
rect 86056 -39269 86066 -39235
rect 86012 -39305 86066 -39269
rect 86012 -39339 86022 -39305
rect 86056 -39339 86066 -39305
rect 86012 -39355 86066 -39339
rect 86096 -39167 86150 -39155
rect 86096 -39201 86106 -39167
rect 86140 -39201 86150 -39167
rect 86096 -39235 86150 -39201
rect 86096 -39269 86106 -39235
rect 86140 -39269 86150 -39235
rect 86096 -39355 86150 -39269
rect 86180 -39167 86234 -39155
rect 86180 -39201 86190 -39167
rect 86224 -39201 86234 -39167
rect 86180 -39235 86234 -39201
rect 86180 -39269 86190 -39235
rect 86224 -39269 86234 -39235
rect 86180 -39305 86234 -39269
rect 86180 -39339 86190 -39305
rect 86224 -39339 86234 -39305
rect 86180 -39355 86234 -39339
rect 86264 -39167 86318 -39155
rect 86264 -39201 86274 -39167
rect 86308 -39201 86318 -39167
rect 86264 -39235 86318 -39201
rect 86264 -39269 86274 -39235
rect 86308 -39269 86318 -39235
rect 86264 -39355 86318 -39269
rect 86348 -39167 86402 -39155
rect 86348 -39201 86358 -39167
rect 86392 -39201 86402 -39167
rect 86348 -39235 86402 -39201
rect 86348 -39269 86358 -39235
rect 86392 -39269 86402 -39235
rect 86348 -39305 86402 -39269
rect 86348 -39339 86358 -39305
rect 86392 -39339 86402 -39305
rect 86348 -39355 86402 -39339
rect 86432 -39167 86486 -39155
rect 86432 -39201 86442 -39167
rect 86476 -39201 86486 -39167
rect 86432 -39235 86486 -39201
rect 86432 -39269 86442 -39235
rect 86476 -39269 86486 -39235
rect 86432 -39355 86486 -39269
rect 86516 -39167 86570 -39155
rect 86516 -39201 86526 -39167
rect 86560 -39201 86570 -39167
rect 86516 -39235 86570 -39201
rect 86516 -39269 86526 -39235
rect 86560 -39269 86570 -39235
rect 86516 -39305 86570 -39269
rect 86516 -39339 86526 -39305
rect 86560 -39339 86570 -39305
rect 86516 -39355 86570 -39339
rect 86600 -39167 86654 -39155
rect 86600 -39201 86610 -39167
rect 86644 -39201 86654 -39167
rect 86600 -39235 86654 -39201
rect 86600 -39269 86610 -39235
rect 86644 -39269 86654 -39235
rect 86600 -39355 86654 -39269
rect 86684 -39167 86738 -39155
rect 86684 -39201 86694 -39167
rect 86728 -39201 86738 -39167
rect 86684 -39235 86738 -39201
rect 86684 -39269 86694 -39235
rect 86728 -39269 86738 -39235
rect 86684 -39305 86738 -39269
rect 86684 -39339 86694 -39305
rect 86728 -39339 86738 -39305
rect 86684 -39355 86738 -39339
rect 86768 -39167 86822 -39155
rect 86768 -39201 86778 -39167
rect 86812 -39201 86822 -39167
rect 86768 -39235 86822 -39201
rect 86768 -39269 86778 -39235
rect 86812 -39269 86822 -39235
rect 86768 -39355 86822 -39269
rect 86852 -39167 86906 -39155
rect 86852 -39201 86862 -39167
rect 86896 -39201 86906 -39167
rect 86852 -39235 86906 -39201
rect 86852 -39269 86862 -39235
rect 86896 -39269 86906 -39235
rect 86852 -39305 86906 -39269
rect 86852 -39339 86862 -39305
rect 86896 -39339 86906 -39305
rect 86852 -39355 86906 -39339
rect 86936 -39167 86990 -39155
rect 86936 -39201 86946 -39167
rect 86980 -39201 86990 -39167
rect 86936 -39235 86990 -39201
rect 86936 -39269 86946 -39235
rect 86980 -39269 86990 -39235
rect 86936 -39355 86990 -39269
rect 87020 -39167 87074 -39155
rect 87020 -39201 87030 -39167
rect 87064 -39201 87074 -39167
rect 87020 -39235 87074 -39201
rect 87020 -39269 87030 -39235
rect 87064 -39269 87074 -39235
rect 87020 -39305 87074 -39269
rect 87020 -39339 87030 -39305
rect 87064 -39339 87074 -39305
rect 87020 -39355 87074 -39339
rect 87104 -39167 87158 -39155
rect 87104 -39201 87114 -39167
rect 87148 -39201 87158 -39167
rect 87104 -39235 87158 -39201
rect 87104 -39269 87114 -39235
rect 87148 -39269 87158 -39235
rect 87104 -39355 87158 -39269
rect 87188 -39167 87242 -39155
rect 87188 -39201 87198 -39167
rect 87232 -39201 87242 -39167
rect 87188 -39235 87242 -39201
rect 87188 -39269 87198 -39235
rect 87232 -39269 87242 -39235
rect 87188 -39305 87242 -39269
rect 87188 -39339 87198 -39305
rect 87232 -39339 87242 -39305
rect 87188 -39355 87242 -39339
rect 87272 -39167 87324 -39155
rect 87272 -39201 87282 -39167
rect 87316 -39201 87324 -39167
rect 87272 -39235 87324 -39201
rect 87272 -39269 87282 -39235
rect 87316 -39269 87324 -39235
rect 87272 -39355 87324 -39269
rect 87402 -39167 87454 -39155
rect 87402 -39201 87410 -39167
rect 87444 -39201 87454 -39167
rect 87402 -39235 87454 -39201
rect 87402 -39269 87410 -39235
rect 87444 -39269 87454 -39235
rect 87402 -39305 87454 -39269
rect 87402 -39339 87410 -39305
rect 87444 -39339 87454 -39305
rect 87402 -39355 87454 -39339
rect 87484 -39167 87538 -39155
rect 87484 -39201 87494 -39167
rect 87528 -39201 87538 -39167
rect 87484 -39235 87538 -39201
rect 87484 -39269 87494 -39235
rect 87528 -39269 87538 -39235
rect 87484 -39305 87538 -39269
rect 87484 -39339 87494 -39305
rect 87528 -39339 87538 -39305
rect 87484 -39355 87538 -39339
rect 87568 -39167 87622 -39155
rect 87568 -39201 87578 -39167
rect 87612 -39201 87622 -39167
rect 87568 -39235 87622 -39201
rect 87568 -39269 87578 -39235
rect 87612 -39269 87622 -39235
rect 87568 -39355 87622 -39269
rect 87652 -39167 87706 -39155
rect 87652 -39201 87662 -39167
rect 87696 -39201 87706 -39167
rect 87652 -39235 87706 -39201
rect 87652 -39269 87662 -39235
rect 87696 -39269 87706 -39235
rect 87652 -39305 87706 -39269
rect 87652 -39339 87662 -39305
rect 87696 -39339 87706 -39305
rect 87652 -39355 87706 -39339
rect 87736 -39167 87790 -39155
rect 87736 -39201 87746 -39167
rect 87780 -39201 87790 -39167
rect 87736 -39235 87790 -39201
rect 87736 -39269 87746 -39235
rect 87780 -39269 87790 -39235
rect 87736 -39355 87790 -39269
rect 87820 -39167 87874 -39155
rect 87820 -39201 87830 -39167
rect 87864 -39201 87874 -39167
rect 87820 -39235 87874 -39201
rect 87820 -39269 87830 -39235
rect 87864 -39269 87874 -39235
rect 87820 -39305 87874 -39269
rect 87820 -39339 87830 -39305
rect 87864 -39339 87874 -39305
rect 87820 -39355 87874 -39339
rect 87904 -39167 87958 -39155
rect 87904 -39201 87914 -39167
rect 87948 -39201 87958 -39167
rect 87904 -39235 87958 -39201
rect 87904 -39269 87914 -39235
rect 87948 -39269 87958 -39235
rect 87904 -39355 87958 -39269
rect 87988 -39167 88042 -39155
rect 87988 -39201 87998 -39167
rect 88032 -39201 88042 -39167
rect 87988 -39235 88042 -39201
rect 87988 -39269 87998 -39235
rect 88032 -39269 88042 -39235
rect 87988 -39305 88042 -39269
rect 87988 -39339 87998 -39305
rect 88032 -39339 88042 -39305
rect 87988 -39355 88042 -39339
rect 88072 -39167 88126 -39155
rect 88072 -39201 88082 -39167
rect 88116 -39201 88126 -39167
rect 88072 -39235 88126 -39201
rect 88072 -39269 88082 -39235
rect 88116 -39269 88126 -39235
rect 88072 -39355 88126 -39269
rect 88156 -39167 88210 -39155
rect 88156 -39201 88166 -39167
rect 88200 -39201 88210 -39167
rect 88156 -39235 88210 -39201
rect 88156 -39269 88166 -39235
rect 88200 -39269 88210 -39235
rect 88156 -39305 88210 -39269
rect 88156 -39339 88166 -39305
rect 88200 -39339 88210 -39305
rect 88156 -39355 88210 -39339
rect 88240 -39167 88294 -39155
rect 88240 -39201 88250 -39167
rect 88284 -39201 88294 -39167
rect 88240 -39235 88294 -39201
rect 88240 -39269 88250 -39235
rect 88284 -39269 88294 -39235
rect 88240 -39355 88294 -39269
rect 88324 -39167 88378 -39155
rect 88324 -39201 88334 -39167
rect 88368 -39201 88378 -39167
rect 88324 -39235 88378 -39201
rect 88324 -39269 88334 -39235
rect 88368 -39269 88378 -39235
rect 88324 -39305 88378 -39269
rect 88324 -39339 88334 -39305
rect 88368 -39339 88378 -39305
rect 88324 -39355 88378 -39339
rect 88408 -39167 88462 -39155
rect 88408 -39201 88418 -39167
rect 88452 -39201 88462 -39167
rect 88408 -39235 88462 -39201
rect 88408 -39269 88418 -39235
rect 88452 -39269 88462 -39235
rect 88408 -39355 88462 -39269
rect 88492 -39167 88546 -39155
rect 88492 -39201 88502 -39167
rect 88536 -39201 88546 -39167
rect 88492 -39235 88546 -39201
rect 88492 -39269 88502 -39235
rect 88536 -39269 88546 -39235
rect 88492 -39305 88546 -39269
rect 88492 -39339 88502 -39305
rect 88536 -39339 88546 -39305
rect 88492 -39355 88546 -39339
rect 88576 -39167 88630 -39155
rect 88576 -39201 88586 -39167
rect 88620 -39201 88630 -39167
rect 88576 -39235 88630 -39201
rect 88576 -39269 88586 -39235
rect 88620 -39269 88630 -39235
rect 88576 -39355 88630 -39269
rect 88660 -39167 88714 -39155
rect 88660 -39201 88670 -39167
rect 88704 -39201 88714 -39167
rect 88660 -39235 88714 -39201
rect 88660 -39269 88670 -39235
rect 88704 -39269 88714 -39235
rect 88660 -39305 88714 -39269
rect 88660 -39339 88670 -39305
rect 88704 -39339 88714 -39305
rect 88660 -39355 88714 -39339
rect 88744 -39167 88796 -39155
rect 88744 -39201 88754 -39167
rect 88788 -39201 88796 -39167
rect 88744 -39235 88796 -39201
rect 88744 -39269 88754 -39235
rect 88788 -39269 88796 -39235
rect 88744 -39355 88796 -39269
rect 54079 -39828 54879 -39816
rect 54079 -39862 54091 -39828
rect 54867 -39862 54879 -39828
rect 54079 -39874 54879 -39862
rect 54079 -39956 54879 -39944
rect 54079 -39990 54091 -39956
rect 54867 -39990 54879 -39956
rect 54079 -40002 54879 -39990
rect 57123 -39929 57175 -39909
rect 57123 -39963 57131 -39929
rect 57165 -39963 57175 -39929
rect 57123 -39997 57175 -39963
rect 57123 -40031 57131 -39997
rect 57165 -40031 57175 -39997
rect 57123 -40067 57175 -40031
rect 57205 -39929 57263 -39909
rect 57205 -39963 57217 -39929
rect 57251 -39963 57263 -39929
rect 57205 -39997 57263 -39963
rect 57205 -40031 57217 -39997
rect 57251 -40031 57263 -39997
rect 57205 -40067 57263 -40031
rect 57293 -39929 57345 -39909
rect 57293 -39963 57303 -39929
rect 57337 -39963 57345 -39929
rect 57293 -40010 57345 -39963
rect 57293 -40044 57303 -40010
rect 57337 -40044 57345 -40010
rect 57293 -40067 57345 -40044
rect 59113 -39847 59513 -39835
rect 59113 -39881 59125 -39847
rect 59501 -39881 59513 -39847
rect 59113 -39893 59513 -39881
rect 59113 -39955 59513 -39943
rect 59113 -39989 59125 -39955
rect 59501 -39989 59513 -39955
rect 59113 -40001 59513 -39989
rect 59113 -40063 59513 -40051
rect 59113 -40097 59125 -40063
rect 59501 -40097 59513 -40063
rect 59113 -40109 59513 -40097
rect 77605 -40008 77657 -39985
rect 77605 -40042 77613 -40008
rect 77647 -40042 77657 -40008
rect 77605 -40069 77657 -40042
rect 77687 -40069 77753 -39985
rect 77783 -40069 77825 -39985
rect 77855 -40069 77921 -39985
rect 77951 -40069 78019 -39985
rect 54069 -41788 54869 -41776
rect 54069 -41822 54081 -41788
rect 54857 -41822 54869 -41788
rect 54069 -41834 54869 -41822
rect 54069 -41916 54869 -41904
rect 54069 -41950 54081 -41916
rect 54857 -41950 54869 -41916
rect 54069 -41962 54869 -41950
rect 56418 -40499 56476 -40487
rect 56418 -41275 56430 -40499
rect 56464 -41275 56476 -40499
rect 56418 -41287 56476 -41275
rect 56546 -40499 56604 -40487
rect 56546 -41275 56558 -40499
rect 56592 -41275 56604 -40499
rect 56546 -41287 56604 -41275
rect 59032 -40371 59090 -40359
rect 59032 -40747 59044 -40371
rect 59078 -40747 59090 -40371
rect 59032 -40759 59090 -40747
rect 59150 -40371 59208 -40359
rect 59150 -40747 59162 -40371
rect 59196 -40747 59208 -40371
rect 59150 -40759 59208 -40747
rect 77966 -40071 78019 -40069
rect 77966 -40105 77974 -40071
rect 78008 -40105 78019 -40071
rect 77966 -40139 78019 -40105
rect 77966 -40173 77974 -40139
rect 78008 -40173 78019 -40139
rect 77966 -40185 78019 -40173
rect 78049 -40040 78103 -39985
rect 78049 -40074 78059 -40040
rect 78093 -40074 78103 -40040
rect 78049 -40108 78103 -40074
rect 78049 -40142 78059 -40108
rect 78093 -40142 78103 -40108
rect 78049 -40185 78103 -40142
rect 80856 -40043 80908 -40025
rect 80856 -40077 80864 -40043
rect 80898 -40077 80908 -40043
rect 80856 -40111 80908 -40077
rect 80856 -40145 80864 -40111
rect 80898 -40145 80908 -40111
rect 80856 -40179 80908 -40145
rect 80856 -40213 80864 -40179
rect 80898 -40213 80908 -40179
rect 80856 -40225 80908 -40213
rect 80938 -40043 80990 -40025
rect 80938 -40077 80948 -40043
rect 80982 -40077 80990 -40043
rect 80938 -40111 80990 -40077
rect 80938 -40145 80948 -40111
rect 80982 -40145 80990 -40111
rect 80938 -40179 80990 -40145
rect 80938 -40213 80948 -40179
rect 80982 -40213 80990 -40179
rect 80938 -40225 80990 -40213
rect 77833 -40367 77885 -40355
rect 77833 -40397 77841 -40367
rect 77637 -40409 77693 -40397
rect 77637 -40443 77649 -40409
rect 77683 -40443 77693 -40409
rect 77637 -40481 77693 -40443
rect 77723 -40409 77777 -40397
rect 77723 -40443 77733 -40409
rect 77767 -40443 77777 -40409
rect 77723 -40481 77777 -40443
rect 77807 -40401 77841 -40397
rect 77875 -40401 77885 -40367
rect 77807 -40435 77885 -40401
rect 77807 -40469 77841 -40435
rect 77875 -40469 77885 -40435
rect 77807 -40481 77885 -40469
rect 77823 -40555 77885 -40481
rect 77915 -40367 78010 -40355
rect 77915 -40401 77945 -40367
rect 77979 -40401 78010 -40367
rect 77915 -40435 78010 -40401
rect 77915 -40469 77945 -40435
rect 77979 -40469 78010 -40435
rect 77915 -40555 78010 -40469
rect 60441 -40773 60641 -40765
rect 60441 -40807 60459 -40773
rect 60493 -40807 60527 -40773
rect 60561 -40807 60595 -40773
rect 60629 -40807 60641 -40773
rect 60441 -40817 60641 -40807
rect 60811 -40773 61011 -40765
rect 60811 -40807 60823 -40773
rect 60857 -40807 60891 -40773
rect 60925 -40807 60959 -40773
rect 60993 -40807 61011 -40773
rect 60811 -40817 61011 -40807
rect 60441 -40857 60641 -40847
rect 60441 -40891 60459 -40857
rect 60493 -40891 60527 -40857
rect 60561 -40891 60595 -40857
rect 60629 -40891 60641 -40857
rect 60441 -40901 60641 -40891
rect 60811 -40857 61011 -40847
rect 60811 -40891 60823 -40857
rect 60857 -40891 60891 -40857
rect 60925 -40891 60959 -40857
rect 60993 -40891 61011 -40857
rect 60811 -40901 61011 -40891
rect 59032 -41101 59090 -41089
rect 59032 -41477 59044 -41101
rect 59078 -41477 59090 -41101
rect 59032 -41489 59090 -41477
rect 59150 -41101 59208 -41089
rect 59150 -41477 59162 -41101
rect 59196 -41477 59208 -41101
rect 59150 -41489 59208 -41477
rect 60441 -40941 60641 -40931
rect 60441 -40975 60527 -40941
rect 60561 -40975 60595 -40941
rect 60629 -40975 60641 -40941
rect 60441 -40985 60641 -40975
rect 60811 -40941 61011 -40931
rect 60811 -40975 60823 -40941
rect 60857 -40975 60891 -40941
rect 60925 -40975 61011 -40941
rect 60811 -40985 61011 -40975
rect 60441 -41025 60641 -41015
rect 60441 -41059 60459 -41025
rect 60493 -41059 60527 -41025
rect 60561 -41059 60595 -41025
rect 60629 -41059 60641 -41025
rect 60441 -41069 60641 -41059
rect 60811 -41025 61011 -41015
rect 60811 -41059 60823 -41025
rect 60857 -41059 60891 -41025
rect 60925 -41059 60959 -41025
rect 60993 -41059 61011 -41025
rect 60811 -41069 61011 -41059
rect 60441 -41109 60641 -41099
rect 60441 -41143 60595 -41109
rect 60629 -41143 60641 -41109
rect 60441 -41151 60641 -41143
rect 60811 -41109 61011 -41099
rect 60811 -41143 60823 -41109
rect 60857 -41143 61011 -41109
rect 60811 -41151 61011 -41143
rect 77823 -41299 77885 -41225
rect 77637 -41337 77693 -41299
rect 77637 -41371 77649 -41337
rect 77683 -41371 77693 -41337
rect 77637 -41383 77693 -41371
rect 77723 -41337 77777 -41299
rect 77723 -41371 77733 -41337
rect 77767 -41371 77777 -41337
rect 77723 -41383 77777 -41371
rect 77807 -41311 77885 -41299
rect 77807 -41345 77841 -41311
rect 77875 -41345 77885 -41311
rect 77807 -41379 77885 -41345
rect 77807 -41383 77841 -41379
rect 77833 -41413 77841 -41383
rect 77875 -41413 77885 -41379
rect 77833 -41425 77885 -41413
rect 77915 -41311 78010 -41225
rect 78065 -41248 78117 -41225
rect 78065 -41282 78073 -41248
rect 78107 -41282 78117 -41248
rect 78065 -41309 78117 -41282
rect 78147 -41309 78213 -41225
rect 78243 -41309 78285 -41225
rect 78315 -41309 78381 -41225
rect 78411 -41309 78479 -41225
rect 77915 -41345 77945 -41311
rect 77979 -41345 78010 -41311
rect 77915 -41379 78010 -41345
rect 78426 -41311 78479 -41309
rect 78426 -41345 78434 -41311
rect 78468 -41345 78479 -41311
rect 77915 -41413 77945 -41379
rect 77979 -41413 78010 -41379
rect 78426 -41379 78479 -41345
rect 77915 -41425 78010 -41413
rect 78426 -41413 78434 -41379
rect 78468 -41413 78479 -41379
rect 78426 -41425 78479 -41413
rect 78509 -41280 78563 -41225
rect 78509 -41314 78519 -41280
rect 78553 -41314 78563 -41280
rect 78509 -41348 78563 -41314
rect 78509 -41382 78519 -41348
rect 78553 -41382 78563 -41348
rect 78509 -41425 78563 -41382
rect 57123 -41757 57175 -41721
rect 57123 -41791 57131 -41757
rect 57165 -41791 57175 -41757
rect 57123 -41825 57175 -41791
rect 57123 -41859 57131 -41825
rect 57165 -41859 57175 -41825
rect 57123 -41879 57175 -41859
rect 57205 -41757 57263 -41721
rect 57205 -41791 57217 -41757
rect 57251 -41791 57263 -41757
rect 57205 -41825 57263 -41791
rect 57205 -41859 57217 -41825
rect 57251 -41859 57263 -41825
rect 57205 -41879 57263 -41859
rect 57293 -41744 57345 -41721
rect 57293 -41778 57303 -41744
rect 57337 -41778 57345 -41744
rect 57293 -41825 57345 -41778
rect 57293 -41859 57303 -41825
rect 57337 -41859 57345 -41825
rect 57293 -41879 57345 -41859
rect 59113 -41754 59513 -41742
rect 59113 -41788 59125 -41754
rect 59501 -41788 59513 -41754
rect 59113 -41800 59513 -41788
rect 59113 -41862 59513 -41850
rect 59113 -41896 59125 -41862
rect 59501 -41896 59513 -41862
rect 59113 -41908 59513 -41896
rect 59113 -41970 59513 -41958
rect 59113 -42004 59125 -41970
rect 59501 -42004 59513 -41970
rect 59113 -42016 59513 -42004
rect 54069 -42144 54869 -42132
rect 54069 -42178 54081 -42144
rect 54857 -42178 54869 -42144
rect 54069 -42190 54869 -42178
rect 54069 -42272 54869 -42260
rect 54069 -42306 54081 -42272
rect 54857 -42306 54869 -42272
rect 54069 -42318 54869 -42306
rect 77833 -41607 77885 -41595
rect 77833 -41637 77841 -41607
rect 77637 -41649 77693 -41637
rect 77637 -41683 77649 -41649
rect 77683 -41683 77693 -41649
rect 77637 -41721 77693 -41683
rect 77723 -41649 77777 -41637
rect 77723 -41683 77733 -41649
rect 77767 -41683 77777 -41649
rect 77723 -41721 77777 -41683
rect 77807 -41641 77841 -41637
rect 77875 -41641 77885 -41607
rect 77807 -41675 77885 -41641
rect 77807 -41709 77841 -41675
rect 77875 -41709 77885 -41675
rect 77807 -41721 77885 -41709
rect 77823 -41795 77885 -41721
rect 77915 -41607 78010 -41595
rect 77915 -41641 77945 -41607
rect 77979 -41641 78010 -41607
rect 77915 -41675 78010 -41641
rect 77915 -41709 77945 -41675
rect 77979 -41709 78010 -41675
rect 77915 -41795 78010 -41709
rect 77825 -42553 77887 -42479
rect 77639 -42591 77695 -42553
rect 77639 -42625 77651 -42591
rect 77685 -42625 77695 -42591
rect 77639 -42637 77695 -42625
rect 77725 -42591 77779 -42553
rect 77725 -42625 77735 -42591
rect 77769 -42625 77779 -42591
rect 77725 -42637 77779 -42625
rect 77809 -42565 77887 -42553
rect 77809 -42599 77843 -42565
rect 77877 -42599 77887 -42565
rect 77809 -42633 77887 -42599
rect 77809 -42637 77843 -42633
rect 77835 -42667 77843 -42637
rect 77877 -42667 77887 -42633
rect 77835 -42679 77887 -42667
rect 77917 -42565 78012 -42479
rect 77917 -42599 77947 -42565
rect 77981 -42599 78012 -42565
rect 77917 -42633 78012 -42599
rect 77917 -42667 77947 -42633
rect 77981 -42667 78012 -42633
rect 77917 -42679 78012 -42667
rect 77605 -42857 77657 -42845
rect 77605 -42891 77613 -42857
rect 77647 -42891 77657 -42857
rect 77605 -42929 77657 -42891
rect 77687 -42865 77757 -42845
rect 77687 -42899 77705 -42865
rect 77739 -42899 77757 -42865
rect 77687 -42929 77757 -42899
rect 77787 -42857 77861 -42845
rect 77787 -42891 77807 -42857
rect 77841 -42891 77861 -42857
rect 77787 -42929 77861 -42891
rect 77891 -42865 77947 -42845
rect 77891 -42899 77902 -42865
rect 77936 -42899 77947 -42865
rect 77891 -42929 77947 -42899
rect 77977 -42857 78113 -42845
rect 77977 -42891 78053 -42857
rect 78087 -42891 78113 -42857
rect 77977 -42925 78113 -42891
rect 77977 -42929 78053 -42925
rect 77996 -42959 78053 -42929
rect 78087 -42959 78113 -42925
rect 77996 -43045 78113 -42959
rect 78143 -42857 78195 -42845
rect 78143 -42891 78153 -42857
rect 78187 -42891 78195 -42857
rect 78710 -42857 78763 -42845
rect 78143 -42925 78195 -42891
rect 78710 -42891 78718 -42857
rect 78752 -42891 78763 -42857
rect 78143 -42959 78153 -42925
rect 78187 -42959 78195 -42925
rect 78143 -42993 78195 -42959
rect 78710 -42925 78763 -42891
rect 78710 -42959 78718 -42925
rect 78752 -42959 78763 -42925
rect 78710 -42961 78763 -42959
rect 78143 -43027 78153 -42993
rect 78187 -43027 78195 -42993
rect 78143 -43045 78195 -43027
rect 78349 -42988 78401 -42961
rect 78349 -43022 78357 -42988
rect 78391 -43022 78401 -42988
rect 78349 -43045 78401 -43022
rect 78431 -43045 78497 -42961
rect 78527 -43045 78569 -42961
rect 78599 -43045 78665 -42961
rect 78695 -43045 78763 -42961
rect 78793 -42888 78847 -42845
rect 78793 -42922 78803 -42888
rect 78837 -42922 78847 -42888
rect 78793 -42956 78847 -42922
rect 78793 -42990 78803 -42956
rect 78837 -42990 78847 -42956
rect 78793 -43045 78847 -42990
rect 83075 -43683 83127 -43655
rect 77996 -43797 78113 -43711
rect 77996 -43827 78053 -43797
rect 77605 -43865 77657 -43827
rect 77605 -43899 77613 -43865
rect 77647 -43899 77657 -43865
rect 77605 -43911 77657 -43899
rect 77687 -43857 77757 -43827
rect 77687 -43891 77705 -43857
rect 77739 -43891 77757 -43857
rect 77687 -43911 77757 -43891
rect 77787 -43865 77861 -43827
rect 77787 -43899 77807 -43865
rect 77841 -43899 77861 -43865
rect 77787 -43911 77861 -43899
rect 77891 -43857 77947 -43827
rect 77891 -43891 77902 -43857
rect 77936 -43891 77947 -43857
rect 77891 -43911 77947 -43891
rect 77977 -43831 78053 -43827
rect 78087 -43831 78113 -43797
rect 77977 -43865 78113 -43831
rect 77977 -43899 78053 -43865
rect 78087 -43899 78113 -43865
rect 77977 -43911 78113 -43899
rect 78143 -43729 78195 -43711
rect 78143 -43763 78153 -43729
rect 78187 -43763 78195 -43729
rect 83075 -43717 83083 -43683
rect 83117 -43717 83127 -43683
rect 78143 -43797 78195 -43763
rect 83075 -43751 83127 -43717
rect 83075 -43771 83083 -43751
rect 78143 -43831 78153 -43797
rect 78187 -43831 78195 -43797
rect 78143 -43865 78195 -43831
rect 82906 -43803 82958 -43771
rect 82906 -43837 82914 -43803
rect 82948 -43837 82958 -43803
rect 82906 -43855 82958 -43837
rect 82988 -43855 83030 -43771
rect 83060 -43785 83083 -43771
rect 83117 -43785 83127 -43751
rect 83060 -43855 83127 -43785
rect 83157 -43667 83225 -43655
rect 83157 -43701 83183 -43667
rect 83217 -43701 83225 -43667
rect 83157 -43735 83225 -43701
rect 83157 -43769 83183 -43735
rect 83217 -43769 83225 -43735
rect 83157 -43855 83225 -43769
rect 83366 -43667 83418 -43655
rect 83366 -43701 83374 -43667
rect 83408 -43701 83418 -43667
rect 83366 -43735 83418 -43701
rect 83366 -43769 83374 -43735
rect 83408 -43769 83418 -43735
rect 83366 -43803 83418 -43769
rect 83366 -43837 83374 -43803
rect 83408 -43837 83418 -43803
rect 83366 -43855 83418 -43837
rect 83448 -43667 83500 -43655
rect 83448 -43701 83458 -43667
rect 83492 -43701 83500 -43667
rect 83448 -43735 83500 -43701
rect 83448 -43769 83458 -43735
rect 83492 -43769 83500 -43735
rect 83448 -43803 83500 -43769
rect 83448 -43837 83458 -43803
rect 83492 -43837 83500 -43803
rect 83448 -43855 83500 -43837
rect 83611 -43667 83663 -43655
rect 83611 -43701 83619 -43667
rect 83653 -43701 83663 -43667
rect 83611 -43735 83663 -43701
rect 83611 -43769 83619 -43735
rect 83653 -43769 83663 -43735
rect 83611 -43803 83663 -43769
rect 83611 -43837 83619 -43803
rect 83653 -43837 83663 -43803
rect 83611 -43855 83663 -43837
rect 83693 -43667 83747 -43655
rect 83693 -43701 83703 -43667
rect 83737 -43701 83747 -43667
rect 83693 -43735 83747 -43701
rect 83693 -43769 83703 -43735
rect 83737 -43769 83747 -43735
rect 83693 -43803 83747 -43769
rect 83693 -43837 83703 -43803
rect 83737 -43837 83747 -43803
rect 83693 -43855 83747 -43837
rect 83777 -43667 83831 -43655
rect 83777 -43701 83787 -43667
rect 83821 -43701 83831 -43667
rect 83777 -43735 83831 -43701
rect 83777 -43769 83787 -43735
rect 83821 -43769 83831 -43735
rect 83777 -43855 83831 -43769
rect 83861 -43667 83915 -43655
rect 83861 -43701 83871 -43667
rect 83905 -43701 83915 -43667
rect 83861 -43735 83915 -43701
rect 83861 -43769 83871 -43735
rect 83905 -43769 83915 -43735
rect 83861 -43803 83915 -43769
rect 83861 -43837 83871 -43803
rect 83905 -43837 83915 -43803
rect 83861 -43855 83915 -43837
rect 83945 -43667 83997 -43655
rect 83945 -43701 83955 -43667
rect 83989 -43701 83997 -43667
rect 83945 -43855 83997 -43701
rect 84074 -43667 84126 -43655
rect 84074 -43701 84082 -43667
rect 84116 -43701 84126 -43667
rect 84074 -43735 84126 -43701
rect 84074 -43769 84082 -43735
rect 84116 -43769 84126 -43735
rect 84074 -43805 84126 -43769
rect 84074 -43839 84082 -43805
rect 84116 -43839 84126 -43805
rect 84074 -43855 84126 -43839
rect 84156 -43667 84210 -43655
rect 84156 -43701 84166 -43667
rect 84200 -43701 84210 -43667
rect 84156 -43735 84210 -43701
rect 84156 -43769 84166 -43735
rect 84200 -43769 84210 -43735
rect 84156 -43805 84210 -43769
rect 84156 -43839 84166 -43805
rect 84200 -43839 84210 -43805
rect 84156 -43855 84210 -43839
rect 84240 -43667 84294 -43655
rect 84240 -43701 84250 -43667
rect 84284 -43701 84294 -43667
rect 84240 -43735 84294 -43701
rect 84240 -43769 84250 -43735
rect 84284 -43769 84294 -43735
rect 84240 -43855 84294 -43769
rect 84324 -43667 84378 -43655
rect 84324 -43701 84334 -43667
rect 84368 -43701 84378 -43667
rect 84324 -43735 84378 -43701
rect 84324 -43769 84334 -43735
rect 84368 -43769 84378 -43735
rect 84324 -43805 84378 -43769
rect 84324 -43839 84334 -43805
rect 84368 -43839 84378 -43805
rect 84324 -43855 84378 -43839
rect 84408 -43667 84462 -43655
rect 84408 -43701 84418 -43667
rect 84452 -43701 84462 -43667
rect 84408 -43735 84462 -43701
rect 84408 -43769 84418 -43735
rect 84452 -43769 84462 -43735
rect 84408 -43855 84462 -43769
rect 84492 -43667 84546 -43655
rect 84492 -43701 84502 -43667
rect 84536 -43701 84546 -43667
rect 84492 -43735 84546 -43701
rect 84492 -43769 84502 -43735
rect 84536 -43769 84546 -43735
rect 84492 -43805 84546 -43769
rect 84492 -43839 84502 -43805
rect 84536 -43839 84546 -43805
rect 84492 -43855 84546 -43839
rect 84576 -43667 84630 -43655
rect 84576 -43701 84586 -43667
rect 84620 -43701 84630 -43667
rect 84576 -43735 84630 -43701
rect 84576 -43769 84586 -43735
rect 84620 -43769 84630 -43735
rect 84576 -43855 84630 -43769
rect 84660 -43667 84714 -43655
rect 84660 -43701 84670 -43667
rect 84704 -43701 84714 -43667
rect 84660 -43735 84714 -43701
rect 84660 -43769 84670 -43735
rect 84704 -43769 84714 -43735
rect 84660 -43805 84714 -43769
rect 84660 -43839 84670 -43805
rect 84704 -43839 84714 -43805
rect 84660 -43855 84714 -43839
rect 84744 -43667 84798 -43655
rect 84744 -43701 84754 -43667
rect 84788 -43701 84798 -43667
rect 84744 -43735 84798 -43701
rect 84744 -43769 84754 -43735
rect 84788 -43769 84798 -43735
rect 84744 -43855 84798 -43769
rect 84828 -43667 84882 -43655
rect 84828 -43701 84838 -43667
rect 84872 -43701 84882 -43667
rect 84828 -43735 84882 -43701
rect 84828 -43769 84838 -43735
rect 84872 -43769 84882 -43735
rect 84828 -43805 84882 -43769
rect 84828 -43839 84838 -43805
rect 84872 -43839 84882 -43805
rect 84828 -43855 84882 -43839
rect 84912 -43667 84966 -43655
rect 84912 -43701 84922 -43667
rect 84956 -43701 84966 -43667
rect 84912 -43735 84966 -43701
rect 84912 -43769 84922 -43735
rect 84956 -43769 84966 -43735
rect 84912 -43855 84966 -43769
rect 84996 -43667 85050 -43655
rect 84996 -43701 85006 -43667
rect 85040 -43701 85050 -43667
rect 84996 -43735 85050 -43701
rect 84996 -43769 85006 -43735
rect 85040 -43769 85050 -43735
rect 84996 -43805 85050 -43769
rect 84996 -43839 85006 -43805
rect 85040 -43839 85050 -43805
rect 84996 -43855 85050 -43839
rect 85080 -43667 85134 -43655
rect 85080 -43701 85090 -43667
rect 85124 -43701 85134 -43667
rect 85080 -43735 85134 -43701
rect 85080 -43769 85090 -43735
rect 85124 -43769 85134 -43735
rect 85080 -43855 85134 -43769
rect 85164 -43667 85218 -43655
rect 85164 -43701 85174 -43667
rect 85208 -43701 85218 -43667
rect 85164 -43735 85218 -43701
rect 85164 -43769 85174 -43735
rect 85208 -43769 85218 -43735
rect 85164 -43805 85218 -43769
rect 85164 -43839 85174 -43805
rect 85208 -43839 85218 -43805
rect 85164 -43855 85218 -43839
rect 85248 -43667 85302 -43655
rect 85248 -43701 85258 -43667
rect 85292 -43701 85302 -43667
rect 85248 -43735 85302 -43701
rect 85248 -43769 85258 -43735
rect 85292 -43769 85302 -43735
rect 85248 -43855 85302 -43769
rect 85332 -43667 85386 -43655
rect 85332 -43701 85342 -43667
rect 85376 -43701 85386 -43667
rect 85332 -43735 85386 -43701
rect 85332 -43769 85342 -43735
rect 85376 -43769 85386 -43735
rect 85332 -43805 85386 -43769
rect 85332 -43839 85342 -43805
rect 85376 -43839 85386 -43805
rect 85332 -43855 85386 -43839
rect 85416 -43667 85468 -43655
rect 85416 -43701 85426 -43667
rect 85460 -43701 85468 -43667
rect 85416 -43735 85468 -43701
rect 85416 -43769 85426 -43735
rect 85460 -43769 85468 -43735
rect 85416 -43855 85468 -43769
rect 85546 -43667 85598 -43655
rect 85546 -43701 85554 -43667
rect 85588 -43701 85598 -43667
rect 85546 -43735 85598 -43701
rect 85546 -43769 85554 -43735
rect 85588 -43769 85598 -43735
rect 85546 -43805 85598 -43769
rect 85546 -43839 85554 -43805
rect 85588 -43839 85598 -43805
rect 85546 -43855 85598 -43839
rect 85628 -43667 85682 -43655
rect 85628 -43701 85638 -43667
rect 85672 -43701 85682 -43667
rect 85628 -43735 85682 -43701
rect 85628 -43769 85638 -43735
rect 85672 -43769 85682 -43735
rect 85628 -43805 85682 -43769
rect 85628 -43839 85638 -43805
rect 85672 -43839 85682 -43805
rect 85628 -43855 85682 -43839
rect 85712 -43667 85766 -43655
rect 85712 -43701 85722 -43667
rect 85756 -43701 85766 -43667
rect 85712 -43735 85766 -43701
rect 85712 -43769 85722 -43735
rect 85756 -43769 85766 -43735
rect 85712 -43855 85766 -43769
rect 85796 -43667 85850 -43655
rect 85796 -43701 85806 -43667
rect 85840 -43701 85850 -43667
rect 85796 -43735 85850 -43701
rect 85796 -43769 85806 -43735
rect 85840 -43769 85850 -43735
rect 85796 -43805 85850 -43769
rect 85796 -43839 85806 -43805
rect 85840 -43839 85850 -43805
rect 85796 -43855 85850 -43839
rect 85880 -43667 85934 -43655
rect 85880 -43701 85890 -43667
rect 85924 -43701 85934 -43667
rect 85880 -43735 85934 -43701
rect 85880 -43769 85890 -43735
rect 85924 -43769 85934 -43735
rect 85880 -43855 85934 -43769
rect 85964 -43667 86018 -43655
rect 85964 -43701 85974 -43667
rect 86008 -43701 86018 -43667
rect 85964 -43735 86018 -43701
rect 85964 -43769 85974 -43735
rect 86008 -43769 86018 -43735
rect 85964 -43805 86018 -43769
rect 85964 -43839 85974 -43805
rect 86008 -43839 86018 -43805
rect 85964 -43855 86018 -43839
rect 86048 -43667 86102 -43655
rect 86048 -43701 86058 -43667
rect 86092 -43701 86102 -43667
rect 86048 -43735 86102 -43701
rect 86048 -43769 86058 -43735
rect 86092 -43769 86102 -43735
rect 86048 -43855 86102 -43769
rect 86132 -43667 86186 -43655
rect 86132 -43701 86142 -43667
rect 86176 -43701 86186 -43667
rect 86132 -43735 86186 -43701
rect 86132 -43769 86142 -43735
rect 86176 -43769 86186 -43735
rect 86132 -43805 86186 -43769
rect 86132 -43839 86142 -43805
rect 86176 -43839 86186 -43805
rect 86132 -43855 86186 -43839
rect 86216 -43667 86270 -43655
rect 86216 -43701 86226 -43667
rect 86260 -43701 86270 -43667
rect 86216 -43735 86270 -43701
rect 86216 -43769 86226 -43735
rect 86260 -43769 86270 -43735
rect 86216 -43855 86270 -43769
rect 86300 -43667 86354 -43655
rect 86300 -43701 86310 -43667
rect 86344 -43701 86354 -43667
rect 86300 -43735 86354 -43701
rect 86300 -43769 86310 -43735
rect 86344 -43769 86354 -43735
rect 86300 -43805 86354 -43769
rect 86300 -43839 86310 -43805
rect 86344 -43839 86354 -43805
rect 86300 -43855 86354 -43839
rect 86384 -43667 86438 -43655
rect 86384 -43701 86394 -43667
rect 86428 -43701 86438 -43667
rect 86384 -43735 86438 -43701
rect 86384 -43769 86394 -43735
rect 86428 -43769 86438 -43735
rect 86384 -43855 86438 -43769
rect 86468 -43667 86522 -43655
rect 86468 -43701 86478 -43667
rect 86512 -43701 86522 -43667
rect 86468 -43735 86522 -43701
rect 86468 -43769 86478 -43735
rect 86512 -43769 86522 -43735
rect 86468 -43805 86522 -43769
rect 86468 -43839 86478 -43805
rect 86512 -43839 86522 -43805
rect 86468 -43855 86522 -43839
rect 86552 -43667 86606 -43655
rect 86552 -43701 86562 -43667
rect 86596 -43701 86606 -43667
rect 86552 -43735 86606 -43701
rect 86552 -43769 86562 -43735
rect 86596 -43769 86606 -43735
rect 86552 -43855 86606 -43769
rect 86636 -43667 86690 -43655
rect 86636 -43701 86646 -43667
rect 86680 -43701 86690 -43667
rect 86636 -43735 86690 -43701
rect 86636 -43769 86646 -43735
rect 86680 -43769 86690 -43735
rect 86636 -43805 86690 -43769
rect 86636 -43839 86646 -43805
rect 86680 -43839 86690 -43805
rect 86636 -43855 86690 -43839
rect 86720 -43667 86774 -43655
rect 86720 -43701 86730 -43667
rect 86764 -43701 86774 -43667
rect 86720 -43735 86774 -43701
rect 86720 -43769 86730 -43735
rect 86764 -43769 86774 -43735
rect 86720 -43855 86774 -43769
rect 86804 -43667 86858 -43655
rect 86804 -43701 86814 -43667
rect 86848 -43701 86858 -43667
rect 86804 -43735 86858 -43701
rect 86804 -43769 86814 -43735
rect 86848 -43769 86858 -43735
rect 86804 -43805 86858 -43769
rect 86804 -43839 86814 -43805
rect 86848 -43839 86858 -43805
rect 86804 -43855 86858 -43839
rect 86888 -43667 86940 -43655
rect 86888 -43701 86898 -43667
rect 86932 -43701 86940 -43667
rect 86888 -43735 86940 -43701
rect 86888 -43769 86898 -43735
rect 86932 -43769 86940 -43735
rect 86888 -43855 86940 -43769
rect 87018 -43667 87070 -43655
rect 87018 -43701 87026 -43667
rect 87060 -43701 87070 -43667
rect 87018 -43735 87070 -43701
rect 87018 -43769 87026 -43735
rect 87060 -43769 87070 -43735
rect 87018 -43805 87070 -43769
rect 87018 -43839 87026 -43805
rect 87060 -43839 87070 -43805
rect 87018 -43855 87070 -43839
rect 87100 -43667 87154 -43655
rect 87100 -43701 87110 -43667
rect 87144 -43701 87154 -43667
rect 87100 -43735 87154 -43701
rect 87100 -43769 87110 -43735
rect 87144 -43769 87154 -43735
rect 87100 -43805 87154 -43769
rect 87100 -43839 87110 -43805
rect 87144 -43839 87154 -43805
rect 87100 -43855 87154 -43839
rect 87184 -43667 87238 -43655
rect 87184 -43701 87194 -43667
rect 87228 -43701 87238 -43667
rect 87184 -43735 87238 -43701
rect 87184 -43769 87194 -43735
rect 87228 -43769 87238 -43735
rect 87184 -43855 87238 -43769
rect 87268 -43667 87322 -43655
rect 87268 -43701 87278 -43667
rect 87312 -43701 87322 -43667
rect 87268 -43735 87322 -43701
rect 87268 -43769 87278 -43735
rect 87312 -43769 87322 -43735
rect 87268 -43805 87322 -43769
rect 87268 -43839 87278 -43805
rect 87312 -43839 87322 -43805
rect 87268 -43855 87322 -43839
rect 87352 -43667 87406 -43655
rect 87352 -43701 87362 -43667
rect 87396 -43701 87406 -43667
rect 87352 -43735 87406 -43701
rect 87352 -43769 87362 -43735
rect 87396 -43769 87406 -43735
rect 87352 -43855 87406 -43769
rect 87436 -43667 87490 -43655
rect 87436 -43701 87446 -43667
rect 87480 -43701 87490 -43667
rect 87436 -43735 87490 -43701
rect 87436 -43769 87446 -43735
rect 87480 -43769 87490 -43735
rect 87436 -43805 87490 -43769
rect 87436 -43839 87446 -43805
rect 87480 -43839 87490 -43805
rect 87436 -43855 87490 -43839
rect 87520 -43667 87574 -43655
rect 87520 -43701 87530 -43667
rect 87564 -43701 87574 -43667
rect 87520 -43735 87574 -43701
rect 87520 -43769 87530 -43735
rect 87564 -43769 87574 -43735
rect 87520 -43855 87574 -43769
rect 87604 -43667 87658 -43655
rect 87604 -43701 87614 -43667
rect 87648 -43701 87658 -43667
rect 87604 -43735 87658 -43701
rect 87604 -43769 87614 -43735
rect 87648 -43769 87658 -43735
rect 87604 -43805 87658 -43769
rect 87604 -43839 87614 -43805
rect 87648 -43839 87658 -43805
rect 87604 -43855 87658 -43839
rect 87688 -43667 87742 -43655
rect 87688 -43701 87698 -43667
rect 87732 -43701 87742 -43667
rect 87688 -43735 87742 -43701
rect 87688 -43769 87698 -43735
rect 87732 -43769 87742 -43735
rect 87688 -43855 87742 -43769
rect 87772 -43667 87826 -43655
rect 87772 -43701 87782 -43667
rect 87816 -43701 87826 -43667
rect 87772 -43735 87826 -43701
rect 87772 -43769 87782 -43735
rect 87816 -43769 87826 -43735
rect 87772 -43805 87826 -43769
rect 87772 -43839 87782 -43805
rect 87816 -43839 87826 -43805
rect 87772 -43855 87826 -43839
rect 87856 -43667 87910 -43655
rect 87856 -43701 87866 -43667
rect 87900 -43701 87910 -43667
rect 87856 -43735 87910 -43701
rect 87856 -43769 87866 -43735
rect 87900 -43769 87910 -43735
rect 87856 -43855 87910 -43769
rect 87940 -43667 87994 -43655
rect 87940 -43701 87950 -43667
rect 87984 -43701 87994 -43667
rect 87940 -43735 87994 -43701
rect 87940 -43769 87950 -43735
rect 87984 -43769 87994 -43735
rect 87940 -43805 87994 -43769
rect 87940 -43839 87950 -43805
rect 87984 -43839 87994 -43805
rect 87940 -43855 87994 -43839
rect 88024 -43667 88078 -43655
rect 88024 -43701 88034 -43667
rect 88068 -43701 88078 -43667
rect 88024 -43735 88078 -43701
rect 88024 -43769 88034 -43735
rect 88068 -43769 88078 -43735
rect 88024 -43855 88078 -43769
rect 88108 -43667 88162 -43655
rect 88108 -43701 88118 -43667
rect 88152 -43701 88162 -43667
rect 88108 -43735 88162 -43701
rect 88108 -43769 88118 -43735
rect 88152 -43769 88162 -43735
rect 88108 -43805 88162 -43769
rect 88108 -43839 88118 -43805
rect 88152 -43839 88162 -43805
rect 88108 -43855 88162 -43839
rect 88192 -43667 88246 -43655
rect 88192 -43701 88202 -43667
rect 88236 -43701 88246 -43667
rect 88192 -43735 88246 -43701
rect 88192 -43769 88202 -43735
rect 88236 -43769 88246 -43735
rect 88192 -43855 88246 -43769
rect 88276 -43667 88330 -43655
rect 88276 -43701 88286 -43667
rect 88320 -43701 88330 -43667
rect 88276 -43735 88330 -43701
rect 88276 -43769 88286 -43735
rect 88320 -43769 88330 -43735
rect 88276 -43805 88330 -43769
rect 88276 -43839 88286 -43805
rect 88320 -43839 88330 -43805
rect 88276 -43855 88330 -43839
rect 88360 -43667 88412 -43655
rect 88360 -43701 88370 -43667
rect 88404 -43701 88412 -43667
rect 88360 -43735 88412 -43701
rect 88360 -43769 88370 -43735
rect 88404 -43769 88412 -43735
rect 88360 -43855 88412 -43769
rect 88490 -43667 88542 -43655
rect 88490 -43701 88498 -43667
rect 88532 -43701 88542 -43667
rect 88490 -43735 88542 -43701
rect 88490 -43769 88498 -43735
rect 88532 -43769 88542 -43735
rect 88490 -43805 88542 -43769
rect 88490 -43839 88498 -43805
rect 88532 -43839 88542 -43805
rect 88490 -43855 88542 -43839
rect 88572 -43667 88626 -43655
rect 88572 -43701 88582 -43667
rect 88616 -43701 88626 -43667
rect 88572 -43735 88626 -43701
rect 88572 -43769 88582 -43735
rect 88616 -43769 88626 -43735
rect 88572 -43805 88626 -43769
rect 88572 -43839 88582 -43805
rect 88616 -43839 88626 -43805
rect 88572 -43855 88626 -43839
rect 88656 -43667 88710 -43655
rect 88656 -43701 88666 -43667
rect 88700 -43701 88710 -43667
rect 88656 -43735 88710 -43701
rect 88656 -43769 88666 -43735
rect 88700 -43769 88710 -43735
rect 88656 -43855 88710 -43769
rect 88740 -43667 88794 -43655
rect 88740 -43701 88750 -43667
rect 88784 -43701 88794 -43667
rect 88740 -43735 88794 -43701
rect 88740 -43769 88750 -43735
rect 88784 -43769 88794 -43735
rect 88740 -43805 88794 -43769
rect 88740 -43839 88750 -43805
rect 88784 -43839 88794 -43805
rect 88740 -43855 88794 -43839
rect 88824 -43667 88878 -43655
rect 88824 -43701 88834 -43667
rect 88868 -43701 88878 -43667
rect 88824 -43735 88878 -43701
rect 88824 -43769 88834 -43735
rect 88868 -43769 88878 -43735
rect 88824 -43855 88878 -43769
rect 88908 -43667 88962 -43655
rect 88908 -43701 88918 -43667
rect 88952 -43701 88962 -43667
rect 88908 -43735 88962 -43701
rect 88908 -43769 88918 -43735
rect 88952 -43769 88962 -43735
rect 88908 -43805 88962 -43769
rect 88908 -43839 88918 -43805
rect 88952 -43839 88962 -43805
rect 88908 -43855 88962 -43839
rect 88992 -43667 89046 -43655
rect 88992 -43701 89002 -43667
rect 89036 -43701 89046 -43667
rect 88992 -43735 89046 -43701
rect 88992 -43769 89002 -43735
rect 89036 -43769 89046 -43735
rect 88992 -43855 89046 -43769
rect 89076 -43667 89130 -43655
rect 89076 -43701 89086 -43667
rect 89120 -43701 89130 -43667
rect 89076 -43735 89130 -43701
rect 89076 -43769 89086 -43735
rect 89120 -43769 89130 -43735
rect 89076 -43805 89130 -43769
rect 89076 -43839 89086 -43805
rect 89120 -43839 89130 -43805
rect 89076 -43855 89130 -43839
rect 89160 -43667 89214 -43655
rect 89160 -43701 89170 -43667
rect 89204 -43701 89214 -43667
rect 89160 -43735 89214 -43701
rect 89160 -43769 89170 -43735
rect 89204 -43769 89214 -43735
rect 89160 -43855 89214 -43769
rect 89244 -43667 89298 -43655
rect 89244 -43701 89254 -43667
rect 89288 -43701 89298 -43667
rect 89244 -43735 89298 -43701
rect 89244 -43769 89254 -43735
rect 89288 -43769 89298 -43735
rect 89244 -43805 89298 -43769
rect 89244 -43839 89254 -43805
rect 89288 -43839 89298 -43805
rect 89244 -43855 89298 -43839
rect 89328 -43667 89382 -43655
rect 89328 -43701 89338 -43667
rect 89372 -43701 89382 -43667
rect 89328 -43735 89382 -43701
rect 89328 -43769 89338 -43735
rect 89372 -43769 89382 -43735
rect 89328 -43855 89382 -43769
rect 89412 -43667 89466 -43655
rect 89412 -43701 89422 -43667
rect 89456 -43701 89466 -43667
rect 89412 -43735 89466 -43701
rect 89412 -43769 89422 -43735
rect 89456 -43769 89466 -43735
rect 89412 -43805 89466 -43769
rect 89412 -43839 89422 -43805
rect 89456 -43839 89466 -43805
rect 89412 -43855 89466 -43839
rect 89496 -43667 89550 -43655
rect 89496 -43701 89506 -43667
rect 89540 -43701 89550 -43667
rect 89496 -43735 89550 -43701
rect 89496 -43769 89506 -43735
rect 89540 -43769 89550 -43735
rect 89496 -43855 89550 -43769
rect 89580 -43667 89634 -43655
rect 89580 -43701 89590 -43667
rect 89624 -43701 89634 -43667
rect 89580 -43735 89634 -43701
rect 89580 -43769 89590 -43735
rect 89624 -43769 89634 -43735
rect 89580 -43805 89634 -43769
rect 89580 -43839 89590 -43805
rect 89624 -43839 89634 -43805
rect 89580 -43855 89634 -43839
rect 89664 -43667 89718 -43655
rect 89664 -43701 89674 -43667
rect 89708 -43701 89718 -43667
rect 89664 -43735 89718 -43701
rect 89664 -43769 89674 -43735
rect 89708 -43769 89718 -43735
rect 89664 -43855 89718 -43769
rect 89748 -43667 89802 -43655
rect 89748 -43701 89758 -43667
rect 89792 -43701 89802 -43667
rect 89748 -43735 89802 -43701
rect 89748 -43769 89758 -43735
rect 89792 -43769 89802 -43735
rect 89748 -43805 89802 -43769
rect 89748 -43839 89758 -43805
rect 89792 -43839 89802 -43805
rect 89748 -43855 89802 -43839
rect 89832 -43667 89884 -43655
rect 89832 -43701 89842 -43667
rect 89876 -43701 89884 -43667
rect 89832 -43735 89884 -43701
rect 89832 -43769 89842 -43735
rect 89876 -43769 89884 -43735
rect 89832 -43855 89884 -43769
rect 89962 -43667 90014 -43655
rect 89962 -43701 89970 -43667
rect 90004 -43701 90014 -43667
rect 89962 -43735 90014 -43701
rect 89962 -43769 89970 -43735
rect 90004 -43769 90014 -43735
rect 89962 -43805 90014 -43769
rect 89962 -43839 89970 -43805
rect 90004 -43839 90014 -43805
rect 89962 -43855 90014 -43839
rect 90044 -43667 90098 -43655
rect 90044 -43701 90054 -43667
rect 90088 -43701 90098 -43667
rect 90044 -43735 90098 -43701
rect 90044 -43769 90054 -43735
rect 90088 -43769 90098 -43735
rect 90044 -43805 90098 -43769
rect 90044 -43839 90054 -43805
rect 90088 -43839 90098 -43805
rect 90044 -43855 90098 -43839
rect 90128 -43667 90182 -43655
rect 90128 -43701 90138 -43667
rect 90172 -43701 90182 -43667
rect 90128 -43735 90182 -43701
rect 90128 -43769 90138 -43735
rect 90172 -43769 90182 -43735
rect 90128 -43855 90182 -43769
rect 90212 -43667 90266 -43655
rect 90212 -43701 90222 -43667
rect 90256 -43701 90266 -43667
rect 90212 -43735 90266 -43701
rect 90212 -43769 90222 -43735
rect 90256 -43769 90266 -43735
rect 90212 -43805 90266 -43769
rect 90212 -43839 90222 -43805
rect 90256 -43839 90266 -43805
rect 90212 -43855 90266 -43839
rect 90296 -43667 90350 -43655
rect 90296 -43701 90306 -43667
rect 90340 -43701 90350 -43667
rect 90296 -43735 90350 -43701
rect 90296 -43769 90306 -43735
rect 90340 -43769 90350 -43735
rect 90296 -43855 90350 -43769
rect 90380 -43667 90434 -43655
rect 90380 -43701 90390 -43667
rect 90424 -43701 90434 -43667
rect 90380 -43735 90434 -43701
rect 90380 -43769 90390 -43735
rect 90424 -43769 90434 -43735
rect 90380 -43805 90434 -43769
rect 90380 -43839 90390 -43805
rect 90424 -43839 90434 -43805
rect 90380 -43855 90434 -43839
rect 90464 -43667 90518 -43655
rect 90464 -43701 90474 -43667
rect 90508 -43701 90518 -43667
rect 90464 -43735 90518 -43701
rect 90464 -43769 90474 -43735
rect 90508 -43769 90518 -43735
rect 90464 -43855 90518 -43769
rect 90548 -43667 90602 -43655
rect 90548 -43701 90558 -43667
rect 90592 -43701 90602 -43667
rect 90548 -43735 90602 -43701
rect 90548 -43769 90558 -43735
rect 90592 -43769 90602 -43735
rect 90548 -43805 90602 -43769
rect 90548 -43839 90558 -43805
rect 90592 -43839 90602 -43805
rect 90548 -43855 90602 -43839
rect 90632 -43667 90686 -43655
rect 90632 -43701 90642 -43667
rect 90676 -43701 90686 -43667
rect 90632 -43735 90686 -43701
rect 90632 -43769 90642 -43735
rect 90676 -43769 90686 -43735
rect 90632 -43855 90686 -43769
rect 90716 -43667 90770 -43655
rect 90716 -43701 90726 -43667
rect 90760 -43701 90770 -43667
rect 90716 -43735 90770 -43701
rect 90716 -43769 90726 -43735
rect 90760 -43769 90770 -43735
rect 90716 -43805 90770 -43769
rect 90716 -43839 90726 -43805
rect 90760 -43839 90770 -43805
rect 90716 -43855 90770 -43839
rect 90800 -43667 90854 -43655
rect 90800 -43701 90810 -43667
rect 90844 -43701 90854 -43667
rect 90800 -43735 90854 -43701
rect 90800 -43769 90810 -43735
rect 90844 -43769 90854 -43735
rect 90800 -43855 90854 -43769
rect 90884 -43667 90938 -43655
rect 90884 -43701 90894 -43667
rect 90928 -43701 90938 -43667
rect 90884 -43735 90938 -43701
rect 90884 -43769 90894 -43735
rect 90928 -43769 90938 -43735
rect 90884 -43805 90938 -43769
rect 90884 -43839 90894 -43805
rect 90928 -43839 90938 -43805
rect 90884 -43855 90938 -43839
rect 90968 -43667 91022 -43655
rect 90968 -43701 90978 -43667
rect 91012 -43701 91022 -43667
rect 90968 -43735 91022 -43701
rect 90968 -43769 90978 -43735
rect 91012 -43769 91022 -43735
rect 90968 -43855 91022 -43769
rect 91052 -43667 91106 -43655
rect 91052 -43701 91062 -43667
rect 91096 -43701 91106 -43667
rect 91052 -43735 91106 -43701
rect 91052 -43769 91062 -43735
rect 91096 -43769 91106 -43735
rect 91052 -43805 91106 -43769
rect 91052 -43839 91062 -43805
rect 91096 -43839 91106 -43805
rect 91052 -43855 91106 -43839
rect 91136 -43667 91190 -43655
rect 91136 -43701 91146 -43667
rect 91180 -43701 91190 -43667
rect 91136 -43735 91190 -43701
rect 91136 -43769 91146 -43735
rect 91180 -43769 91190 -43735
rect 91136 -43855 91190 -43769
rect 91220 -43667 91274 -43655
rect 91220 -43701 91230 -43667
rect 91264 -43701 91274 -43667
rect 91220 -43735 91274 -43701
rect 91220 -43769 91230 -43735
rect 91264 -43769 91274 -43735
rect 91220 -43805 91274 -43769
rect 91220 -43839 91230 -43805
rect 91264 -43839 91274 -43805
rect 91220 -43855 91274 -43839
rect 91304 -43667 91356 -43655
rect 91304 -43701 91314 -43667
rect 91348 -43701 91356 -43667
rect 91304 -43735 91356 -43701
rect 91304 -43769 91314 -43735
rect 91348 -43769 91356 -43735
rect 91304 -43855 91356 -43769
rect 78143 -43899 78153 -43865
rect 78187 -43899 78195 -43865
rect 78143 -43911 78195 -43899
rect 77605 -44089 77657 -44077
rect 77605 -44123 77613 -44089
rect 77647 -44123 77657 -44089
rect 77605 -44161 77657 -44123
rect 77687 -44097 77757 -44077
rect 77687 -44131 77705 -44097
rect 77739 -44131 77757 -44097
rect 77687 -44161 77757 -44131
rect 77787 -44089 77861 -44077
rect 77787 -44123 77807 -44089
rect 77841 -44123 77861 -44089
rect 77787 -44161 77861 -44123
rect 77891 -44097 77947 -44077
rect 77891 -44131 77902 -44097
rect 77936 -44131 77947 -44097
rect 77891 -44161 77947 -44131
rect 77977 -44089 78113 -44077
rect 77977 -44123 78053 -44089
rect 78087 -44123 78113 -44089
rect 77977 -44157 78113 -44123
rect 77977 -44161 78053 -44157
rect 77996 -44191 78053 -44161
rect 78087 -44191 78113 -44157
rect 77996 -44277 78113 -44191
rect 78143 -44089 78195 -44077
rect 78143 -44123 78153 -44089
rect 78187 -44123 78195 -44089
rect 78143 -44157 78195 -44123
rect 78143 -44191 78153 -44157
rect 78187 -44191 78195 -44157
rect 78143 -44225 78195 -44191
rect 78143 -44259 78153 -44225
rect 78187 -44259 78195 -44225
rect 78143 -44277 78195 -44259
rect 54079 -44872 54879 -44860
rect 54079 -44906 54091 -44872
rect 54867 -44906 54879 -44872
rect 54079 -44918 54879 -44906
rect 54079 -45000 54879 -44988
rect 54079 -45034 54091 -45000
rect 54867 -45034 54879 -45000
rect 54079 -45046 54879 -45034
rect 77996 -45031 78113 -44945
rect 77996 -45061 78053 -45031
rect 54079 -45228 54879 -45216
rect 54079 -45262 54091 -45228
rect 54867 -45262 54879 -45228
rect 54079 -45274 54879 -45262
rect 54079 -45356 54879 -45344
rect 54079 -45390 54091 -45356
rect 54867 -45390 54879 -45356
rect 54079 -45402 54879 -45390
rect 77605 -45099 77657 -45061
rect 77605 -45133 77613 -45099
rect 77647 -45133 77657 -45099
rect 77605 -45145 77657 -45133
rect 77687 -45091 77757 -45061
rect 77687 -45125 77705 -45091
rect 77739 -45125 77757 -45091
rect 77687 -45145 77757 -45125
rect 77787 -45099 77861 -45061
rect 77787 -45133 77807 -45099
rect 77841 -45133 77861 -45099
rect 77787 -45145 77861 -45133
rect 77891 -45091 77947 -45061
rect 77891 -45125 77902 -45091
rect 77936 -45125 77947 -45091
rect 77891 -45145 77947 -45125
rect 77977 -45065 78053 -45061
rect 78087 -45065 78113 -45031
rect 77977 -45099 78113 -45065
rect 77977 -45133 78053 -45099
rect 78087 -45133 78113 -45099
rect 77977 -45145 78113 -45133
rect 78143 -44963 78195 -44945
rect 78143 -44997 78153 -44963
rect 78187 -44997 78195 -44963
rect 78143 -45031 78195 -44997
rect 78143 -45065 78153 -45031
rect 78187 -45065 78195 -45031
rect 78143 -45099 78195 -45065
rect 78143 -45133 78153 -45099
rect 78187 -45133 78195 -45099
rect 78143 -45145 78195 -45133
rect 57123 -45329 57175 -45309
rect 57123 -45363 57131 -45329
rect 57165 -45363 57175 -45329
rect 57123 -45397 57175 -45363
rect 57123 -45431 57131 -45397
rect 57165 -45431 57175 -45397
rect 57123 -45467 57175 -45431
rect 57205 -45329 57263 -45309
rect 57205 -45363 57217 -45329
rect 57251 -45363 57263 -45329
rect 57205 -45397 57263 -45363
rect 57205 -45431 57217 -45397
rect 57251 -45431 57263 -45397
rect 57205 -45467 57263 -45431
rect 57293 -45329 57345 -45309
rect 57293 -45363 57303 -45329
rect 57337 -45363 57345 -45329
rect 57293 -45410 57345 -45363
rect 57293 -45444 57303 -45410
rect 57337 -45444 57345 -45410
rect 57293 -45467 57345 -45444
rect 59113 -45247 59513 -45235
rect 59113 -45281 59125 -45247
rect 59501 -45281 59513 -45247
rect 59113 -45293 59513 -45281
rect 59113 -45355 59513 -45343
rect 59113 -45389 59125 -45355
rect 59501 -45389 59513 -45355
rect 59113 -45401 59513 -45389
rect 59113 -45463 59513 -45451
rect 59113 -45497 59125 -45463
rect 59501 -45497 59513 -45463
rect 59113 -45509 59513 -45497
rect 77877 -45327 77929 -45315
rect 77877 -45361 77885 -45327
rect 77919 -45361 77929 -45327
rect 77877 -45374 77929 -45361
rect 77879 -45428 77929 -45374
rect 54069 -47188 54869 -47176
rect 54069 -47222 54081 -47188
rect 54857 -47222 54869 -47188
rect 54069 -47234 54869 -47222
rect 54069 -47316 54869 -47304
rect 54069 -47350 54081 -47316
rect 54857 -47350 54869 -47316
rect 54069 -47362 54869 -47350
rect 56418 -45899 56476 -45887
rect 56418 -46675 56430 -45899
rect 56464 -46675 56476 -45899
rect 56418 -46687 56476 -46675
rect 56546 -45899 56604 -45887
rect 56546 -46675 56558 -45899
rect 56592 -46675 56604 -45899
rect 56546 -46687 56604 -46675
rect 59032 -45771 59090 -45759
rect 59032 -46147 59044 -45771
rect 59078 -46147 59090 -45771
rect 59032 -46159 59090 -46147
rect 59150 -45771 59208 -45759
rect 59150 -46147 59162 -45771
rect 59196 -46147 59208 -45771
rect 59150 -46159 59208 -46147
rect 77605 -45466 77657 -45428
rect 77605 -45500 77613 -45466
rect 77647 -45500 77657 -45466
rect 77605 -45512 77657 -45500
rect 77687 -45436 77741 -45428
rect 77687 -45470 77697 -45436
rect 77731 -45470 77741 -45436
rect 77687 -45512 77741 -45470
rect 77771 -45455 77834 -45428
rect 77771 -45489 77790 -45455
rect 77824 -45489 77834 -45455
rect 77771 -45512 77834 -45489
rect 77864 -45512 77929 -45428
rect 77879 -45515 77929 -45512
rect 77959 -45341 78011 -45315
rect 78293 -45327 78345 -45315
rect 77959 -45375 77969 -45341
rect 78003 -45375 78011 -45341
rect 78293 -45357 78301 -45327
rect 77959 -45409 78011 -45375
rect 77959 -45443 77969 -45409
rect 78003 -45443 78011 -45409
rect 78097 -45369 78153 -45357
rect 78097 -45403 78109 -45369
rect 78143 -45403 78153 -45369
rect 78097 -45441 78153 -45403
rect 78183 -45369 78237 -45357
rect 78183 -45403 78193 -45369
rect 78227 -45403 78237 -45369
rect 78183 -45441 78237 -45403
rect 78267 -45361 78301 -45357
rect 78335 -45361 78345 -45327
rect 78267 -45395 78345 -45361
rect 78267 -45429 78301 -45395
rect 78335 -45429 78345 -45395
rect 78267 -45441 78345 -45429
rect 77959 -45515 78011 -45443
rect 78283 -45515 78345 -45441
rect 78375 -45327 78470 -45315
rect 78375 -45361 78405 -45327
rect 78439 -45361 78470 -45327
rect 78886 -45327 78939 -45315
rect 78375 -45395 78470 -45361
rect 78886 -45361 78894 -45327
rect 78928 -45361 78939 -45327
rect 78375 -45429 78405 -45395
rect 78439 -45429 78470 -45395
rect 78375 -45515 78470 -45429
rect 78886 -45395 78939 -45361
rect 78886 -45429 78894 -45395
rect 78928 -45429 78939 -45395
rect 78886 -45431 78939 -45429
rect 78525 -45458 78577 -45431
rect 78525 -45492 78533 -45458
rect 78567 -45492 78577 -45458
rect 78525 -45515 78577 -45492
rect 78607 -45515 78673 -45431
rect 78703 -45515 78745 -45431
rect 78775 -45515 78841 -45431
rect 78871 -45515 78939 -45431
rect 78969 -45358 79023 -45315
rect 78969 -45392 78979 -45358
rect 79013 -45392 79023 -45358
rect 78969 -45426 79023 -45392
rect 78969 -45460 78979 -45426
rect 79013 -45460 79023 -45426
rect 78969 -45515 79023 -45460
rect 60441 -46173 60641 -46165
rect 60441 -46207 60459 -46173
rect 60493 -46207 60527 -46173
rect 60561 -46207 60595 -46173
rect 60629 -46207 60641 -46173
rect 60441 -46217 60641 -46207
rect 60811 -46173 61011 -46165
rect 60811 -46207 60823 -46173
rect 60857 -46207 60891 -46173
rect 60925 -46207 60959 -46173
rect 60993 -46207 61011 -46173
rect 60811 -46217 61011 -46207
rect 60441 -46257 60641 -46247
rect 60441 -46291 60459 -46257
rect 60493 -46291 60527 -46257
rect 60561 -46291 60595 -46257
rect 60629 -46291 60641 -46257
rect 60441 -46301 60641 -46291
rect 60811 -46257 61011 -46247
rect 60811 -46291 60823 -46257
rect 60857 -46291 60891 -46257
rect 60925 -46291 60959 -46257
rect 60993 -46291 61011 -46257
rect 60811 -46301 61011 -46291
rect 59032 -46501 59090 -46489
rect 59032 -46877 59044 -46501
rect 59078 -46877 59090 -46501
rect 59032 -46889 59090 -46877
rect 59150 -46501 59208 -46489
rect 59150 -46877 59162 -46501
rect 59196 -46877 59208 -46501
rect 59150 -46889 59208 -46877
rect 60441 -46341 60641 -46331
rect 60441 -46375 60527 -46341
rect 60561 -46375 60595 -46341
rect 60629 -46375 60641 -46341
rect 60441 -46385 60641 -46375
rect 60811 -46341 61011 -46331
rect 60811 -46375 60823 -46341
rect 60857 -46375 60891 -46341
rect 60925 -46375 61011 -46341
rect 60811 -46385 61011 -46375
rect 60441 -46425 60641 -46415
rect 60441 -46459 60459 -46425
rect 60493 -46459 60527 -46425
rect 60561 -46459 60595 -46425
rect 60629 -46459 60641 -46425
rect 60441 -46469 60641 -46459
rect 60811 -46425 61011 -46415
rect 60811 -46459 60823 -46425
rect 60857 -46459 60891 -46425
rect 60925 -46459 60959 -46425
rect 60993 -46459 61011 -46425
rect 60811 -46469 61011 -46459
rect 60441 -46509 60641 -46499
rect 60441 -46543 60595 -46509
rect 60629 -46543 60641 -46509
rect 60441 -46551 60641 -46543
rect 60811 -46509 61011 -46499
rect 60811 -46543 60823 -46509
rect 60857 -46543 61011 -46509
rect 60811 -46551 61011 -46543
rect 75574 -46743 75626 -46725
rect 75574 -46777 75582 -46743
rect 75616 -46777 75626 -46743
rect 75574 -46811 75626 -46777
rect 57123 -47157 57175 -47121
rect 57123 -47191 57131 -47157
rect 57165 -47191 57175 -47157
rect 57123 -47225 57175 -47191
rect 57123 -47259 57131 -47225
rect 57165 -47259 57175 -47225
rect 57123 -47279 57175 -47259
rect 57205 -47157 57263 -47121
rect 57205 -47191 57217 -47157
rect 57251 -47191 57263 -47157
rect 57205 -47225 57263 -47191
rect 57205 -47259 57217 -47225
rect 57251 -47259 57263 -47225
rect 57205 -47279 57263 -47259
rect 57293 -47144 57345 -47121
rect 57293 -47178 57303 -47144
rect 57337 -47178 57345 -47144
rect 57293 -47225 57345 -47178
rect 57293 -47259 57303 -47225
rect 57337 -47259 57345 -47225
rect 57293 -47279 57345 -47259
rect 59113 -47154 59513 -47142
rect 59113 -47188 59125 -47154
rect 59501 -47188 59513 -47154
rect 59113 -47200 59513 -47188
rect 59113 -47262 59513 -47250
rect 59113 -47296 59125 -47262
rect 59501 -47296 59513 -47262
rect 59113 -47308 59513 -47296
rect 59113 -47370 59513 -47358
rect 59113 -47404 59125 -47370
rect 59501 -47404 59513 -47370
rect 59113 -47416 59513 -47404
rect 54069 -47544 54869 -47532
rect 54069 -47578 54081 -47544
rect 54857 -47578 54869 -47544
rect 54069 -47590 54869 -47578
rect 54069 -47672 54869 -47660
rect 54069 -47706 54081 -47672
rect 54857 -47706 54869 -47672
rect 54069 -47718 54869 -47706
rect 75574 -46845 75582 -46811
rect 75616 -46845 75626 -46811
rect 75574 -46879 75626 -46845
rect 75574 -46913 75582 -46879
rect 75616 -46913 75626 -46879
rect 75574 -46925 75626 -46913
rect 75656 -46743 75708 -46725
rect 75656 -46777 75666 -46743
rect 75700 -46777 75708 -46743
rect 75656 -46811 75708 -46777
rect 75656 -46845 75666 -46811
rect 75700 -46845 75708 -46811
rect 75656 -46879 75708 -46845
rect 75656 -46913 75666 -46879
rect 75700 -46913 75708 -46879
rect 75656 -46925 75708 -46913
rect 75850 -46743 75902 -46725
rect 75850 -46777 75858 -46743
rect 75892 -46777 75902 -46743
rect 75850 -46811 75902 -46777
rect 75850 -46845 75858 -46811
rect 75892 -46845 75902 -46811
rect 75850 -46879 75902 -46845
rect 75850 -46913 75858 -46879
rect 75892 -46913 75902 -46879
rect 75850 -46925 75902 -46913
rect 75932 -46743 75984 -46725
rect 75932 -46777 75942 -46743
rect 75976 -46777 75984 -46743
rect 75932 -46811 75984 -46777
rect 75932 -46845 75942 -46811
rect 75976 -46845 75984 -46811
rect 75932 -46879 75984 -46845
rect 75932 -46913 75942 -46879
rect 75976 -46913 75984 -46879
rect 75932 -46925 75984 -46913
rect 76124 -46743 76176 -46725
rect 76124 -46777 76132 -46743
rect 76166 -46777 76176 -46743
rect 76124 -46811 76176 -46777
rect 76124 -46845 76132 -46811
rect 76166 -46845 76176 -46811
rect 76124 -46879 76176 -46845
rect 76124 -46913 76132 -46879
rect 76166 -46913 76176 -46879
rect 76124 -46925 76176 -46913
rect 76206 -46743 76258 -46725
rect 76206 -46777 76216 -46743
rect 76250 -46777 76258 -46743
rect 76206 -46811 76258 -46777
rect 76206 -46845 76216 -46811
rect 76250 -46845 76258 -46811
rect 76206 -46879 76258 -46845
rect 76206 -46913 76216 -46879
rect 76250 -46913 76258 -46879
rect 76206 -46925 76258 -46913
rect 76400 -46743 76452 -46725
rect 76400 -46777 76408 -46743
rect 76442 -46777 76452 -46743
rect 76400 -46811 76452 -46777
rect 76400 -46845 76408 -46811
rect 76442 -46845 76452 -46811
rect 76400 -46879 76452 -46845
rect 76400 -46913 76408 -46879
rect 76442 -46913 76452 -46879
rect 76400 -46925 76452 -46913
rect 76482 -46743 76534 -46725
rect 76482 -46777 76492 -46743
rect 76526 -46777 76534 -46743
rect 76482 -46811 76534 -46777
rect 76482 -46845 76492 -46811
rect 76526 -46845 76534 -46811
rect 76482 -46879 76534 -46845
rect 76482 -46913 76492 -46879
rect 76526 -46913 76534 -46879
rect 76482 -46925 76534 -46913
rect 76676 -46743 76728 -46725
rect 76676 -46777 76684 -46743
rect 76718 -46777 76728 -46743
rect 76676 -46811 76728 -46777
rect 76676 -46845 76684 -46811
rect 76718 -46845 76728 -46811
rect 76676 -46879 76728 -46845
rect 76676 -46913 76684 -46879
rect 76718 -46913 76728 -46879
rect 76676 -46925 76728 -46913
rect 76758 -46743 76810 -46725
rect 76758 -46777 76768 -46743
rect 76802 -46777 76810 -46743
rect 76758 -46811 76810 -46777
rect 76758 -46845 76768 -46811
rect 76802 -46845 76810 -46811
rect 76758 -46879 76810 -46845
rect 76758 -46913 76768 -46879
rect 76802 -46913 76810 -46879
rect 76758 -46925 76810 -46913
rect 77966 -47157 78019 -47145
rect 77966 -47191 77974 -47157
rect 78008 -47191 78019 -47157
rect 77966 -47225 78019 -47191
rect 77966 -47259 77974 -47225
rect 78008 -47259 78019 -47225
rect 77966 -47261 78019 -47259
rect 77605 -47288 77657 -47261
rect 77605 -47322 77613 -47288
rect 77647 -47322 77657 -47288
rect 77605 -47345 77657 -47322
rect 77687 -47345 77753 -47261
rect 77783 -47345 77825 -47261
rect 77855 -47345 77921 -47261
rect 77951 -47345 78019 -47261
rect 78049 -47188 78103 -47145
rect 78424 -47157 78477 -47145
rect 78049 -47222 78059 -47188
rect 78093 -47222 78103 -47188
rect 78424 -47191 78432 -47157
rect 78466 -47191 78477 -47157
rect 78049 -47256 78103 -47222
rect 78049 -47290 78059 -47256
rect 78093 -47290 78103 -47256
rect 78424 -47225 78477 -47191
rect 78424 -47259 78432 -47225
rect 78466 -47259 78477 -47225
rect 78424 -47261 78477 -47259
rect 78049 -47345 78103 -47290
rect 78159 -47288 78211 -47261
rect 78159 -47322 78167 -47288
rect 78201 -47322 78211 -47288
rect 78159 -47345 78211 -47322
rect 78241 -47345 78283 -47261
rect 78313 -47345 78379 -47261
rect 78409 -47345 78477 -47261
rect 78507 -47188 78563 -47145
rect 78845 -47157 78897 -47145
rect 78845 -47187 78853 -47157
rect 78507 -47222 78517 -47188
rect 78551 -47222 78563 -47188
rect 78507 -47256 78563 -47222
rect 78507 -47290 78517 -47256
rect 78551 -47290 78563 -47256
rect 78649 -47199 78705 -47187
rect 78649 -47233 78661 -47199
rect 78695 -47233 78705 -47199
rect 78649 -47271 78705 -47233
rect 78735 -47199 78789 -47187
rect 78735 -47233 78745 -47199
rect 78779 -47233 78789 -47199
rect 78735 -47271 78789 -47233
rect 78819 -47191 78853 -47187
rect 78887 -47191 78897 -47157
rect 78819 -47225 78897 -47191
rect 78819 -47259 78853 -47225
rect 78887 -47259 78897 -47225
rect 78819 -47271 78897 -47259
rect 78507 -47345 78563 -47290
rect 78835 -47345 78897 -47271
rect 78927 -47157 79022 -47145
rect 78927 -47191 78957 -47157
rect 78991 -47191 79022 -47157
rect 78927 -47225 79022 -47191
rect 78927 -47259 78957 -47225
rect 78991 -47259 79022 -47225
rect 78927 -47345 79022 -47259
rect 83075 -47823 83127 -47795
rect 83075 -47857 83083 -47823
rect 83117 -47857 83127 -47823
rect 83075 -47891 83127 -47857
rect 83075 -47911 83083 -47891
rect 82906 -47943 82958 -47911
rect 82906 -47977 82914 -47943
rect 82948 -47977 82958 -47943
rect 82906 -47995 82958 -47977
rect 82988 -47995 83030 -47911
rect 83060 -47925 83083 -47911
rect 83117 -47925 83127 -47891
rect 83060 -47995 83127 -47925
rect 83157 -47807 83225 -47795
rect 83157 -47841 83183 -47807
rect 83217 -47841 83225 -47807
rect 83157 -47875 83225 -47841
rect 83157 -47909 83183 -47875
rect 83217 -47909 83225 -47875
rect 83157 -47995 83225 -47909
rect 83366 -47807 83418 -47795
rect 83366 -47841 83374 -47807
rect 83408 -47841 83418 -47807
rect 83366 -47875 83418 -47841
rect 83366 -47909 83374 -47875
rect 83408 -47909 83418 -47875
rect 83366 -47943 83418 -47909
rect 83366 -47977 83374 -47943
rect 83408 -47977 83418 -47943
rect 83366 -47995 83418 -47977
rect 83448 -47807 83500 -47795
rect 83448 -47841 83458 -47807
rect 83492 -47841 83500 -47807
rect 83448 -47875 83500 -47841
rect 83448 -47909 83458 -47875
rect 83492 -47909 83500 -47875
rect 83448 -47943 83500 -47909
rect 83448 -47977 83458 -47943
rect 83492 -47977 83500 -47943
rect 83448 -47995 83500 -47977
rect 83611 -47807 83663 -47795
rect 83611 -47841 83619 -47807
rect 83653 -47841 83663 -47807
rect 83611 -47875 83663 -47841
rect 83611 -47909 83619 -47875
rect 83653 -47909 83663 -47875
rect 83611 -47943 83663 -47909
rect 83611 -47977 83619 -47943
rect 83653 -47977 83663 -47943
rect 83611 -47995 83663 -47977
rect 83693 -47807 83747 -47795
rect 83693 -47841 83703 -47807
rect 83737 -47841 83747 -47807
rect 83693 -47875 83747 -47841
rect 83693 -47909 83703 -47875
rect 83737 -47909 83747 -47875
rect 83693 -47943 83747 -47909
rect 83693 -47977 83703 -47943
rect 83737 -47977 83747 -47943
rect 83693 -47995 83747 -47977
rect 83777 -47807 83831 -47795
rect 83777 -47841 83787 -47807
rect 83821 -47841 83831 -47807
rect 83777 -47875 83831 -47841
rect 83777 -47909 83787 -47875
rect 83821 -47909 83831 -47875
rect 83777 -47995 83831 -47909
rect 83861 -47807 83915 -47795
rect 83861 -47841 83871 -47807
rect 83905 -47841 83915 -47807
rect 83861 -47875 83915 -47841
rect 83861 -47909 83871 -47875
rect 83905 -47909 83915 -47875
rect 83861 -47943 83915 -47909
rect 83861 -47977 83871 -47943
rect 83905 -47977 83915 -47943
rect 83861 -47995 83915 -47977
rect 83945 -47807 83997 -47795
rect 83945 -47841 83955 -47807
rect 83989 -47841 83997 -47807
rect 83945 -47995 83997 -47841
rect 84074 -47807 84126 -47795
rect 84074 -47841 84082 -47807
rect 84116 -47841 84126 -47807
rect 84074 -47875 84126 -47841
rect 84074 -47909 84082 -47875
rect 84116 -47909 84126 -47875
rect 84074 -47945 84126 -47909
rect 84074 -47979 84082 -47945
rect 84116 -47979 84126 -47945
rect 84074 -47995 84126 -47979
rect 84156 -47807 84210 -47795
rect 84156 -47841 84166 -47807
rect 84200 -47841 84210 -47807
rect 84156 -47875 84210 -47841
rect 84156 -47909 84166 -47875
rect 84200 -47909 84210 -47875
rect 84156 -47945 84210 -47909
rect 84156 -47979 84166 -47945
rect 84200 -47979 84210 -47945
rect 84156 -47995 84210 -47979
rect 84240 -47807 84294 -47795
rect 84240 -47841 84250 -47807
rect 84284 -47841 84294 -47807
rect 84240 -47875 84294 -47841
rect 84240 -47909 84250 -47875
rect 84284 -47909 84294 -47875
rect 84240 -47995 84294 -47909
rect 84324 -47807 84378 -47795
rect 84324 -47841 84334 -47807
rect 84368 -47841 84378 -47807
rect 84324 -47875 84378 -47841
rect 84324 -47909 84334 -47875
rect 84368 -47909 84378 -47875
rect 84324 -47945 84378 -47909
rect 84324 -47979 84334 -47945
rect 84368 -47979 84378 -47945
rect 84324 -47995 84378 -47979
rect 84408 -47807 84462 -47795
rect 84408 -47841 84418 -47807
rect 84452 -47841 84462 -47807
rect 84408 -47875 84462 -47841
rect 84408 -47909 84418 -47875
rect 84452 -47909 84462 -47875
rect 84408 -47995 84462 -47909
rect 84492 -47807 84546 -47795
rect 84492 -47841 84502 -47807
rect 84536 -47841 84546 -47807
rect 84492 -47875 84546 -47841
rect 84492 -47909 84502 -47875
rect 84536 -47909 84546 -47875
rect 84492 -47945 84546 -47909
rect 84492 -47979 84502 -47945
rect 84536 -47979 84546 -47945
rect 84492 -47995 84546 -47979
rect 84576 -47807 84630 -47795
rect 84576 -47841 84586 -47807
rect 84620 -47841 84630 -47807
rect 84576 -47875 84630 -47841
rect 84576 -47909 84586 -47875
rect 84620 -47909 84630 -47875
rect 84576 -47995 84630 -47909
rect 84660 -47807 84714 -47795
rect 84660 -47841 84670 -47807
rect 84704 -47841 84714 -47807
rect 84660 -47875 84714 -47841
rect 84660 -47909 84670 -47875
rect 84704 -47909 84714 -47875
rect 84660 -47945 84714 -47909
rect 84660 -47979 84670 -47945
rect 84704 -47979 84714 -47945
rect 84660 -47995 84714 -47979
rect 84744 -47807 84798 -47795
rect 84744 -47841 84754 -47807
rect 84788 -47841 84798 -47807
rect 84744 -47875 84798 -47841
rect 84744 -47909 84754 -47875
rect 84788 -47909 84798 -47875
rect 84744 -47995 84798 -47909
rect 84828 -47807 84882 -47795
rect 84828 -47841 84838 -47807
rect 84872 -47841 84882 -47807
rect 84828 -47875 84882 -47841
rect 84828 -47909 84838 -47875
rect 84872 -47909 84882 -47875
rect 84828 -47945 84882 -47909
rect 84828 -47979 84838 -47945
rect 84872 -47979 84882 -47945
rect 84828 -47995 84882 -47979
rect 84912 -47807 84966 -47795
rect 84912 -47841 84922 -47807
rect 84956 -47841 84966 -47807
rect 84912 -47875 84966 -47841
rect 84912 -47909 84922 -47875
rect 84956 -47909 84966 -47875
rect 84912 -47995 84966 -47909
rect 84996 -47807 85050 -47795
rect 84996 -47841 85006 -47807
rect 85040 -47841 85050 -47807
rect 84996 -47875 85050 -47841
rect 84996 -47909 85006 -47875
rect 85040 -47909 85050 -47875
rect 84996 -47945 85050 -47909
rect 84996 -47979 85006 -47945
rect 85040 -47979 85050 -47945
rect 84996 -47995 85050 -47979
rect 85080 -47807 85134 -47795
rect 85080 -47841 85090 -47807
rect 85124 -47841 85134 -47807
rect 85080 -47875 85134 -47841
rect 85080 -47909 85090 -47875
rect 85124 -47909 85134 -47875
rect 85080 -47995 85134 -47909
rect 85164 -47807 85218 -47795
rect 85164 -47841 85174 -47807
rect 85208 -47841 85218 -47807
rect 85164 -47875 85218 -47841
rect 85164 -47909 85174 -47875
rect 85208 -47909 85218 -47875
rect 85164 -47945 85218 -47909
rect 85164 -47979 85174 -47945
rect 85208 -47979 85218 -47945
rect 85164 -47995 85218 -47979
rect 85248 -47807 85302 -47795
rect 85248 -47841 85258 -47807
rect 85292 -47841 85302 -47807
rect 85248 -47875 85302 -47841
rect 85248 -47909 85258 -47875
rect 85292 -47909 85302 -47875
rect 85248 -47995 85302 -47909
rect 85332 -47807 85386 -47795
rect 85332 -47841 85342 -47807
rect 85376 -47841 85386 -47807
rect 85332 -47875 85386 -47841
rect 85332 -47909 85342 -47875
rect 85376 -47909 85386 -47875
rect 85332 -47945 85386 -47909
rect 85332 -47979 85342 -47945
rect 85376 -47979 85386 -47945
rect 85332 -47995 85386 -47979
rect 85416 -47807 85468 -47795
rect 85416 -47841 85426 -47807
rect 85460 -47841 85468 -47807
rect 85416 -47875 85468 -47841
rect 85416 -47909 85426 -47875
rect 85460 -47909 85468 -47875
rect 85416 -47995 85468 -47909
rect 85546 -47807 85598 -47795
rect 85546 -47841 85554 -47807
rect 85588 -47841 85598 -47807
rect 85546 -47875 85598 -47841
rect 85546 -47909 85554 -47875
rect 85588 -47909 85598 -47875
rect 85546 -47945 85598 -47909
rect 85546 -47979 85554 -47945
rect 85588 -47979 85598 -47945
rect 85546 -47995 85598 -47979
rect 85628 -47807 85682 -47795
rect 85628 -47841 85638 -47807
rect 85672 -47841 85682 -47807
rect 85628 -47875 85682 -47841
rect 85628 -47909 85638 -47875
rect 85672 -47909 85682 -47875
rect 85628 -47945 85682 -47909
rect 85628 -47979 85638 -47945
rect 85672 -47979 85682 -47945
rect 85628 -47995 85682 -47979
rect 85712 -47807 85766 -47795
rect 85712 -47841 85722 -47807
rect 85756 -47841 85766 -47807
rect 85712 -47875 85766 -47841
rect 85712 -47909 85722 -47875
rect 85756 -47909 85766 -47875
rect 85712 -47995 85766 -47909
rect 85796 -47807 85850 -47795
rect 85796 -47841 85806 -47807
rect 85840 -47841 85850 -47807
rect 85796 -47875 85850 -47841
rect 85796 -47909 85806 -47875
rect 85840 -47909 85850 -47875
rect 85796 -47945 85850 -47909
rect 85796 -47979 85806 -47945
rect 85840 -47979 85850 -47945
rect 85796 -47995 85850 -47979
rect 85880 -47807 85934 -47795
rect 85880 -47841 85890 -47807
rect 85924 -47841 85934 -47807
rect 85880 -47875 85934 -47841
rect 85880 -47909 85890 -47875
rect 85924 -47909 85934 -47875
rect 85880 -47995 85934 -47909
rect 85964 -47807 86018 -47795
rect 85964 -47841 85974 -47807
rect 86008 -47841 86018 -47807
rect 85964 -47875 86018 -47841
rect 85964 -47909 85974 -47875
rect 86008 -47909 86018 -47875
rect 85964 -47945 86018 -47909
rect 85964 -47979 85974 -47945
rect 86008 -47979 86018 -47945
rect 85964 -47995 86018 -47979
rect 86048 -47807 86102 -47795
rect 86048 -47841 86058 -47807
rect 86092 -47841 86102 -47807
rect 86048 -47875 86102 -47841
rect 86048 -47909 86058 -47875
rect 86092 -47909 86102 -47875
rect 86048 -47995 86102 -47909
rect 86132 -47807 86186 -47795
rect 86132 -47841 86142 -47807
rect 86176 -47841 86186 -47807
rect 86132 -47875 86186 -47841
rect 86132 -47909 86142 -47875
rect 86176 -47909 86186 -47875
rect 86132 -47945 86186 -47909
rect 86132 -47979 86142 -47945
rect 86176 -47979 86186 -47945
rect 86132 -47995 86186 -47979
rect 86216 -47807 86270 -47795
rect 86216 -47841 86226 -47807
rect 86260 -47841 86270 -47807
rect 86216 -47875 86270 -47841
rect 86216 -47909 86226 -47875
rect 86260 -47909 86270 -47875
rect 86216 -47995 86270 -47909
rect 86300 -47807 86354 -47795
rect 86300 -47841 86310 -47807
rect 86344 -47841 86354 -47807
rect 86300 -47875 86354 -47841
rect 86300 -47909 86310 -47875
rect 86344 -47909 86354 -47875
rect 86300 -47945 86354 -47909
rect 86300 -47979 86310 -47945
rect 86344 -47979 86354 -47945
rect 86300 -47995 86354 -47979
rect 86384 -47807 86438 -47795
rect 86384 -47841 86394 -47807
rect 86428 -47841 86438 -47807
rect 86384 -47875 86438 -47841
rect 86384 -47909 86394 -47875
rect 86428 -47909 86438 -47875
rect 86384 -47995 86438 -47909
rect 86468 -47807 86522 -47795
rect 86468 -47841 86478 -47807
rect 86512 -47841 86522 -47807
rect 86468 -47875 86522 -47841
rect 86468 -47909 86478 -47875
rect 86512 -47909 86522 -47875
rect 86468 -47945 86522 -47909
rect 86468 -47979 86478 -47945
rect 86512 -47979 86522 -47945
rect 86468 -47995 86522 -47979
rect 86552 -47807 86606 -47795
rect 86552 -47841 86562 -47807
rect 86596 -47841 86606 -47807
rect 86552 -47875 86606 -47841
rect 86552 -47909 86562 -47875
rect 86596 -47909 86606 -47875
rect 86552 -47995 86606 -47909
rect 86636 -47807 86690 -47795
rect 86636 -47841 86646 -47807
rect 86680 -47841 86690 -47807
rect 86636 -47875 86690 -47841
rect 86636 -47909 86646 -47875
rect 86680 -47909 86690 -47875
rect 86636 -47945 86690 -47909
rect 86636 -47979 86646 -47945
rect 86680 -47979 86690 -47945
rect 86636 -47995 86690 -47979
rect 86720 -47807 86774 -47795
rect 86720 -47841 86730 -47807
rect 86764 -47841 86774 -47807
rect 86720 -47875 86774 -47841
rect 86720 -47909 86730 -47875
rect 86764 -47909 86774 -47875
rect 86720 -47995 86774 -47909
rect 86804 -47807 86858 -47795
rect 86804 -47841 86814 -47807
rect 86848 -47841 86858 -47807
rect 86804 -47875 86858 -47841
rect 86804 -47909 86814 -47875
rect 86848 -47909 86858 -47875
rect 86804 -47945 86858 -47909
rect 86804 -47979 86814 -47945
rect 86848 -47979 86858 -47945
rect 86804 -47995 86858 -47979
rect 86888 -47807 86940 -47795
rect 86888 -47841 86898 -47807
rect 86932 -47841 86940 -47807
rect 86888 -47875 86940 -47841
rect 86888 -47909 86898 -47875
rect 86932 -47909 86940 -47875
rect 86888 -47995 86940 -47909
rect 87018 -47807 87070 -47795
rect 87018 -47841 87026 -47807
rect 87060 -47841 87070 -47807
rect 87018 -47875 87070 -47841
rect 87018 -47909 87026 -47875
rect 87060 -47909 87070 -47875
rect 87018 -47945 87070 -47909
rect 87018 -47979 87026 -47945
rect 87060 -47979 87070 -47945
rect 87018 -47995 87070 -47979
rect 87100 -47807 87154 -47795
rect 87100 -47841 87110 -47807
rect 87144 -47841 87154 -47807
rect 87100 -47875 87154 -47841
rect 87100 -47909 87110 -47875
rect 87144 -47909 87154 -47875
rect 87100 -47945 87154 -47909
rect 87100 -47979 87110 -47945
rect 87144 -47979 87154 -47945
rect 87100 -47995 87154 -47979
rect 87184 -47807 87238 -47795
rect 87184 -47841 87194 -47807
rect 87228 -47841 87238 -47807
rect 87184 -47875 87238 -47841
rect 87184 -47909 87194 -47875
rect 87228 -47909 87238 -47875
rect 87184 -47995 87238 -47909
rect 87268 -47807 87322 -47795
rect 87268 -47841 87278 -47807
rect 87312 -47841 87322 -47807
rect 87268 -47875 87322 -47841
rect 87268 -47909 87278 -47875
rect 87312 -47909 87322 -47875
rect 87268 -47945 87322 -47909
rect 87268 -47979 87278 -47945
rect 87312 -47979 87322 -47945
rect 87268 -47995 87322 -47979
rect 87352 -47807 87406 -47795
rect 87352 -47841 87362 -47807
rect 87396 -47841 87406 -47807
rect 87352 -47875 87406 -47841
rect 87352 -47909 87362 -47875
rect 87396 -47909 87406 -47875
rect 87352 -47995 87406 -47909
rect 87436 -47807 87490 -47795
rect 87436 -47841 87446 -47807
rect 87480 -47841 87490 -47807
rect 87436 -47875 87490 -47841
rect 87436 -47909 87446 -47875
rect 87480 -47909 87490 -47875
rect 87436 -47945 87490 -47909
rect 87436 -47979 87446 -47945
rect 87480 -47979 87490 -47945
rect 87436 -47995 87490 -47979
rect 87520 -47807 87574 -47795
rect 87520 -47841 87530 -47807
rect 87564 -47841 87574 -47807
rect 87520 -47875 87574 -47841
rect 87520 -47909 87530 -47875
rect 87564 -47909 87574 -47875
rect 87520 -47995 87574 -47909
rect 87604 -47807 87658 -47795
rect 87604 -47841 87614 -47807
rect 87648 -47841 87658 -47807
rect 87604 -47875 87658 -47841
rect 87604 -47909 87614 -47875
rect 87648 -47909 87658 -47875
rect 87604 -47945 87658 -47909
rect 87604 -47979 87614 -47945
rect 87648 -47979 87658 -47945
rect 87604 -47995 87658 -47979
rect 87688 -47807 87742 -47795
rect 87688 -47841 87698 -47807
rect 87732 -47841 87742 -47807
rect 87688 -47875 87742 -47841
rect 87688 -47909 87698 -47875
rect 87732 -47909 87742 -47875
rect 87688 -47995 87742 -47909
rect 87772 -47807 87826 -47795
rect 87772 -47841 87782 -47807
rect 87816 -47841 87826 -47807
rect 87772 -47875 87826 -47841
rect 87772 -47909 87782 -47875
rect 87816 -47909 87826 -47875
rect 87772 -47945 87826 -47909
rect 87772 -47979 87782 -47945
rect 87816 -47979 87826 -47945
rect 87772 -47995 87826 -47979
rect 87856 -47807 87910 -47795
rect 87856 -47841 87866 -47807
rect 87900 -47841 87910 -47807
rect 87856 -47875 87910 -47841
rect 87856 -47909 87866 -47875
rect 87900 -47909 87910 -47875
rect 87856 -47995 87910 -47909
rect 87940 -47807 87994 -47795
rect 87940 -47841 87950 -47807
rect 87984 -47841 87994 -47807
rect 87940 -47875 87994 -47841
rect 87940 -47909 87950 -47875
rect 87984 -47909 87994 -47875
rect 87940 -47945 87994 -47909
rect 87940 -47979 87950 -47945
rect 87984 -47979 87994 -47945
rect 87940 -47995 87994 -47979
rect 88024 -47807 88078 -47795
rect 88024 -47841 88034 -47807
rect 88068 -47841 88078 -47807
rect 88024 -47875 88078 -47841
rect 88024 -47909 88034 -47875
rect 88068 -47909 88078 -47875
rect 88024 -47995 88078 -47909
rect 88108 -47807 88162 -47795
rect 88108 -47841 88118 -47807
rect 88152 -47841 88162 -47807
rect 88108 -47875 88162 -47841
rect 88108 -47909 88118 -47875
rect 88152 -47909 88162 -47875
rect 88108 -47945 88162 -47909
rect 88108 -47979 88118 -47945
rect 88152 -47979 88162 -47945
rect 88108 -47995 88162 -47979
rect 88192 -47807 88246 -47795
rect 88192 -47841 88202 -47807
rect 88236 -47841 88246 -47807
rect 88192 -47875 88246 -47841
rect 88192 -47909 88202 -47875
rect 88236 -47909 88246 -47875
rect 88192 -47995 88246 -47909
rect 88276 -47807 88330 -47795
rect 88276 -47841 88286 -47807
rect 88320 -47841 88330 -47807
rect 88276 -47875 88330 -47841
rect 88276 -47909 88286 -47875
rect 88320 -47909 88330 -47875
rect 88276 -47945 88330 -47909
rect 88276 -47979 88286 -47945
rect 88320 -47979 88330 -47945
rect 88276 -47995 88330 -47979
rect 88360 -47807 88412 -47795
rect 88360 -47841 88370 -47807
rect 88404 -47841 88412 -47807
rect 88360 -47875 88412 -47841
rect 88360 -47909 88370 -47875
rect 88404 -47909 88412 -47875
rect 88360 -47995 88412 -47909
rect 88490 -47807 88542 -47795
rect 88490 -47841 88498 -47807
rect 88532 -47841 88542 -47807
rect 88490 -47875 88542 -47841
rect 88490 -47909 88498 -47875
rect 88532 -47909 88542 -47875
rect 88490 -47945 88542 -47909
rect 88490 -47979 88498 -47945
rect 88532 -47979 88542 -47945
rect 88490 -47995 88542 -47979
rect 88572 -47807 88626 -47795
rect 88572 -47841 88582 -47807
rect 88616 -47841 88626 -47807
rect 88572 -47875 88626 -47841
rect 88572 -47909 88582 -47875
rect 88616 -47909 88626 -47875
rect 88572 -47945 88626 -47909
rect 88572 -47979 88582 -47945
rect 88616 -47979 88626 -47945
rect 88572 -47995 88626 -47979
rect 88656 -47807 88710 -47795
rect 88656 -47841 88666 -47807
rect 88700 -47841 88710 -47807
rect 88656 -47875 88710 -47841
rect 88656 -47909 88666 -47875
rect 88700 -47909 88710 -47875
rect 88656 -47995 88710 -47909
rect 88740 -47807 88794 -47795
rect 88740 -47841 88750 -47807
rect 88784 -47841 88794 -47807
rect 88740 -47875 88794 -47841
rect 88740 -47909 88750 -47875
rect 88784 -47909 88794 -47875
rect 88740 -47945 88794 -47909
rect 88740 -47979 88750 -47945
rect 88784 -47979 88794 -47945
rect 88740 -47995 88794 -47979
rect 88824 -47807 88878 -47795
rect 88824 -47841 88834 -47807
rect 88868 -47841 88878 -47807
rect 88824 -47875 88878 -47841
rect 88824 -47909 88834 -47875
rect 88868 -47909 88878 -47875
rect 88824 -47995 88878 -47909
rect 88908 -47807 88962 -47795
rect 88908 -47841 88918 -47807
rect 88952 -47841 88962 -47807
rect 88908 -47875 88962 -47841
rect 88908 -47909 88918 -47875
rect 88952 -47909 88962 -47875
rect 88908 -47945 88962 -47909
rect 88908 -47979 88918 -47945
rect 88952 -47979 88962 -47945
rect 88908 -47995 88962 -47979
rect 88992 -47807 89046 -47795
rect 88992 -47841 89002 -47807
rect 89036 -47841 89046 -47807
rect 88992 -47875 89046 -47841
rect 88992 -47909 89002 -47875
rect 89036 -47909 89046 -47875
rect 88992 -47995 89046 -47909
rect 89076 -47807 89130 -47795
rect 89076 -47841 89086 -47807
rect 89120 -47841 89130 -47807
rect 89076 -47875 89130 -47841
rect 89076 -47909 89086 -47875
rect 89120 -47909 89130 -47875
rect 89076 -47945 89130 -47909
rect 89076 -47979 89086 -47945
rect 89120 -47979 89130 -47945
rect 89076 -47995 89130 -47979
rect 89160 -47807 89214 -47795
rect 89160 -47841 89170 -47807
rect 89204 -47841 89214 -47807
rect 89160 -47875 89214 -47841
rect 89160 -47909 89170 -47875
rect 89204 -47909 89214 -47875
rect 89160 -47995 89214 -47909
rect 89244 -47807 89298 -47795
rect 89244 -47841 89254 -47807
rect 89288 -47841 89298 -47807
rect 89244 -47875 89298 -47841
rect 89244 -47909 89254 -47875
rect 89288 -47909 89298 -47875
rect 89244 -47945 89298 -47909
rect 89244 -47979 89254 -47945
rect 89288 -47979 89298 -47945
rect 89244 -47995 89298 -47979
rect 89328 -47807 89382 -47795
rect 89328 -47841 89338 -47807
rect 89372 -47841 89382 -47807
rect 89328 -47875 89382 -47841
rect 89328 -47909 89338 -47875
rect 89372 -47909 89382 -47875
rect 89328 -47995 89382 -47909
rect 89412 -47807 89466 -47795
rect 89412 -47841 89422 -47807
rect 89456 -47841 89466 -47807
rect 89412 -47875 89466 -47841
rect 89412 -47909 89422 -47875
rect 89456 -47909 89466 -47875
rect 89412 -47945 89466 -47909
rect 89412 -47979 89422 -47945
rect 89456 -47979 89466 -47945
rect 89412 -47995 89466 -47979
rect 89496 -47807 89550 -47795
rect 89496 -47841 89506 -47807
rect 89540 -47841 89550 -47807
rect 89496 -47875 89550 -47841
rect 89496 -47909 89506 -47875
rect 89540 -47909 89550 -47875
rect 89496 -47995 89550 -47909
rect 89580 -47807 89634 -47795
rect 89580 -47841 89590 -47807
rect 89624 -47841 89634 -47807
rect 89580 -47875 89634 -47841
rect 89580 -47909 89590 -47875
rect 89624 -47909 89634 -47875
rect 89580 -47945 89634 -47909
rect 89580 -47979 89590 -47945
rect 89624 -47979 89634 -47945
rect 89580 -47995 89634 -47979
rect 89664 -47807 89718 -47795
rect 89664 -47841 89674 -47807
rect 89708 -47841 89718 -47807
rect 89664 -47875 89718 -47841
rect 89664 -47909 89674 -47875
rect 89708 -47909 89718 -47875
rect 89664 -47995 89718 -47909
rect 89748 -47807 89802 -47795
rect 89748 -47841 89758 -47807
rect 89792 -47841 89802 -47807
rect 89748 -47875 89802 -47841
rect 89748 -47909 89758 -47875
rect 89792 -47909 89802 -47875
rect 89748 -47945 89802 -47909
rect 89748 -47979 89758 -47945
rect 89792 -47979 89802 -47945
rect 89748 -47995 89802 -47979
rect 89832 -47807 89884 -47795
rect 89832 -47841 89842 -47807
rect 89876 -47841 89884 -47807
rect 89832 -47875 89884 -47841
rect 89832 -47909 89842 -47875
rect 89876 -47909 89884 -47875
rect 89832 -47995 89884 -47909
rect 89962 -47807 90014 -47795
rect 89962 -47841 89970 -47807
rect 90004 -47841 90014 -47807
rect 89962 -47875 90014 -47841
rect 89962 -47909 89970 -47875
rect 90004 -47909 90014 -47875
rect 89962 -47945 90014 -47909
rect 89962 -47979 89970 -47945
rect 90004 -47979 90014 -47945
rect 89962 -47995 90014 -47979
rect 90044 -47807 90098 -47795
rect 90044 -47841 90054 -47807
rect 90088 -47841 90098 -47807
rect 90044 -47875 90098 -47841
rect 90044 -47909 90054 -47875
rect 90088 -47909 90098 -47875
rect 90044 -47945 90098 -47909
rect 90044 -47979 90054 -47945
rect 90088 -47979 90098 -47945
rect 90044 -47995 90098 -47979
rect 90128 -47807 90182 -47795
rect 90128 -47841 90138 -47807
rect 90172 -47841 90182 -47807
rect 90128 -47875 90182 -47841
rect 90128 -47909 90138 -47875
rect 90172 -47909 90182 -47875
rect 90128 -47995 90182 -47909
rect 90212 -47807 90266 -47795
rect 90212 -47841 90222 -47807
rect 90256 -47841 90266 -47807
rect 90212 -47875 90266 -47841
rect 90212 -47909 90222 -47875
rect 90256 -47909 90266 -47875
rect 90212 -47945 90266 -47909
rect 90212 -47979 90222 -47945
rect 90256 -47979 90266 -47945
rect 90212 -47995 90266 -47979
rect 90296 -47807 90350 -47795
rect 90296 -47841 90306 -47807
rect 90340 -47841 90350 -47807
rect 90296 -47875 90350 -47841
rect 90296 -47909 90306 -47875
rect 90340 -47909 90350 -47875
rect 90296 -47995 90350 -47909
rect 90380 -47807 90434 -47795
rect 90380 -47841 90390 -47807
rect 90424 -47841 90434 -47807
rect 90380 -47875 90434 -47841
rect 90380 -47909 90390 -47875
rect 90424 -47909 90434 -47875
rect 90380 -47945 90434 -47909
rect 90380 -47979 90390 -47945
rect 90424 -47979 90434 -47945
rect 90380 -47995 90434 -47979
rect 90464 -47807 90518 -47795
rect 90464 -47841 90474 -47807
rect 90508 -47841 90518 -47807
rect 90464 -47875 90518 -47841
rect 90464 -47909 90474 -47875
rect 90508 -47909 90518 -47875
rect 90464 -47995 90518 -47909
rect 90548 -47807 90602 -47795
rect 90548 -47841 90558 -47807
rect 90592 -47841 90602 -47807
rect 90548 -47875 90602 -47841
rect 90548 -47909 90558 -47875
rect 90592 -47909 90602 -47875
rect 90548 -47945 90602 -47909
rect 90548 -47979 90558 -47945
rect 90592 -47979 90602 -47945
rect 90548 -47995 90602 -47979
rect 90632 -47807 90686 -47795
rect 90632 -47841 90642 -47807
rect 90676 -47841 90686 -47807
rect 90632 -47875 90686 -47841
rect 90632 -47909 90642 -47875
rect 90676 -47909 90686 -47875
rect 90632 -47995 90686 -47909
rect 90716 -47807 90770 -47795
rect 90716 -47841 90726 -47807
rect 90760 -47841 90770 -47807
rect 90716 -47875 90770 -47841
rect 90716 -47909 90726 -47875
rect 90760 -47909 90770 -47875
rect 90716 -47945 90770 -47909
rect 90716 -47979 90726 -47945
rect 90760 -47979 90770 -47945
rect 90716 -47995 90770 -47979
rect 90800 -47807 90854 -47795
rect 90800 -47841 90810 -47807
rect 90844 -47841 90854 -47807
rect 90800 -47875 90854 -47841
rect 90800 -47909 90810 -47875
rect 90844 -47909 90854 -47875
rect 90800 -47995 90854 -47909
rect 90884 -47807 90938 -47795
rect 90884 -47841 90894 -47807
rect 90928 -47841 90938 -47807
rect 90884 -47875 90938 -47841
rect 90884 -47909 90894 -47875
rect 90928 -47909 90938 -47875
rect 90884 -47945 90938 -47909
rect 90884 -47979 90894 -47945
rect 90928 -47979 90938 -47945
rect 90884 -47995 90938 -47979
rect 90968 -47807 91022 -47795
rect 90968 -47841 90978 -47807
rect 91012 -47841 91022 -47807
rect 90968 -47875 91022 -47841
rect 90968 -47909 90978 -47875
rect 91012 -47909 91022 -47875
rect 90968 -47995 91022 -47909
rect 91052 -47807 91106 -47795
rect 91052 -47841 91062 -47807
rect 91096 -47841 91106 -47807
rect 91052 -47875 91106 -47841
rect 91052 -47909 91062 -47875
rect 91096 -47909 91106 -47875
rect 91052 -47945 91106 -47909
rect 91052 -47979 91062 -47945
rect 91096 -47979 91106 -47945
rect 91052 -47995 91106 -47979
rect 91136 -47807 91190 -47795
rect 91136 -47841 91146 -47807
rect 91180 -47841 91190 -47807
rect 91136 -47875 91190 -47841
rect 91136 -47909 91146 -47875
rect 91180 -47909 91190 -47875
rect 91136 -47995 91190 -47909
rect 91220 -47807 91274 -47795
rect 91220 -47841 91230 -47807
rect 91264 -47841 91274 -47807
rect 91220 -47875 91274 -47841
rect 91220 -47909 91230 -47875
rect 91264 -47909 91274 -47875
rect 91220 -47945 91274 -47909
rect 91220 -47979 91230 -47945
rect 91264 -47979 91274 -47945
rect 91220 -47995 91274 -47979
rect 91304 -47807 91356 -47795
rect 91304 -47841 91314 -47807
rect 91348 -47841 91356 -47807
rect 91304 -47875 91356 -47841
rect 91304 -47909 91314 -47875
rect 91348 -47909 91356 -47875
rect 91304 -47995 91356 -47909
rect 77605 -48048 77657 -48025
rect 77605 -48082 77613 -48048
rect 77647 -48082 77657 -48048
rect 77605 -48109 77657 -48082
rect 77687 -48109 77753 -48025
rect 77783 -48109 77825 -48025
rect 77855 -48109 77921 -48025
rect 77951 -48109 78019 -48025
rect 77966 -48111 78019 -48109
rect 77966 -48145 77974 -48111
rect 78008 -48145 78019 -48111
rect 77966 -48179 78019 -48145
rect 77966 -48213 77974 -48179
rect 78008 -48213 78019 -48179
rect 77966 -48225 78019 -48213
rect 78049 -48080 78103 -48025
rect 78049 -48114 78059 -48080
rect 78093 -48114 78103 -48080
rect 78049 -48148 78103 -48114
rect 78049 -48182 78059 -48148
rect 78093 -48182 78103 -48148
rect 78049 -48225 78103 -48182
rect 77833 -48407 77885 -48395
rect 77833 -48437 77841 -48407
rect 77637 -48449 77693 -48437
rect 77637 -48483 77649 -48449
rect 77683 -48483 77693 -48449
rect 77637 -48521 77693 -48483
rect 77723 -48449 77777 -48437
rect 77723 -48483 77733 -48449
rect 77767 -48483 77777 -48449
rect 77723 -48521 77777 -48483
rect 77807 -48441 77841 -48437
rect 77875 -48441 77885 -48407
rect 77807 -48475 77885 -48441
rect 77807 -48509 77841 -48475
rect 77875 -48509 77885 -48475
rect 77807 -48521 77885 -48509
rect 77823 -48595 77885 -48521
rect 77915 -48407 78010 -48395
rect 77915 -48441 77945 -48407
rect 77979 -48441 78010 -48407
rect 77915 -48475 78010 -48441
rect 77915 -48509 77945 -48475
rect 77979 -48509 78010 -48475
rect 77915 -48595 78010 -48509
rect 77823 -49339 77885 -49265
rect 77637 -49377 77693 -49339
rect 77637 -49411 77649 -49377
rect 77683 -49411 77693 -49377
rect 77637 -49423 77693 -49411
rect 77723 -49377 77777 -49339
rect 77723 -49411 77733 -49377
rect 77767 -49411 77777 -49377
rect 77723 -49423 77777 -49411
rect 77807 -49351 77885 -49339
rect 77807 -49385 77841 -49351
rect 77875 -49385 77885 -49351
rect 77807 -49419 77885 -49385
rect 77807 -49423 77841 -49419
rect 77833 -49453 77841 -49423
rect 77875 -49453 77885 -49419
rect 77833 -49465 77885 -49453
rect 77915 -49351 78010 -49265
rect 78065 -49288 78117 -49265
rect 78065 -49322 78073 -49288
rect 78107 -49322 78117 -49288
rect 78065 -49349 78117 -49322
rect 78147 -49349 78213 -49265
rect 78243 -49349 78285 -49265
rect 78315 -49349 78381 -49265
rect 78411 -49349 78479 -49265
rect 77915 -49385 77945 -49351
rect 77979 -49385 78010 -49351
rect 77915 -49419 78010 -49385
rect 78426 -49351 78479 -49349
rect 78426 -49385 78434 -49351
rect 78468 -49385 78479 -49351
rect 77915 -49453 77945 -49419
rect 77979 -49453 78010 -49419
rect 78426 -49419 78479 -49385
rect 77915 -49465 78010 -49453
rect 78426 -49453 78434 -49419
rect 78468 -49453 78479 -49419
rect 78426 -49465 78479 -49453
rect 78509 -49320 78563 -49265
rect 78509 -49354 78519 -49320
rect 78553 -49354 78563 -49320
rect 78509 -49388 78563 -49354
rect 78509 -49422 78519 -49388
rect 78553 -49422 78563 -49388
rect 78509 -49465 78563 -49422
rect 77833 -49647 77885 -49635
rect 77833 -49677 77841 -49647
rect 77637 -49689 77693 -49677
rect 77637 -49723 77649 -49689
rect 77683 -49723 77693 -49689
rect 77637 -49761 77693 -49723
rect 77723 -49689 77777 -49677
rect 77723 -49723 77733 -49689
rect 77767 -49723 77777 -49689
rect 77723 -49761 77777 -49723
rect 77807 -49681 77841 -49677
rect 77875 -49681 77885 -49647
rect 77807 -49715 77885 -49681
rect 77807 -49749 77841 -49715
rect 77875 -49749 77885 -49715
rect 77807 -49761 77885 -49749
rect 77823 -49835 77885 -49761
rect 77915 -49647 78010 -49635
rect 77915 -49681 77945 -49647
rect 77979 -49681 78010 -49647
rect 77915 -49715 78010 -49681
rect 77915 -49749 77945 -49715
rect 77979 -49749 78010 -49715
rect 77915 -49835 78010 -49749
rect 54079 -50272 54879 -50260
rect 54079 -50306 54091 -50272
rect 54867 -50306 54879 -50272
rect 54079 -50318 54879 -50306
rect 54079 -50400 54879 -50388
rect 54079 -50434 54091 -50400
rect 54867 -50434 54879 -50400
rect 54079 -50446 54879 -50434
rect 54079 -50628 54879 -50616
rect 54079 -50662 54091 -50628
rect 54867 -50662 54879 -50628
rect 54079 -50674 54879 -50662
rect 54079 -50756 54879 -50744
rect 54079 -50790 54091 -50756
rect 54867 -50790 54879 -50756
rect 54079 -50802 54879 -50790
rect 57123 -50729 57175 -50709
rect 57123 -50763 57131 -50729
rect 57165 -50763 57175 -50729
rect 57123 -50797 57175 -50763
rect 57123 -50831 57131 -50797
rect 57165 -50831 57175 -50797
rect 57123 -50867 57175 -50831
rect 57205 -50729 57263 -50709
rect 57205 -50763 57217 -50729
rect 57251 -50763 57263 -50729
rect 57205 -50797 57263 -50763
rect 57205 -50831 57217 -50797
rect 57251 -50831 57263 -50797
rect 57205 -50867 57263 -50831
rect 57293 -50729 57345 -50709
rect 57293 -50763 57303 -50729
rect 57337 -50763 57345 -50729
rect 57293 -50810 57345 -50763
rect 57293 -50844 57303 -50810
rect 57337 -50844 57345 -50810
rect 57293 -50867 57345 -50844
rect 77825 -50593 77887 -50519
rect 59113 -50647 59513 -50635
rect 59113 -50681 59125 -50647
rect 59501 -50681 59513 -50647
rect 59113 -50693 59513 -50681
rect 59113 -50755 59513 -50743
rect 59113 -50789 59125 -50755
rect 59501 -50789 59513 -50755
rect 59113 -50801 59513 -50789
rect 59113 -50863 59513 -50851
rect 59113 -50897 59125 -50863
rect 59501 -50897 59513 -50863
rect 59113 -50909 59513 -50897
rect 77639 -50631 77695 -50593
rect 77639 -50665 77651 -50631
rect 77685 -50665 77695 -50631
rect 77639 -50677 77695 -50665
rect 77725 -50631 77779 -50593
rect 77725 -50665 77735 -50631
rect 77769 -50665 77779 -50631
rect 77725 -50677 77779 -50665
rect 77809 -50605 77887 -50593
rect 77809 -50639 77843 -50605
rect 77877 -50639 77887 -50605
rect 77809 -50673 77887 -50639
rect 77809 -50677 77843 -50673
rect 77835 -50707 77843 -50677
rect 77877 -50707 77887 -50673
rect 77835 -50719 77887 -50707
rect 77917 -50605 78012 -50519
rect 77917 -50639 77947 -50605
rect 77981 -50639 78012 -50605
rect 77917 -50673 78012 -50639
rect 77917 -50707 77947 -50673
rect 77981 -50707 78012 -50673
rect 77917 -50719 78012 -50707
rect 54069 -52588 54869 -52576
rect 54069 -52622 54081 -52588
rect 54857 -52622 54869 -52588
rect 54069 -52634 54869 -52622
rect 54069 -52716 54869 -52704
rect 54069 -52750 54081 -52716
rect 54857 -52750 54869 -52716
rect 54069 -52762 54869 -52750
rect 56418 -51299 56476 -51287
rect 56418 -52075 56430 -51299
rect 56464 -52075 56476 -51299
rect 56418 -52087 56476 -52075
rect 56546 -51299 56604 -51287
rect 56546 -52075 56558 -51299
rect 56592 -52075 56604 -51299
rect 56546 -52087 56604 -52075
rect 59032 -51171 59090 -51159
rect 59032 -51547 59044 -51171
rect 59078 -51547 59090 -51171
rect 59032 -51559 59090 -51547
rect 59150 -51171 59208 -51159
rect 59150 -51547 59162 -51171
rect 59196 -51547 59208 -51171
rect 59150 -51559 59208 -51547
rect 77605 -50897 77657 -50885
rect 77605 -50931 77613 -50897
rect 77647 -50931 77657 -50897
rect 77605 -50969 77657 -50931
rect 77687 -50905 77757 -50885
rect 77687 -50939 77705 -50905
rect 77739 -50939 77757 -50905
rect 77687 -50969 77757 -50939
rect 77787 -50897 77861 -50885
rect 77787 -50931 77807 -50897
rect 77841 -50931 77861 -50897
rect 77787 -50969 77861 -50931
rect 77891 -50905 77947 -50885
rect 77891 -50939 77902 -50905
rect 77936 -50939 77947 -50905
rect 77891 -50969 77947 -50939
rect 77977 -50897 78113 -50885
rect 77977 -50931 78053 -50897
rect 78087 -50931 78113 -50897
rect 77977 -50965 78113 -50931
rect 77977 -50969 78053 -50965
rect 77996 -50999 78053 -50969
rect 78087 -50999 78113 -50965
rect 77996 -51085 78113 -50999
rect 78143 -50897 78195 -50885
rect 78143 -50931 78153 -50897
rect 78187 -50931 78195 -50897
rect 78710 -50897 78763 -50885
rect 78143 -50965 78195 -50931
rect 78710 -50931 78718 -50897
rect 78752 -50931 78763 -50897
rect 78143 -50999 78153 -50965
rect 78187 -50999 78195 -50965
rect 78143 -51033 78195 -50999
rect 78710 -50965 78763 -50931
rect 78710 -50999 78718 -50965
rect 78752 -50999 78763 -50965
rect 78710 -51001 78763 -50999
rect 78143 -51067 78153 -51033
rect 78187 -51067 78195 -51033
rect 78143 -51085 78195 -51067
rect 78349 -51028 78401 -51001
rect 78349 -51062 78357 -51028
rect 78391 -51062 78401 -51028
rect 78349 -51085 78401 -51062
rect 78431 -51085 78497 -51001
rect 78527 -51085 78569 -51001
rect 78599 -51085 78665 -51001
rect 78695 -51085 78763 -51001
rect 78793 -50928 78847 -50885
rect 78793 -50962 78803 -50928
rect 78837 -50962 78847 -50928
rect 78793 -50996 78847 -50962
rect 78793 -51030 78803 -50996
rect 78837 -51030 78847 -50996
rect 78793 -51085 78847 -51030
rect 83075 -51473 83127 -51445
rect 60441 -51573 60641 -51565
rect 60441 -51607 60459 -51573
rect 60493 -51607 60527 -51573
rect 60561 -51607 60595 -51573
rect 60629 -51607 60641 -51573
rect 60441 -51617 60641 -51607
rect 60811 -51573 61011 -51565
rect 60811 -51607 60823 -51573
rect 60857 -51607 60891 -51573
rect 60925 -51607 60959 -51573
rect 60993 -51607 61011 -51573
rect 60811 -51617 61011 -51607
rect 60441 -51657 60641 -51647
rect 60441 -51691 60459 -51657
rect 60493 -51691 60527 -51657
rect 60561 -51691 60595 -51657
rect 60629 -51691 60641 -51657
rect 60441 -51701 60641 -51691
rect 60811 -51657 61011 -51647
rect 60811 -51691 60823 -51657
rect 60857 -51691 60891 -51657
rect 60925 -51691 60959 -51657
rect 60993 -51691 61011 -51657
rect 60811 -51701 61011 -51691
rect 59032 -51901 59090 -51889
rect 59032 -52277 59044 -51901
rect 59078 -52277 59090 -51901
rect 59032 -52289 59090 -52277
rect 59150 -51901 59208 -51889
rect 59150 -52277 59162 -51901
rect 59196 -52277 59208 -51901
rect 59150 -52289 59208 -52277
rect 83075 -51507 83083 -51473
rect 83117 -51507 83127 -51473
rect 83075 -51541 83127 -51507
rect 83075 -51561 83083 -51541
rect 82906 -51593 82958 -51561
rect 82906 -51627 82914 -51593
rect 82948 -51627 82958 -51593
rect 82906 -51645 82958 -51627
rect 82988 -51645 83030 -51561
rect 83060 -51575 83083 -51561
rect 83117 -51575 83127 -51541
rect 83060 -51645 83127 -51575
rect 83157 -51457 83225 -51445
rect 83157 -51491 83183 -51457
rect 83217 -51491 83225 -51457
rect 83157 -51525 83225 -51491
rect 83157 -51559 83183 -51525
rect 83217 -51559 83225 -51525
rect 83157 -51645 83225 -51559
rect 83366 -51457 83418 -51445
rect 83366 -51491 83374 -51457
rect 83408 -51491 83418 -51457
rect 83366 -51525 83418 -51491
rect 83366 -51559 83374 -51525
rect 83408 -51559 83418 -51525
rect 83366 -51593 83418 -51559
rect 83366 -51627 83374 -51593
rect 83408 -51627 83418 -51593
rect 83366 -51645 83418 -51627
rect 83448 -51457 83500 -51445
rect 83448 -51491 83458 -51457
rect 83492 -51491 83500 -51457
rect 83448 -51525 83500 -51491
rect 83448 -51559 83458 -51525
rect 83492 -51559 83500 -51525
rect 83448 -51593 83500 -51559
rect 83448 -51627 83458 -51593
rect 83492 -51627 83500 -51593
rect 83448 -51645 83500 -51627
rect 83611 -51457 83663 -51445
rect 83611 -51491 83619 -51457
rect 83653 -51491 83663 -51457
rect 83611 -51525 83663 -51491
rect 83611 -51559 83619 -51525
rect 83653 -51559 83663 -51525
rect 83611 -51593 83663 -51559
rect 83611 -51627 83619 -51593
rect 83653 -51627 83663 -51593
rect 83611 -51645 83663 -51627
rect 83693 -51457 83747 -51445
rect 83693 -51491 83703 -51457
rect 83737 -51491 83747 -51457
rect 83693 -51525 83747 -51491
rect 83693 -51559 83703 -51525
rect 83737 -51559 83747 -51525
rect 83693 -51593 83747 -51559
rect 83693 -51627 83703 -51593
rect 83737 -51627 83747 -51593
rect 83693 -51645 83747 -51627
rect 83777 -51457 83831 -51445
rect 83777 -51491 83787 -51457
rect 83821 -51491 83831 -51457
rect 83777 -51525 83831 -51491
rect 83777 -51559 83787 -51525
rect 83821 -51559 83831 -51525
rect 83777 -51645 83831 -51559
rect 83861 -51457 83915 -51445
rect 83861 -51491 83871 -51457
rect 83905 -51491 83915 -51457
rect 83861 -51525 83915 -51491
rect 83861 -51559 83871 -51525
rect 83905 -51559 83915 -51525
rect 83861 -51593 83915 -51559
rect 83861 -51627 83871 -51593
rect 83905 -51627 83915 -51593
rect 83861 -51645 83915 -51627
rect 83945 -51457 83997 -51445
rect 83945 -51491 83955 -51457
rect 83989 -51491 83997 -51457
rect 83945 -51645 83997 -51491
rect 84074 -51457 84126 -51445
rect 84074 -51491 84082 -51457
rect 84116 -51491 84126 -51457
rect 84074 -51525 84126 -51491
rect 84074 -51559 84082 -51525
rect 84116 -51559 84126 -51525
rect 84074 -51595 84126 -51559
rect 84074 -51629 84082 -51595
rect 84116 -51629 84126 -51595
rect 84074 -51645 84126 -51629
rect 84156 -51457 84210 -51445
rect 84156 -51491 84166 -51457
rect 84200 -51491 84210 -51457
rect 84156 -51525 84210 -51491
rect 84156 -51559 84166 -51525
rect 84200 -51559 84210 -51525
rect 84156 -51595 84210 -51559
rect 84156 -51629 84166 -51595
rect 84200 -51629 84210 -51595
rect 84156 -51645 84210 -51629
rect 84240 -51457 84294 -51445
rect 84240 -51491 84250 -51457
rect 84284 -51491 84294 -51457
rect 84240 -51525 84294 -51491
rect 84240 -51559 84250 -51525
rect 84284 -51559 84294 -51525
rect 84240 -51645 84294 -51559
rect 84324 -51457 84378 -51445
rect 84324 -51491 84334 -51457
rect 84368 -51491 84378 -51457
rect 84324 -51525 84378 -51491
rect 84324 -51559 84334 -51525
rect 84368 -51559 84378 -51525
rect 84324 -51595 84378 -51559
rect 84324 -51629 84334 -51595
rect 84368 -51629 84378 -51595
rect 84324 -51645 84378 -51629
rect 84408 -51457 84462 -51445
rect 84408 -51491 84418 -51457
rect 84452 -51491 84462 -51457
rect 84408 -51525 84462 -51491
rect 84408 -51559 84418 -51525
rect 84452 -51559 84462 -51525
rect 84408 -51645 84462 -51559
rect 84492 -51457 84546 -51445
rect 84492 -51491 84502 -51457
rect 84536 -51491 84546 -51457
rect 84492 -51525 84546 -51491
rect 84492 -51559 84502 -51525
rect 84536 -51559 84546 -51525
rect 84492 -51595 84546 -51559
rect 84492 -51629 84502 -51595
rect 84536 -51629 84546 -51595
rect 84492 -51645 84546 -51629
rect 84576 -51457 84630 -51445
rect 84576 -51491 84586 -51457
rect 84620 -51491 84630 -51457
rect 84576 -51525 84630 -51491
rect 84576 -51559 84586 -51525
rect 84620 -51559 84630 -51525
rect 84576 -51645 84630 -51559
rect 84660 -51457 84714 -51445
rect 84660 -51491 84670 -51457
rect 84704 -51491 84714 -51457
rect 84660 -51525 84714 -51491
rect 84660 -51559 84670 -51525
rect 84704 -51559 84714 -51525
rect 84660 -51595 84714 -51559
rect 84660 -51629 84670 -51595
rect 84704 -51629 84714 -51595
rect 84660 -51645 84714 -51629
rect 84744 -51457 84798 -51445
rect 84744 -51491 84754 -51457
rect 84788 -51491 84798 -51457
rect 84744 -51525 84798 -51491
rect 84744 -51559 84754 -51525
rect 84788 -51559 84798 -51525
rect 84744 -51645 84798 -51559
rect 84828 -51457 84882 -51445
rect 84828 -51491 84838 -51457
rect 84872 -51491 84882 -51457
rect 84828 -51525 84882 -51491
rect 84828 -51559 84838 -51525
rect 84872 -51559 84882 -51525
rect 84828 -51595 84882 -51559
rect 84828 -51629 84838 -51595
rect 84872 -51629 84882 -51595
rect 84828 -51645 84882 -51629
rect 84912 -51457 84966 -51445
rect 84912 -51491 84922 -51457
rect 84956 -51491 84966 -51457
rect 84912 -51525 84966 -51491
rect 84912 -51559 84922 -51525
rect 84956 -51559 84966 -51525
rect 84912 -51645 84966 -51559
rect 84996 -51457 85050 -51445
rect 84996 -51491 85006 -51457
rect 85040 -51491 85050 -51457
rect 84996 -51525 85050 -51491
rect 84996 -51559 85006 -51525
rect 85040 -51559 85050 -51525
rect 84996 -51595 85050 -51559
rect 84996 -51629 85006 -51595
rect 85040 -51629 85050 -51595
rect 84996 -51645 85050 -51629
rect 85080 -51457 85134 -51445
rect 85080 -51491 85090 -51457
rect 85124 -51491 85134 -51457
rect 85080 -51525 85134 -51491
rect 85080 -51559 85090 -51525
rect 85124 -51559 85134 -51525
rect 85080 -51645 85134 -51559
rect 85164 -51457 85218 -51445
rect 85164 -51491 85174 -51457
rect 85208 -51491 85218 -51457
rect 85164 -51525 85218 -51491
rect 85164 -51559 85174 -51525
rect 85208 -51559 85218 -51525
rect 85164 -51595 85218 -51559
rect 85164 -51629 85174 -51595
rect 85208 -51629 85218 -51595
rect 85164 -51645 85218 -51629
rect 85248 -51457 85302 -51445
rect 85248 -51491 85258 -51457
rect 85292 -51491 85302 -51457
rect 85248 -51525 85302 -51491
rect 85248 -51559 85258 -51525
rect 85292 -51559 85302 -51525
rect 85248 -51645 85302 -51559
rect 85332 -51457 85386 -51445
rect 85332 -51491 85342 -51457
rect 85376 -51491 85386 -51457
rect 85332 -51525 85386 -51491
rect 85332 -51559 85342 -51525
rect 85376 -51559 85386 -51525
rect 85332 -51595 85386 -51559
rect 85332 -51629 85342 -51595
rect 85376 -51629 85386 -51595
rect 85332 -51645 85386 -51629
rect 85416 -51457 85468 -51445
rect 85416 -51491 85426 -51457
rect 85460 -51491 85468 -51457
rect 85416 -51525 85468 -51491
rect 85416 -51559 85426 -51525
rect 85460 -51559 85468 -51525
rect 85416 -51645 85468 -51559
rect 85546 -51457 85598 -51445
rect 85546 -51491 85554 -51457
rect 85588 -51491 85598 -51457
rect 85546 -51525 85598 -51491
rect 85546 -51559 85554 -51525
rect 85588 -51559 85598 -51525
rect 85546 -51595 85598 -51559
rect 85546 -51629 85554 -51595
rect 85588 -51629 85598 -51595
rect 85546 -51645 85598 -51629
rect 85628 -51457 85682 -51445
rect 85628 -51491 85638 -51457
rect 85672 -51491 85682 -51457
rect 85628 -51525 85682 -51491
rect 85628 -51559 85638 -51525
rect 85672 -51559 85682 -51525
rect 85628 -51595 85682 -51559
rect 85628 -51629 85638 -51595
rect 85672 -51629 85682 -51595
rect 85628 -51645 85682 -51629
rect 85712 -51457 85766 -51445
rect 85712 -51491 85722 -51457
rect 85756 -51491 85766 -51457
rect 85712 -51525 85766 -51491
rect 85712 -51559 85722 -51525
rect 85756 -51559 85766 -51525
rect 85712 -51645 85766 -51559
rect 85796 -51457 85850 -51445
rect 85796 -51491 85806 -51457
rect 85840 -51491 85850 -51457
rect 85796 -51525 85850 -51491
rect 85796 -51559 85806 -51525
rect 85840 -51559 85850 -51525
rect 85796 -51595 85850 -51559
rect 85796 -51629 85806 -51595
rect 85840 -51629 85850 -51595
rect 85796 -51645 85850 -51629
rect 85880 -51457 85934 -51445
rect 85880 -51491 85890 -51457
rect 85924 -51491 85934 -51457
rect 85880 -51525 85934 -51491
rect 85880 -51559 85890 -51525
rect 85924 -51559 85934 -51525
rect 85880 -51645 85934 -51559
rect 85964 -51457 86018 -51445
rect 85964 -51491 85974 -51457
rect 86008 -51491 86018 -51457
rect 85964 -51525 86018 -51491
rect 85964 -51559 85974 -51525
rect 86008 -51559 86018 -51525
rect 85964 -51595 86018 -51559
rect 85964 -51629 85974 -51595
rect 86008 -51629 86018 -51595
rect 85964 -51645 86018 -51629
rect 86048 -51457 86102 -51445
rect 86048 -51491 86058 -51457
rect 86092 -51491 86102 -51457
rect 86048 -51525 86102 -51491
rect 86048 -51559 86058 -51525
rect 86092 -51559 86102 -51525
rect 86048 -51645 86102 -51559
rect 86132 -51457 86186 -51445
rect 86132 -51491 86142 -51457
rect 86176 -51491 86186 -51457
rect 86132 -51525 86186 -51491
rect 86132 -51559 86142 -51525
rect 86176 -51559 86186 -51525
rect 86132 -51595 86186 -51559
rect 86132 -51629 86142 -51595
rect 86176 -51629 86186 -51595
rect 86132 -51645 86186 -51629
rect 86216 -51457 86270 -51445
rect 86216 -51491 86226 -51457
rect 86260 -51491 86270 -51457
rect 86216 -51525 86270 -51491
rect 86216 -51559 86226 -51525
rect 86260 -51559 86270 -51525
rect 86216 -51645 86270 -51559
rect 86300 -51457 86354 -51445
rect 86300 -51491 86310 -51457
rect 86344 -51491 86354 -51457
rect 86300 -51525 86354 -51491
rect 86300 -51559 86310 -51525
rect 86344 -51559 86354 -51525
rect 86300 -51595 86354 -51559
rect 86300 -51629 86310 -51595
rect 86344 -51629 86354 -51595
rect 86300 -51645 86354 -51629
rect 86384 -51457 86438 -51445
rect 86384 -51491 86394 -51457
rect 86428 -51491 86438 -51457
rect 86384 -51525 86438 -51491
rect 86384 -51559 86394 -51525
rect 86428 -51559 86438 -51525
rect 86384 -51645 86438 -51559
rect 86468 -51457 86522 -51445
rect 86468 -51491 86478 -51457
rect 86512 -51491 86522 -51457
rect 86468 -51525 86522 -51491
rect 86468 -51559 86478 -51525
rect 86512 -51559 86522 -51525
rect 86468 -51595 86522 -51559
rect 86468 -51629 86478 -51595
rect 86512 -51629 86522 -51595
rect 86468 -51645 86522 -51629
rect 86552 -51457 86606 -51445
rect 86552 -51491 86562 -51457
rect 86596 -51491 86606 -51457
rect 86552 -51525 86606 -51491
rect 86552 -51559 86562 -51525
rect 86596 -51559 86606 -51525
rect 86552 -51645 86606 -51559
rect 86636 -51457 86690 -51445
rect 86636 -51491 86646 -51457
rect 86680 -51491 86690 -51457
rect 86636 -51525 86690 -51491
rect 86636 -51559 86646 -51525
rect 86680 -51559 86690 -51525
rect 86636 -51595 86690 -51559
rect 86636 -51629 86646 -51595
rect 86680 -51629 86690 -51595
rect 86636 -51645 86690 -51629
rect 86720 -51457 86774 -51445
rect 86720 -51491 86730 -51457
rect 86764 -51491 86774 -51457
rect 86720 -51525 86774 -51491
rect 86720 -51559 86730 -51525
rect 86764 -51559 86774 -51525
rect 86720 -51645 86774 -51559
rect 86804 -51457 86858 -51445
rect 86804 -51491 86814 -51457
rect 86848 -51491 86858 -51457
rect 86804 -51525 86858 -51491
rect 86804 -51559 86814 -51525
rect 86848 -51559 86858 -51525
rect 86804 -51595 86858 -51559
rect 86804 -51629 86814 -51595
rect 86848 -51629 86858 -51595
rect 86804 -51645 86858 -51629
rect 86888 -51457 86940 -51445
rect 86888 -51491 86898 -51457
rect 86932 -51491 86940 -51457
rect 86888 -51525 86940 -51491
rect 86888 -51559 86898 -51525
rect 86932 -51559 86940 -51525
rect 86888 -51645 86940 -51559
rect 87018 -51457 87070 -51445
rect 87018 -51491 87026 -51457
rect 87060 -51491 87070 -51457
rect 87018 -51525 87070 -51491
rect 87018 -51559 87026 -51525
rect 87060 -51559 87070 -51525
rect 87018 -51595 87070 -51559
rect 87018 -51629 87026 -51595
rect 87060 -51629 87070 -51595
rect 87018 -51645 87070 -51629
rect 87100 -51457 87154 -51445
rect 87100 -51491 87110 -51457
rect 87144 -51491 87154 -51457
rect 87100 -51525 87154 -51491
rect 87100 -51559 87110 -51525
rect 87144 -51559 87154 -51525
rect 87100 -51595 87154 -51559
rect 87100 -51629 87110 -51595
rect 87144 -51629 87154 -51595
rect 87100 -51645 87154 -51629
rect 87184 -51457 87238 -51445
rect 87184 -51491 87194 -51457
rect 87228 -51491 87238 -51457
rect 87184 -51525 87238 -51491
rect 87184 -51559 87194 -51525
rect 87228 -51559 87238 -51525
rect 87184 -51645 87238 -51559
rect 87268 -51457 87322 -51445
rect 87268 -51491 87278 -51457
rect 87312 -51491 87322 -51457
rect 87268 -51525 87322 -51491
rect 87268 -51559 87278 -51525
rect 87312 -51559 87322 -51525
rect 87268 -51595 87322 -51559
rect 87268 -51629 87278 -51595
rect 87312 -51629 87322 -51595
rect 87268 -51645 87322 -51629
rect 87352 -51457 87406 -51445
rect 87352 -51491 87362 -51457
rect 87396 -51491 87406 -51457
rect 87352 -51525 87406 -51491
rect 87352 -51559 87362 -51525
rect 87396 -51559 87406 -51525
rect 87352 -51645 87406 -51559
rect 87436 -51457 87490 -51445
rect 87436 -51491 87446 -51457
rect 87480 -51491 87490 -51457
rect 87436 -51525 87490 -51491
rect 87436 -51559 87446 -51525
rect 87480 -51559 87490 -51525
rect 87436 -51595 87490 -51559
rect 87436 -51629 87446 -51595
rect 87480 -51629 87490 -51595
rect 87436 -51645 87490 -51629
rect 87520 -51457 87574 -51445
rect 87520 -51491 87530 -51457
rect 87564 -51491 87574 -51457
rect 87520 -51525 87574 -51491
rect 87520 -51559 87530 -51525
rect 87564 -51559 87574 -51525
rect 87520 -51645 87574 -51559
rect 87604 -51457 87658 -51445
rect 87604 -51491 87614 -51457
rect 87648 -51491 87658 -51457
rect 87604 -51525 87658 -51491
rect 87604 -51559 87614 -51525
rect 87648 -51559 87658 -51525
rect 87604 -51595 87658 -51559
rect 87604 -51629 87614 -51595
rect 87648 -51629 87658 -51595
rect 87604 -51645 87658 -51629
rect 87688 -51457 87742 -51445
rect 87688 -51491 87698 -51457
rect 87732 -51491 87742 -51457
rect 87688 -51525 87742 -51491
rect 87688 -51559 87698 -51525
rect 87732 -51559 87742 -51525
rect 87688 -51645 87742 -51559
rect 87772 -51457 87826 -51445
rect 87772 -51491 87782 -51457
rect 87816 -51491 87826 -51457
rect 87772 -51525 87826 -51491
rect 87772 -51559 87782 -51525
rect 87816 -51559 87826 -51525
rect 87772 -51595 87826 -51559
rect 87772 -51629 87782 -51595
rect 87816 -51629 87826 -51595
rect 87772 -51645 87826 -51629
rect 87856 -51457 87910 -51445
rect 87856 -51491 87866 -51457
rect 87900 -51491 87910 -51457
rect 87856 -51525 87910 -51491
rect 87856 -51559 87866 -51525
rect 87900 -51559 87910 -51525
rect 87856 -51645 87910 -51559
rect 87940 -51457 87994 -51445
rect 87940 -51491 87950 -51457
rect 87984 -51491 87994 -51457
rect 87940 -51525 87994 -51491
rect 87940 -51559 87950 -51525
rect 87984 -51559 87994 -51525
rect 87940 -51595 87994 -51559
rect 87940 -51629 87950 -51595
rect 87984 -51629 87994 -51595
rect 87940 -51645 87994 -51629
rect 88024 -51457 88078 -51445
rect 88024 -51491 88034 -51457
rect 88068 -51491 88078 -51457
rect 88024 -51525 88078 -51491
rect 88024 -51559 88034 -51525
rect 88068 -51559 88078 -51525
rect 88024 -51645 88078 -51559
rect 88108 -51457 88162 -51445
rect 88108 -51491 88118 -51457
rect 88152 -51491 88162 -51457
rect 88108 -51525 88162 -51491
rect 88108 -51559 88118 -51525
rect 88152 -51559 88162 -51525
rect 88108 -51595 88162 -51559
rect 88108 -51629 88118 -51595
rect 88152 -51629 88162 -51595
rect 88108 -51645 88162 -51629
rect 88192 -51457 88246 -51445
rect 88192 -51491 88202 -51457
rect 88236 -51491 88246 -51457
rect 88192 -51525 88246 -51491
rect 88192 -51559 88202 -51525
rect 88236 -51559 88246 -51525
rect 88192 -51645 88246 -51559
rect 88276 -51457 88330 -51445
rect 88276 -51491 88286 -51457
rect 88320 -51491 88330 -51457
rect 88276 -51525 88330 -51491
rect 88276 -51559 88286 -51525
rect 88320 -51559 88330 -51525
rect 88276 -51595 88330 -51559
rect 88276 -51629 88286 -51595
rect 88320 -51629 88330 -51595
rect 88276 -51645 88330 -51629
rect 88360 -51457 88412 -51445
rect 88360 -51491 88370 -51457
rect 88404 -51491 88412 -51457
rect 88360 -51525 88412 -51491
rect 88360 -51559 88370 -51525
rect 88404 -51559 88412 -51525
rect 88360 -51645 88412 -51559
rect 88490 -51457 88542 -51445
rect 88490 -51491 88498 -51457
rect 88532 -51491 88542 -51457
rect 88490 -51525 88542 -51491
rect 88490 -51559 88498 -51525
rect 88532 -51559 88542 -51525
rect 88490 -51595 88542 -51559
rect 88490 -51629 88498 -51595
rect 88532 -51629 88542 -51595
rect 88490 -51645 88542 -51629
rect 88572 -51457 88626 -51445
rect 88572 -51491 88582 -51457
rect 88616 -51491 88626 -51457
rect 88572 -51525 88626 -51491
rect 88572 -51559 88582 -51525
rect 88616 -51559 88626 -51525
rect 88572 -51595 88626 -51559
rect 88572 -51629 88582 -51595
rect 88616 -51629 88626 -51595
rect 88572 -51645 88626 -51629
rect 88656 -51457 88710 -51445
rect 88656 -51491 88666 -51457
rect 88700 -51491 88710 -51457
rect 88656 -51525 88710 -51491
rect 88656 -51559 88666 -51525
rect 88700 -51559 88710 -51525
rect 88656 -51645 88710 -51559
rect 88740 -51457 88794 -51445
rect 88740 -51491 88750 -51457
rect 88784 -51491 88794 -51457
rect 88740 -51525 88794 -51491
rect 88740 -51559 88750 -51525
rect 88784 -51559 88794 -51525
rect 88740 -51595 88794 -51559
rect 88740 -51629 88750 -51595
rect 88784 -51629 88794 -51595
rect 88740 -51645 88794 -51629
rect 88824 -51457 88878 -51445
rect 88824 -51491 88834 -51457
rect 88868 -51491 88878 -51457
rect 88824 -51525 88878 -51491
rect 88824 -51559 88834 -51525
rect 88868 -51559 88878 -51525
rect 88824 -51645 88878 -51559
rect 88908 -51457 88962 -51445
rect 88908 -51491 88918 -51457
rect 88952 -51491 88962 -51457
rect 88908 -51525 88962 -51491
rect 88908 -51559 88918 -51525
rect 88952 -51559 88962 -51525
rect 88908 -51595 88962 -51559
rect 88908 -51629 88918 -51595
rect 88952 -51629 88962 -51595
rect 88908 -51645 88962 -51629
rect 88992 -51457 89046 -51445
rect 88992 -51491 89002 -51457
rect 89036 -51491 89046 -51457
rect 88992 -51525 89046 -51491
rect 88992 -51559 89002 -51525
rect 89036 -51559 89046 -51525
rect 88992 -51645 89046 -51559
rect 89076 -51457 89130 -51445
rect 89076 -51491 89086 -51457
rect 89120 -51491 89130 -51457
rect 89076 -51525 89130 -51491
rect 89076 -51559 89086 -51525
rect 89120 -51559 89130 -51525
rect 89076 -51595 89130 -51559
rect 89076 -51629 89086 -51595
rect 89120 -51629 89130 -51595
rect 89076 -51645 89130 -51629
rect 89160 -51457 89214 -51445
rect 89160 -51491 89170 -51457
rect 89204 -51491 89214 -51457
rect 89160 -51525 89214 -51491
rect 89160 -51559 89170 -51525
rect 89204 -51559 89214 -51525
rect 89160 -51645 89214 -51559
rect 89244 -51457 89298 -51445
rect 89244 -51491 89254 -51457
rect 89288 -51491 89298 -51457
rect 89244 -51525 89298 -51491
rect 89244 -51559 89254 -51525
rect 89288 -51559 89298 -51525
rect 89244 -51595 89298 -51559
rect 89244 -51629 89254 -51595
rect 89288 -51629 89298 -51595
rect 89244 -51645 89298 -51629
rect 89328 -51457 89382 -51445
rect 89328 -51491 89338 -51457
rect 89372 -51491 89382 -51457
rect 89328 -51525 89382 -51491
rect 89328 -51559 89338 -51525
rect 89372 -51559 89382 -51525
rect 89328 -51645 89382 -51559
rect 89412 -51457 89466 -51445
rect 89412 -51491 89422 -51457
rect 89456 -51491 89466 -51457
rect 89412 -51525 89466 -51491
rect 89412 -51559 89422 -51525
rect 89456 -51559 89466 -51525
rect 89412 -51595 89466 -51559
rect 89412 -51629 89422 -51595
rect 89456 -51629 89466 -51595
rect 89412 -51645 89466 -51629
rect 89496 -51457 89550 -51445
rect 89496 -51491 89506 -51457
rect 89540 -51491 89550 -51457
rect 89496 -51525 89550 -51491
rect 89496 -51559 89506 -51525
rect 89540 -51559 89550 -51525
rect 89496 -51645 89550 -51559
rect 89580 -51457 89634 -51445
rect 89580 -51491 89590 -51457
rect 89624 -51491 89634 -51457
rect 89580 -51525 89634 -51491
rect 89580 -51559 89590 -51525
rect 89624 -51559 89634 -51525
rect 89580 -51595 89634 -51559
rect 89580 -51629 89590 -51595
rect 89624 -51629 89634 -51595
rect 89580 -51645 89634 -51629
rect 89664 -51457 89718 -51445
rect 89664 -51491 89674 -51457
rect 89708 -51491 89718 -51457
rect 89664 -51525 89718 -51491
rect 89664 -51559 89674 -51525
rect 89708 -51559 89718 -51525
rect 89664 -51645 89718 -51559
rect 89748 -51457 89802 -51445
rect 89748 -51491 89758 -51457
rect 89792 -51491 89802 -51457
rect 89748 -51525 89802 -51491
rect 89748 -51559 89758 -51525
rect 89792 -51559 89802 -51525
rect 89748 -51595 89802 -51559
rect 89748 -51629 89758 -51595
rect 89792 -51629 89802 -51595
rect 89748 -51645 89802 -51629
rect 89832 -51457 89884 -51445
rect 89832 -51491 89842 -51457
rect 89876 -51491 89884 -51457
rect 89832 -51525 89884 -51491
rect 89832 -51559 89842 -51525
rect 89876 -51559 89884 -51525
rect 89832 -51645 89884 -51559
rect 89962 -51457 90014 -51445
rect 89962 -51491 89970 -51457
rect 90004 -51491 90014 -51457
rect 89962 -51525 90014 -51491
rect 89962 -51559 89970 -51525
rect 90004 -51559 90014 -51525
rect 89962 -51595 90014 -51559
rect 89962 -51629 89970 -51595
rect 90004 -51629 90014 -51595
rect 89962 -51645 90014 -51629
rect 90044 -51457 90098 -51445
rect 90044 -51491 90054 -51457
rect 90088 -51491 90098 -51457
rect 90044 -51525 90098 -51491
rect 90044 -51559 90054 -51525
rect 90088 -51559 90098 -51525
rect 90044 -51595 90098 -51559
rect 90044 -51629 90054 -51595
rect 90088 -51629 90098 -51595
rect 90044 -51645 90098 -51629
rect 90128 -51457 90182 -51445
rect 90128 -51491 90138 -51457
rect 90172 -51491 90182 -51457
rect 90128 -51525 90182 -51491
rect 90128 -51559 90138 -51525
rect 90172 -51559 90182 -51525
rect 90128 -51645 90182 -51559
rect 90212 -51457 90266 -51445
rect 90212 -51491 90222 -51457
rect 90256 -51491 90266 -51457
rect 90212 -51525 90266 -51491
rect 90212 -51559 90222 -51525
rect 90256 -51559 90266 -51525
rect 90212 -51595 90266 -51559
rect 90212 -51629 90222 -51595
rect 90256 -51629 90266 -51595
rect 90212 -51645 90266 -51629
rect 90296 -51457 90350 -51445
rect 90296 -51491 90306 -51457
rect 90340 -51491 90350 -51457
rect 90296 -51525 90350 -51491
rect 90296 -51559 90306 -51525
rect 90340 -51559 90350 -51525
rect 90296 -51645 90350 -51559
rect 90380 -51457 90434 -51445
rect 90380 -51491 90390 -51457
rect 90424 -51491 90434 -51457
rect 90380 -51525 90434 -51491
rect 90380 -51559 90390 -51525
rect 90424 -51559 90434 -51525
rect 90380 -51595 90434 -51559
rect 90380 -51629 90390 -51595
rect 90424 -51629 90434 -51595
rect 90380 -51645 90434 -51629
rect 90464 -51457 90518 -51445
rect 90464 -51491 90474 -51457
rect 90508 -51491 90518 -51457
rect 90464 -51525 90518 -51491
rect 90464 -51559 90474 -51525
rect 90508 -51559 90518 -51525
rect 90464 -51645 90518 -51559
rect 90548 -51457 90602 -51445
rect 90548 -51491 90558 -51457
rect 90592 -51491 90602 -51457
rect 90548 -51525 90602 -51491
rect 90548 -51559 90558 -51525
rect 90592 -51559 90602 -51525
rect 90548 -51595 90602 -51559
rect 90548 -51629 90558 -51595
rect 90592 -51629 90602 -51595
rect 90548 -51645 90602 -51629
rect 90632 -51457 90686 -51445
rect 90632 -51491 90642 -51457
rect 90676 -51491 90686 -51457
rect 90632 -51525 90686 -51491
rect 90632 -51559 90642 -51525
rect 90676 -51559 90686 -51525
rect 90632 -51645 90686 -51559
rect 90716 -51457 90770 -51445
rect 90716 -51491 90726 -51457
rect 90760 -51491 90770 -51457
rect 90716 -51525 90770 -51491
rect 90716 -51559 90726 -51525
rect 90760 -51559 90770 -51525
rect 90716 -51595 90770 -51559
rect 90716 -51629 90726 -51595
rect 90760 -51629 90770 -51595
rect 90716 -51645 90770 -51629
rect 90800 -51457 90854 -51445
rect 90800 -51491 90810 -51457
rect 90844 -51491 90854 -51457
rect 90800 -51525 90854 -51491
rect 90800 -51559 90810 -51525
rect 90844 -51559 90854 -51525
rect 90800 -51645 90854 -51559
rect 90884 -51457 90938 -51445
rect 90884 -51491 90894 -51457
rect 90928 -51491 90938 -51457
rect 90884 -51525 90938 -51491
rect 90884 -51559 90894 -51525
rect 90928 -51559 90938 -51525
rect 90884 -51595 90938 -51559
rect 90884 -51629 90894 -51595
rect 90928 -51629 90938 -51595
rect 90884 -51645 90938 -51629
rect 90968 -51457 91022 -51445
rect 90968 -51491 90978 -51457
rect 91012 -51491 91022 -51457
rect 90968 -51525 91022 -51491
rect 90968 -51559 90978 -51525
rect 91012 -51559 91022 -51525
rect 90968 -51645 91022 -51559
rect 91052 -51457 91106 -51445
rect 91052 -51491 91062 -51457
rect 91096 -51491 91106 -51457
rect 91052 -51525 91106 -51491
rect 91052 -51559 91062 -51525
rect 91096 -51559 91106 -51525
rect 91052 -51595 91106 -51559
rect 91052 -51629 91062 -51595
rect 91096 -51629 91106 -51595
rect 91052 -51645 91106 -51629
rect 91136 -51457 91190 -51445
rect 91136 -51491 91146 -51457
rect 91180 -51491 91190 -51457
rect 91136 -51525 91190 -51491
rect 91136 -51559 91146 -51525
rect 91180 -51559 91190 -51525
rect 91136 -51645 91190 -51559
rect 91220 -51457 91274 -51445
rect 91220 -51491 91230 -51457
rect 91264 -51491 91274 -51457
rect 91220 -51525 91274 -51491
rect 91220 -51559 91230 -51525
rect 91264 -51559 91274 -51525
rect 91220 -51595 91274 -51559
rect 91220 -51629 91230 -51595
rect 91264 -51629 91274 -51595
rect 91220 -51645 91274 -51629
rect 91304 -51457 91356 -51445
rect 91304 -51491 91314 -51457
rect 91348 -51491 91356 -51457
rect 91304 -51525 91356 -51491
rect 91304 -51559 91314 -51525
rect 91348 -51559 91356 -51525
rect 91304 -51645 91356 -51559
rect 60441 -51741 60641 -51731
rect 60441 -51775 60527 -51741
rect 60561 -51775 60595 -51741
rect 60629 -51775 60641 -51741
rect 60441 -51785 60641 -51775
rect 60811 -51741 61011 -51731
rect 60811 -51775 60823 -51741
rect 60857 -51775 60891 -51741
rect 60925 -51775 61011 -51741
rect 60811 -51785 61011 -51775
rect 60441 -51825 60641 -51815
rect 60441 -51859 60459 -51825
rect 60493 -51859 60527 -51825
rect 60561 -51859 60595 -51825
rect 60629 -51859 60641 -51825
rect 60441 -51869 60641 -51859
rect 60811 -51825 61011 -51815
rect 60811 -51859 60823 -51825
rect 60857 -51859 60891 -51825
rect 60925 -51859 60959 -51825
rect 60993 -51859 61011 -51825
rect 60811 -51869 61011 -51859
rect 77996 -51837 78113 -51751
rect 77996 -51867 78053 -51837
rect 60441 -51909 60641 -51899
rect 60441 -51943 60595 -51909
rect 60629 -51943 60641 -51909
rect 60441 -51951 60641 -51943
rect 60811 -51909 61011 -51899
rect 60811 -51943 60823 -51909
rect 60857 -51943 61011 -51909
rect 60811 -51951 61011 -51943
rect 77605 -51905 77657 -51867
rect 77605 -51939 77613 -51905
rect 77647 -51939 77657 -51905
rect 77605 -51951 77657 -51939
rect 77687 -51897 77757 -51867
rect 77687 -51931 77705 -51897
rect 77739 -51931 77757 -51897
rect 77687 -51951 77757 -51931
rect 77787 -51905 77861 -51867
rect 77787 -51939 77807 -51905
rect 77841 -51939 77861 -51905
rect 77787 -51951 77861 -51939
rect 77891 -51897 77947 -51867
rect 77891 -51931 77902 -51897
rect 77936 -51931 77947 -51897
rect 77891 -51951 77947 -51931
rect 77977 -51871 78053 -51867
rect 78087 -51871 78113 -51837
rect 77977 -51905 78113 -51871
rect 77977 -51939 78053 -51905
rect 78087 -51939 78113 -51905
rect 77977 -51951 78113 -51939
rect 78143 -51769 78195 -51751
rect 78143 -51803 78153 -51769
rect 78187 -51803 78195 -51769
rect 78143 -51837 78195 -51803
rect 78143 -51871 78153 -51837
rect 78187 -51871 78195 -51837
rect 78143 -51905 78195 -51871
rect 78143 -51939 78153 -51905
rect 78187 -51939 78195 -51905
rect 78143 -51951 78195 -51939
rect 77605 -52129 77657 -52117
rect 77605 -52163 77613 -52129
rect 77647 -52163 77657 -52129
rect 77605 -52201 77657 -52163
rect 77687 -52137 77757 -52117
rect 77687 -52171 77705 -52137
rect 77739 -52171 77757 -52137
rect 77687 -52201 77757 -52171
rect 77787 -52129 77861 -52117
rect 77787 -52163 77807 -52129
rect 77841 -52163 77861 -52129
rect 77787 -52201 77861 -52163
rect 77891 -52137 77947 -52117
rect 77891 -52171 77902 -52137
rect 77936 -52171 77947 -52137
rect 77891 -52201 77947 -52171
rect 77977 -52129 78113 -52117
rect 77977 -52163 78053 -52129
rect 78087 -52163 78113 -52129
rect 77977 -52197 78113 -52163
rect 77977 -52201 78053 -52197
rect 57123 -52557 57175 -52521
rect 57123 -52591 57131 -52557
rect 57165 -52591 57175 -52557
rect 57123 -52625 57175 -52591
rect 57123 -52659 57131 -52625
rect 57165 -52659 57175 -52625
rect 57123 -52679 57175 -52659
rect 57205 -52557 57263 -52521
rect 57205 -52591 57217 -52557
rect 57251 -52591 57263 -52557
rect 57205 -52625 57263 -52591
rect 57205 -52659 57217 -52625
rect 57251 -52659 57263 -52625
rect 57205 -52679 57263 -52659
rect 57293 -52544 57345 -52521
rect 57293 -52578 57303 -52544
rect 57337 -52578 57345 -52544
rect 57293 -52625 57345 -52578
rect 57293 -52659 57303 -52625
rect 57337 -52659 57345 -52625
rect 57293 -52679 57345 -52659
rect 59113 -52554 59513 -52542
rect 59113 -52588 59125 -52554
rect 59501 -52588 59513 -52554
rect 59113 -52600 59513 -52588
rect 59113 -52662 59513 -52650
rect 59113 -52696 59125 -52662
rect 59501 -52696 59513 -52662
rect 59113 -52708 59513 -52696
rect 59113 -52770 59513 -52758
rect 59113 -52804 59125 -52770
rect 59501 -52804 59513 -52770
rect 59113 -52816 59513 -52804
rect 54069 -52944 54869 -52932
rect 54069 -52978 54081 -52944
rect 54857 -52978 54869 -52944
rect 54069 -52990 54869 -52978
rect 54069 -53072 54869 -53060
rect 54069 -53106 54081 -53072
rect 54857 -53106 54869 -53072
rect 54069 -53118 54869 -53106
rect 77996 -52231 78053 -52201
rect 78087 -52231 78113 -52197
rect 77996 -52317 78113 -52231
rect 78143 -52129 78195 -52117
rect 78143 -52163 78153 -52129
rect 78187 -52163 78195 -52129
rect 78143 -52197 78195 -52163
rect 78143 -52231 78153 -52197
rect 78187 -52231 78195 -52197
rect 78143 -52265 78195 -52231
rect 78143 -52299 78153 -52265
rect 78187 -52299 78195 -52265
rect 78143 -52317 78195 -52299
rect 77996 -53071 78113 -52985
rect 77996 -53101 78053 -53071
rect 77605 -53139 77657 -53101
rect 77605 -53173 77613 -53139
rect 77647 -53173 77657 -53139
rect 77605 -53185 77657 -53173
rect 77687 -53131 77757 -53101
rect 77687 -53165 77705 -53131
rect 77739 -53165 77757 -53131
rect 77687 -53185 77757 -53165
rect 77787 -53139 77861 -53101
rect 77787 -53173 77807 -53139
rect 77841 -53173 77861 -53139
rect 77787 -53185 77861 -53173
rect 77891 -53131 77947 -53101
rect 77891 -53165 77902 -53131
rect 77936 -53165 77947 -53131
rect 77891 -53185 77947 -53165
rect 77977 -53105 78053 -53101
rect 78087 -53105 78113 -53071
rect 77977 -53139 78113 -53105
rect 77977 -53173 78053 -53139
rect 78087 -53173 78113 -53139
rect 77977 -53185 78113 -53173
rect 78143 -53003 78195 -52985
rect 78143 -53037 78153 -53003
rect 78187 -53037 78195 -53003
rect 78143 -53071 78195 -53037
rect 78143 -53105 78153 -53071
rect 78187 -53105 78195 -53071
rect 78143 -53139 78195 -53105
rect 78143 -53173 78153 -53139
rect 78187 -53173 78195 -53139
rect 78143 -53185 78195 -53173
rect 77877 -53367 77929 -53355
rect 77877 -53401 77885 -53367
rect 77919 -53401 77929 -53367
rect 77877 -53414 77929 -53401
rect 77879 -53468 77929 -53414
rect 77605 -53506 77657 -53468
rect 77605 -53540 77613 -53506
rect 77647 -53540 77657 -53506
rect 77605 -53552 77657 -53540
rect 77687 -53476 77741 -53468
rect 77687 -53510 77697 -53476
rect 77731 -53510 77741 -53476
rect 77687 -53552 77741 -53510
rect 77771 -53495 77834 -53468
rect 77771 -53529 77790 -53495
rect 77824 -53529 77834 -53495
rect 77771 -53552 77834 -53529
rect 77864 -53552 77929 -53468
rect 77879 -53555 77929 -53552
rect 77959 -53381 78011 -53355
rect 78293 -53367 78345 -53355
rect 77959 -53415 77969 -53381
rect 78003 -53415 78011 -53381
rect 78293 -53397 78301 -53367
rect 77959 -53449 78011 -53415
rect 77959 -53483 77969 -53449
rect 78003 -53483 78011 -53449
rect 78097 -53409 78153 -53397
rect 78097 -53443 78109 -53409
rect 78143 -53443 78153 -53409
rect 78097 -53481 78153 -53443
rect 78183 -53409 78237 -53397
rect 78183 -53443 78193 -53409
rect 78227 -53443 78237 -53409
rect 78183 -53481 78237 -53443
rect 78267 -53401 78301 -53397
rect 78335 -53401 78345 -53367
rect 78267 -53435 78345 -53401
rect 78267 -53469 78301 -53435
rect 78335 -53469 78345 -53435
rect 78267 -53481 78345 -53469
rect 77959 -53555 78011 -53483
rect 78283 -53555 78345 -53481
rect 78375 -53367 78470 -53355
rect 78375 -53401 78405 -53367
rect 78439 -53401 78470 -53367
rect 78886 -53367 78939 -53355
rect 78375 -53435 78470 -53401
rect 78886 -53401 78894 -53367
rect 78928 -53401 78939 -53367
rect 78375 -53469 78405 -53435
rect 78439 -53469 78470 -53435
rect 78375 -53555 78470 -53469
rect 78886 -53435 78939 -53401
rect 78886 -53469 78894 -53435
rect 78928 -53469 78939 -53435
rect 78886 -53471 78939 -53469
rect 78525 -53498 78577 -53471
rect 78525 -53532 78533 -53498
rect 78567 -53532 78577 -53498
rect 78525 -53555 78577 -53532
rect 78607 -53555 78673 -53471
rect 78703 -53555 78745 -53471
rect 78775 -53555 78841 -53471
rect 78871 -53555 78939 -53471
rect 78969 -53398 79023 -53355
rect 78969 -53432 78979 -53398
rect 79013 -53432 79023 -53398
rect 78969 -53466 79023 -53432
rect 78969 -53500 78979 -53466
rect 79013 -53500 79023 -53466
rect 78969 -53555 79023 -53500
rect 54079 -55672 54879 -55660
rect 54079 -55706 54091 -55672
rect 54867 -55706 54879 -55672
rect 54079 -55718 54879 -55706
rect 54079 -55800 54879 -55788
rect 54079 -55834 54091 -55800
rect 54867 -55834 54879 -55800
rect 54079 -55846 54879 -55834
rect 54079 -56028 54879 -56016
rect 54079 -56062 54091 -56028
rect 54867 -56062 54879 -56028
rect 54079 -56074 54879 -56062
rect 54079 -56156 54879 -56144
rect 54079 -56190 54091 -56156
rect 54867 -56190 54879 -56156
rect 54079 -56202 54879 -56190
rect 57123 -56129 57175 -56109
rect 57123 -56163 57131 -56129
rect 57165 -56163 57175 -56129
rect 57123 -56197 57175 -56163
rect 57123 -56231 57131 -56197
rect 57165 -56231 57175 -56197
rect 57123 -56267 57175 -56231
rect 57205 -56129 57263 -56109
rect 57205 -56163 57217 -56129
rect 57251 -56163 57263 -56129
rect 57205 -56197 57263 -56163
rect 57205 -56231 57217 -56197
rect 57251 -56231 57263 -56197
rect 57205 -56267 57263 -56231
rect 57293 -56129 57345 -56109
rect 57293 -56163 57303 -56129
rect 57337 -56163 57345 -56129
rect 57293 -56210 57345 -56163
rect 57293 -56244 57303 -56210
rect 57337 -56244 57345 -56210
rect 57293 -56267 57345 -56244
rect 59113 -56047 59513 -56035
rect 59113 -56081 59125 -56047
rect 59501 -56081 59513 -56047
rect 59113 -56093 59513 -56081
rect 59113 -56155 59513 -56143
rect 59113 -56189 59125 -56155
rect 59501 -56189 59513 -56155
rect 59113 -56201 59513 -56189
rect 59113 -56263 59513 -56251
rect 59113 -56297 59125 -56263
rect 59501 -56297 59513 -56263
rect 59113 -56309 59513 -56297
rect 54069 -57988 54869 -57976
rect 54069 -58022 54081 -57988
rect 54857 -58022 54869 -57988
rect 54069 -58034 54869 -58022
rect 54069 -58116 54869 -58104
rect 54069 -58150 54081 -58116
rect 54857 -58150 54869 -58116
rect 54069 -58162 54869 -58150
rect 56418 -56699 56476 -56687
rect 56418 -57475 56430 -56699
rect 56464 -57475 56476 -56699
rect 56418 -57487 56476 -57475
rect 56546 -56699 56604 -56687
rect 56546 -57475 56558 -56699
rect 56592 -57475 56604 -56699
rect 56546 -57487 56604 -57475
rect 59032 -56571 59090 -56559
rect 59032 -56947 59044 -56571
rect 59078 -56947 59090 -56571
rect 59032 -56959 59090 -56947
rect 59150 -56571 59208 -56559
rect 59150 -56947 59162 -56571
rect 59196 -56947 59208 -56571
rect 59150 -56959 59208 -56947
rect 60441 -56973 60641 -56965
rect 60441 -57007 60459 -56973
rect 60493 -57007 60527 -56973
rect 60561 -57007 60595 -56973
rect 60629 -57007 60641 -56973
rect 60441 -57017 60641 -57007
rect 60811 -56973 61011 -56965
rect 60811 -57007 60823 -56973
rect 60857 -57007 60891 -56973
rect 60925 -57007 60959 -56973
rect 60993 -57007 61011 -56973
rect 60811 -57017 61011 -57007
rect 60441 -57057 60641 -57047
rect 60441 -57091 60459 -57057
rect 60493 -57091 60527 -57057
rect 60561 -57091 60595 -57057
rect 60629 -57091 60641 -57057
rect 60441 -57101 60641 -57091
rect 60811 -57057 61011 -57047
rect 60811 -57091 60823 -57057
rect 60857 -57091 60891 -57057
rect 60925 -57091 60959 -57057
rect 60993 -57091 61011 -57057
rect 60811 -57101 61011 -57091
rect 59032 -57301 59090 -57289
rect 59032 -57677 59044 -57301
rect 59078 -57677 59090 -57301
rect 59032 -57689 59090 -57677
rect 59150 -57301 59208 -57289
rect 59150 -57677 59162 -57301
rect 59196 -57677 59208 -57301
rect 59150 -57689 59208 -57677
rect 60441 -57141 60641 -57131
rect 60441 -57175 60527 -57141
rect 60561 -57175 60595 -57141
rect 60629 -57175 60641 -57141
rect 60441 -57185 60641 -57175
rect 60811 -57141 61011 -57131
rect 60811 -57175 60823 -57141
rect 60857 -57175 60891 -57141
rect 60925 -57175 61011 -57141
rect 60811 -57185 61011 -57175
rect 60441 -57225 60641 -57215
rect 60441 -57259 60459 -57225
rect 60493 -57259 60527 -57225
rect 60561 -57259 60595 -57225
rect 60629 -57259 60641 -57225
rect 60441 -57269 60641 -57259
rect 60811 -57225 61011 -57215
rect 60811 -57259 60823 -57225
rect 60857 -57259 60891 -57225
rect 60925 -57259 60959 -57225
rect 60993 -57259 61011 -57225
rect 60811 -57269 61011 -57259
rect 60441 -57309 60641 -57299
rect 60441 -57343 60595 -57309
rect 60629 -57343 60641 -57309
rect 60441 -57351 60641 -57343
rect 60811 -57309 61011 -57299
rect 60811 -57343 60823 -57309
rect 60857 -57343 61011 -57309
rect 60811 -57351 61011 -57343
rect 57123 -57957 57175 -57921
rect 57123 -57991 57131 -57957
rect 57165 -57991 57175 -57957
rect 57123 -58025 57175 -57991
rect 57123 -58059 57131 -58025
rect 57165 -58059 57175 -58025
rect 57123 -58079 57175 -58059
rect 57205 -57957 57263 -57921
rect 57205 -57991 57217 -57957
rect 57251 -57991 57263 -57957
rect 57205 -58025 57263 -57991
rect 57205 -58059 57217 -58025
rect 57251 -58059 57263 -58025
rect 57205 -58079 57263 -58059
rect 57293 -57944 57345 -57921
rect 57293 -57978 57303 -57944
rect 57337 -57978 57345 -57944
rect 57293 -58025 57345 -57978
rect 57293 -58059 57303 -58025
rect 57337 -58059 57345 -58025
rect 57293 -58079 57345 -58059
rect 59113 -57954 59513 -57942
rect 59113 -57988 59125 -57954
rect 59501 -57988 59513 -57954
rect 59113 -58000 59513 -57988
rect 59113 -58062 59513 -58050
rect 59113 -58096 59125 -58062
rect 59501 -58096 59513 -58062
rect 59113 -58108 59513 -58096
rect 59113 -58170 59513 -58158
rect 59113 -58204 59125 -58170
rect 59501 -58204 59513 -58170
rect 59113 -58216 59513 -58204
rect 54069 -58344 54869 -58332
rect 54069 -58378 54081 -58344
rect 54857 -58378 54869 -58344
rect 54069 -58390 54869 -58378
rect 54069 -58472 54869 -58460
rect 54069 -58506 54081 -58472
rect 54857 -58506 54869 -58472
rect 54069 -58518 54869 -58506
rect 54079 -61072 54879 -61060
rect 54079 -61106 54091 -61072
rect 54867 -61106 54879 -61072
rect 54079 -61118 54879 -61106
rect 54079 -61200 54879 -61188
rect 54079 -61234 54091 -61200
rect 54867 -61234 54879 -61200
rect 54079 -61246 54879 -61234
rect 54079 -61428 54879 -61416
rect 54079 -61462 54091 -61428
rect 54867 -61462 54879 -61428
rect 54079 -61474 54879 -61462
rect 54079 -61556 54879 -61544
rect 54079 -61590 54091 -61556
rect 54867 -61590 54879 -61556
rect 54079 -61602 54879 -61590
rect 57123 -61529 57175 -61509
rect 57123 -61563 57131 -61529
rect 57165 -61563 57175 -61529
rect 57123 -61597 57175 -61563
rect 57123 -61631 57131 -61597
rect 57165 -61631 57175 -61597
rect 57123 -61667 57175 -61631
rect 57205 -61529 57263 -61509
rect 57205 -61563 57217 -61529
rect 57251 -61563 57263 -61529
rect 57205 -61597 57263 -61563
rect 57205 -61631 57217 -61597
rect 57251 -61631 57263 -61597
rect 57205 -61667 57263 -61631
rect 57293 -61529 57345 -61509
rect 57293 -61563 57303 -61529
rect 57337 -61563 57345 -61529
rect 57293 -61610 57345 -61563
rect 57293 -61644 57303 -61610
rect 57337 -61644 57345 -61610
rect 57293 -61667 57345 -61644
rect 59113 -61447 59513 -61435
rect 59113 -61481 59125 -61447
rect 59501 -61481 59513 -61447
rect 59113 -61493 59513 -61481
rect 59113 -61555 59513 -61543
rect 59113 -61589 59125 -61555
rect 59501 -61589 59513 -61555
rect 59113 -61601 59513 -61589
rect 59113 -61663 59513 -61651
rect 59113 -61697 59125 -61663
rect 59501 -61697 59513 -61663
rect 59113 -61709 59513 -61697
rect 54069 -63388 54869 -63376
rect 54069 -63422 54081 -63388
rect 54857 -63422 54869 -63388
rect 54069 -63434 54869 -63422
rect 54069 -63516 54869 -63504
rect 54069 -63550 54081 -63516
rect 54857 -63550 54869 -63516
rect 54069 -63562 54869 -63550
rect 56418 -62099 56476 -62087
rect 56418 -62875 56430 -62099
rect 56464 -62875 56476 -62099
rect 56418 -62887 56476 -62875
rect 56546 -62099 56604 -62087
rect 56546 -62875 56558 -62099
rect 56592 -62875 56604 -62099
rect 56546 -62887 56604 -62875
rect 59032 -61971 59090 -61959
rect 59032 -62347 59044 -61971
rect 59078 -62347 59090 -61971
rect 59032 -62359 59090 -62347
rect 59150 -61971 59208 -61959
rect 59150 -62347 59162 -61971
rect 59196 -62347 59208 -61971
rect 59150 -62359 59208 -62347
rect 60441 -62373 60641 -62365
rect 60441 -62407 60459 -62373
rect 60493 -62407 60527 -62373
rect 60561 -62407 60595 -62373
rect 60629 -62407 60641 -62373
rect 60441 -62417 60641 -62407
rect 60811 -62373 61011 -62365
rect 60811 -62407 60823 -62373
rect 60857 -62407 60891 -62373
rect 60925 -62407 60959 -62373
rect 60993 -62407 61011 -62373
rect 60811 -62417 61011 -62407
rect 60441 -62457 60641 -62447
rect 60441 -62491 60459 -62457
rect 60493 -62491 60527 -62457
rect 60561 -62491 60595 -62457
rect 60629 -62491 60641 -62457
rect 60441 -62501 60641 -62491
rect 60811 -62457 61011 -62447
rect 60811 -62491 60823 -62457
rect 60857 -62491 60891 -62457
rect 60925 -62491 60959 -62457
rect 60993 -62491 61011 -62457
rect 60811 -62501 61011 -62491
rect 59032 -62701 59090 -62689
rect 59032 -63077 59044 -62701
rect 59078 -63077 59090 -62701
rect 59032 -63089 59090 -63077
rect 59150 -62701 59208 -62689
rect 59150 -63077 59162 -62701
rect 59196 -63077 59208 -62701
rect 59150 -63089 59208 -63077
rect 60441 -62541 60641 -62531
rect 60441 -62575 60527 -62541
rect 60561 -62575 60595 -62541
rect 60629 -62575 60641 -62541
rect 60441 -62585 60641 -62575
rect 60811 -62541 61011 -62531
rect 60811 -62575 60823 -62541
rect 60857 -62575 60891 -62541
rect 60925 -62575 61011 -62541
rect 60811 -62585 61011 -62575
rect 60441 -62625 60641 -62615
rect 60441 -62659 60459 -62625
rect 60493 -62659 60527 -62625
rect 60561 -62659 60595 -62625
rect 60629 -62659 60641 -62625
rect 60441 -62669 60641 -62659
rect 60811 -62625 61011 -62615
rect 60811 -62659 60823 -62625
rect 60857 -62659 60891 -62625
rect 60925 -62659 60959 -62625
rect 60993 -62659 61011 -62625
rect 60811 -62669 61011 -62659
rect 60441 -62709 60641 -62699
rect 60441 -62743 60595 -62709
rect 60629 -62743 60641 -62709
rect 60441 -62751 60641 -62743
rect 60811 -62709 61011 -62699
rect 60811 -62743 60823 -62709
rect 60857 -62743 61011 -62709
rect 60811 -62751 61011 -62743
rect 57123 -63357 57175 -63321
rect 57123 -63391 57131 -63357
rect 57165 -63391 57175 -63357
rect 57123 -63425 57175 -63391
rect 57123 -63459 57131 -63425
rect 57165 -63459 57175 -63425
rect 57123 -63479 57175 -63459
rect 57205 -63357 57263 -63321
rect 57205 -63391 57217 -63357
rect 57251 -63391 57263 -63357
rect 57205 -63425 57263 -63391
rect 57205 -63459 57217 -63425
rect 57251 -63459 57263 -63425
rect 57205 -63479 57263 -63459
rect 57293 -63344 57345 -63321
rect 57293 -63378 57303 -63344
rect 57337 -63378 57345 -63344
rect 57293 -63425 57345 -63378
rect 57293 -63459 57303 -63425
rect 57337 -63459 57345 -63425
rect 57293 -63479 57345 -63459
rect 59113 -63354 59513 -63342
rect 59113 -63388 59125 -63354
rect 59501 -63388 59513 -63354
rect 59113 -63400 59513 -63388
rect 59113 -63462 59513 -63450
rect 59113 -63496 59125 -63462
rect 59501 -63496 59513 -63462
rect 59113 -63508 59513 -63496
rect 59113 -63570 59513 -63558
rect 59113 -63604 59125 -63570
rect 59501 -63604 59513 -63570
rect 59113 -63616 59513 -63604
rect 54069 -63744 54869 -63732
rect 54069 -63778 54081 -63744
rect 54857 -63778 54869 -63744
rect 54069 -63790 54869 -63778
rect 54069 -63872 54869 -63860
rect 54069 -63906 54081 -63872
rect 54857 -63906 54869 -63872
rect 54069 -63918 54869 -63906
rect 54079 -66472 54879 -66460
rect 54079 -66506 54091 -66472
rect 54867 -66506 54879 -66472
rect 54079 -66518 54879 -66506
rect 54079 -66600 54879 -66588
rect 54079 -66634 54091 -66600
rect 54867 -66634 54879 -66600
rect 54079 -66646 54879 -66634
rect 54079 -66828 54879 -66816
rect 54079 -66862 54091 -66828
rect 54867 -66862 54879 -66828
rect 54079 -66874 54879 -66862
rect 54079 -66956 54879 -66944
rect 54079 -66990 54091 -66956
rect 54867 -66990 54879 -66956
rect 54079 -67002 54879 -66990
rect 57123 -66929 57175 -66909
rect 57123 -66963 57131 -66929
rect 57165 -66963 57175 -66929
rect 57123 -66997 57175 -66963
rect 57123 -67031 57131 -66997
rect 57165 -67031 57175 -66997
rect 57123 -67067 57175 -67031
rect 57205 -66929 57263 -66909
rect 57205 -66963 57217 -66929
rect 57251 -66963 57263 -66929
rect 57205 -66997 57263 -66963
rect 57205 -67031 57217 -66997
rect 57251 -67031 57263 -66997
rect 57205 -67067 57263 -67031
rect 57293 -66929 57345 -66909
rect 57293 -66963 57303 -66929
rect 57337 -66963 57345 -66929
rect 57293 -67010 57345 -66963
rect 57293 -67044 57303 -67010
rect 57337 -67044 57345 -67010
rect 57293 -67067 57345 -67044
rect 59113 -66847 59513 -66835
rect 59113 -66881 59125 -66847
rect 59501 -66881 59513 -66847
rect 59113 -66893 59513 -66881
rect 59113 -66955 59513 -66943
rect 59113 -66989 59125 -66955
rect 59501 -66989 59513 -66955
rect 59113 -67001 59513 -66989
rect 59113 -67063 59513 -67051
rect 59113 -67097 59125 -67063
rect 59501 -67097 59513 -67063
rect 59113 -67109 59513 -67097
rect 54069 -68788 54869 -68776
rect 54069 -68822 54081 -68788
rect 54857 -68822 54869 -68788
rect 54069 -68834 54869 -68822
rect 54069 -68916 54869 -68904
rect 54069 -68950 54081 -68916
rect 54857 -68950 54869 -68916
rect 54069 -68962 54869 -68950
rect 56418 -67499 56476 -67487
rect 56418 -68275 56430 -67499
rect 56464 -68275 56476 -67499
rect 56418 -68287 56476 -68275
rect 56546 -67499 56604 -67487
rect 56546 -68275 56558 -67499
rect 56592 -68275 56604 -67499
rect 56546 -68287 56604 -68275
rect 59032 -67371 59090 -67359
rect 59032 -67747 59044 -67371
rect 59078 -67747 59090 -67371
rect 59032 -67759 59090 -67747
rect 59150 -67371 59208 -67359
rect 59150 -67747 59162 -67371
rect 59196 -67747 59208 -67371
rect 59150 -67759 59208 -67747
rect 60441 -67773 60641 -67765
rect 60441 -67807 60459 -67773
rect 60493 -67807 60527 -67773
rect 60561 -67807 60595 -67773
rect 60629 -67807 60641 -67773
rect 60441 -67817 60641 -67807
rect 60811 -67773 61011 -67765
rect 60811 -67807 60823 -67773
rect 60857 -67807 60891 -67773
rect 60925 -67807 60959 -67773
rect 60993 -67807 61011 -67773
rect 60811 -67817 61011 -67807
rect 60441 -67857 60641 -67847
rect 60441 -67891 60459 -67857
rect 60493 -67891 60527 -67857
rect 60561 -67891 60595 -67857
rect 60629 -67891 60641 -67857
rect 60441 -67901 60641 -67891
rect 60811 -67857 61011 -67847
rect 60811 -67891 60823 -67857
rect 60857 -67891 60891 -67857
rect 60925 -67891 60959 -67857
rect 60993 -67891 61011 -67857
rect 60811 -67901 61011 -67891
rect 59032 -68101 59090 -68089
rect 59032 -68477 59044 -68101
rect 59078 -68477 59090 -68101
rect 59032 -68489 59090 -68477
rect 59150 -68101 59208 -68089
rect 59150 -68477 59162 -68101
rect 59196 -68477 59208 -68101
rect 59150 -68489 59208 -68477
rect 60441 -67941 60641 -67931
rect 60441 -67975 60527 -67941
rect 60561 -67975 60595 -67941
rect 60629 -67975 60641 -67941
rect 60441 -67985 60641 -67975
rect 60811 -67941 61011 -67931
rect 60811 -67975 60823 -67941
rect 60857 -67975 60891 -67941
rect 60925 -67975 61011 -67941
rect 60811 -67985 61011 -67975
rect 60441 -68025 60641 -68015
rect 60441 -68059 60459 -68025
rect 60493 -68059 60527 -68025
rect 60561 -68059 60595 -68025
rect 60629 -68059 60641 -68025
rect 60441 -68069 60641 -68059
rect 60811 -68025 61011 -68015
rect 60811 -68059 60823 -68025
rect 60857 -68059 60891 -68025
rect 60925 -68059 60959 -68025
rect 60993 -68059 61011 -68025
rect 60811 -68069 61011 -68059
rect 60441 -68109 60641 -68099
rect 60441 -68143 60595 -68109
rect 60629 -68143 60641 -68109
rect 60441 -68151 60641 -68143
rect 60811 -68109 61011 -68099
rect 60811 -68143 60823 -68109
rect 60857 -68143 61011 -68109
rect 60811 -68151 61011 -68143
rect 57123 -68757 57175 -68721
rect 57123 -68791 57131 -68757
rect 57165 -68791 57175 -68757
rect 57123 -68825 57175 -68791
rect 57123 -68859 57131 -68825
rect 57165 -68859 57175 -68825
rect 57123 -68879 57175 -68859
rect 57205 -68757 57263 -68721
rect 57205 -68791 57217 -68757
rect 57251 -68791 57263 -68757
rect 57205 -68825 57263 -68791
rect 57205 -68859 57217 -68825
rect 57251 -68859 57263 -68825
rect 57205 -68879 57263 -68859
rect 57293 -68744 57345 -68721
rect 57293 -68778 57303 -68744
rect 57337 -68778 57345 -68744
rect 57293 -68825 57345 -68778
rect 57293 -68859 57303 -68825
rect 57337 -68859 57345 -68825
rect 57293 -68879 57345 -68859
rect 59113 -68754 59513 -68742
rect 59113 -68788 59125 -68754
rect 59501 -68788 59513 -68754
rect 59113 -68800 59513 -68788
rect 59113 -68862 59513 -68850
rect 59113 -68896 59125 -68862
rect 59501 -68896 59513 -68862
rect 59113 -68908 59513 -68896
rect 59113 -68970 59513 -68958
rect 59113 -69004 59125 -68970
rect 59501 -69004 59513 -68970
rect 59113 -69016 59513 -69004
rect 54069 -69144 54869 -69132
rect 54069 -69178 54081 -69144
rect 54857 -69178 54869 -69144
rect 54069 -69190 54869 -69178
rect 54069 -69272 54869 -69260
rect 54069 -69306 54081 -69272
rect 54857 -69306 54869 -69272
rect 54069 -69318 54869 -69306
rect 54079 -71872 54879 -71860
rect 54079 -71906 54091 -71872
rect 54867 -71906 54879 -71872
rect 54079 -71918 54879 -71906
rect 54079 -72000 54879 -71988
rect 54079 -72034 54091 -72000
rect 54867 -72034 54879 -72000
rect 54079 -72046 54879 -72034
rect 54079 -72228 54879 -72216
rect 54079 -72262 54091 -72228
rect 54867 -72262 54879 -72228
rect 54079 -72274 54879 -72262
rect 54079 -72356 54879 -72344
rect 54079 -72390 54091 -72356
rect 54867 -72390 54879 -72356
rect 54079 -72402 54879 -72390
rect 57123 -72329 57175 -72309
rect 57123 -72363 57131 -72329
rect 57165 -72363 57175 -72329
rect 57123 -72397 57175 -72363
rect 57123 -72431 57131 -72397
rect 57165 -72431 57175 -72397
rect 57123 -72467 57175 -72431
rect 57205 -72329 57263 -72309
rect 57205 -72363 57217 -72329
rect 57251 -72363 57263 -72329
rect 57205 -72397 57263 -72363
rect 57205 -72431 57217 -72397
rect 57251 -72431 57263 -72397
rect 57205 -72467 57263 -72431
rect 57293 -72329 57345 -72309
rect 57293 -72363 57303 -72329
rect 57337 -72363 57345 -72329
rect 57293 -72410 57345 -72363
rect 57293 -72444 57303 -72410
rect 57337 -72444 57345 -72410
rect 57293 -72467 57345 -72444
rect 59113 -72247 59513 -72235
rect 59113 -72281 59125 -72247
rect 59501 -72281 59513 -72247
rect 59113 -72293 59513 -72281
rect 59113 -72355 59513 -72343
rect 59113 -72389 59125 -72355
rect 59501 -72389 59513 -72355
rect 59113 -72401 59513 -72389
rect 59113 -72463 59513 -72451
rect 59113 -72497 59125 -72463
rect 59501 -72497 59513 -72463
rect 59113 -72509 59513 -72497
rect 54069 -74188 54869 -74176
rect 54069 -74222 54081 -74188
rect 54857 -74222 54869 -74188
rect 54069 -74234 54869 -74222
rect 54069 -74316 54869 -74304
rect 54069 -74350 54081 -74316
rect 54857 -74350 54869 -74316
rect 54069 -74362 54869 -74350
rect 56418 -72899 56476 -72887
rect 56418 -73675 56430 -72899
rect 56464 -73675 56476 -72899
rect 56418 -73687 56476 -73675
rect 56546 -72899 56604 -72887
rect 56546 -73675 56558 -72899
rect 56592 -73675 56604 -72899
rect 56546 -73687 56604 -73675
rect 59032 -72771 59090 -72759
rect 59032 -73147 59044 -72771
rect 59078 -73147 59090 -72771
rect 59032 -73159 59090 -73147
rect 59150 -72771 59208 -72759
rect 59150 -73147 59162 -72771
rect 59196 -73147 59208 -72771
rect 59150 -73159 59208 -73147
rect 60441 -73173 60641 -73165
rect 60441 -73207 60459 -73173
rect 60493 -73207 60527 -73173
rect 60561 -73207 60595 -73173
rect 60629 -73207 60641 -73173
rect 60441 -73217 60641 -73207
rect 60811 -73173 61011 -73165
rect 60811 -73207 60823 -73173
rect 60857 -73207 60891 -73173
rect 60925 -73207 60959 -73173
rect 60993 -73207 61011 -73173
rect 60811 -73217 61011 -73207
rect 60441 -73257 60641 -73247
rect 60441 -73291 60459 -73257
rect 60493 -73291 60527 -73257
rect 60561 -73291 60595 -73257
rect 60629 -73291 60641 -73257
rect 60441 -73301 60641 -73291
rect 60811 -73257 61011 -73247
rect 60811 -73291 60823 -73257
rect 60857 -73291 60891 -73257
rect 60925 -73291 60959 -73257
rect 60993 -73291 61011 -73257
rect 60811 -73301 61011 -73291
rect 59032 -73501 59090 -73489
rect 59032 -73877 59044 -73501
rect 59078 -73877 59090 -73501
rect 59032 -73889 59090 -73877
rect 59150 -73501 59208 -73489
rect 59150 -73877 59162 -73501
rect 59196 -73877 59208 -73501
rect 59150 -73889 59208 -73877
rect 60441 -73341 60641 -73331
rect 60441 -73375 60527 -73341
rect 60561 -73375 60595 -73341
rect 60629 -73375 60641 -73341
rect 60441 -73385 60641 -73375
rect 60811 -73341 61011 -73331
rect 60811 -73375 60823 -73341
rect 60857 -73375 60891 -73341
rect 60925 -73375 61011 -73341
rect 60811 -73385 61011 -73375
rect 60441 -73425 60641 -73415
rect 60441 -73459 60459 -73425
rect 60493 -73459 60527 -73425
rect 60561 -73459 60595 -73425
rect 60629 -73459 60641 -73425
rect 60441 -73469 60641 -73459
rect 60811 -73425 61011 -73415
rect 60811 -73459 60823 -73425
rect 60857 -73459 60891 -73425
rect 60925 -73459 60959 -73425
rect 60993 -73459 61011 -73425
rect 60811 -73469 61011 -73459
rect 60441 -73509 60641 -73499
rect 60441 -73543 60595 -73509
rect 60629 -73543 60641 -73509
rect 60441 -73551 60641 -73543
rect 60811 -73509 61011 -73499
rect 60811 -73543 60823 -73509
rect 60857 -73543 61011 -73509
rect 60811 -73551 61011 -73543
rect 57123 -74157 57175 -74121
rect 57123 -74191 57131 -74157
rect 57165 -74191 57175 -74157
rect 57123 -74225 57175 -74191
rect 57123 -74259 57131 -74225
rect 57165 -74259 57175 -74225
rect 57123 -74279 57175 -74259
rect 57205 -74157 57263 -74121
rect 57205 -74191 57217 -74157
rect 57251 -74191 57263 -74157
rect 57205 -74225 57263 -74191
rect 57205 -74259 57217 -74225
rect 57251 -74259 57263 -74225
rect 57205 -74279 57263 -74259
rect 57293 -74144 57345 -74121
rect 57293 -74178 57303 -74144
rect 57337 -74178 57345 -74144
rect 57293 -74225 57345 -74178
rect 57293 -74259 57303 -74225
rect 57337 -74259 57345 -74225
rect 57293 -74279 57345 -74259
rect 59113 -74154 59513 -74142
rect 59113 -74188 59125 -74154
rect 59501 -74188 59513 -74154
rect 59113 -74200 59513 -74188
rect 59113 -74262 59513 -74250
rect 59113 -74296 59125 -74262
rect 59501 -74296 59513 -74262
rect 59113 -74308 59513 -74296
rect 59113 -74370 59513 -74358
rect 59113 -74404 59125 -74370
rect 59501 -74404 59513 -74370
rect 59113 -74416 59513 -74404
rect 54069 -74544 54869 -74532
rect 54069 -74578 54081 -74544
rect 54857 -74578 54869 -74544
rect 54069 -74590 54869 -74578
rect 54069 -74672 54869 -74660
rect 54069 -74706 54081 -74672
rect 54857 -74706 54869 -74672
rect 54069 -74718 54869 -74706
rect 54079 -77272 54879 -77260
rect 54079 -77306 54091 -77272
rect 54867 -77306 54879 -77272
rect 54079 -77318 54879 -77306
rect 54079 -77400 54879 -77388
rect 54079 -77434 54091 -77400
rect 54867 -77434 54879 -77400
rect 54079 -77446 54879 -77434
rect 54079 -77628 54879 -77616
rect 54079 -77662 54091 -77628
rect 54867 -77662 54879 -77628
rect 54079 -77674 54879 -77662
rect 54079 -77756 54879 -77744
rect 54079 -77790 54091 -77756
rect 54867 -77790 54879 -77756
rect 54079 -77802 54879 -77790
rect 57123 -77729 57175 -77709
rect 57123 -77763 57131 -77729
rect 57165 -77763 57175 -77729
rect 57123 -77797 57175 -77763
rect 57123 -77831 57131 -77797
rect 57165 -77831 57175 -77797
rect 57123 -77867 57175 -77831
rect 57205 -77729 57263 -77709
rect 57205 -77763 57217 -77729
rect 57251 -77763 57263 -77729
rect 57205 -77797 57263 -77763
rect 57205 -77831 57217 -77797
rect 57251 -77831 57263 -77797
rect 57205 -77867 57263 -77831
rect 57293 -77729 57345 -77709
rect 57293 -77763 57303 -77729
rect 57337 -77763 57345 -77729
rect 57293 -77810 57345 -77763
rect 57293 -77844 57303 -77810
rect 57337 -77844 57345 -77810
rect 57293 -77867 57345 -77844
rect 59113 -77647 59513 -77635
rect 59113 -77681 59125 -77647
rect 59501 -77681 59513 -77647
rect 59113 -77693 59513 -77681
rect 59113 -77755 59513 -77743
rect 59113 -77789 59125 -77755
rect 59501 -77789 59513 -77755
rect 59113 -77801 59513 -77789
rect 59113 -77863 59513 -77851
rect 59113 -77897 59125 -77863
rect 59501 -77897 59513 -77863
rect 59113 -77909 59513 -77897
rect 54069 -79588 54869 -79576
rect 54069 -79622 54081 -79588
rect 54857 -79622 54869 -79588
rect 54069 -79634 54869 -79622
rect 54069 -79716 54869 -79704
rect 54069 -79750 54081 -79716
rect 54857 -79750 54869 -79716
rect 54069 -79762 54869 -79750
rect 56418 -78299 56476 -78287
rect 56418 -79075 56430 -78299
rect 56464 -79075 56476 -78299
rect 56418 -79087 56476 -79075
rect 56546 -78299 56604 -78287
rect 56546 -79075 56558 -78299
rect 56592 -79075 56604 -78299
rect 56546 -79087 56604 -79075
rect 59032 -78171 59090 -78159
rect 59032 -78547 59044 -78171
rect 59078 -78547 59090 -78171
rect 59032 -78559 59090 -78547
rect 59150 -78171 59208 -78159
rect 59150 -78547 59162 -78171
rect 59196 -78547 59208 -78171
rect 59150 -78559 59208 -78547
rect 60441 -78573 60641 -78565
rect 60441 -78607 60459 -78573
rect 60493 -78607 60527 -78573
rect 60561 -78607 60595 -78573
rect 60629 -78607 60641 -78573
rect 60441 -78617 60641 -78607
rect 60811 -78573 61011 -78565
rect 60811 -78607 60823 -78573
rect 60857 -78607 60891 -78573
rect 60925 -78607 60959 -78573
rect 60993 -78607 61011 -78573
rect 60811 -78617 61011 -78607
rect 60441 -78657 60641 -78647
rect 60441 -78691 60459 -78657
rect 60493 -78691 60527 -78657
rect 60561 -78691 60595 -78657
rect 60629 -78691 60641 -78657
rect 60441 -78701 60641 -78691
rect 60811 -78657 61011 -78647
rect 60811 -78691 60823 -78657
rect 60857 -78691 60891 -78657
rect 60925 -78691 60959 -78657
rect 60993 -78691 61011 -78657
rect 60811 -78701 61011 -78691
rect 59032 -78901 59090 -78889
rect 59032 -79277 59044 -78901
rect 59078 -79277 59090 -78901
rect 59032 -79289 59090 -79277
rect 59150 -78901 59208 -78889
rect 59150 -79277 59162 -78901
rect 59196 -79277 59208 -78901
rect 59150 -79289 59208 -79277
rect 60441 -78741 60641 -78731
rect 60441 -78775 60527 -78741
rect 60561 -78775 60595 -78741
rect 60629 -78775 60641 -78741
rect 60441 -78785 60641 -78775
rect 60811 -78741 61011 -78731
rect 60811 -78775 60823 -78741
rect 60857 -78775 60891 -78741
rect 60925 -78775 61011 -78741
rect 60811 -78785 61011 -78775
rect 60441 -78825 60641 -78815
rect 60441 -78859 60459 -78825
rect 60493 -78859 60527 -78825
rect 60561 -78859 60595 -78825
rect 60629 -78859 60641 -78825
rect 60441 -78869 60641 -78859
rect 60811 -78825 61011 -78815
rect 60811 -78859 60823 -78825
rect 60857 -78859 60891 -78825
rect 60925 -78859 60959 -78825
rect 60993 -78859 61011 -78825
rect 60811 -78869 61011 -78859
rect 60441 -78909 60641 -78899
rect 60441 -78943 60595 -78909
rect 60629 -78943 60641 -78909
rect 60441 -78951 60641 -78943
rect 60811 -78909 61011 -78899
rect 60811 -78943 60823 -78909
rect 60857 -78943 61011 -78909
rect 60811 -78951 61011 -78943
rect 57123 -79557 57175 -79521
rect 57123 -79591 57131 -79557
rect 57165 -79591 57175 -79557
rect 57123 -79625 57175 -79591
rect 57123 -79659 57131 -79625
rect 57165 -79659 57175 -79625
rect 57123 -79679 57175 -79659
rect 57205 -79557 57263 -79521
rect 57205 -79591 57217 -79557
rect 57251 -79591 57263 -79557
rect 57205 -79625 57263 -79591
rect 57205 -79659 57217 -79625
rect 57251 -79659 57263 -79625
rect 57205 -79679 57263 -79659
rect 57293 -79544 57345 -79521
rect 57293 -79578 57303 -79544
rect 57337 -79578 57345 -79544
rect 57293 -79625 57345 -79578
rect 57293 -79659 57303 -79625
rect 57337 -79659 57345 -79625
rect 57293 -79679 57345 -79659
rect 59113 -79554 59513 -79542
rect 59113 -79588 59125 -79554
rect 59501 -79588 59513 -79554
rect 59113 -79600 59513 -79588
rect 59113 -79662 59513 -79650
rect 59113 -79696 59125 -79662
rect 59501 -79696 59513 -79662
rect 59113 -79708 59513 -79696
rect 59113 -79770 59513 -79758
rect 59113 -79804 59125 -79770
rect 59501 -79804 59513 -79770
rect 59113 -79816 59513 -79804
rect 54069 -79944 54869 -79932
rect 54069 -79978 54081 -79944
rect 54857 -79978 54869 -79944
rect 54069 -79990 54869 -79978
rect 54069 -80072 54869 -80060
rect 54069 -80106 54081 -80072
rect 54857 -80106 54869 -80072
rect 54069 -80118 54869 -80106
rect 54079 -82672 54879 -82660
rect 54079 -82706 54091 -82672
rect 54867 -82706 54879 -82672
rect 54079 -82718 54879 -82706
rect 54079 -82800 54879 -82788
rect 54079 -82834 54091 -82800
rect 54867 -82834 54879 -82800
rect 54079 -82846 54879 -82834
rect 54079 -83028 54879 -83016
rect 54079 -83062 54091 -83028
rect 54867 -83062 54879 -83028
rect 54079 -83074 54879 -83062
rect 54079 -83156 54879 -83144
rect 54079 -83190 54091 -83156
rect 54867 -83190 54879 -83156
rect 54079 -83202 54879 -83190
rect 57123 -83129 57175 -83109
rect 57123 -83163 57131 -83129
rect 57165 -83163 57175 -83129
rect 57123 -83197 57175 -83163
rect 57123 -83231 57131 -83197
rect 57165 -83231 57175 -83197
rect 57123 -83267 57175 -83231
rect 57205 -83129 57263 -83109
rect 57205 -83163 57217 -83129
rect 57251 -83163 57263 -83129
rect 57205 -83197 57263 -83163
rect 57205 -83231 57217 -83197
rect 57251 -83231 57263 -83197
rect 57205 -83267 57263 -83231
rect 57293 -83129 57345 -83109
rect 57293 -83163 57303 -83129
rect 57337 -83163 57345 -83129
rect 57293 -83210 57345 -83163
rect 57293 -83244 57303 -83210
rect 57337 -83244 57345 -83210
rect 57293 -83267 57345 -83244
rect 59113 -83047 59513 -83035
rect 59113 -83081 59125 -83047
rect 59501 -83081 59513 -83047
rect 59113 -83093 59513 -83081
rect 59113 -83155 59513 -83143
rect 59113 -83189 59125 -83155
rect 59501 -83189 59513 -83155
rect 59113 -83201 59513 -83189
rect 59113 -83263 59513 -83251
rect 59113 -83297 59125 -83263
rect 59501 -83297 59513 -83263
rect 59113 -83309 59513 -83297
rect 54069 -84988 54869 -84976
rect 54069 -85022 54081 -84988
rect 54857 -85022 54869 -84988
rect 54069 -85034 54869 -85022
rect 54069 -85116 54869 -85104
rect 54069 -85150 54081 -85116
rect 54857 -85150 54869 -85116
rect 54069 -85162 54869 -85150
rect 56418 -83699 56476 -83687
rect 56418 -84475 56430 -83699
rect 56464 -84475 56476 -83699
rect 56418 -84487 56476 -84475
rect 56546 -83699 56604 -83687
rect 56546 -84475 56558 -83699
rect 56592 -84475 56604 -83699
rect 56546 -84487 56604 -84475
rect 59032 -83571 59090 -83559
rect 59032 -83947 59044 -83571
rect 59078 -83947 59090 -83571
rect 59032 -83959 59090 -83947
rect 59150 -83571 59208 -83559
rect 59150 -83947 59162 -83571
rect 59196 -83947 59208 -83571
rect 59150 -83959 59208 -83947
rect 60441 -83973 60641 -83965
rect 60441 -84007 60459 -83973
rect 60493 -84007 60527 -83973
rect 60561 -84007 60595 -83973
rect 60629 -84007 60641 -83973
rect 60441 -84017 60641 -84007
rect 60811 -83973 61011 -83965
rect 60811 -84007 60823 -83973
rect 60857 -84007 60891 -83973
rect 60925 -84007 60959 -83973
rect 60993 -84007 61011 -83973
rect 60811 -84017 61011 -84007
rect 60441 -84057 60641 -84047
rect 60441 -84091 60459 -84057
rect 60493 -84091 60527 -84057
rect 60561 -84091 60595 -84057
rect 60629 -84091 60641 -84057
rect 60441 -84101 60641 -84091
rect 60811 -84057 61011 -84047
rect 60811 -84091 60823 -84057
rect 60857 -84091 60891 -84057
rect 60925 -84091 60959 -84057
rect 60993 -84091 61011 -84057
rect 60811 -84101 61011 -84091
rect 59032 -84301 59090 -84289
rect 59032 -84677 59044 -84301
rect 59078 -84677 59090 -84301
rect 59032 -84689 59090 -84677
rect 59150 -84301 59208 -84289
rect 59150 -84677 59162 -84301
rect 59196 -84677 59208 -84301
rect 59150 -84689 59208 -84677
rect 60441 -84141 60641 -84131
rect 60441 -84175 60527 -84141
rect 60561 -84175 60595 -84141
rect 60629 -84175 60641 -84141
rect 60441 -84185 60641 -84175
rect 60811 -84141 61011 -84131
rect 60811 -84175 60823 -84141
rect 60857 -84175 60891 -84141
rect 60925 -84175 61011 -84141
rect 60811 -84185 61011 -84175
rect 60441 -84225 60641 -84215
rect 60441 -84259 60459 -84225
rect 60493 -84259 60527 -84225
rect 60561 -84259 60595 -84225
rect 60629 -84259 60641 -84225
rect 60441 -84269 60641 -84259
rect 60811 -84225 61011 -84215
rect 60811 -84259 60823 -84225
rect 60857 -84259 60891 -84225
rect 60925 -84259 60959 -84225
rect 60993 -84259 61011 -84225
rect 60811 -84269 61011 -84259
rect 60441 -84309 60641 -84299
rect 60441 -84343 60595 -84309
rect 60629 -84343 60641 -84309
rect 60441 -84351 60641 -84343
rect 60811 -84309 61011 -84299
rect 60811 -84343 60823 -84309
rect 60857 -84343 61011 -84309
rect 60811 -84351 61011 -84343
rect 57123 -84957 57175 -84921
rect 57123 -84991 57131 -84957
rect 57165 -84991 57175 -84957
rect 57123 -85025 57175 -84991
rect 57123 -85059 57131 -85025
rect 57165 -85059 57175 -85025
rect 57123 -85079 57175 -85059
rect 57205 -84957 57263 -84921
rect 57205 -84991 57217 -84957
rect 57251 -84991 57263 -84957
rect 57205 -85025 57263 -84991
rect 57205 -85059 57217 -85025
rect 57251 -85059 57263 -85025
rect 57205 -85079 57263 -85059
rect 57293 -84944 57345 -84921
rect 57293 -84978 57303 -84944
rect 57337 -84978 57345 -84944
rect 57293 -85025 57345 -84978
rect 57293 -85059 57303 -85025
rect 57337 -85059 57345 -85025
rect 57293 -85079 57345 -85059
rect 59113 -84954 59513 -84942
rect 59113 -84988 59125 -84954
rect 59501 -84988 59513 -84954
rect 59113 -85000 59513 -84988
rect 59113 -85062 59513 -85050
rect 59113 -85096 59125 -85062
rect 59501 -85096 59513 -85062
rect 59113 -85108 59513 -85096
rect 59113 -85170 59513 -85158
rect 59113 -85204 59125 -85170
rect 59501 -85204 59513 -85170
rect 59113 -85216 59513 -85204
rect 54069 -85344 54869 -85332
rect 54069 -85378 54081 -85344
rect 54857 -85378 54869 -85344
rect 54069 -85390 54869 -85378
rect 54069 -85472 54869 -85460
rect 54069 -85506 54081 -85472
rect 54857 -85506 54869 -85472
rect 54069 -85518 54869 -85506
<< ndiffc >>
rect 53464 -2966 53498 -2190
rect 53642 -2966 53676 -2190
rect 55290 -2428 55324 -2252
rect 55378 -2428 55412 -2252
rect 53942 -2812 54718 -2778
rect 53942 -2990 54718 -2956
rect 55820 -2916 55854 -2140
rect 55998 -2916 56032 -2140
rect 53464 -3984 53498 -3208
rect 53642 -3984 53676 -3208
rect 53942 -3218 54718 -3184
rect 53942 -3396 54718 -3362
rect 55280 -3924 55314 -3748
rect 55368 -3924 55402 -3748
rect 55820 -4030 55854 -3254
rect 55998 -4030 56032 -3254
rect 57131 -2534 57165 -2500
rect 57217 -2547 57251 -2513
rect 57303 -2517 57337 -2483
rect 59958 -2408 60334 -2374
rect 59958 -2516 60334 -2482
rect 59502 -2958 59536 -2782
rect 59590 -2958 59624 -2782
rect 59818 -2958 59852 -2782
rect 59906 -2958 59940 -2782
rect 60203 -3007 60237 -2973
rect 61215 -3007 61249 -2973
rect 60211 -3091 60245 -3057
rect 61207 -3091 61241 -3057
rect 57131 -3688 57165 -3654
rect 57217 -3675 57251 -3641
rect 57303 -3705 57337 -3671
rect 59501 -3471 59535 -3295
rect 59589 -3471 59623 -3295
rect 60203 -3175 60237 -3141
rect 61215 -3175 61249 -3141
rect 59817 -3471 59851 -3295
rect 59905 -3471 59939 -3295
rect 60211 -3259 60245 -3225
rect 61207 -3259 61241 -3225
rect 60204 -3343 60238 -3309
rect 61214 -3343 61248 -3309
rect 59958 -3774 60334 -3740
rect 59958 -3882 60334 -3848
rect 55300 -4592 55476 -4558
rect 55300 -4680 55476 -4646
rect 53464 -8366 53498 -7590
rect 53642 -8366 53676 -7590
rect 55290 -7828 55324 -7652
rect 55378 -7828 55412 -7652
rect 53942 -8212 54718 -8178
rect 53942 -8390 54718 -8356
rect 55820 -8316 55854 -7540
rect 55998 -8316 56032 -7540
rect 53464 -9384 53498 -8608
rect 53642 -9384 53676 -8608
rect 53942 -8618 54718 -8584
rect 53942 -8796 54718 -8762
rect 55280 -9324 55314 -9148
rect 55368 -9324 55402 -9148
rect 55820 -9430 55854 -8654
rect 55998 -9430 56032 -8654
rect 57131 -7934 57165 -7900
rect 57217 -7947 57251 -7913
rect 57303 -7917 57337 -7883
rect 59958 -7808 60334 -7774
rect 59958 -7916 60334 -7882
rect 59502 -8358 59536 -8182
rect 59590 -8358 59624 -8182
rect 59818 -8358 59852 -8182
rect 59906 -8358 59940 -8182
rect 60203 -8407 60237 -8373
rect 61215 -8407 61249 -8373
rect 60211 -8491 60245 -8457
rect 61207 -8491 61241 -8457
rect 57131 -9088 57165 -9054
rect 57217 -9075 57251 -9041
rect 57303 -9105 57337 -9071
rect 59501 -8871 59535 -8695
rect 59589 -8871 59623 -8695
rect 60203 -8575 60237 -8541
rect 61215 -8575 61249 -8541
rect 59817 -8871 59851 -8695
rect 59905 -8871 59939 -8695
rect 60211 -8659 60245 -8625
rect 61207 -8659 61241 -8625
rect 60204 -8743 60238 -8709
rect 61214 -8743 61248 -8709
rect 59958 -9174 60334 -9140
rect 59958 -9282 60334 -9248
rect 55300 -9992 55476 -9958
rect 55300 -10080 55476 -10046
rect 20280 -11964 20340 -11930
rect 20280 -12052 20340 -12018
rect 16553 -13105 16587 -12329
rect 16731 -13105 16765 -12329
rect 16959 -13105 16993 -12329
rect 17137 -13105 17171 -12329
rect 17365 -13105 17399 -12329
rect 17543 -13105 17577 -12329
rect 17771 -13105 17805 -12329
rect 17949 -13105 17983 -12329
rect 18177 -13105 18211 -12329
rect 18355 -13105 18389 -12329
rect 18583 -13105 18617 -12329
rect 18761 -13105 18795 -12329
rect 18989 -13105 19023 -12329
rect 19167 -13105 19201 -12329
rect 19395 -13105 19429 -12329
rect 19573 -13105 19607 -12329
rect 19801 -13105 19835 -12329
rect 19979 -13105 20013 -12329
rect 20207 -13105 20241 -12329
rect 20385 -13105 20419 -12329
rect 20613 -13105 20647 -12329
rect 20791 -13105 20825 -12329
rect 21019 -13105 21053 -12329
rect 21197 -13105 21231 -12329
rect 21425 -13105 21459 -12329
rect 21603 -13105 21637 -12329
rect 21831 -13105 21865 -12329
rect 22009 -13105 22043 -12329
rect 22237 -13105 22271 -12329
rect 22415 -13105 22449 -12329
rect 22643 -13105 22677 -12329
rect 22821 -13105 22855 -12329
rect 23049 -13105 23083 -12329
rect 23227 -13105 23261 -12329
rect 23455 -13105 23489 -12329
rect 23633 -13105 23667 -12329
rect 23861 -13105 23895 -12329
rect 24039 -13105 24073 -12329
rect 24267 -13105 24301 -12329
rect 24445 -13105 24479 -12329
rect 24673 -13105 24707 -12329
rect 24851 -13105 24885 -12329
rect 25079 -13105 25113 -12329
rect 25257 -13105 25291 -12329
rect 53464 -13766 53498 -12990
rect 53642 -13766 53676 -12990
rect 55290 -13228 55324 -13052
rect 55378 -13228 55412 -13052
rect 53942 -13612 54718 -13578
rect 53942 -13790 54718 -13756
rect 55820 -13716 55854 -12940
rect 55998 -13716 56032 -12940
rect 53464 -14784 53498 -14008
rect 53642 -14784 53676 -14008
rect 53942 -14018 54718 -13984
rect 53942 -14196 54718 -14162
rect 55280 -14724 55314 -14548
rect 55368 -14724 55402 -14548
rect 55820 -14830 55854 -14054
rect 55998 -14830 56032 -14054
rect 57131 -13334 57165 -13300
rect 57217 -13347 57251 -13313
rect 57303 -13317 57337 -13283
rect 59958 -13208 60334 -13174
rect 59958 -13316 60334 -13282
rect 59502 -13758 59536 -13582
rect 59590 -13758 59624 -13582
rect 59818 -13758 59852 -13582
rect 59906 -13758 59940 -13582
rect 60203 -13807 60237 -13773
rect 61215 -13807 61249 -13773
rect 60211 -13891 60245 -13857
rect 61207 -13891 61241 -13857
rect 57131 -14488 57165 -14454
rect 57217 -14475 57251 -14441
rect 57303 -14505 57337 -14471
rect 59501 -14271 59535 -14095
rect 59589 -14271 59623 -14095
rect 60203 -13975 60237 -13941
rect 61215 -13975 61249 -13941
rect 59817 -14271 59851 -14095
rect 59905 -14271 59939 -14095
rect 60211 -14059 60245 -14025
rect 61207 -14059 61241 -14025
rect 60204 -14143 60238 -14109
rect 61214 -14143 61248 -14109
rect 59958 -14574 60334 -14540
rect 59958 -14682 60334 -14648
rect 55300 -15392 55476 -15358
rect 55300 -15480 55476 -15446
rect 53464 -19166 53498 -18390
rect 53642 -19166 53676 -18390
rect 55290 -18628 55324 -18452
rect 55378 -18628 55412 -18452
rect 53942 -19012 54718 -18978
rect 53942 -19190 54718 -19156
rect 55820 -19116 55854 -18340
rect 55998 -19116 56032 -18340
rect 53464 -20184 53498 -19408
rect 53642 -20184 53676 -19408
rect 53942 -19418 54718 -19384
rect 53942 -19596 54718 -19562
rect 55280 -20124 55314 -19948
rect 55368 -20124 55402 -19948
rect 55820 -20230 55854 -19454
rect 55998 -20230 56032 -19454
rect 57131 -18734 57165 -18700
rect 57217 -18747 57251 -18713
rect 57303 -18717 57337 -18683
rect 59958 -18608 60334 -18574
rect 59958 -18716 60334 -18682
rect 59502 -19158 59536 -18982
rect 59590 -19158 59624 -18982
rect 59818 -19158 59852 -18982
rect 59906 -19158 59940 -18982
rect 60203 -19207 60237 -19173
rect 61215 -19207 61249 -19173
rect 60211 -19291 60245 -19257
rect 61207 -19291 61241 -19257
rect 57131 -19888 57165 -19854
rect 57217 -19875 57251 -19841
rect 57303 -19905 57337 -19871
rect 59501 -19671 59535 -19495
rect 59589 -19671 59623 -19495
rect 60203 -19375 60237 -19341
rect 61215 -19375 61249 -19341
rect 59817 -19671 59851 -19495
rect 59905 -19671 59939 -19495
rect 60211 -19459 60245 -19425
rect 61207 -19459 61241 -19425
rect 60204 -19543 60238 -19509
rect 61214 -19543 61248 -19509
rect 59958 -19974 60334 -19940
rect 59958 -20082 60334 -20048
rect 55300 -20792 55476 -20758
rect 55300 -20880 55476 -20846
rect 53464 -24566 53498 -23790
rect 53642 -24566 53676 -23790
rect 55290 -24028 55324 -23852
rect 55378 -24028 55412 -23852
rect 53942 -24412 54718 -24378
rect 53942 -24590 54718 -24556
rect 55820 -24516 55854 -23740
rect 55998 -24516 56032 -23740
rect 53464 -25584 53498 -24808
rect 53642 -25584 53676 -24808
rect 53942 -24818 54718 -24784
rect 53942 -24996 54718 -24962
rect 55280 -25524 55314 -25348
rect 55368 -25524 55402 -25348
rect 55820 -25630 55854 -24854
rect 55998 -25630 56032 -24854
rect 57131 -24134 57165 -24100
rect 57217 -24147 57251 -24113
rect 57303 -24117 57337 -24083
rect 59958 -24008 60334 -23974
rect 59958 -24116 60334 -24082
rect 59502 -24558 59536 -24382
rect 59590 -24558 59624 -24382
rect 59818 -24558 59852 -24382
rect 59906 -24558 59940 -24382
rect 60203 -24607 60237 -24573
rect 61215 -24607 61249 -24573
rect 60211 -24691 60245 -24657
rect 61207 -24691 61241 -24657
rect 57131 -25288 57165 -25254
rect 57217 -25275 57251 -25241
rect 57303 -25305 57337 -25271
rect 59501 -25071 59535 -24895
rect 59589 -25071 59623 -24895
rect 60203 -24775 60237 -24741
rect 61215 -24775 61249 -24741
rect 59817 -25071 59851 -24895
rect 59905 -25071 59939 -24895
rect 60211 -24859 60245 -24825
rect 61207 -24859 61241 -24825
rect 60204 -24943 60238 -24909
rect 61214 -24943 61248 -24909
rect 59958 -25374 60334 -25340
rect 59958 -25482 60334 -25448
rect 55300 -26192 55476 -26158
rect 55300 -26280 55476 -26246
rect 53464 -29966 53498 -29190
rect 53642 -29966 53676 -29190
rect 55290 -29428 55324 -29252
rect 55378 -29428 55412 -29252
rect 53942 -29812 54718 -29778
rect 53942 -29990 54718 -29956
rect 55820 -29916 55854 -29140
rect 55998 -29916 56032 -29140
rect 53464 -30984 53498 -30208
rect 53642 -30984 53676 -30208
rect 53942 -30218 54718 -30184
rect 53942 -30396 54718 -30362
rect 55280 -30924 55314 -30748
rect 55368 -30924 55402 -30748
rect 55820 -31030 55854 -30254
rect 55998 -31030 56032 -30254
rect 57131 -29534 57165 -29500
rect 57217 -29547 57251 -29513
rect 57303 -29517 57337 -29483
rect 59958 -29408 60334 -29374
rect 59958 -29516 60334 -29482
rect 59502 -29958 59536 -29782
rect 59590 -29958 59624 -29782
rect 59818 -29958 59852 -29782
rect 59906 -29958 59940 -29782
rect 60203 -30007 60237 -29973
rect 61215 -30007 61249 -29973
rect 60211 -30091 60245 -30057
rect 61207 -30091 61241 -30057
rect 57131 -30688 57165 -30654
rect 57217 -30675 57251 -30641
rect 57303 -30705 57337 -30671
rect 59501 -30471 59535 -30295
rect 59589 -30471 59623 -30295
rect 60203 -30175 60237 -30141
rect 61215 -30175 61249 -30141
rect 59817 -30471 59851 -30295
rect 59905 -30471 59939 -30295
rect 60211 -30259 60245 -30225
rect 61207 -30259 61241 -30225
rect 60204 -30343 60238 -30309
rect 61214 -30343 61248 -30309
rect 59958 -30774 60334 -30740
rect 59958 -30882 60334 -30848
rect 55300 -31592 55476 -31558
rect 55300 -31680 55476 -31646
rect 53464 -35366 53498 -34590
rect 53642 -35366 53676 -34590
rect 55290 -34828 55324 -34652
rect 55378 -34828 55412 -34652
rect 53942 -35212 54718 -35178
rect 53942 -35390 54718 -35356
rect 55820 -35316 55854 -34540
rect 55998 -35316 56032 -34540
rect 53464 -36384 53498 -35608
rect 53642 -36384 53676 -35608
rect 53942 -35618 54718 -35584
rect 53942 -35796 54718 -35762
rect 55280 -36324 55314 -36148
rect 55368 -36324 55402 -36148
rect 55820 -36430 55854 -35654
rect 55998 -36430 56032 -35654
rect 57131 -34934 57165 -34900
rect 57217 -34947 57251 -34913
rect 57303 -34917 57337 -34883
rect 59958 -34808 60334 -34774
rect 59958 -34916 60334 -34882
rect 59502 -35358 59536 -35182
rect 59590 -35358 59624 -35182
rect 59818 -35358 59852 -35182
rect 59906 -35358 59940 -35182
rect 60203 -35407 60237 -35373
rect 61215 -35407 61249 -35373
rect 60211 -35491 60245 -35457
rect 61207 -35491 61241 -35457
rect 57131 -36088 57165 -36054
rect 57217 -36075 57251 -36041
rect 57303 -36105 57337 -36071
rect 59501 -35871 59535 -35695
rect 59589 -35871 59623 -35695
rect 60203 -35575 60237 -35541
rect 61215 -35575 61249 -35541
rect 59817 -35871 59851 -35695
rect 59905 -35871 59939 -35695
rect 60211 -35659 60245 -35625
rect 61207 -35659 61241 -35625
rect 60204 -35743 60238 -35709
rect 61214 -35743 61248 -35709
rect 59958 -36174 60334 -36140
rect 59958 -36282 60334 -36248
rect 55300 -36992 55476 -36958
rect 55300 -37080 55476 -37046
rect 75582 -38485 75616 -38451
rect 75582 -38553 75616 -38519
rect 75666 -38485 75700 -38451
rect 75666 -38553 75700 -38519
rect 75858 -38485 75892 -38451
rect 75858 -38553 75892 -38519
rect 75942 -38485 75976 -38451
rect 75942 -38553 75976 -38519
rect 76132 -38485 76166 -38451
rect 76132 -38553 76166 -38519
rect 76216 -38485 76250 -38451
rect 76216 -38553 76250 -38519
rect 76408 -38485 76442 -38451
rect 76408 -38553 76442 -38519
rect 76492 -38485 76526 -38451
rect 76492 -38553 76526 -38519
rect 76684 -38485 76718 -38451
rect 76684 -38553 76718 -38519
rect 76768 -38485 76802 -38451
rect 76768 -38553 76802 -38519
rect 77613 -39519 77647 -39485
rect 77703 -39525 77737 -39491
rect 77793 -39539 77827 -39505
rect 77877 -39525 77911 -39491
rect 77971 -39539 78005 -39505
rect 78059 -39501 78093 -39467
rect 78167 -39525 78201 -39491
rect 78251 -39539 78285 -39505
rect 78335 -39525 78369 -39491
rect 78429 -39539 78463 -39505
rect 78517 -39501 78551 -39467
rect 78661 -39515 78695 -39481
rect 78853 -39543 78887 -39509
rect 78937 -39543 78971 -39509
rect 80814 -39521 80848 -39487
rect 80814 -39589 80848 -39555
rect 80898 -39521 80932 -39487
rect 80898 -39589 80932 -39555
rect 81059 -39593 81093 -39559
rect 81143 -39585 81177 -39551
rect 81227 -39593 81261 -39559
rect 81311 -39585 81345 -39551
rect 81395 -39592 81429 -39558
rect 81522 -39525 81556 -39491
rect 81522 -39593 81556 -39559
rect 81606 -39525 81640 -39491
rect 81606 -39593 81640 -39559
rect 81690 -39593 81724 -39559
rect 81774 -39525 81808 -39491
rect 81774 -39593 81808 -39559
rect 81858 -39593 81892 -39559
rect 81942 -39525 81976 -39491
rect 81942 -39593 81976 -39559
rect 82026 -39593 82060 -39559
rect 82110 -39525 82144 -39491
rect 82110 -39593 82144 -39559
rect 82194 -39593 82228 -39559
rect 82278 -39525 82312 -39491
rect 82278 -39593 82312 -39559
rect 82362 -39593 82396 -39559
rect 82446 -39525 82480 -39491
rect 82446 -39593 82480 -39559
rect 82530 -39593 82564 -39559
rect 82614 -39525 82648 -39491
rect 82614 -39593 82648 -39559
rect 82698 -39593 82732 -39559
rect 82782 -39525 82816 -39491
rect 82782 -39593 82816 -39559
rect 82866 -39525 82900 -39491
rect 82866 -39593 82900 -39559
rect 82994 -39525 83028 -39491
rect 82994 -39593 83028 -39559
rect 83078 -39525 83112 -39491
rect 83078 -39593 83112 -39559
rect 83162 -39593 83196 -39559
rect 83246 -39525 83280 -39491
rect 83246 -39593 83280 -39559
rect 83330 -39593 83364 -39559
rect 83414 -39525 83448 -39491
rect 83414 -39593 83448 -39559
rect 83498 -39593 83532 -39559
rect 83582 -39525 83616 -39491
rect 83582 -39593 83616 -39559
rect 83666 -39593 83700 -39559
rect 83750 -39525 83784 -39491
rect 83750 -39593 83784 -39559
rect 83834 -39593 83868 -39559
rect 83918 -39525 83952 -39491
rect 83918 -39593 83952 -39559
rect 84002 -39593 84036 -39559
rect 84086 -39525 84120 -39491
rect 84086 -39593 84120 -39559
rect 84170 -39593 84204 -39559
rect 84254 -39525 84288 -39491
rect 84254 -39593 84288 -39559
rect 84338 -39525 84372 -39491
rect 84338 -39593 84372 -39559
rect 84466 -39525 84500 -39491
rect 84466 -39593 84500 -39559
rect 84550 -39525 84584 -39491
rect 84550 -39593 84584 -39559
rect 84634 -39593 84668 -39559
rect 84718 -39525 84752 -39491
rect 84718 -39593 84752 -39559
rect 84802 -39593 84836 -39559
rect 84886 -39525 84920 -39491
rect 84886 -39593 84920 -39559
rect 84970 -39593 85004 -39559
rect 85054 -39525 85088 -39491
rect 85054 -39593 85088 -39559
rect 85138 -39593 85172 -39559
rect 85222 -39525 85256 -39491
rect 85222 -39593 85256 -39559
rect 85306 -39593 85340 -39559
rect 85390 -39525 85424 -39491
rect 85390 -39593 85424 -39559
rect 85474 -39593 85508 -39559
rect 85558 -39525 85592 -39491
rect 85558 -39593 85592 -39559
rect 85642 -39593 85676 -39559
rect 85726 -39525 85760 -39491
rect 85726 -39593 85760 -39559
rect 85810 -39525 85844 -39491
rect 85810 -39593 85844 -39559
rect 85938 -39525 85972 -39491
rect 85938 -39593 85972 -39559
rect 86022 -39525 86056 -39491
rect 86022 -39593 86056 -39559
rect 86106 -39593 86140 -39559
rect 86190 -39525 86224 -39491
rect 86190 -39593 86224 -39559
rect 86274 -39593 86308 -39559
rect 86358 -39525 86392 -39491
rect 86358 -39593 86392 -39559
rect 86442 -39593 86476 -39559
rect 86526 -39525 86560 -39491
rect 86526 -39593 86560 -39559
rect 86610 -39593 86644 -39559
rect 86694 -39525 86728 -39491
rect 86694 -39593 86728 -39559
rect 86778 -39593 86812 -39559
rect 86862 -39525 86896 -39491
rect 86862 -39593 86896 -39559
rect 86946 -39593 86980 -39559
rect 87030 -39525 87064 -39491
rect 87030 -39593 87064 -39559
rect 87114 -39593 87148 -39559
rect 87198 -39525 87232 -39491
rect 87198 -39593 87232 -39559
rect 87282 -39525 87316 -39491
rect 87282 -39593 87316 -39559
rect 87410 -39525 87444 -39491
rect 87410 -39593 87444 -39559
rect 87494 -39525 87528 -39491
rect 87494 -39593 87528 -39559
rect 87578 -39593 87612 -39559
rect 87662 -39525 87696 -39491
rect 87662 -39593 87696 -39559
rect 87746 -39593 87780 -39559
rect 87830 -39525 87864 -39491
rect 87830 -39593 87864 -39559
rect 87914 -39593 87948 -39559
rect 87998 -39525 88032 -39491
rect 87998 -39593 88032 -39559
rect 88082 -39593 88116 -39559
rect 88166 -39525 88200 -39491
rect 88166 -39593 88200 -39559
rect 88250 -39593 88284 -39559
rect 88334 -39525 88368 -39491
rect 88334 -39593 88368 -39559
rect 88418 -39593 88452 -39559
rect 88502 -39525 88536 -39491
rect 88502 -39593 88536 -39559
rect 88586 -39593 88620 -39559
rect 88670 -39525 88704 -39491
rect 88670 -39593 88704 -39559
rect 88754 -39525 88788 -39491
rect 88754 -39593 88788 -39559
rect 53464 -40766 53498 -39990
rect 53642 -40766 53676 -39990
rect 55290 -40228 55324 -40052
rect 55378 -40228 55412 -40052
rect 53942 -40612 54718 -40578
rect 53942 -40790 54718 -40756
rect 55820 -40716 55854 -39940
rect 55998 -40716 56032 -39940
rect 77613 -39805 77647 -39771
rect 77703 -39799 77737 -39765
rect 77793 -39785 77827 -39751
rect 77877 -39799 77911 -39765
rect 77971 -39785 78005 -39751
rect 78059 -39823 78093 -39789
rect 80864 -39825 80898 -39791
rect 80864 -39893 80898 -39859
rect 80948 -39825 80982 -39791
rect 80948 -39893 80982 -39859
rect 53464 -41784 53498 -41008
rect 53642 -41784 53676 -41008
rect 53942 -41018 54718 -40984
rect 53942 -41196 54718 -41162
rect 55280 -41724 55314 -41548
rect 55368 -41724 55402 -41548
rect 55820 -41830 55854 -41054
rect 55998 -41830 56032 -41054
rect 57131 -40334 57165 -40300
rect 57217 -40347 57251 -40313
rect 57303 -40317 57337 -40283
rect 59958 -40208 60334 -40174
rect 59958 -40316 60334 -40282
rect 59502 -40758 59536 -40582
rect 59590 -40758 59624 -40582
rect 59818 -40758 59852 -40582
rect 59906 -40758 59940 -40582
rect 60203 -40807 60237 -40773
rect 61215 -40807 61249 -40773
rect 77649 -40765 77683 -40731
rect 77841 -40793 77875 -40759
rect 77925 -40793 77959 -40759
rect 60211 -40891 60245 -40857
rect 61207 -40891 61241 -40857
rect 57131 -41488 57165 -41454
rect 57217 -41475 57251 -41441
rect 57303 -41505 57337 -41471
rect 59501 -41271 59535 -41095
rect 59589 -41271 59623 -41095
rect 60203 -40975 60237 -40941
rect 61215 -40975 61249 -40941
rect 59817 -41271 59851 -41095
rect 59905 -41271 59939 -41095
rect 60211 -41059 60245 -41025
rect 61207 -41059 61241 -41025
rect 77649 -41049 77683 -41015
rect 77841 -41021 77875 -40987
rect 60204 -41143 60238 -41109
rect 61214 -41143 61248 -41109
rect 77925 -41021 77959 -40987
rect 78073 -41045 78107 -41011
rect 78163 -41039 78197 -41005
rect 78253 -41025 78287 -40991
rect 78337 -41039 78371 -41005
rect 78431 -41025 78465 -40991
rect 78519 -41063 78553 -41029
rect 59958 -41574 60334 -41540
rect 59958 -41682 60334 -41648
rect 77649 -42005 77683 -41971
rect 77841 -42033 77875 -41999
rect 77925 -42033 77959 -41999
rect 55300 -42392 55476 -42358
rect 55300 -42480 55476 -42446
rect 77651 -42303 77685 -42269
rect 77843 -42275 77877 -42241
rect 77927 -42275 77961 -42241
rect 77613 -43275 77647 -43241
rect 78054 -43215 78088 -43181
rect 78054 -43283 78088 -43249
rect 78153 -43215 78187 -43181
rect 78153 -43283 78187 -43249
rect 78357 -43259 78391 -43225
rect 78447 -43265 78481 -43231
rect 78537 -43279 78571 -43245
rect 78621 -43265 78655 -43231
rect 78715 -43279 78749 -43245
rect 78803 -43241 78837 -43207
rect 77613 -43515 77647 -43481
rect 78054 -43507 78088 -43473
rect 78054 -43575 78088 -43541
rect 78153 -43507 78187 -43473
rect 78153 -43575 78187 -43541
rect 82902 -44083 82936 -44049
rect 82986 -44083 83020 -44049
rect 83082 -44083 83116 -44049
rect 83167 -44023 83201 -43989
rect 83167 -44091 83201 -44057
rect 83374 -44021 83408 -43987
rect 83374 -44089 83408 -44055
rect 83458 -44021 83492 -43987
rect 83458 -44089 83492 -44055
rect 83619 -44093 83653 -44059
rect 83703 -44085 83737 -44051
rect 83787 -44093 83821 -44059
rect 83871 -44085 83905 -44051
rect 83955 -44092 83989 -44058
rect 84082 -44025 84116 -43991
rect 84082 -44093 84116 -44059
rect 84166 -44025 84200 -43991
rect 84166 -44093 84200 -44059
rect 84250 -44093 84284 -44059
rect 84334 -44025 84368 -43991
rect 84334 -44093 84368 -44059
rect 84418 -44093 84452 -44059
rect 84502 -44025 84536 -43991
rect 84502 -44093 84536 -44059
rect 84586 -44093 84620 -44059
rect 84670 -44025 84704 -43991
rect 84670 -44093 84704 -44059
rect 84754 -44093 84788 -44059
rect 84838 -44025 84872 -43991
rect 84838 -44093 84872 -44059
rect 84922 -44093 84956 -44059
rect 85006 -44025 85040 -43991
rect 85006 -44093 85040 -44059
rect 85090 -44093 85124 -44059
rect 85174 -44025 85208 -43991
rect 85174 -44093 85208 -44059
rect 85258 -44093 85292 -44059
rect 85342 -44025 85376 -43991
rect 85342 -44093 85376 -44059
rect 85426 -44025 85460 -43991
rect 85426 -44093 85460 -44059
rect 85554 -44025 85588 -43991
rect 85554 -44093 85588 -44059
rect 85638 -44025 85672 -43991
rect 85638 -44093 85672 -44059
rect 85722 -44093 85756 -44059
rect 85806 -44025 85840 -43991
rect 85806 -44093 85840 -44059
rect 85890 -44093 85924 -44059
rect 85974 -44025 86008 -43991
rect 85974 -44093 86008 -44059
rect 86058 -44093 86092 -44059
rect 86142 -44025 86176 -43991
rect 86142 -44093 86176 -44059
rect 86226 -44093 86260 -44059
rect 86310 -44025 86344 -43991
rect 86310 -44093 86344 -44059
rect 86394 -44093 86428 -44059
rect 86478 -44025 86512 -43991
rect 86478 -44093 86512 -44059
rect 86562 -44093 86596 -44059
rect 86646 -44025 86680 -43991
rect 86646 -44093 86680 -44059
rect 86730 -44093 86764 -44059
rect 86814 -44025 86848 -43991
rect 86814 -44093 86848 -44059
rect 86898 -44025 86932 -43991
rect 86898 -44093 86932 -44059
rect 87026 -44025 87060 -43991
rect 87026 -44093 87060 -44059
rect 87110 -44025 87144 -43991
rect 87110 -44093 87144 -44059
rect 87194 -44093 87228 -44059
rect 87278 -44025 87312 -43991
rect 87278 -44093 87312 -44059
rect 87362 -44093 87396 -44059
rect 87446 -44025 87480 -43991
rect 87446 -44093 87480 -44059
rect 87530 -44093 87564 -44059
rect 87614 -44025 87648 -43991
rect 87614 -44093 87648 -44059
rect 87698 -44093 87732 -44059
rect 87782 -44025 87816 -43991
rect 87782 -44093 87816 -44059
rect 87866 -44093 87900 -44059
rect 87950 -44025 87984 -43991
rect 87950 -44093 87984 -44059
rect 88034 -44093 88068 -44059
rect 88118 -44025 88152 -43991
rect 88118 -44093 88152 -44059
rect 88202 -44093 88236 -44059
rect 88286 -44025 88320 -43991
rect 88286 -44093 88320 -44059
rect 88370 -44025 88404 -43991
rect 88370 -44093 88404 -44059
rect 88498 -44025 88532 -43991
rect 88498 -44093 88532 -44059
rect 88582 -44025 88616 -43991
rect 88582 -44093 88616 -44059
rect 88666 -44093 88700 -44059
rect 88750 -44025 88784 -43991
rect 88750 -44093 88784 -44059
rect 88834 -44093 88868 -44059
rect 88918 -44025 88952 -43991
rect 88918 -44093 88952 -44059
rect 89002 -44093 89036 -44059
rect 89086 -44025 89120 -43991
rect 89086 -44093 89120 -44059
rect 89170 -44093 89204 -44059
rect 89254 -44025 89288 -43991
rect 89254 -44093 89288 -44059
rect 89338 -44093 89372 -44059
rect 89422 -44025 89456 -43991
rect 89422 -44093 89456 -44059
rect 89506 -44093 89540 -44059
rect 89590 -44025 89624 -43991
rect 89590 -44093 89624 -44059
rect 89674 -44093 89708 -44059
rect 89758 -44025 89792 -43991
rect 89758 -44093 89792 -44059
rect 89842 -44025 89876 -43991
rect 89842 -44093 89876 -44059
rect 89970 -44025 90004 -43991
rect 89970 -44093 90004 -44059
rect 90054 -44025 90088 -43991
rect 90054 -44093 90088 -44059
rect 90138 -44093 90172 -44059
rect 90222 -44025 90256 -43991
rect 90222 -44093 90256 -44059
rect 90306 -44093 90340 -44059
rect 90390 -44025 90424 -43991
rect 90390 -44093 90424 -44059
rect 90474 -44093 90508 -44059
rect 90558 -44025 90592 -43991
rect 90558 -44093 90592 -44059
rect 90642 -44093 90676 -44059
rect 90726 -44025 90760 -43991
rect 90726 -44093 90760 -44059
rect 90810 -44093 90844 -44059
rect 90894 -44025 90928 -43991
rect 90894 -44093 90928 -44059
rect 90978 -44093 91012 -44059
rect 91062 -44025 91096 -43991
rect 91062 -44093 91096 -44059
rect 91146 -44093 91180 -44059
rect 91230 -44025 91264 -43991
rect 91230 -44093 91264 -44059
rect 91314 -44025 91348 -43991
rect 91314 -44093 91348 -44059
rect 77613 -44507 77647 -44473
rect 78054 -44447 78088 -44413
rect 78054 -44515 78088 -44481
rect 78153 -44447 78187 -44413
rect 78153 -44515 78187 -44481
rect 77613 -44749 77647 -44715
rect 78054 -44741 78088 -44707
rect 78054 -44809 78088 -44775
rect 78153 -44741 78187 -44707
rect 78153 -44809 78187 -44775
rect 53464 -46166 53498 -45390
rect 53642 -46166 53676 -45390
rect 55290 -45628 55324 -45452
rect 55378 -45628 55412 -45452
rect 53942 -46012 54718 -45978
rect 53942 -46190 54718 -46156
rect 55820 -46116 55854 -45340
rect 55998 -46116 56032 -45340
rect 53464 -47184 53498 -46408
rect 53642 -47184 53676 -46408
rect 53942 -46418 54718 -46384
rect 53942 -46596 54718 -46562
rect 55280 -47124 55314 -46948
rect 55368 -47124 55402 -46948
rect 55820 -47230 55854 -46454
rect 55998 -47230 56032 -46454
rect 57131 -45734 57165 -45700
rect 57217 -45747 57251 -45713
rect 57303 -45717 57337 -45683
rect 59958 -45608 60334 -45574
rect 59958 -45716 60334 -45682
rect 77613 -45753 77647 -45719
rect 77885 -45737 77919 -45703
rect 77969 -45727 78003 -45693
rect 78109 -45725 78143 -45691
rect 78301 -45753 78335 -45719
rect 78385 -45753 78419 -45719
rect 78533 -45729 78567 -45695
rect 78623 -45735 78657 -45701
rect 78713 -45749 78747 -45715
rect 78797 -45735 78831 -45701
rect 78891 -45749 78925 -45715
rect 78979 -45711 79013 -45677
rect 59502 -46158 59536 -45982
rect 59590 -46158 59624 -45982
rect 59818 -46158 59852 -45982
rect 59906 -46158 59940 -45982
rect 60203 -46207 60237 -46173
rect 61215 -46207 61249 -46173
rect 60211 -46291 60245 -46257
rect 61207 -46291 61241 -46257
rect 57131 -46888 57165 -46854
rect 57217 -46875 57251 -46841
rect 57303 -46905 57337 -46871
rect 59501 -46671 59535 -46495
rect 59589 -46671 59623 -46495
rect 60203 -46375 60237 -46341
rect 61215 -46375 61249 -46341
rect 59817 -46671 59851 -46495
rect 59905 -46671 59939 -46495
rect 60211 -46459 60245 -46425
rect 61207 -46459 61241 -46425
rect 60204 -46543 60238 -46509
rect 61214 -46543 61248 -46509
rect 75582 -46525 75616 -46491
rect 75582 -46593 75616 -46559
rect 75666 -46525 75700 -46491
rect 75666 -46593 75700 -46559
rect 75858 -46525 75892 -46491
rect 75858 -46593 75892 -46559
rect 75942 -46525 75976 -46491
rect 75942 -46593 75976 -46559
rect 76132 -46525 76166 -46491
rect 76132 -46593 76166 -46559
rect 76216 -46525 76250 -46491
rect 76216 -46593 76250 -46559
rect 76408 -46525 76442 -46491
rect 76408 -46593 76442 -46559
rect 76492 -46525 76526 -46491
rect 76492 -46593 76526 -46559
rect 76684 -46525 76718 -46491
rect 76684 -46593 76718 -46559
rect 76768 -46525 76802 -46491
rect 76768 -46593 76802 -46559
rect 59958 -46974 60334 -46940
rect 59958 -47082 60334 -47048
rect 77613 -47559 77647 -47525
rect 77703 -47565 77737 -47531
rect 77793 -47579 77827 -47545
rect 77877 -47565 77911 -47531
rect 77971 -47579 78005 -47545
rect 78059 -47541 78093 -47507
rect 78167 -47565 78201 -47531
rect 78251 -47579 78285 -47545
rect 78335 -47565 78369 -47531
rect 78429 -47579 78463 -47545
rect 78517 -47541 78551 -47507
rect 78661 -47555 78695 -47521
rect 78853 -47583 78887 -47549
rect 78937 -47583 78971 -47549
rect 55300 -47792 55476 -47758
rect 55300 -47880 55476 -47846
rect 77613 -47845 77647 -47811
rect 77703 -47839 77737 -47805
rect 77793 -47825 77827 -47791
rect 77877 -47839 77911 -47805
rect 77971 -47825 78005 -47791
rect 78059 -47863 78093 -47829
rect 82902 -48223 82936 -48189
rect 82986 -48223 83020 -48189
rect 83082 -48223 83116 -48189
rect 83167 -48163 83201 -48129
rect 83167 -48231 83201 -48197
rect 83374 -48161 83408 -48127
rect 83374 -48229 83408 -48195
rect 83458 -48161 83492 -48127
rect 83458 -48229 83492 -48195
rect 83619 -48233 83653 -48199
rect 83703 -48225 83737 -48191
rect 83787 -48233 83821 -48199
rect 83871 -48225 83905 -48191
rect 83955 -48232 83989 -48198
rect 84082 -48165 84116 -48131
rect 84082 -48233 84116 -48199
rect 84166 -48165 84200 -48131
rect 84166 -48233 84200 -48199
rect 84250 -48233 84284 -48199
rect 84334 -48165 84368 -48131
rect 84334 -48233 84368 -48199
rect 84418 -48233 84452 -48199
rect 84502 -48165 84536 -48131
rect 84502 -48233 84536 -48199
rect 84586 -48233 84620 -48199
rect 84670 -48165 84704 -48131
rect 84670 -48233 84704 -48199
rect 84754 -48233 84788 -48199
rect 84838 -48165 84872 -48131
rect 84838 -48233 84872 -48199
rect 84922 -48233 84956 -48199
rect 85006 -48165 85040 -48131
rect 85006 -48233 85040 -48199
rect 85090 -48233 85124 -48199
rect 85174 -48165 85208 -48131
rect 85174 -48233 85208 -48199
rect 85258 -48233 85292 -48199
rect 85342 -48165 85376 -48131
rect 85342 -48233 85376 -48199
rect 85426 -48165 85460 -48131
rect 85426 -48233 85460 -48199
rect 85554 -48165 85588 -48131
rect 85554 -48233 85588 -48199
rect 85638 -48165 85672 -48131
rect 85638 -48233 85672 -48199
rect 85722 -48233 85756 -48199
rect 85806 -48165 85840 -48131
rect 85806 -48233 85840 -48199
rect 85890 -48233 85924 -48199
rect 85974 -48165 86008 -48131
rect 85974 -48233 86008 -48199
rect 86058 -48233 86092 -48199
rect 86142 -48165 86176 -48131
rect 86142 -48233 86176 -48199
rect 86226 -48233 86260 -48199
rect 86310 -48165 86344 -48131
rect 86310 -48233 86344 -48199
rect 86394 -48233 86428 -48199
rect 86478 -48165 86512 -48131
rect 86478 -48233 86512 -48199
rect 86562 -48233 86596 -48199
rect 86646 -48165 86680 -48131
rect 86646 -48233 86680 -48199
rect 86730 -48233 86764 -48199
rect 86814 -48165 86848 -48131
rect 86814 -48233 86848 -48199
rect 86898 -48165 86932 -48131
rect 86898 -48233 86932 -48199
rect 87026 -48165 87060 -48131
rect 87026 -48233 87060 -48199
rect 87110 -48165 87144 -48131
rect 87110 -48233 87144 -48199
rect 87194 -48233 87228 -48199
rect 87278 -48165 87312 -48131
rect 87278 -48233 87312 -48199
rect 87362 -48233 87396 -48199
rect 87446 -48165 87480 -48131
rect 87446 -48233 87480 -48199
rect 87530 -48233 87564 -48199
rect 87614 -48165 87648 -48131
rect 87614 -48233 87648 -48199
rect 87698 -48233 87732 -48199
rect 87782 -48165 87816 -48131
rect 87782 -48233 87816 -48199
rect 87866 -48233 87900 -48199
rect 87950 -48165 87984 -48131
rect 87950 -48233 87984 -48199
rect 88034 -48233 88068 -48199
rect 88118 -48165 88152 -48131
rect 88118 -48233 88152 -48199
rect 88202 -48233 88236 -48199
rect 88286 -48165 88320 -48131
rect 88286 -48233 88320 -48199
rect 88370 -48165 88404 -48131
rect 88370 -48233 88404 -48199
rect 88498 -48165 88532 -48131
rect 88498 -48233 88532 -48199
rect 88582 -48165 88616 -48131
rect 88582 -48233 88616 -48199
rect 88666 -48233 88700 -48199
rect 88750 -48165 88784 -48131
rect 88750 -48233 88784 -48199
rect 88834 -48233 88868 -48199
rect 88918 -48165 88952 -48131
rect 88918 -48233 88952 -48199
rect 89002 -48233 89036 -48199
rect 89086 -48165 89120 -48131
rect 89086 -48233 89120 -48199
rect 89170 -48233 89204 -48199
rect 89254 -48165 89288 -48131
rect 89254 -48233 89288 -48199
rect 89338 -48233 89372 -48199
rect 89422 -48165 89456 -48131
rect 89422 -48233 89456 -48199
rect 89506 -48233 89540 -48199
rect 89590 -48165 89624 -48131
rect 89590 -48233 89624 -48199
rect 89674 -48233 89708 -48199
rect 89758 -48165 89792 -48131
rect 89758 -48233 89792 -48199
rect 89842 -48165 89876 -48131
rect 89842 -48233 89876 -48199
rect 89970 -48165 90004 -48131
rect 89970 -48233 90004 -48199
rect 90054 -48165 90088 -48131
rect 90054 -48233 90088 -48199
rect 90138 -48233 90172 -48199
rect 90222 -48165 90256 -48131
rect 90222 -48233 90256 -48199
rect 90306 -48233 90340 -48199
rect 90390 -48165 90424 -48131
rect 90390 -48233 90424 -48199
rect 90474 -48233 90508 -48199
rect 90558 -48165 90592 -48131
rect 90558 -48233 90592 -48199
rect 90642 -48233 90676 -48199
rect 90726 -48165 90760 -48131
rect 90726 -48233 90760 -48199
rect 90810 -48233 90844 -48199
rect 90894 -48165 90928 -48131
rect 90894 -48233 90928 -48199
rect 90978 -48233 91012 -48199
rect 91062 -48165 91096 -48131
rect 91062 -48233 91096 -48199
rect 91146 -48233 91180 -48199
rect 91230 -48165 91264 -48131
rect 91230 -48233 91264 -48199
rect 91314 -48165 91348 -48131
rect 91314 -48233 91348 -48199
rect 77649 -48805 77683 -48771
rect 77841 -48833 77875 -48799
rect 77925 -48833 77959 -48799
rect 77649 -49089 77683 -49055
rect 77841 -49061 77875 -49027
rect 77925 -49061 77959 -49027
rect 78073 -49085 78107 -49051
rect 78163 -49079 78197 -49045
rect 78253 -49065 78287 -49031
rect 78337 -49079 78371 -49045
rect 78431 -49065 78465 -49031
rect 78519 -49103 78553 -49069
rect 77649 -50045 77683 -50011
rect 77841 -50073 77875 -50039
rect 77925 -50073 77959 -50039
rect 77651 -50343 77685 -50309
rect 77843 -50315 77877 -50281
rect 53464 -51566 53498 -50790
rect 53642 -51566 53676 -50790
rect 55290 -51028 55324 -50852
rect 55378 -51028 55412 -50852
rect 53942 -51412 54718 -51378
rect 53942 -51590 54718 -51556
rect 55820 -51516 55854 -50740
rect 55998 -51516 56032 -50740
rect 77927 -50315 77961 -50281
rect 53464 -52584 53498 -51808
rect 53642 -52584 53676 -51808
rect 53942 -51818 54718 -51784
rect 53942 -51996 54718 -51962
rect 55280 -52524 55314 -52348
rect 55368 -52524 55402 -52348
rect 55820 -52630 55854 -51854
rect 55998 -52630 56032 -51854
rect 57131 -51134 57165 -51100
rect 57217 -51147 57251 -51113
rect 57303 -51117 57337 -51083
rect 59958 -51008 60334 -50974
rect 59958 -51116 60334 -51082
rect 59502 -51558 59536 -51382
rect 59590 -51558 59624 -51382
rect 59818 -51558 59852 -51382
rect 59906 -51558 59940 -51382
rect 77613 -51315 77647 -51281
rect 78054 -51255 78088 -51221
rect 78054 -51323 78088 -51289
rect 78153 -51255 78187 -51221
rect 78153 -51323 78187 -51289
rect 78357 -51299 78391 -51265
rect 78447 -51305 78481 -51271
rect 78537 -51319 78571 -51285
rect 78621 -51305 78655 -51271
rect 78715 -51319 78749 -51285
rect 78803 -51281 78837 -51247
rect 77613 -51555 77647 -51521
rect 60203 -51607 60237 -51573
rect 61215 -51607 61249 -51573
rect 78054 -51547 78088 -51513
rect 60211 -51691 60245 -51657
rect 61207 -51691 61241 -51657
rect 57131 -52288 57165 -52254
rect 57217 -52275 57251 -52241
rect 57303 -52305 57337 -52271
rect 78054 -51615 78088 -51581
rect 78153 -51547 78187 -51513
rect 78153 -51615 78187 -51581
rect 59501 -52071 59535 -51895
rect 59589 -52071 59623 -51895
rect 60203 -51775 60237 -51741
rect 61215 -51775 61249 -51741
rect 59817 -52071 59851 -51895
rect 59905 -52071 59939 -51895
rect 60211 -51859 60245 -51825
rect 61207 -51859 61241 -51825
rect 60204 -51943 60238 -51909
rect 61214 -51943 61248 -51909
rect 82902 -51873 82936 -51839
rect 82986 -51873 83020 -51839
rect 83082 -51873 83116 -51839
rect 83167 -51813 83201 -51779
rect 83167 -51881 83201 -51847
rect 83374 -51811 83408 -51777
rect 83374 -51879 83408 -51845
rect 83458 -51811 83492 -51777
rect 83458 -51879 83492 -51845
rect 83619 -51883 83653 -51849
rect 83703 -51875 83737 -51841
rect 83787 -51883 83821 -51849
rect 83871 -51875 83905 -51841
rect 83955 -51882 83989 -51848
rect 84082 -51815 84116 -51781
rect 84082 -51883 84116 -51849
rect 84166 -51815 84200 -51781
rect 84166 -51883 84200 -51849
rect 84250 -51883 84284 -51849
rect 84334 -51815 84368 -51781
rect 84334 -51883 84368 -51849
rect 84418 -51883 84452 -51849
rect 84502 -51815 84536 -51781
rect 84502 -51883 84536 -51849
rect 84586 -51883 84620 -51849
rect 84670 -51815 84704 -51781
rect 84670 -51883 84704 -51849
rect 84754 -51883 84788 -51849
rect 84838 -51815 84872 -51781
rect 84838 -51883 84872 -51849
rect 84922 -51883 84956 -51849
rect 85006 -51815 85040 -51781
rect 85006 -51883 85040 -51849
rect 85090 -51883 85124 -51849
rect 85174 -51815 85208 -51781
rect 85174 -51883 85208 -51849
rect 85258 -51883 85292 -51849
rect 85342 -51815 85376 -51781
rect 85342 -51883 85376 -51849
rect 85426 -51815 85460 -51781
rect 85426 -51883 85460 -51849
rect 85554 -51815 85588 -51781
rect 85554 -51883 85588 -51849
rect 85638 -51815 85672 -51781
rect 85638 -51883 85672 -51849
rect 85722 -51883 85756 -51849
rect 85806 -51815 85840 -51781
rect 85806 -51883 85840 -51849
rect 85890 -51883 85924 -51849
rect 85974 -51815 86008 -51781
rect 85974 -51883 86008 -51849
rect 86058 -51883 86092 -51849
rect 86142 -51815 86176 -51781
rect 86142 -51883 86176 -51849
rect 86226 -51883 86260 -51849
rect 86310 -51815 86344 -51781
rect 86310 -51883 86344 -51849
rect 86394 -51883 86428 -51849
rect 86478 -51815 86512 -51781
rect 86478 -51883 86512 -51849
rect 86562 -51883 86596 -51849
rect 86646 -51815 86680 -51781
rect 86646 -51883 86680 -51849
rect 86730 -51883 86764 -51849
rect 86814 -51815 86848 -51781
rect 86814 -51883 86848 -51849
rect 86898 -51815 86932 -51781
rect 86898 -51883 86932 -51849
rect 87026 -51815 87060 -51781
rect 87026 -51883 87060 -51849
rect 87110 -51815 87144 -51781
rect 87110 -51883 87144 -51849
rect 87194 -51883 87228 -51849
rect 87278 -51815 87312 -51781
rect 87278 -51883 87312 -51849
rect 87362 -51883 87396 -51849
rect 87446 -51815 87480 -51781
rect 87446 -51883 87480 -51849
rect 87530 -51883 87564 -51849
rect 87614 -51815 87648 -51781
rect 87614 -51883 87648 -51849
rect 87698 -51883 87732 -51849
rect 87782 -51815 87816 -51781
rect 87782 -51883 87816 -51849
rect 87866 -51883 87900 -51849
rect 87950 -51815 87984 -51781
rect 87950 -51883 87984 -51849
rect 88034 -51883 88068 -51849
rect 88118 -51815 88152 -51781
rect 88118 -51883 88152 -51849
rect 88202 -51883 88236 -51849
rect 88286 -51815 88320 -51781
rect 88286 -51883 88320 -51849
rect 88370 -51815 88404 -51781
rect 88370 -51883 88404 -51849
rect 88498 -51815 88532 -51781
rect 88498 -51883 88532 -51849
rect 88582 -51815 88616 -51781
rect 88582 -51883 88616 -51849
rect 88666 -51883 88700 -51849
rect 88750 -51815 88784 -51781
rect 88750 -51883 88784 -51849
rect 88834 -51883 88868 -51849
rect 88918 -51815 88952 -51781
rect 88918 -51883 88952 -51849
rect 89002 -51883 89036 -51849
rect 89086 -51815 89120 -51781
rect 89086 -51883 89120 -51849
rect 89170 -51883 89204 -51849
rect 89254 -51815 89288 -51781
rect 89254 -51883 89288 -51849
rect 89338 -51883 89372 -51849
rect 89422 -51815 89456 -51781
rect 89422 -51883 89456 -51849
rect 89506 -51883 89540 -51849
rect 89590 -51815 89624 -51781
rect 89590 -51883 89624 -51849
rect 89674 -51883 89708 -51849
rect 89758 -51815 89792 -51781
rect 89758 -51883 89792 -51849
rect 89842 -51815 89876 -51781
rect 89842 -51883 89876 -51849
rect 89970 -51815 90004 -51781
rect 89970 -51883 90004 -51849
rect 90054 -51815 90088 -51781
rect 90054 -51883 90088 -51849
rect 90138 -51883 90172 -51849
rect 90222 -51815 90256 -51781
rect 90222 -51883 90256 -51849
rect 90306 -51883 90340 -51849
rect 90390 -51815 90424 -51781
rect 90390 -51883 90424 -51849
rect 90474 -51883 90508 -51849
rect 90558 -51815 90592 -51781
rect 90558 -51883 90592 -51849
rect 90642 -51883 90676 -51849
rect 90726 -51815 90760 -51781
rect 90726 -51883 90760 -51849
rect 90810 -51883 90844 -51849
rect 90894 -51815 90928 -51781
rect 90894 -51883 90928 -51849
rect 90978 -51883 91012 -51849
rect 91062 -51815 91096 -51781
rect 91062 -51883 91096 -51849
rect 91146 -51883 91180 -51849
rect 91230 -51815 91264 -51781
rect 91230 -51883 91264 -51849
rect 91314 -51815 91348 -51781
rect 91314 -51883 91348 -51849
rect 59958 -52374 60334 -52340
rect 59958 -52482 60334 -52448
rect 77613 -52547 77647 -52513
rect 78054 -52487 78088 -52453
rect 78054 -52555 78088 -52521
rect 78153 -52487 78187 -52453
rect 78153 -52555 78187 -52521
rect 77613 -52789 77647 -52755
rect 78054 -52781 78088 -52747
rect 78054 -52849 78088 -52815
rect 78153 -52781 78187 -52747
rect 78153 -52849 78187 -52815
rect 55300 -53192 55476 -53158
rect 55300 -53280 55476 -53246
rect 77613 -53793 77647 -53759
rect 77885 -53777 77919 -53743
rect 77969 -53767 78003 -53733
rect 78109 -53765 78143 -53731
rect 78301 -53793 78335 -53759
rect 78385 -53793 78419 -53759
rect 78533 -53769 78567 -53735
rect 78623 -53775 78657 -53741
rect 78713 -53789 78747 -53755
rect 78797 -53775 78831 -53741
rect 78891 -53789 78925 -53755
rect 78979 -53751 79013 -53717
rect 53464 -56966 53498 -56190
rect 53642 -56966 53676 -56190
rect 55290 -56428 55324 -56252
rect 55378 -56428 55412 -56252
rect 53942 -56812 54718 -56778
rect 53942 -56990 54718 -56956
rect 55820 -56916 55854 -56140
rect 55998 -56916 56032 -56140
rect 53464 -57984 53498 -57208
rect 53642 -57984 53676 -57208
rect 53942 -57218 54718 -57184
rect 53942 -57396 54718 -57362
rect 55280 -57924 55314 -57748
rect 55368 -57924 55402 -57748
rect 55820 -58030 55854 -57254
rect 55998 -58030 56032 -57254
rect 57131 -56534 57165 -56500
rect 57217 -56547 57251 -56513
rect 57303 -56517 57337 -56483
rect 59958 -56408 60334 -56374
rect 59958 -56516 60334 -56482
rect 59502 -56958 59536 -56782
rect 59590 -56958 59624 -56782
rect 59818 -56958 59852 -56782
rect 59906 -56958 59940 -56782
rect 60203 -57007 60237 -56973
rect 61215 -57007 61249 -56973
rect 60211 -57091 60245 -57057
rect 61207 -57091 61241 -57057
rect 57131 -57688 57165 -57654
rect 57217 -57675 57251 -57641
rect 57303 -57705 57337 -57671
rect 59501 -57471 59535 -57295
rect 59589 -57471 59623 -57295
rect 60203 -57175 60237 -57141
rect 61215 -57175 61249 -57141
rect 59817 -57471 59851 -57295
rect 59905 -57471 59939 -57295
rect 60211 -57259 60245 -57225
rect 61207 -57259 61241 -57225
rect 60204 -57343 60238 -57309
rect 61214 -57343 61248 -57309
rect 59958 -57774 60334 -57740
rect 59958 -57882 60334 -57848
rect 55300 -58592 55476 -58558
rect 55300 -58680 55476 -58646
rect 53464 -62366 53498 -61590
rect 53642 -62366 53676 -61590
rect 55290 -61828 55324 -61652
rect 55378 -61828 55412 -61652
rect 53942 -62212 54718 -62178
rect 53942 -62390 54718 -62356
rect 55820 -62316 55854 -61540
rect 55998 -62316 56032 -61540
rect 53464 -63384 53498 -62608
rect 53642 -63384 53676 -62608
rect 53942 -62618 54718 -62584
rect 53942 -62796 54718 -62762
rect 55280 -63324 55314 -63148
rect 55368 -63324 55402 -63148
rect 55820 -63430 55854 -62654
rect 55998 -63430 56032 -62654
rect 57131 -61934 57165 -61900
rect 57217 -61947 57251 -61913
rect 57303 -61917 57337 -61883
rect 59958 -61808 60334 -61774
rect 59958 -61916 60334 -61882
rect 59502 -62358 59536 -62182
rect 59590 -62358 59624 -62182
rect 59818 -62358 59852 -62182
rect 59906 -62358 59940 -62182
rect 60203 -62407 60237 -62373
rect 61215 -62407 61249 -62373
rect 60211 -62491 60245 -62457
rect 61207 -62491 61241 -62457
rect 57131 -63088 57165 -63054
rect 57217 -63075 57251 -63041
rect 57303 -63105 57337 -63071
rect 59501 -62871 59535 -62695
rect 59589 -62871 59623 -62695
rect 60203 -62575 60237 -62541
rect 61215 -62575 61249 -62541
rect 59817 -62871 59851 -62695
rect 59905 -62871 59939 -62695
rect 60211 -62659 60245 -62625
rect 61207 -62659 61241 -62625
rect 60204 -62743 60238 -62709
rect 61214 -62743 61248 -62709
rect 59958 -63174 60334 -63140
rect 59958 -63282 60334 -63248
rect 55300 -63992 55476 -63958
rect 55300 -64080 55476 -64046
rect 53464 -67766 53498 -66990
rect 53642 -67766 53676 -66990
rect 55290 -67228 55324 -67052
rect 55378 -67228 55412 -67052
rect 53942 -67612 54718 -67578
rect 53942 -67790 54718 -67756
rect 55820 -67716 55854 -66940
rect 55998 -67716 56032 -66940
rect 53464 -68784 53498 -68008
rect 53642 -68784 53676 -68008
rect 53942 -68018 54718 -67984
rect 53942 -68196 54718 -68162
rect 55280 -68724 55314 -68548
rect 55368 -68724 55402 -68548
rect 55820 -68830 55854 -68054
rect 55998 -68830 56032 -68054
rect 57131 -67334 57165 -67300
rect 57217 -67347 57251 -67313
rect 57303 -67317 57337 -67283
rect 59958 -67208 60334 -67174
rect 59958 -67316 60334 -67282
rect 59502 -67758 59536 -67582
rect 59590 -67758 59624 -67582
rect 59818 -67758 59852 -67582
rect 59906 -67758 59940 -67582
rect 60203 -67807 60237 -67773
rect 61215 -67807 61249 -67773
rect 60211 -67891 60245 -67857
rect 61207 -67891 61241 -67857
rect 57131 -68488 57165 -68454
rect 57217 -68475 57251 -68441
rect 57303 -68505 57337 -68471
rect 59501 -68271 59535 -68095
rect 59589 -68271 59623 -68095
rect 60203 -67975 60237 -67941
rect 61215 -67975 61249 -67941
rect 59817 -68271 59851 -68095
rect 59905 -68271 59939 -68095
rect 60211 -68059 60245 -68025
rect 61207 -68059 61241 -68025
rect 60204 -68143 60238 -68109
rect 61214 -68143 61248 -68109
rect 59958 -68574 60334 -68540
rect 59958 -68682 60334 -68648
rect 55300 -69392 55476 -69358
rect 55300 -69480 55476 -69446
rect 53464 -73166 53498 -72390
rect 53642 -73166 53676 -72390
rect 55290 -72628 55324 -72452
rect 55378 -72628 55412 -72452
rect 53942 -73012 54718 -72978
rect 53942 -73190 54718 -73156
rect 55820 -73116 55854 -72340
rect 55998 -73116 56032 -72340
rect 53464 -74184 53498 -73408
rect 53642 -74184 53676 -73408
rect 53942 -73418 54718 -73384
rect 53942 -73596 54718 -73562
rect 55280 -74124 55314 -73948
rect 55368 -74124 55402 -73948
rect 55820 -74230 55854 -73454
rect 55998 -74230 56032 -73454
rect 57131 -72734 57165 -72700
rect 57217 -72747 57251 -72713
rect 57303 -72717 57337 -72683
rect 59958 -72608 60334 -72574
rect 59958 -72716 60334 -72682
rect 59502 -73158 59536 -72982
rect 59590 -73158 59624 -72982
rect 59818 -73158 59852 -72982
rect 59906 -73158 59940 -72982
rect 60203 -73207 60237 -73173
rect 61215 -73207 61249 -73173
rect 60211 -73291 60245 -73257
rect 61207 -73291 61241 -73257
rect 57131 -73888 57165 -73854
rect 57217 -73875 57251 -73841
rect 57303 -73905 57337 -73871
rect 59501 -73671 59535 -73495
rect 59589 -73671 59623 -73495
rect 60203 -73375 60237 -73341
rect 61215 -73375 61249 -73341
rect 59817 -73671 59851 -73495
rect 59905 -73671 59939 -73495
rect 60211 -73459 60245 -73425
rect 61207 -73459 61241 -73425
rect 60204 -73543 60238 -73509
rect 61214 -73543 61248 -73509
rect 59958 -73974 60334 -73940
rect 59958 -74082 60334 -74048
rect 55300 -74792 55476 -74758
rect 55300 -74880 55476 -74846
rect 53464 -78566 53498 -77790
rect 53642 -78566 53676 -77790
rect 55290 -78028 55324 -77852
rect 55378 -78028 55412 -77852
rect 53942 -78412 54718 -78378
rect 53942 -78590 54718 -78556
rect 55820 -78516 55854 -77740
rect 55998 -78516 56032 -77740
rect 53464 -79584 53498 -78808
rect 53642 -79584 53676 -78808
rect 53942 -78818 54718 -78784
rect 53942 -78996 54718 -78962
rect 55280 -79524 55314 -79348
rect 55368 -79524 55402 -79348
rect 55820 -79630 55854 -78854
rect 55998 -79630 56032 -78854
rect 57131 -78134 57165 -78100
rect 57217 -78147 57251 -78113
rect 57303 -78117 57337 -78083
rect 59958 -78008 60334 -77974
rect 59958 -78116 60334 -78082
rect 59502 -78558 59536 -78382
rect 59590 -78558 59624 -78382
rect 59818 -78558 59852 -78382
rect 59906 -78558 59940 -78382
rect 60203 -78607 60237 -78573
rect 61215 -78607 61249 -78573
rect 60211 -78691 60245 -78657
rect 61207 -78691 61241 -78657
rect 57131 -79288 57165 -79254
rect 57217 -79275 57251 -79241
rect 57303 -79305 57337 -79271
rect 59501 -79071 59535 -78895
rect 59589 -79071 59623 -78895
rect 60203 -78775 60237 -78741
rect 61215 -78775 61249 -78741
rect 59817 -79071 59851 -78895
rect 59905 -79071 59939 -78895
rect 60211 -78859 60245 -78825
rect 61207 -78859 61241 -78825
rect 60204 -78943 60238 -78909
rect 61214 -78943 61248 -78909
rect 59958 -79374 60334 -79340
rect 59958 -79482 60334 -79448
rect 55300 -80192 55476 -80158
rect 55300 -80280 55476 -80246
rect 53464 -83966 53498 -83190
rect 53642 -83966 53676 -83190
rect 55290 -83428 55324 -83252
rect 55378 -83428 55412 -83252
rect 53942 -83812 54718 -83778
rect 53942 -83990 54718 -83956
rect 55820 -83916 55854 -83140
rect 55998 -83916 56032 -83140
rect 53464 -84984 53498 -84208
rect 53642 -84984 53676 -84208
rect 53942 -84218 54718 -84184
rect 53942 -84396 54718 -84362
rect 55280 -84924 55314 -84748
rect 55368 -84924 55402 -84748
rect 55820 -85030 55854 -84254
rect 55998 -85030 56032 -84254
rect 57131 -83534 57165 -83500
rect 57217 -83547 57251 -83513
rect 57303 -83517 57337 -83483
rect 59958 -83408 60334 -83374
rect 59958 -83516 60334 -83482
rect 59502 -83958 59536 -83782
rect 59590 -83958 59624 -83782
rect 59818 -83958 59852 -83782
rect 59906 -83958 59940 -83782
rect 60203 -84007 60237 -83973
rect 61215 -84007 61249 -83973
rect 60211 -84091 60245 -84057
rect 61207 -84091 61241 -84057
rect 57131 -84688 57165 -84654
rect 57217 -84675 57251 -84641
rect 57303 -84705 57337 -84671
rect 59501 -84471 59535 -84295
rect 59589 -84471 59623 -84295
rect 60203 -84175 60237 -84141
rect 61215 -84175 61249 -84141
rect 59817 -84471 59851 -84295
rect 59905 -84471 59939 -84295
rect 60211 -84259 60245 -84225
rect 61207 -84259 61241 -84225
rect 60204 -84343 60238 -84309
rect 61214 -84343 61248 -84309
rect 59958 -84774 60334 -84740
rect 59958 -84882 60334 -84848
rect 55300 -85592 55476 -85558
rect 55300 -85680 55476 -85646
<< pdiffc >>
rect 54091 -1706 54867 -1672
rect 54091 -1834 54867 -1800
rect 54091 -2062 54867 -2028
rect 54091 -2190 54867 -2156
rect 57131 -2163 57165 -2129
rect 57131 -2231 57165 -2197
rect 57217 -2163 57251 -2129
rect 57217 -2231 57251 -2197
rect 57303 -2163 57337 -2129
rect 57303 -2244 57337 -2210
rect 59125 -2081 59501 -2047
rect 59125 -2189 59501 -2155
rect 59125 -2297 59501 -2263
rect 54081 -4022 54857 -3988
rect 54081 -4150 54857 -4116
rect 56430 -3475 56464 -2699
rect 56558 -3475 56592 -2699
rect 59044 -2947 59078 -2571
rect 59162 -2947 59196 -2571
rect 60459 -3007 60493 -2973
rect 60527 -3007 60561 -2973
rect 60595 -3007 60629 -2973
rect 60823 -3007 60857 -2973
rect 60891 -3007 60925 -2973
rect 60959 -3007 60993 -2973
rect 60459 -3091 60493 -3057
rect 60527 -3091 60561 -3057
rect 60595 -3091 60629 -3057
rect 60823 -3091 60857 -3057
rect 60891 -3091 60925 -3057
rect 60959 -3091 60993 -3057
rect 59044 -3677 59078 -3301
rect 59162 -3677 59196 -3301
rect 60527 -3175 60561 -3141
rect 60595 -3175 60629 -3141
rect 60823 -3175 60857 -3141
rect 60891 -3175 60925 -3141
rect 60459 -3259 60493 -3225
rect 60527 -3259 60561 -3225
rect 60595 -3259 60629 -3225
rect 60823 -3259 60857 -3225
rect 60891 -3259 60925 -3225
rect 60959 -3259 60993 -3225
rect 60595 -3343 60629 -3309
rect 60823 -3343 60857 -3309
rect 57131 -3991 57165 -3957
rect 57131 -4059 57165 -4025
rect 57217 -3991 57251 -3957
rect 57217 -4059 57251 -4025
rect 57303 -3978 57337 -3944
rect 57303 -4059 57337 -4025
rect 59125 -3988 59501 -3954
rect 59125 -4096 59501 -4062
rect 59125 -4204 59501 -4170
rect 54081 -4378 54857 -4344
rect 54081 -4506 54857 -4472
rect 54091 -7106 54867 -7072
rect 54091 -7234 54867 -7200
rect 20846 -11644 20880 -7868
rect 21104 -11644 21138 -7868
rect 21332 -11644 21366 -7868
rect 21590 -11644 21624 -7868
rect 21818 -11644 21852 -7868
rect 22076 -11644 22110 -7868
rect 54091 -7462 54867 -7428
rect 54091 -7590 54867 -7556
rect 57131 -7563 57165 -7529
rect 57131 -7631 57165 -7597
rect 57217 -7563 57251 -7529
rect 57217 -7631 57251 -7597
rect 57303 -7563 57337 -7529
rect 57303 -7644 57337 -7610
rect 59125 -7481 59501 -7447
rect 59125 -7589 59501 -7555
rect 59125 -7697 59501 -7663
rect 54081 -9422 54857 -9388
rect 54081 -9550 54857 -9516
rect 56430 -8875 56464 -8099
rect 56558 -8875 56592 -8099
rect 59044 -8347 59078 -7971
rect 59162 -8347 59196 -7971
rect 60459 -8407 60493 -8373
rect 60527 -8407 60561 -8373
rect 60595 -8407 60629 -8373
rect 60823 -8407 60857 -8373
rect 60891 -8407 60925 -8373
rect 60959 -8407 60993 -8373
rect 60459 -8491 60493 -8457
rect 60527 -8491 60561 -8457
rect 60595 -8491 60629 -8457
rect 60823 -8491 60857 -8457
rect 60891 -8491 60925 -8457
rect 60959 -8491 60993 -8457
rect 59044 -9077 59078 -8701
rect 59162 -9077 59196 -8701
rect 60527 -8575 60561 -8541
rect 60595 -8575 60629 -8541
rect 60823 -8575 60857 -8541
rect 60891 -8575 60925 -8541
rect 60459 -8659 60493 -8625
rect 60527 -8659 60561 -8625
rect 60595 -8659 60629 -8625
rect 60823 -8659 60857 -8625
rect 60891 -8659 60925 -8625
rect 60959 -8659 60993 -8625
rect 60595 -8743 60629 -8709
rect 60823 -8743 60857 -8709
rect 57131 -9391 57165 -9357
rect 57131 -9459 57165 -9425
rect 57217 -9391 57251 -9357
rect 57217 -9459 57251 -9425
rect 57303 -9378 57337 -9344
rect 57303 -9459 57337 -9425
rect 59125 -9388 59501 -9354
rect 59125 -9496 59501 -9462
rect 59125 -9604 59501 -9570
rect 54081 -9778 54857 -9744
rect 54081 -9906 54857 -9872
rect 54091 -12506 54867 -12472
rect 54091 -12634 54867 -12600
rect 54091 -12862 54867 -12828
rect 54091 -12990 54867 -12956
rect 57131 -12963 57165 -12929
rect 57131 -13031 57165 -12997
rect 57217 -12963 57251 -12929
rect 57217 -13031 57251 -12997
rect 57303 -12963 57337 -12929
rect 57303 -13044 57337 -13010
rect 59125 -12881 59501 -12847
rect 59125 -12989 59501 -12955
rect 59125 -13097 59501 -13063
rect 54081 -14822 54857 -14788
rect 54081 -14950 54857 -14916
rect 56430 -14275 56464 -13499
rect 56558 -14275 56592 -13499
rect 59044 -13747 59078 -13371
rect 59162 -13747 59196 -13371
rect 60459 -13807 60493 -13773
rect 60527 -13807 60561 -13773
rect 60595 -13807 60629 -13773
rect 60823 -13807 60857 -13773
rect 60891 -13807 60925 -13773
rect 60959 -13807 60993 -13773
rect 60459 -13891 60493 -13857
rect 60527 -13891 60561 -13857
rect 60595 -13891 60629 -13857
rect 60823 -13891 60857 -13857
rect 60891 -13891 60925 -13857
rect 60959 -13891 60993 -13857
rect 59044 -14477 59078 -14101
rect 59162 -14477 59196 -14101
rect 60527 -13975 60561 -13941
rect 60595 -13975 60629 -13941
rect 60823 -13975 60857 -13941
rect 60891 -13975 60925 -13941
rect 60459 -14059 60493 -14025
rect 60527 -14059 60561 -14025
rect 60595 -14059 60629 -14025
rect 60823 -14059 60857 -14025
rect 60891 -14059 60925 -14025
rect 60959 -14059 60993 -14025
rect 60595 -14143 60629 -14109
rect 60823 -14143 60857 -14109
rect 57131 -14791 57165 -14757
rect 57131 -14859 57165 -14825
rect 57217 -14791 57251 -14757
rect 57217 -14859 57251 -14825
rect 57303 -14778 57337 -14744
rect 57303 -14859 57337 -14825
rect 59125 -14788 59501 -14754
rect 59125 -14896 59501 -14862
rect 59125 -15004 59501 -14970
rect 54081 -15178 54857 -15144
rect 54081 -15306 54857 -15272
rect 54091 -17906 54867 -17872
rect 54091 -18034 54867 -18000
rect 54091 -18262 54867 -18228
rect 54091 -18390 54867 -18356
rect 57131 -18363 57165 -18329
rect 57131 -18431 57165 -18397
rect 57217 -18363 57251 -18329
rect 57217 -18431 57251 -18397
rect 57303 -18363 57337 -18329
rect 57303 -18444 57337 -18410
rect 59125 -18281 59501 -18247
rect 59125 -18389 59501 -18355
rect 59125 -18497 59501 -18463
rect 54081 -20222 54857 -20188
rect 54081 -20350 54857 -20316
rect 56430 -19675 56464 -18899
rect 56558 -19675 56592 -18899
rect 59044 -19147 59078 -18771
rect 59162 -19147 59196 -18771
rect 60459 -19207 60493 -19173
rect 60527 -19207 60561 -19173
rect 60595 -19207 60629 -19173
rect 60823 -19207 60857 -19173
rect 60891 -19207 60925 -19173
rect 60959 -19207 60993 -19173
rect 60459 -19291 60493 -19257
rect 60527 -19291 60561 -19257
rect 60595 -19291 60629 -19257
rect 60823 -19291 60857 -19257
rect 60891 -19291 60925 -19257
rect 60959 -19291 60993 -19257
rect 59044 -19877 59078 -19501
rect 59162 -19877 59196 -19501
rect 60527 -19375 60561 -19341
rect 60595 -19375 60629 -19341
rect 60823 -19375 60857 -19341
rect 60891 -19375 60925 -19341
rect 60459 -19459 60493 -19425
rect 60527 -19459 60561 -19425
rect 60595 -19459 60629 -19425
rect 60823 -19459 60857 -19425
rect 60891 -19459 60925 -19425
rect 60959 -19459 60993 -19425
rect 60595 -19543 60629 -19509
rect 60823 -19543 60857 -19509
rect 57131 -20191 57165 -20157
rect 57131 -20259 57165 -20225
rect 57217 -20191 57251 -20157
rect 57217 -20259 57251 -20225
rect 57303 -20178 57337 -20144
rect 57303 -20259 57337 -20225
rect 59125 -20188 59501 -20154
rect 59125 -20296 59501 -20262
rect 59125 -20404 59501 -20370
rect 54081 -20578 54857 -20544
rect 54081 -20706 54857 -20672
rect 54091 -23306 54867 -23272
rect 54091 -23434 54867 -23400
rect 54091 -23662 54867 -23628
rect 54091 -23790 54867 -23756
rect 57131 -23763 57165 -23729
rect 57131 -23831 57165 -23797
rect 57217 -23763 57251 -23729
rect 57217 -23831 57251 -23797
rect 57303 -23763 57337 -23729
rect 57303 -23844 57337 -23810
rect 59125 -23681 59501 -23647
rect 59125 -23789 59501 -23755
rect 59125 -23897 59501 -23863
rect 54081 -25622 54857 -25588
rect 54081 -25750 54857 -25716
rect 56430 -25075 56464 -24299
rect 56558 -25075 56592 -24299
rect 59044 -24547 59078 -24171
rect 59162 -24547 59196 -24171
rect 60459 -24607 60493 -24573
rect 60527 -24607 60561 -24573
rect 60595 -24607 60629 -24573
rect 60823 -24607 60857 -24573
rect 60891 -24607 60925 -24573
rect 60959 -24607 60993 -24573
rect 60459 -24691 60493 -24657
rect 60527 -24691 60561 -24657
rect 60595 -24691 60629 -24657
rect 60823 -24691 60857 -24657
rect 60891 -24691 60925 -24657
rect 60959 -24691 60993 -24657
rect 59044 -25277 59078 -24901
rect 59162 -25277 59196 -24901
rect 60527 -24775 60561 -24741
rect 60595 -24775 60629 -24741
rect 60823 -24775 60857 -24741
rect 60891 -24775 60925 -24741
rect 60459 -24859 60493 -24825
rect 60527 -24859 60561 -24825
rect 60595 -24859 60629 -24825
rect 60823 -24859 60857 -24825
rect 60891 -24859 60925 -24825
rect 60959 -24859 60993 -24825
rect 60595 -24943 60629 -24909
rect 60823 -24943 60857 -24909
rect 57131 -25591 57165 -25557
rect 57131 -25659 57165 -25625
rect 57217 -25591 57251 -25557
rect 57217 -25659 57251 -25625
rect 57303 -25578 57337 -25544
rect 57303 -25659 57337 -25625
rect 59125 -25588 59501 -25554
rect 59125 -25696 59501 -25662
rect 59125 -25804 59501 -25770
rect 54081 -25978 54857 -25944
rect 54081 -26106 54857 -26072
rect 54091 -28706 54867 -28672
rect 54091 -28834 54867 -28800
rect 54091 -29062 54867 -29028
rect 54091 -29190 54867 -29156
rect 57131 -29163 57165 -29129
rect 57131 -29231 57165 -29197
rect 57217 -29163 57251 -29129
rect 57217 -29231 57251 -29197
rect 57303 -29163 57337 -29129
rect 57303 -29244 57337 -29210
rect 59125 -29081 59501 -29047
rect 59125 -29189 59501 -29155
rect 59125 -29297 59501 -29263
rect 54081 -31022 54857 -30988
rect 54081 -31150 54857 -31116
rect 56430 -30475 56464 -29699
rect 56558 -30475 56592 -29699
rect 59044 -29947 59078 -29571
rect 59162 -29947 59196 -29571
rect 60459 -30007 60493 -29973
rect 60527 -30007 60561 -29973
rect 60595 -30007 60629 -29973
rect 60823 -30007 60857 -29973
rect 60891 -30007 60925 -29973
rect 60959 -30007 60993 -29973
rect 60459 -30091 60493 -30057
rect 60527 -30091 60561 -30057
rect 60595 -30091 60629 -30057
rect 60823 -30091 60857 -30057
rect 60891 -30091 60925 -30057
rect 60959 -30091 60993 -30057
rect 59044 -30677 59078 -30301
rect 59162 -30677 59196 -30301
rect 60527 -30175 60561 -30141
rect 60595 -30175 60629 -30141
rect 60823 -30175 60857 -30141
rect 60891 -30175 60925 -30141
rect 60459 -30259 60493 -30225
rect 60527 -30259 60561 -30225
rect 60595 -30259 60629 -30225
rect 60823 -30259 60857 -30225
rect 60891 -30259 60925 -30225
rect 60959 -30259 60993 -30225
rect 60595 -30343 60629 -30309
rect 60823 -30343 60857 -30309
rect 57131 -30991 57165 -30957
rect 57131 -31059 57165 -31025
rect 57217 -30991 57251 -30957
rect 57217 -31059 57251 -31025
rect 57303 -30978 57337 -30944
rect 57303 -31059 57337 -31025
rect 59125 -30988 59501 -30954
rect 59125 -31096 59501 -31062
rect 59125 -31204 59501 -31170
rect 54081 -31378 54857 -31344
rect 54081 -31506 54857 -31472
rect 54091 -34106 54867 -34072
rect 54091 -34234 54867 -34200
rect 54091 -34462 54867 -34428
rect 54091 -34590 54867 -34556
rect 57131 -34563 57165 -34529
rect 57131 -34631 57165 -34597
rect 57217 -34563 57251 -34529
rect 57217 -34631 57251 -34597
rect 57303 -34563 57337 -34529
rect 57303 -34644 57337 -34610
rect 59125 -34481 59501 -34447
rect 59125 -34589 59501 -34555
rect 59125 -34697 59501 -34663
rect 54081 -36422 54857 -36388
rect 54081 -36550 54857 -36516
rect 56430 -35875 56464 -35099
rect 56558 -35875 56592 -35099
rect 59044 -35347 59078 -34971
rect 59162 -35347 59196 -34971
rect 60459 -35407 60493 -35373
rect 60527 -35407 60561 -35373
rect 60595 -35407 60629 -35373
rect 60823 -35407 60857 -35373
rect 60891 -35407 60925 -35373
rect 60959 -35407 60993 -35373
rect 60459 -35491 60493 -35457
rect 60527 -35491 60561 -35457
rect 60595 -35491 60629 -35457
rect 60823 -35491 60857 -35457
rect 60891 -35491 60925 -35457
rect 60959 -35491 60993 -35457
rect 59044 -36077 59078 -35701
rect 59162 -36077 59196 -35701
rect 60527 -35575 60561 -35541
rect 60595 -35575 60629 -35541
rect 60823 -35575 60857 -35541
rect 60891 -35575 60925 -35541
rect 60459 -35659 60493 -35625
rect 60527 -35659 60561 -35625
rect 60595 -35659 60629 -35625
rect 60823 -35659 60857 -35625
rect 60891 -35659 60925 -35625
rect 60959 -35659 60993 -35625
rect 60595 -35743 60629 -35709
rect 60823 -35743 60857 -35709
rect 57131 -36391 57165 -36357
rect 57131 -36459 57165 -36425
rect 57217 -36391 57251 -36357
rect 57217 -36459 57251 -36425
rect 57303 -36378 57337 -36344
rect 57303 -36459 57337 -36425
rect 59125 -36388 59501 -36354
rect 59125 -36496 59501 -36462
rect 59125 -36604 59501 -36570
rect 54081 -36778 54857 -36744
rect 54081 -36906 54857 -36872
rect 75582 -38737 75616 -38703
rect 75582 -38805 75616 -38771
rect 75582 -38873 75616 -38839
rect 75666 -38737 75700 -38703
rect 75666 -38805 75700 -38771
rect 75666 -38873 75700 -38839
rect 75858 -38737 75892 -38703
rect 75858 -38805 75892 -38771
rect 75858 -38873 75892 -38839
rect 75942 -38737 75976 -38703
rect 75942 -38805 75976 -38771
rect 75942 -38873 75976 -38839
rect 76132 -38737 76166 -38703
rect 76132 -38805 76166 -38771
rect 76132 -38873 76166 -38839
rect 76216 -38737 76250 -38703
rect 76216 -38805 76250 -38771
rect 76216 -38873 76250 -38839
rect 76408 -38737 76442 -38703
rect 76408 -38805 76442 -38771
rect 76408 -38873 76442 -38839
rect 76492 -38737 76526 -38703
rect 76492 -38805 76526 -38771
rect 76492 -38873 76526 -38839
rect 76684 -38737 76718 -38703
rect 76684 -38805 76718 -38771
rect 76684 -38873 76718 -38839
rect 76768 -38737 76802 -38703
rect 76768 -38805 76802 -38771
rect 76768 -38873 76802 -38839
rect 77974 -39151 78008 -39117
rect 77974 -39219 78008 -39185
rect 77613 -39282 77647 -39248
rect 78059 -39182 78093 -39148
rect 78432 -39151 78466 -39117
rect 78059 -39250 78093 -39216
rect 78432 -39219 78466 -39185
rect 78167 -39282 78201 -39248
rect 78517 -39182 78551 -39148
rect 78517 -39250 78551 -39216
rect 78661 -39193 78695 -39159
rect 78745 -39193 78779 -39159
rect 78853 -39151 78887 -39117
rect 78853 -39219 78887 -39185
rect 54091 -39506 54867 -39472
rect 54091 -39634 54867 -39600
rect 78957 -39151 78991 -39117
rect 78957 -39219 78991 -39185
rect 80814 -39201 80848 -39167
rect 80814 -39269 80848 -39235
rect 80814 -39337 80848 -39303
rect 80898 -39201 80932 -39167
rect 80898 -39269 80932 -39235
rect 80898 -39337 80932 -39303
rect 81059 -39201 81093 -39167
rect 81059 -39269 81093 -39235
rect 81059 -39337 81093 -39303
rect 81143 -39201 81177 -39167
rect 81143 -39269 81177 -39235
rect 81143 -39337 81177 -39303
rect 81227 -39201 81261 -39167
rect 81227 -39269 81261 -39235
rect 81311 -39201 81345 -39167
rect 81311 -39269 81345 -39235
rect 81311 -39337 81345 -39303
rect 81395 -39201 81429 -39167
rect 81522 -39201 81556 -39167
rect 81522 -39269 81556 -39235
rect 81522 -39339 81556 -39305
rect 81606 -39201 81640 -39167
rect 81606 -39269 81640 -39235
rect 81606 -39339 81640 -39305
rect 81690 -39201 81724 -39167
rect 81690 -39269 81724 -39235
rect 81774 -39201 81808 -39167
rect 81774 -39269 81808 -39235
rect 81774 -39339 81808 -39305
rect 81858 -39201 81892 -39167
rect 81858 -39269 81892 -39235
rect 81942 -39201 81976 -39167
rect 81942 -39269 81976 -39235
rect 81942 -39339 81976 -39305
rect 82026 -39201 82060 -39167
rect 82026 -39269 82060 -39235
rect 82110 -39201 82144 -39167
rect 82110 -39269 82144 -39235
rect 82110 -39339 82144 -39305
rect 82194 -39201 82228 -39167
rect 82194 -39269 82228 -39235
rect 82278 -39201 82312 -39167
rect 82278 -39269 82312 -39235
rect 82278 -39339 82312 -39305
rect 82362 -39201 82396 -39167
rect 82362 -39269 82396 -39235
rect 82446 -39201 82480 -39167
rect 82446 -39269 82480 -39235
rect 82446 -39339 82480 -39305
rect 82530 -39201 82564 -39167
rect 82530 -39269 82564 -39235
rect 82614 -39201 82648 -39167
rect 82614 -39269 82648 -39235
rect 82614 -39339 82648 -39305
rect 82698 -39201 82732 -39167
rect 82698 -39269 82732 -39235
rect 82782 -39201 82816 -39167
rect 82782 -39269 82816 -39235
rect 82782 -39339 82816 -39305
rect 82866 -39201 82900 -39167
rect 82866 -39269 82900 -39235
rect 82994 -39201 83028 -39167
rect 82994 -39269 83028 -39235
rect 82994 -39339 83028 -39305
rect 83078 -39201 83112 -39167
rect 83078 -39269 83112 -39235
rect 83078 -39339 83112 -39305
rect 83162 -39201 83196 -39167
rect 83162 -39269 83196 -39235
rect 83246 -39201 83280 -39167
rect 83246 -39269 83280 -39235
rect 83246 -39339 83280 -39305
rect 83330 -39201 83364 -39167
rect 83330 -39269 83364 -39235
rect 83414 -39201 83448 -39167
rect 83414 -39269 83448 -39235
rect 83414 -39339 83448 -39305
rect 83498 -39201 83532 -39167
rect 83498 -39269 83532 -39235
rect 83582 -39201 83616 -39167
rect 83582 -39269 83616 -39235
rect 83582 -39339 83616 -39305
rect 83666 -39201 83700 -39167
rect 83666 -39269 83700 -39235
rect 83750 -39201 83784 -39167
rect 83750 -39269 83784 -39235
rect 83750 -39339 83784 -39305
rect 83834 -39201 83868 -39167
rect 83834 -39269 83868 -39235
rect 83918 -39201 83952 -39167
rect 83918 -39269 83952 -39235
rect 83918 -39339 83952 -39305
rect 84002 -39201 84036 -39167
rect 84002 -39269 84036 -39235
rect 84086 -39201 84120 -39167
rect 84086 -39269 84120 -39235
rect 84086 -39339 84120 -39305
rect 84170 -39201 84204 -39167
rect 84170 -39269 84204 -39235
rect 84254 -39201 84288 -39167
rect 84254 -39269 84288 -39235
rect 84254 -39339 84288 -39305
rect 84338 -39201 84372 -39167
rect 84338 -39269 84372 -39235
rect 84466 -39201 84500 -39167
rect 84466 -39269 84500 -39235
rect 84466 -39339 84500 -39305
rect 84550 -39201 84584 -39167
rect 84550 -39269 84584 -39235
rect 84550 -39339 84584 -39305
rect 84634 -39201 84668 -39167
rect 84634 -39269 84668 -39235
rect 84718 -39201 84752 -39167
rect 84718 -39269 84752 -39235
rect 84718 -39339 84752 -39305
rect 84802 -39201 84836 -39167
rect 84802 -39269 84836 -39235
rect 84886 -39201 84920 -39167
rect 84886 -39269 84920 -39235
rect 84886 -39339 84920 -39305
rect 84970 -39201 85004 -39167
rect 84970 -39269 85004 -39235
rect 85054 -39201 85088 -39167
rect 85054 -39269 85088 -39235
rect 85054 -39339 85088 -39305
rect 85138 -39201 85172 -39167
rect 85138 -39269 85172 -39235
rect 85222 -39201 85256 -39167
rect 85222 -39269 85256 -39235
rect 85222 -39339 85256 -39305
rect 85306 -39201 85340 -39167
rect 85306 -39269 85340 -39235
rect 85390 -39201 85424 -39167
rect 85390 -39269 85424 -39235
rect 85390 -39339 85424 -39305
rect 85474 -39201 85508 -39167
rect 85474 -39269 85508 -39235
rect 85558 -39201 85592 -39167
rect 85558 -39269 85592 -39235
rect 85558 -39339 85592 -39305
rect 85642 -39201 85676 -39167
rect 85642 -39269 85676 -39235
rect 85726 -39201 85760 -39167
rect 85726 -39269 85760 -39235
rect 85726 -39339 85760 -39305
rect 85810 -39201 85844 -39167
rect 85810 -39269 85844 -39235
rect 85938 -39201 85972 -39167
rect 85938 -39269 85972 -39235
rect 85938 -39339 85972 -39305
rect 86022 -39201 86056 -39167
rect 86022 -39269 86056 -39235
rect 86022 -39339 86056 -39305
rect 86106 -39201 86140 -39167
rect 86106 -39269 86140 -39235
rect 86190 -39201 86224 -39167
rect 86190 -39269 86224 -39235
rect 86190 -39339 86224 -39305
rect 86274 -39201 86308 -39167
rect 86274 -39269 86308 -39235
rect 86358 -39201 86392 -39167
rect 86358 -39269 86392 -39235
rect 86358 -39339 86392 -39305
rect 86442 -39201 86476 -39167
rect 86442 -39269 86476 -39235
rect 86526 -39201 86560 -39167
rect 86526 -39269 86560 -39235
rect 86526 -39339 86560 -39305
rect 86610 -39201 86644 -39167
rect 86610 -39269 86644 -39235
rect 86694 -39201 86728 -39167
rect 86694 -39269 86728 -39235
rect 86694 -39339 86728 -39305
rect 86778 -39201 86812 -39167
rect 86778 -39269 86812 -39235
rect 86862 -39201 86896 -39167
rect 86862 -39269 86896 -39235
rect 86862 -39339 86896 -39305
rect 86946 -39201 86980 -39167
rect 86946 -39269 86980 -39235
rect 87030 -39201 87064 -39167
rect 87030 -39269 87064 -39235
rect 87030 -39339 87064 -39305
rect 87114 -39201 87148 -39167
rect 87114 -39269 87148 -39235
rect 87198 -39201 87232 -39167
rect 87198 -39269 87232 -39235
rect 87198 -39339 87232 -39305
rect 87282 -39201 87316 -39167
rect 87282 -39269 87316 -39235
rect 87410 -39201 87444 -39167
rect 87410 -39269 87444 -39235
rect 87410 -39339 87444 -39305
rect 87494 -39201 87528 -39167
rect 87494 -39269 87528 -39235
rect 87494 -39339 87528 -39305
rect 87578 -39201 87612 -39167
rect 87578 -39269 87612 -39235
rect 87662 -39201 87696 -39167
rect 87662 -39269 87696 -39235
rect 87662 -39339 87696 -39305
rect 87746 -39201 87780 -39167
rect 87746 -39269 87780 -39235
rect 87830 -39201 87864 -39167
rect 87830 -39269 87864 -39235
rect 87830 -39339 87864 -39305
rect 87914 -39201 87948 -39167
rect 87914 -39269 87948 -39235
rect 87998 -39201 88032 -39167
rect 87998 -39269 88032 -39235
rect 87998 -39339 88032 -39305
rect 88082 -39201 88116 -39167
rect 88082 -39269 88116 -39235
rect 88166 -39201 88200 -39167
rect 88166 -39269 88200 -39235
rect 88166 -39339 88200 -39305
rect 88250 -39201 88284 -39167
rect 88250 -39269 88284 -39235
rect 88334 -39201 88368 -39167
rect 88334 -39269 88368 -39235
rect 88334 -39339 88368 -39305
rect 88418 -39201 88452 -39167
rect 88418 -39269 88452 -39235
rect 88502 -39201 88536 -39167
rect 88502 -39269 88536 -39235
rect 88502 -39339 88536 -39305
rect 88586 -39201 88620 -39167
rect 88586 -39269 88620 -39235
rect 88670 -39201 88704 -39167
rect 88670 -39269 88704 -39235
rect 88670 -39339 88704 -39305
rect 88754 -39201 88788 -39167
rect 88754 -39269 88788 -39235
rect 54091 -39862 54867 -39828
rect 54091 -39990 54867 -39956
rect 57131 -39963 57165 -39929
rect 57131 -40031 57165 -39997
rect 57217 -39963 57251 -39929
rect 57217 -40031 57251 -39997
rect 57303 -39963 57337 -39929
rect 57303 -40044 57337 -40010
rect 59125 -39881 59501 -39847
rect 59125 -39989 59501 -39955
rect 59125 -40097 59501 -40063
rect 77613 -40042 77647 -40008
rect 54081 -41822 54857 -41788
rect 54081 -41950 54857 -41916
rect 56430 -41275 56464 -40499
rect 56558 -41275 56592 -40499
rect 59044 -40747 59078 -40371
rect 59162 -40747 59196 -40371
rect 77974 -40105 78008 -40071
rect 77974 -40173 78008 -40139
rect 78059 -40074 78093 -40040
rect 78059 -40142 78093 -40108
rect 80864 -40077 80898 -40043
rect 80864 -40145 80898 -40111
rect 80864 -40213 80898 -40179
rect 80948 -40077 80982 -40043
rect 80948 -40145 80982 -40111
rect 80948 -40213 80982 -40179
rect 77649 -40443 77683 -40409
rect 77733 -40443 77767 -40409
rect 77841 -40401 77875 -40367
rect 77841 -40469 77875 -40435
rect 77945 -40401 77979 -40367
rect 77945 -40469 77979 -40435
rect 60459 -40807 60493 -40773
rect 60527 -40807 60561 -40773
rect 60595 -40807 60629 -40773
rect 60823 -40807 60857 -40773
rect 60891 -40807 60925 -40773
rect 60959 -40807 60993 -40773
rect 60459 -40891 60493 -40857
rect 60527 -40891 60561 -40857
rect 60595 -40891 60629 -40857
rect 60823 -40891 60857 -40857
rect 60891 -40891 60925 -40857
rect 60959 -40891 60993 -40857
rect 59044 -41477 59078 -41101
rect 59162 -41477 59196 -41101
rect 60527 -40975 60561 -40941
rect 60595 -40975 60629 -40941
rect 60823 -40975 60857 -40941
rect 60891 -40975 60925 -40941
rect 60459 -41059 60493 -41025
rect 60527 -41059 60561 -41025
rect 60595 -41059 60629 -41025
rect 60823 -41059 60857 -41025
rect 60891 -41059 60925 -41025
rect 60959 -41059 60993 -41025
rect 60595 -41143 60629 -41109
rect 60823 -41143 60857 -41109
rect 77649 -41371 77683 -41337
rect 77733 -41371 77767 -41337
rect 77841 -41345 77875 -41311
rect 77841 -41413 77875 -41379
rect 78073 -41282 78107 -41248
rect 77945 -41345 77979 -41311
rect 78434 -41345 78468 -41311
rect 77945 -41413 77979 -41379
rect 78434 -41413 78468 -41379
rect 78519 -41314 78553 -41280
rect 78519 -41382 78553 -41348
rect 57131 -41791 57165 -41757
rect 57131 -41859 57165 -41825
rect 57217 -41791 57251 -41757
rect 57217 -41859 57251 -41825
rect 57303 -41778 57337 -41744
rect 57303 -41859 57337 -41825
rect 59125 -41788 59501 -41754
rect 59125 -41896 59501 -41862
rect 59125 -42004 59501 -41970
rect 54081 -42178 54857 -42144
rect 54081 -42306 54857 -42272
rect 77649 -41683 77683 -41649
rect 77733 -41683 77767 -41649
rect 77841 -41641 77875 -41607
rect 77841 -41709 77875 -41675
rect 77945 -41641 77979 -41607
rect 77945 -41709 77979 -41675
rect 77651 -42625 77685 -42591
rect 77735 -42625 77769 -42591
rect 77843 -42599 77877 -42565
rect 77843 -42667 77877 -42633
rect 77947 -42599 77981 -42565
rect 77947 -42667 77981 -42633
rect 77613 -42891 77647 -42857
rect 77705 -42899 77739 -42865
rect 77807 -42891 77841 -42857
rect 77902 -42899 77936 -42865
rect 78053 -42891 78087 -42857
rect 78053 -42959 78087 -42925
rect 78153 -42891 78187 -42857
rect 78718 -42891 78752 -42857
rect 78153 -42959 78187 -42925
rect 78718 -42959 78752 -42925
rect 78153 -43027 78187 -42993
rect 78357 -43022 78391 -42988
rect 78803 -42922 78837 -42888
rect 78803 -42990 78837 -42956
rect 77613 -43899 77647 -43865
rect 77705 -43891 77739 -43857
rect 77807 -43899 77841 -43865
rect 77902 -43891 77936 -43857
rect 78053 -43831 78087 -43797
rect 78053 -43899 78087 -43865
rect 78153 -43763 78187 -43729
rect 83083 -43717 83117 -43683
rect 78153 -43831 78187 -43797
rect 82914 -43837 82948 -43803
rect 83083 -43785 83117 -43751
rect 83183 -43701 83217 -43667
rect 83183 -43769 83217 -43735
rect 83374 -43701 83408 -43667
rect 83374 -43769 83408 -43735
rect 83374 -43837 83408 -43803
rect 83458 -43701 83492 -43667
rect 83458 -43769 83492 -43735
rect 83458 -43837 83492 -43803
rect 83619 -43701 83653 -43667
rect 83619 -43769 83653 -43735
rect 83619 -43837 83653 -43803
rect 83703 -43701 83737 -43667
rect 83703 -43769 83737 -43735
rect 83703 -43837 83737 -43803
rect 83787 -43701 83821 -43667
rect 83787 -43769 83821 -43735
rect 83871 -43701 83905 -43667
rect 83871 -43769 83905 -43735
rect 83871 -43837 83905 -43803
rect 83955 -43701 83989 -43667
rect 84082 -43701 84116 -43667
rect 84082 -43769 84116 -43735
rect 84082 -43839 84116 -43805
rect 84166 -43701 84200 -43667
rect 84166 -43769 84200 -43735
rect 84166 -43839 84200 -43805
rect 84250 -43701 84284 -43667
rect 84250 -43769 84284 -43735
rect 84334 -43701 84368 -43667
rect 84334 -43769 84368 -43735
rect 84334 -43839 84368 -43805
rect 84418 -43701 84452 -43667
rect 84418 -43769 84452 -43735
rect 84502 -43701 84536 -43667
rect 84502 -43769 84536 -43735
rect 84502 -43839 84536 -43805
rect 84586 -43701 84620 -43667
rect 84586 -43769 84620 -43735
rect 84670 -43701 84704 -43667
rect 84670 -43769 84704 -43735
rect 84670 -43839 84704 -43805
rect 84754 -43701 84788 -43667
rect 84754 -43769 84788 -43735
rect 84838 -43701 84872 -43667
rect 84838 -43769 84872 -43735
rect 84838 -43839 84872 -43805
rect 84922 -43701 84956 -43667
rect 84922 -43769 84956 -43735
rect 85006 -43701 85040 -43667
rect 85006 -43769 85040 -43735
rect 85006 -43839 85040 -43805
rect 85090 -43701 85124 -43667
rect 85090 -43769 85124 -43735
rect 85174 -43701 85208 -43667
rect 85174 -43769 85208 -43735
rect 85174 -43839 85208 -43805
rect 85258 -43701 85292 -43667
rect 85258 -43769 85292 -43735
rect 85342 -43701 85376 -43667
rect 85342 -43769 85376 -43735
rect 85342 -43839 85376 -43805
rect 85426 -43701 85460 -43667
rect 85426 -43769 85460 -43735
rect 85554 -43701 85588 -43667
rect 85554 -43769 85588 -43735
rect 85554 -43839 85588 -43805
rect 85638 -43701 85672 -43667
rect 85638 -43769 85672 -43735
rect 85638 -43839 85672 -43805
rect 85722 -43701 85756 -43667
rect 85722 -43769 85756 -43735
rect 85806 -43701 85840 -43667
rect 85806 -43769 85840 -43735
rect 85806 -43839 85840 -43805
rect 85890 -43701 85924 -43667
rect 85890 -43769 85924 -43735
rect 85974 -43701 86008 -43667
rect 85974 -43769 86008 -43735
rect 85974 -43839 86008 -43805
rect 86058 -43701 86092 -43667
rect 86058 -43769 86092 -43735
rect 86142 -43701 86176 -43667
rect 86142 -43769 86176 -43735
rect 86142 -43839 86176 -43805
rect 86226 -43701 86260 -43667
rect 86226 -43769 86260 -43735
rect 86310 -43701 86344 -43667
rect 86310 -43769 86344 -43735
rect 86310 -43839 86344 -43805
rect 86394 -43701 86428 -43667
rect 86394 -43769 86428 -43735
rect 86478 -43701 86512 -43667
rect 86478 -43769 86512 -43735
rect 86478 -43839 86512 -43805
rect 86562 -43701 86596 -43667
rect 86562 -43769 86596 -43735
rect 86646 -43701 86680 -43667
rect 86646 -43769 86680 -43735
rect 86646 -43839 86680 -43805
rect 86730 -43701 86764 -43667
rect 86730 -43769 86764 -43735
rect 86814 -43701 86848 -43667
rect 86814 -43769 86848 -43735
rect 86814 -43839 86848 -43805
rect 86898 -43701 86932 -43667
rect 86898 -43769 86932 -43735
rect 87026 -43701 87060 -43667
rect 87026 -43769 87060 -43735
rect 87026 -43839 87060 -43805
rect 87110 -43701 87144 -43667
rect 87110 -43769 87144 -43735
rect 87110 -43839 87144 -43805
rect 87194 -43701 87228 -43667
rect 87194 -43769 87228 -43735
rect 87278 -43701 87312 -43667
rect 87278 -43769 87312 -43735
rect 87278 -43839 87312 -43805
rect 87362 -43701 87396 -43667
rect 87362 -43769 87396 -43735
rect 87446 -43701 87480 -43667
rect 87446 -43769 87480 -43735
rect 87446 -43839 87480 -43805
rect 87530 -43701 87564 -43667
rect 87530 -43769 87564 -43735
rect 87614 -43701 87648 -43667
rect 87614 -43769 87648 -43735
rect 87614 -43839 87648 -43805
rect 87698 -43701 87732 -43667
rect 87698 -43769 87732 -43735
rect 87782 -43701 87816 -43667
rect 87782 -43769 87816 -43735
rect 87782 -43839 87816 -43805
rect 87866 -43701 87900 -43667
rect 87866 -43769 87900 -43735
rect 87950 -43701 87984 -43667
rect 87950 -43769 87984 -43735
rect 87950 -43839 87984 -43805
rect 88034 -43701 88068 -43667
rect 88034 -43769 88068 -43735
rect 88118 -43701 88152 -43667
rect 88118 -43769 88152 -43735
rect 88118 -43839 88152 -43805
rect 88202 -43701 88236 -43667
rect 88202 -43769 88236 -43735
rect 88286 -43701 88320 -43667
rect 88286 -43769 88320 -43735
rect 88286 -43839 88320 -43805
rect 88370 -43701 88404 -43667
rect 88370 -43769 88404 -43735
rect 88498 -43701 88532 -43667
rect 88498 -43769 88532 -43735
rect 88498 -43839 88532 -43805
rect 88582 -43701 88616 -43667
rect 88582 -43769 88616 -43735
rect 88582 -43839 88616 -43805
rect 88666 -43701 88700 -43667
rect 88666 -43769 88700 -43735
rect 88750 -43701 88784 -43667
rect 88750 -43769 88784 -43735
rect 88750 -43839 88784 -43805
rect 88834 -43701 88868 -43667
rect 88834 -43769 88868 -43735
rect 88918 -43701 88952 -43667
rect 88918 -43769 88952 -43735
rect 88918 -43839 88952 -43805
rect 89002 -43701 89036 -43667
rect 89002 -43769 89036 -43735
rect 89086 -43701 89120 -43667
rect 89086 -43769 89120 -43735
rect 89086 -43839 89120 -43805
rect 89170 -43701 89204 -43667
rect 89170 -43769 89204 -43735
rect 89254 -43701 89288 -43667
rect 89254 -43769 89288 -43735
rect 89254 -43839 89288 -43805
rect 89338 -43701 89372 -43667
rect 89338 -43769 89372 -43735
rect 89422 -43701 89456 -43667
rect 89422 -43769 89456 -43735
rect 89422 -43839 89456 -43805
rect 89506 -43701 89540 -43667
rect 89506 -43769 89540 -43735
rect 89590 -43701 89624 -43667
rect 89590 -43769 89624 -43735
rect 89590 -43839 89624 -43805
rect 89674 -43701 89708 -43667
rect 89674 -43769 89708 -43735
rect 89758 -43701 89792 -43667
rect 89758 -43769 89792 -43735
rect 89758 -43839 89792 -43805
rect 89842 -43701 89876 -43667
rect 89842 -43769 89876 -43735
rect 89970 -43701 90004 -43667
rect 89970 -43769 90004 -43735
rect 89970 -43839 90004 -43805
rect 90054 -43701 90088 -43667
rect 90054 -43769 90088 -43735
rect 90054 -43839 90088 -43805
rect 90138 -43701 90172 -43667
rect 90138 -43769 90172 -43735
rect 90222 -43701 90256 -43667
rect 90222 -43769 90256 -43735
rect 90222 -43839 90256 -43805
rect 90306 -43701 90340 -43667
rect 90306 -43769 90340 -43735
rect 90390 -43701 90424 -43667
rect 90390 -43769 90424 -43735
rect 90390 -43839 90424 -43805
rect 90474 -43701 90508 -43667
rect 90474 -43769 90508 -43735
rect 90558 -43701 90592 -43667
rect 90558 -43769 90592 -43735
rect 90558 -43839 90592 -43805
rect 90642 -43701 90676 -43667
rect 90642 -43769 90676 -43735
rect 90726 -43701 90760 -43667
rect 90726 -43769 90760 -43735
rect 90726 -43839 90760 -43805
rect 90810 -43701 90844 -43667
rect 90810 -43769 90844 -43735
rect 90894 -43701 90928 -43667
rect 90894 -43769 90928 -43735
rect 90894 -43839 90928 -43805
rect 90978 -43701 91012 -43667
rect 90978 -43769 91012 -43735
rect 91062 -43701 91096 -43667
rect 91062 -43769 91096 -43735
rect 91062 -43839 91096 -43805
rect 91146 -43701 91180 -43667
rect 91146 -43769 91180 -43735
rect 91230 -43701 91264 -43667
rect 91230 -43769 91264 -43735
rect 91230 -43839 91264 -43805
rect 91314 -43701 91348 -43667
rect 91314 -43769 91348 -43735
rect 78153 -43899 78187 -43865
rect 77613 -44123 77647 -44089
rect 77705 -44131 77739 -44097
rect 77807 -44123 77841 -44089
rect 77902 -44131 77936 -44097
rect 78053 -44123 78087 -44089
rect 78053 -44191 78087 -44157
rect 78153 -44123 78187 -44089
rect 78153 -44191 78187 -44157
rect 78153 -44259 78187 -44225
rect 54091 -44906 54867 -44872
rect 54091 -45034 54867 -45000
rect 54091 -45262 54867 -45228
rect 54091 -45390 54867 -45356
rect 77613 -45133 77647 -45099
rect 77705 -45125 77739 -45091
rect 77807 -45133 77841 -45099
rect 77902 -45125 77936 -45091
rect 78053 -45065 78087 -45031
rect 78053 -45133 78087 -45099
rect 78153 -44997 78187 -44963
rect 78153 -45065 78187 -45031
rect 78153 -45133 78187 -45099
rect 57131 -45363 57165 -45329
rect 57131 -45431 57165 -45397
rect 57217 -45363 57251 -45329
rect 57217 -45431 57251 -45397
rect 57303 -45363 57337 -45329
rect 57303 -45444 57337 -45410
rect 59125 -45281 59501 -45247
rect 59125 -45389 59501 -45355
rect 59125 -45497 59501 -45463
rect 77885 -45361 77919 -45327
rect 54081 -47222 54857 -47188
rect 54081 -47350 54857 -47316
rect 56430 -46675 56464 -45899
rect 56558 -46675 56592 -45899
rect 59044 -46147 59078 -45771
rect 59162 -46147 59196 -45771
rect 77613 -45500 77647 -45466
rect 77697 -45470 77731 -45436
rect 77790 -45489 77824 -45455
rect 77969 -45375 78003 -45341
rect 77969 -45443 78003 -45409
rect 78109 -45403 78143 -45369
rect 78193 -45403 78227 -45369
rect 78301 -45361 78335 -45327
rect 78301 -45429 78335 -45395
rect 78405 -45361 78439 -45327
rect 78894 -45361 78928 -45327
rect 78405 -45429 78439 -45395
rect 78894 -45429 78928 -45395
rect 78533 -45492 78567 -45458
rect 78979 -45392 79013 -45358
rect 78979 -45460 79013 -45426
rect 60459 -46207 60493 -46173
rect 60527 -46207 60561 -46173
rect 60595 -46207 60629 -46173
rect 60823 -46207 60857 -46173
rect 60891 -46207 60925 -46173
rect 60959 -46207 60993 -46173
rect 60459 -46291 60493 -46257
rect 60527 -46291 60561 -46257
rect 60595 -46291 60629 -46257
rect 60823 -46291 60857 -46257
rect 60891 -46291 60925 -46257
rect 60959 -46291 60993 -46257
rect 59044 -46877 59078 -46501
rect 59162 -46877 59196 -46501
rect 60527 -46375 60561 -46341
rect 60595 -46375 60629 -46341
rect 60823 -46375 60857 -46341
rect 60891 -46375 60925 -46341
rect 60459 -46459 60493 -46425
rect 60527 -46459 60561 -46425
rect 60595 -46459 60629 -46425
rect 60823 -46459 60857 -46425
rect 60891 -46459 60925 -46425
rect 60959 -46459 60993 -46425
rect 60595 -46543 60629 -46509
rect 60823 -46543 60857 -46509
rect 75582 -46777 75616 -46743
rect 57131 -47191 57165 -47157
rect 57131 -47259 57165 -47225
rect 57217 -47191 57251 -47157
rect 57217 -47259 57251 -47225
rect 57303 -47178 57337 -47144
rect 57303 -47259 57337 -47225
rect 59125 -47188 59501 -47154
rect 59125 -47296 59501 -47262
rect 59125 -47404 59501 -47370
rect 54081 -47578 54857 -47544
rect 54081 -47706 54857 -47672
rect 75582 -46845 75616 -46811
rect 75582 -46913 75616 -46879
rect 75666 -46777 75700 -46743
rect 75666 -46845 75700 -46811
rect 75666 -46913 75700 -46879
rect 75858 -46777 75892 -46743
rect 75858 -46845 75892 -46811
rect 75858 -46913 75892 -46879
rect 75942 -46777 75976 -46743
rect 75942 -46845 75976 -46811
rect 75942 -46913 75976 -46879
rect 76132 -46777 76166 -46743
rect 76132 -46845 76166 -46811
rect 76132 -46913 76166 -46879
rect 76216 -46777 76250 -46743
rect 76216 -46845 76250 -46811
rect 76216 -46913 76250 -46879
rect 76408 -46777 76442 -46743
rect 76408 -46845 76442 -46811
rect 76408 -46913 76442 -46879
rect 76492 -46777 76526 -46743
rect 76492 -46845 76526 -46811
rect 76492 -46913 76526 -46879
rect 76684 -46777 76718 -46743
rect 76684 -46845 76718 -46811
rect 76684 -46913 76718 -46879
rect 76768 -46777 76802 -46743
rect 76768 -46845 76802 -46811
rect 76768 -46913 76802 -46879
rect 77974 -47191 78008 -47157
rect 77974 -47259 78008 -47225
rect 77613 -47322 77647 -47288
rect 78059 -47222 78093 -47188
rect 78432 -47191 78466 -47157
rect 78059 -47290 78093 -47256
rect 78432 -47259 78466 -47225
rect 78167 -47322 78201 -47288
rect 78517 -47222 78551 -47188
rect 78517 -47290 78551 -47256
rect 78661 -47233 78695 -47199
rect 78745 -47233 78779 -47199
rect 78853 -47191 78887 -47157
rect 78853 -47259 78887 -47225
rect 78957 -47191 78991 -47157
rect 78957 -47259 78991 -47225
rect 83083 -47857 83117 -47823
rect 82914 -47977 82948 -47943
rect 83083 -47925 83117 -47891
rect 83183 -47841 83217 -47807
rect 83183 -47909 83217 -47875
rect 83374 -47841 83408 -47807
rect 83374 -47909 83408 -47875
rect 83374 -47977 83408 -47943
rect 83458 -47841 83492 -47807
rect 83458 -47909 83492 -47875
rect 83458 -47977 83492 -47943
rect 83619 -47841 83653 -47807
rect 83619 -47909 83653 -47875
rect 83619 -47977 83653 -47943
rect 83703 -47841 83737 -47807
rect 83703 -47909 83737 -47875
rect 83703 -47977 83737 -47943
rect 83787 -47841 83821 -47807
rect 83787 -47909 83821 -47875
rect 83871 -47841 83905 -47807
rect 83871 -47909 83905 -47875
rect 83871 -47977 83905 -47943
rect 83955 -47841 83989 -47807
rect 84082 -47841 84116 -47807
rect 84082 -47909 84116 -47875
rect 84082 -47979 84116 -47945
rect 84166 -47841 84200 -47807
rect 84166 -47909 84200 -47875
rect 84166 -47979 84200 -47945
rect 84250 -47841 84284 -47807
rect 84250 -47909 84284 -47875
rect 84334 -47841 84368 -47807
rect 84334 -47909 84368 -47875
rect 84334 -47979 84368 -47945
rect 84418 -47841 84452 -47807
rect 84418 -47909 84452 -47875
rect 84502 -47841 84536 -47807
rect 84502 -47909 84536 -47875
rect 84502 -47979 84536 -47945
rect 84586 -47841 84620 -47807
rect 84586 -47909 84620 -47875
rect 84670 -47841 84704 -47807
rect 84670 -47909 84704 -47875
rect 84670 -47979 84704 -47945
rect 84754 -47841 84788 -47807
rect 84754 -47909 84788 -47875
rect 84838 -47841 84872 -47807
rect 84838 -47909 84872 -47875
rect 84838 -47979 84872 -47945
rect 84922 -47841 84956 -47807
rect 84922 -47909 84956 -47875
rect 85006 -47841 85040 -47807
rect 85006 -47909 85040 -47875
rect 85006 -47979 85040 -47945
rect 85090 -47841 85124 -47807
rect 85090 -47909 85124 -47875
rect 85174 -47841 85208 -47807
rect 85174 -47909 85208 -47875
rect 85174 -47979 85208 -47945
rect 85258 -47841 85292 -47807
rect 85258 -47909 85292 -47875
rect 85342 -47841 85376 -47807
rect 85342 -47909 85376 -47875
rect 85342 -47979 85376 -47945
rect 85426 -47841 85460 -47807
rect 85426 -47909 85460 -47875
rect 85554 -47841 85588 -47807
rect 85554 -47909 85588 -47875
rect 85554 -47979 85588 -47945
rect 85638 -47841 85672 -47807
rect 85638 -47909 85672 -47875
rect 85638 -47979 85672 -47945
rect 85722 -47841 85756 -47807
rect 85722 -47909 85756 -47875
rect 85806 -47841 85840 -47807
rect 85806 -47909 85840 -47875
rect 85806 -47979 85840 -47945
rect 85890 -47841 85924 -47807
rect 85890 -47909 85924 -47875
rect 85974 -47841 86008 -47807
rect 85974 -47909 86008 -47875
rect 85974 -47979 86008 -47945
rect 86058 -47841 86092 -47807
rect 86058 -47909 86092 -47875
rect 86142 -47841 86176 -47807
rect 86142 -47909 86176 -47875
rect 86142 -47979 86176 -47945
rect 86226 -47841 86260 -47807
rect 86226 -47909 86260 -47875
rect 86310 -47841 86344 -47807
rect 86310 -47909 86344 -47875
rect 86310 -47979 86344 -47945
rect 86394 -47841 86428 -47807
rect 86394 -47909 86428 -47875
rect 86478 -47841 86512 -47807
rect 86478 -47909 86512 -47875
rect 86478 -47979 86512 -47945
rect 86562 -47841 86596 -47807
rect 86562 -47909 86596 -47875
rect 86646 -47841 86680 -47807
rect 86646 -47909 86680 -47875
rect 86646 -47979 86680 -47945
rect 86730 -47841 86764 -47807
rect 86730 -47909 86764 -47875
rect 86814 -47841 86848 -47807
rect 86814 -47909 86848 -47875
rect 86814 -47979 86848 -47945
rect 86898 -47841 86932 -47807
rect 86898 -47909 86932 -47875
rect 87026 -47841 87060 -47807
rect 87026 -47909 87060 -47875
rect 87026 -47979 87060 -47945
rect 87110 -47841 87144 -47807
rect 87110 -47909 87144 -47875
rect 87110 -47979 87144 -47945
rect 87194 -47841 87228 -47807
rect 87194 -47909 87228 -47875
rect 87278 -47841 87312 -47807
rect 87278 -47909 87312 -47875
rect 87278 -47979 87312 -47945
rect 87362 -47841 87396 -47807
rect 87362 -47909 87396 -47875
rect 87446 -47841 87480 -47807
rect 87446 -47909 87480 -47875
rect 87446 -47979 87480 -47945
rect 87530 -47841 87564 -47807
rect 87530 -47909 87564 -47875
rect 87614 -47841 87648 -47807
rect 87614 -47909 87648 -47875
rect 87614 -47979 87648 -47945
rect 87698 -47841 87732 -47807
rect 87698 -47909 87732 -47875
rect 87782 -47841 87816 -47807
rect 87782 -47909 87816 -47875
rect 87782 -47979 87816 -47945
rect 87866 -47841 87900 -47807
rect 87866 -47909 87900 -47875
rect 87950 -47841 87984 -47807
rect 87950 -47909 87984 -47875
rect 87950 -47979 87984 -47945
rect 88034 -47841 88068 -47807
rect 88034 -47909 88068 -47875
rect 88118 -47841 88152 -47807
rect 88118 -47909 88152 -47875
rect 88118 -47979 88152 -47945
rect 88202 -47841 88236 -47807
rect 88202 -47909 88236 -47875
rect 88286 -47841 88320 -47807
rect 88286 -47909 88320 -47875
rect 88286 -47979 88320 -47945
rect 88370 -47841 88404 -47807
rect 88370 -47909 88404 -47875
rect 88498 -47841 88532 -47807
rect 88498 -47909 88532 -47875
rect 88498 -47979 88532 -47945
rect 88582 -47841 88616 -47807
rect 88582 -47909 88616 -47875
rect 88582 -47979 88616 -47945
rect 88666 -47841 88700 -47807
rect 88666 -47909 88700 -47875
rect 88750 -47841 88784 -47807
rect 88750 -47909 88784 -47875
rect 88750 -47979 88784 -47945
rect 88834 -47841 88868 -47807
rect 88834 -47909 88868 -47875
rect 88918 -47841 88952 -47807
rect 88918 -47909 88952 -47875
rect 88918 -47979 88952 -47945
rect 89002 -47841 89036 -47807
rect 89002 -47909 89036 -47875
rect 89086 -47841 89120 -47807
rect 89086 -47909 89120 -47875
rect 89086 -47979 89120 -47945
rect 89170 -47841 89204 -47807
rect 89170 -47909 89204 -47875
rect 89254 -47841 89288 -47807
rect 89254 -47909 89288 -47875
rect 89254 -47979 89288 -47945
rect 89338 -47841 89372 -47807
rect 89338 -47909 89372 -47875
rect 89422 -47841 89456 -47807
rect 89422 -47909 89456 -47875
rect 89422 -47979 89456 -47945
rect 89506 -47841 89540 -47807
rect 89506 -47909 89540 -47875
rect 89590 -47841 89624 -47807
rect 89590 -47909 89624 -47875
rect 89590 -47979 89624 -47945
rect 89674 -47841 89708 -47807
rect 89674 -47909 89708 -47875
rect 89758 -47841 89792 -47807
rect 89758 -47909 89792 -47875
rect 89758 -47979 89792 -47945
rect 89842 -47841 89876 -47807
rect 89842 -47909 89876 -47875
rect 89970 -47841 90004 -47807
rect 89970 -47909 90004 -47875
rect 89970 -47979 90004 -47945
rect 90054 -47841 90088 -47807
rect 90054 -47909 90088 -47875
rect 90054 -47979 90088 -47945
rect 90138 -47841 90172 -47807
rect 90138 -47909 90172 -47875
rect 90222 -47841 90256 -47807
rect 90222 -47909 90256 -47875
rect 90222 -47979 90256 -47945
rect 90306 -47841 90340 -47807
rect 90306 -47909 90340 -47875
rect 90390 -47841 90424 -47807
rect 90390 -47909 90424 -47875
rect 90390 -47979 90424 -47945
rect 90474 -47841 90508 -47807
rect 90474 -47909 90508 -47875
rect 90558 -47841 90592 -47807
rect 90558 -47909 90592 -47875
rect 90558 -47979 90592 -47945
rect 90642 -47841 90676 -47807
rect 90642 -47909 90676 -47875
rect 90726 -47841 90760 -47807
rect 90726 -47909 90760 -47875
rect 90726 -47979 90760 -47945
rect 90810 -47841 90844 -47807
rect 90810 -47909 90844 -47875
rect 90894 -47841 90928 -47807
rect 90894 -47909 90928 -47875
rect 90894 -47979 90928 -47945
rect 90978 -47841 91012 -47807
rect 90978 -47909 91012 -47875
rect 91062 -47841 91096 -47807
rect 91062 -47909 91096 -47875
rect 91062 -47979 91096 -47945
rect 91146 -47841 91180 -47807
rect 91146 -47909 91180 -47875
rect 91230 -47841 91264 -47807
rect 91230 -47909 91264 -47875
rect 91230 -47979 91264 -47945
rect 91314 -47841 91348 -47807
rect 91314 -47909 91348 -47875
rect 77613 -48082 77647 -48048
rect 77974 -48145 78008 -48111
rect 77974 -48213 78008 -48179
rect 78059 -48114 78093 -48080
rect 78059 -48182 78093 -48148
rect 77649 -48483 77683 -48449
rect 77733 -48483 77767 -48449
rect 77841 -48441 77875 -48407
rect 77841 -48509 77875 -48475
rect 77945 -48441 77979 -48407
rect 77945 -48509 77979 -48475
rect 77649 -49411 77683 -49377
rect 77733 -49411 77767 -49377
rect 77841 -49385 77875 -49351
rect 77841 -49453 77875 -49419
rect 78073 -49322 78107 -49288
rect 77945 -49385 77979 -49351
rect 78434 -49385 78468 -49351
rect 77945 -49453 77979 -49419
rect 78434 -49453 78468 -49419
rect 78519 -49354 78553 -49320
rect 78519 -49422 78553 -49388
rect 77649 -49723 77683 -49689
rect 77733 -49723 77767 -49689
rect 77841 -49681 77875 -49647
rect 77841 -49749 77875 -49715
rect 77945 -49681 77979 -49647
rect 77945 -49749 77979 -49715
rect 54091 -50306 54867 -50272
rect 54091 -50434 54867 -50400
rect 54091 -50662 54867 -50628
rect 54091 -50790 54867 -50756
rect 57131 -50763 57165 -50729
rect 57131 -50831 57165 -50797
rect 57217 -50763 57251 -50729
rect 57217 -50831 57251 -50797
rect 57303 -50763 57337 -50729
rect 57303 -50844 57337 -50810
rect 59125 -50681 59501 -50647
rect 59125 -50789 59501 -50755
rect 59125 -50897 59501 -50863
rect 77651 -50665 77685 -50631
rect 77735 -50665 77769 -50631
rect 77843 -50639 77877 -50605
rect 77843 -50707 77877 -50673
rect 77947 -50639 77981 -50605
rect 77947 -50707 77981 -50673
rect 54081 -52622 54857 -52588
rect 54081 -52750 54857 -52716
rect 56430 -52075 56464 -51299
rect 56558 -52075 56592 -51299
rect 59044 -51547 59078 -51171
rect 59162 -51547 59196 -51171
rect 77613 -50931 77647 -50897
rect 77705 -50939 77739 -50905
rect 77807 -50931 77841 -50897
rect 77902 -50939 77936 -50905
rect 78053 -50931 78087 -50897
rect 78053 -50999 78087 -50965
rect 78153 -50931 78187 -50897
rect 78718 -50931 78752 -50897
rect 78153 -50999 78187 -50965
rect 78718 -50999 78752 -50965
rect 78153 -51067 78187 -51033
rect 78357 -51062 78391 -51028
rect 78803 -50962 78837 -50928
rect 78803 -51030 78837 -50996
rect 60459 -51607 60493 -51573
rect 60527 -51607 60561 -51573
rect 60595 -51607 60629 -51573
rect 60823 -51607 60857 -51573
rect 60891 -51607 60925 -51573
rect 60959 -51607 60993 -51573
rect 60459 -51691 60493 -51657
rect 60527 -51691 60561 -51657
rect 60595 -51691 60629 -51657
rect 60823 -51691 60857 -51657
rect 60891 -51691 60925 -51657
rect 60959 -51691 60993 -51657
rect 59044 -52277 59078 -51901
rect 59162 -52277 59196 -51901
rect 83083 -51507 83117 -51473
rect 82914 -51627 82948 -51593
rect 83083 -51575 83117 -51541
rect 83183 -51491 83217 -51457
rect 83183 -51559 83217 -51525
rect 83374 -51491 83408 -51457
rect 83374 -51559 83408 -51525
rect 83374 -51627 83408 -51593
rect 83458 -51491 83492 -51457
rect 83458 -51559 83492 -51525
rect 83458 -51627 83492 -51593
rect 83619 -51491 83653 -51457
rect 83619 -51559 83653 -51525
rect 83619 -51627 83653 -51593
rect 83703 -51491 83737 -51457
rect 83703 -51559 83737 -51525
rect 83703 -51627 83737 -51593
rect 83787 -51491 83821 -51457
rect 83787 -51559 83821 -51525
rect 83871 -51491 83905 -51457
rect 83871 -51559 83905 -51525
rect 83871 -51627 83905 -51593
rect 83955 -51491 83989 -51457
rect 84082 -51491 84116 -51457
rect 84082 -51559 84116 -51525
rect 84082 -51629 84116 -51595
rect 84166 -51491 84200 -51457
rect 84166 -51559 84200 -51525
rect 84166 -51629 84200 -51595
rect 84250 -51491 84284 -51457
rect 84250 -51559 84284 -51525
rect 84334 -51491 84368 -51457
rect 84334 -51559 84368 -51525
rect 84334 -51629 84368 -51595
rect 84418 -51491 84452 -51457
rect 84418 -51559 84452 -51525
rect 84502 -51491 84536 -51457
rect 84502 -51559 84536 -51525
rect 84502 -51629 84536 -51595
rect 84586 -51491 84620 -51457
rect 84586 -51559 84620 -51525
rect 84670 -51491 84704 -51457
rect 84670 -51559 84704 -51525
rect 84670 -51629 84704 -51595
rect 84754 -51491 84788 -51457
rect 84754 -51559 84788 -51525
rect 84838 -51491 84872 -51457
rect 84838 -51559 84872 -51525
rect 84838 -51629 84872 -51595
rect 84922 -51491 84956 -51457
rect 84922 -51559 84956 -51525
rect 85006 -51491 85040 -51457
rect 85006 -51559 85040 -51525
rect 85006 -51629 85040 -51595
rect 85090 -51491 85124 -51457
rect 85090 -51559 85124 -51525
rect 85174 -51491 85208 -51457
rect 85174 -51559 85208 -51525
rect 85174 -51629 85208 -51595
rect 85258 -51491 85292 -51457
rect 85258 -51559 85292 -51525
rect 85342 -51491 85376 -51457
rect 85342 -51559 85376 -51525
rect 85342 -51629 85376 -51595
rect 85426 -51491 85460 -51457
rect 85426 -51559 85460 -51525
rect 85554 -51491 85588 -51457
rect 85554 -51559 85588 -51525
rect 85554 -51629 85588 -51595
rect 85638 -51491 85672 -51457
rect 85638 -51559 85672 -51525
rect 85638 -51629 85672 -51595
rect 85722 -51491 85756 -51457
rect 85722 -51559 85756 -51525
rect 85806 -51491 85840 -51457
rect 85806 -51559 85840 -51525
rect 85806 -51629 85840 -51595
rect 85890 -51491 85924 -51457
rect 85890 -51559 85924 -51525
rect 85974 -51491 86008 -51457
rect 85974 -51559 86008 -51525
rect 85974 -51629 86008 -51595
rect 86058 -51491 86092 -51457
rect 86058 -51559 86092 -51525
rect 86142 -51491 86176 -51457
rect 86142 -51559 86176 -51525
rect 86142 -51629 86176 -51595
rect 86226 -51491 86260 -51457
rect 86226 -51559 86260 -51525
rect 86310 -51491 86344 -51457
rect 86310 -51559 86344 -51525
rect 86310 -51629 86344 -51595
rect 86394 -51491 86428 -51457
rect 86394 -51559 86428 -51525
rect 86478 -51491 86512 -51457
rect 86478 -51559 86512 -51525
rect 86478 -51629 86512 -51595
rect 86562 -51491 86596 -51457
rect 86562 -51559 86596 -51525
rect 86646 -51491 86680 -51457
rect 86646 -51559 86680 -51525
rect 86646 -51629 86680 -51595
rect 86730 -51491 86764 -51457
rect 86730 -51559 86764 -51525
rect 86814 -51491 86848 -51457
rect 86814 -51559 86848 -51525
rect 86814 -51629 86848 -51595
rect 86898 -51491 86932 -51457
rect 86898 -51559 86932 -51525
rect 87026 -51491 87060 -51457
rect 87026 -51559 87060 -51525
rect 87026 -51629 87060 -51595
rect 87110 -51491 87144 -51457
rect 87110 -51559 87144 -51525
rect 87110 -51629 87144 -51595
rect 87194 -51491 87228 -51457
rect 87194 -51559 87228 -51525
rect 87278 -51491 87312 -51457
rect 87278 -51559 87312 -51525
rect 87278 -51629 87312 -51595
rect 87362 -51491 87396 -51457
rect 87362 -51559 87396 -51525
rect 87446 -51491 87480 -51457
rect 87446 -51559 87480 -51525
rect 87446 -51629 87480 -51595
rect 87530 -51491 87564 -51457
rect 87530 -51559 87564 -51525
rect 87614 -51491 87648 -51457
rect 87614 -51559 87648 -51525
rect 87614 -51629 87648 -51595
rect 87698 -51491 87732 -51457
rect 87698 -51559 87732 -51525
rect 87782 -51491 87816 -51457
rect 87782 -51559 87816 -51525
rect 87782 -51629 87816 -51595
rect 87866 -51491 87900 -51457
rect 87866 -51559 87900 -51525
rect 87950 -51491 87984 -51457
rect 87950 -51559 87984 -51525
rect 87950 -51629 87984 -51595
rect 88034 -51491 88068 -51457
rect 88034 -51559 88068 -51525
rect 88118 -51491 88152 -51457
rect 88118 -51559 88152 -51525
rect 88118 -51629 88152 -51595
rect 88202 -51491 88236 -51457
rect 88202 -51559 88236 -51525
rect 88286 -51491 88320 -51457
rect 88286 -51559 88320 -51525
rect 88286 -51629 88320 -51595
rect 88370 -51491 88404 -51457
rect 88370 -51559 88404 -51525
rect 88498 -51491 88532 -51457
rect 88498 -51559 88532 -51525
rect 88498 -51629 88532 -51595
rect 88582 -51491 88616 -51457
rect 88582 -51559 88616 -51525
rect 88582 -51629 88616 -51595
rect 88666 -51491 88700 -51457
rect 88666 -51559 88700 -51525
rect 88750 -51491 88784 -51457
rect 88750 -51559 88784 -51525
rect 88750 -51629 88784 -51595
rect 88834 -51491 88868 -51457
rect 88834 -51559 88868 -51525
rect 88918 -51491 88952 -51457
rect 88918 -51559 88952 -51525
rect 88918 -51629 88952 -51595
rect 89002 -51491 89036 -51457
rect 89002 -51559 89036 -51525
rect 89086 -51491 89120 -51457
rect 89086 -51559 89120 -51525
rect 89086 -51629 89120 -51595
rect 89170 -51491 89204 -51457
rect 89170 -51559 89204 -51525
rect 89254 -51491 89288 -51457
rect 89254 -51559 89288 -51525
rect 89254 -51629 89288 -51595
rect 89338 -51491 89372 -51457
rect 89338 -51559 89372 -51525
rect 89422 -51491 89456 -51457
rect 89422 -51559 89456 -51525
rect 89422 -51629 89456 -51595
rect 89506 -51491 89540 -51457
rect 89506 -51559 89540 -51525
rect 89590 -51491 89624 -51457
rect 89590 -51559 89624 -51525
rect 89590 -51629 89624 -51595
rect 89674 -51491 89708 -51457
rect 89674 -51559 89708 -51525
rect 89758 -51491 89792 -51457
rect 89758 -51559 89792 -51525
rect 89758 -51629 89792 -51595
rect 89842 -51491 89876 -51457
rect 89842 -51559 89876 -51525
rect 89970 -51491 90004 -51457
rect 89970 -51559 90004 -51525
rect 89970 -51629 90004 -51595
rect 90054 -51491 90088 -51457
rect 90054 -51559 90088 -51525
rect 90054 -51629 90088 -51595
rect 90138 -51491 90172 -51457
rect 90138 -51559 90172 -51525
rect 90222 -51491 90256 -51457
rect 90222 -51559 90256 -51525
rect 90222 -51629 90256 -51595
rect 90306 -51491 90340 -51457
rect 90306 -51559 90340 -51525
rect 90390 -51491 90424 -51457
rect 90390 -51559 90424 -51525
rect 90390 -51629 90424 -51595
rect 90474 -51491 90508 -51457
rect 90474 -51559 90508 -51525
rect 90558 -51491 90592 -51457
rect 90558 -51559 90592 -51525
rect 90558 -51629 90592 -51595
rect 90642 -51491 90676 -51457
rect 90642 -51559 90676 -51525
rect 90726 -51491 90760 -51457
rect 90726 -51559 90760 -51525
rect 90726 -51629 90760 -51595
rect 90810 -51491 90844 -51457
rect 90810 -51559 90844 -51525
rect 90894 -51491 90928 -51457
rect 90894 -51559 90928 -51525
rect 90894 -51629 90928 -51595
rect 90978 -51491 91012 -51457
rect 90978 -51559 91012 -51525
rect 91062 -51491 91096 -51457
rect 91062 -51559 91096 -51525
rect 91062 -51629 91096 -51595
rect 91146 -51491 91180 -51457
rect 91146 -51559 91180 -51525
rect 91230 -51491 91264 -51457
rect 91230 -51559 91264 -51525
rect 91230 -51629 91264 -51595
rect 91314 -51491 91348 -51457
rect 91314 -51559 91348 -51525
rect 60527 -51775 60561 -51741
rect 60595 -51775 60629 -51741
rect 60823 -51775 60857 -51741
rect 60891 -51775 60925 -51741
rect 60459 -51859 60493 -51825
rect 60527 -51859 60561 -51825
rect 60595 -51859 60629 -51825
rect 60823 -51859 60857 -51825
rect 60891 -51859 60925 -51825
rect 60959 -51859 60993 -51825
rect 60595 -51943 60629 -51909
rect 60823 -51943 60857 -51909
rect 77613 -51939 77647 -51905
rect 77705 -51931 77739 -51897
rect 77807 -51939 77841 -51905
rect 77902 -51931 77936 -51897
rect 78053 -51871 78087 -51837
rect 78053 -51939 78087 -51905
rect 78153 -51803 78187 -51769
rect 78153 -51871 78187 -51837
rect 78153 -51939 78187 -51905
rect 77613 -52163 77647 -52129
rect 77705 -52171 77739 -52137
rect 77807 -52163 77841 -52129
rect 77902 -52171 77936 -52137
rect 78053 -52163 78087 -52129
rect 57131 -52591 57165 -52557
rect 57131 -52659 57165 -52625
rect 57217 -52591 57251 -52557
rect 57217 -52659 57251 -52625
rect 57303 -52578 57337 -52544
rect 57303 -52659 57337 -52625
rect 59125 -52588 59501 -52554
rect 59125 -52696 59501 -52662
rect 59125 -52804 59501 -52770
rect 54081 -52978 54857 -52944
rect 54081 -53106 54857 -53072
rect 78053 -52231 78087 -52197
rect 78153 -52163 78187 -52129
rect 78153 -52231 78187 -52197
rect 78153 -52299 78187 -52265
rect 77613 -53173 77647 -53139
rect 77705 -53165 77739 -53131
rect 77807 -53173 77841 -53139
rect 77902 -53165 77936 -53131
rect 78053 -53105 78087 -53071
rect 78053 -53173 78087 -53139
rect 78153 -53037 78187 -53003
rect 78153 -53105 78187 -53071
rect 78153 -53173 78187 -53139
rect 77885 -53401 77919 -53367
rect 77613 -53540 77647 -53506
rect 77697 -53510 77731 -53476
rect 77790 -53529 77824 -53495
rect 77969 -53415 78003 -53381
rect 77969 -53483 78003 -53449
rect 78109 -53443 78143 -53409
rect 78193 -53443 78227 -53409
rect 78301 -53401 78335 -53367
rect 78301 -53469 78335 -53435
rect 78405 -53401 78439 -53367
rect 78894 -53401 78928 -53367
rect 78405 -53469 78439 -53435
rect 78894 -53469 78928 -53435
rect 78533 -53532 78567 -53498
rect 78979 -53432 79013 -53398
rect 78979 -53500 79013 -53466
rect 54091 -55706 54867 -55672
rect 54091 -55834 54867 -55800
rect 54091 -56062 54867 -56028
rect 54091 -56190 54867 -56156
rect 57131 -56163 57165 -56129
rect 57131 -56231 57165 -56197
rect 57217 -56163 57251 -56129
rect 57217 -56231 57251 -56197
rect 57303 -56163 57337 -56129
rect 57303 -56244 57337 -56210
rect 59125 -56081 59501 -56047
rect 59125 -56189 59501 -56155
rect 59125 -56297 59501 -56263
rect 54081 -58022 54857 -57988
rect 54081 -58150 54857 -58116
rect 56430 -57475 56464 -56699
rect 56558 -57475 56592 -56699
rect 59044 -56947 59078 -56571
rect 59162 -56947 59196 -56571
rect 60459 -57007 60493 -56973
rect 60527 -57007 60561 -56973
rect 60595 -57007 60629 -56973
rect 60823 -57007 60857 -56973
rect 60891 -57007 60925 -56973
rect 60959 -57007 60993 -56973
rect 60459 -57091 60493 -57057
rect 60527 -57091 60561 -57057
rect 60595 -57091 60629 -57057
rect 60823 -57091 60857 -57057
rect 60891 -57091 60925 -57057
rect 60959 -57091 60993 -57057
rect 59044 -57677 59078 -57301
rect 59162 -57677 59196 -57301
rect 60527 -57175 60561 -57141
rect 60595 -57175 60629 -57141
rect 60823 -57175 60857 -57141
rect 60891 -57175 60925 -57141
rect 60459 -57259 60493 -57225
rect 60527 -57259 60561 -57225
rect 60595 -57259 60629 -57225
rect 60823 -57259 60857 -57225
rect 60891 -57259 60925 -57225
rect 60959 -57259 60993 -57225
rect 60595 -57343 60629 -57309
rect 60823 -57343 60857 -57309
rect 57131 -57991 57165 -57957
rect 57131 -58059 57165 -58025
rect 57217 -57991 57251 -57957
rect 57217 -58059 57251 -58025
rect 57303 -57978 57337 -57944
rect 57303 -58059 57337 -58025
rect 59125 -57988 59501 -57954
rect 59125 -58096 59501 -58062
rect 59125 -58204 59501 -58170
rect 54081 -58378 54857 -58344
rect 54081 -58506 54857 -58472
rect 54091 -61106 54867 -61072
rect 54091 -61234 54867 -61200
rect 54091 -61462 54867 -61428
rect 54091 -61590 54867 -61556
rect 57131 -61563 57165 -61529
rect 57131 -61631 57165 -61597
rect 57217 -61563 57251 -61529
rect 57217 -61631 57251 -61597
rect 57303 -61563 57337 -61529
rect 57303 -61644 57337 -61610
rect 59125 -61481 59501 -61447
rect 59125 -61589 59501 -61555
rect 59125 -61697 59501 -61663
rect 54081 -63422 54857 -63388
rect 54081 -63550 54857 -63516
rect 56430 -62875 56464 -62099
rect 56558 -62875 56592 -62099
rect 59044 -62347 59078 -61971
rect 59162 -62347 59196 -61971
rect 60459 -62407 60493 -62373
rect 60527 -62407 60561 -62373
rect 60595 -62407 60629 -62373
rect 60823 -62407 60857 -62373
rect 60891 -62407 60925 -62373
rect 60959 -62407 60993 -62373
rect 60459 -62491 60493 -62457
rect 60527 -62491 60561 -62457
rect 60595 -62491 60629 -62457
rect 60823 -62491 60857 -62457
rect 60891 -62491 60925 -62457
rect 60959 -62491 60993 -62457
rect 59044 -63077 59078 -62701
rect 59162 -63077 59196 -62701
rect 60527 -62575 60561 -62541
rect 60595 -62575 60629 -62541
rect 60823 -62575 60857 -62541
rect 60891 -62575 60925 -62541
rect 60459 -62659 60493 -62625
rect 60527 -62659 60561 -62625
rect 60595 -62659 60629 -62625
rect 60823 -62659 60857 -62625
rect 60891 -62659 60925 -62625
rect 60959 -62659 60993 -62625
rect 60595 -62743 60629 -62709
rect 60823 -62743 60857 -62709
rect 57131 -63391 57165 -63357
rect 57131 -63459 57165 -63425
rect 57217 -63391 57251 -63357
rect 57217 -63459 57251 -63425
rect 57303 -63378 57337 -63344
rect 57303 -63459 57337 -63425
rect 59125 -63388 59501 -63354
rect 59125 -63496 59501 -63462
rect 59125 -63604 59501 -63570
rect 54081 -63778 54857 -63744
rect 54081 -63906 54857 -63872
rect 54091 -66506 54867 -66472
rect 54091 -66634 54867 -66600
rect 54091 -66862 54867 -66828
rect 54091 -66990 54867 -66956
rect 57131 -66963 57165 -66929
rect 57131 -67031 57165 -66997
rect 57217 -66963 57251 -66929
rect 57217 -67031 57251 -66997
rect 57303 -66963 57337 -66929
rect 57303 -67044 57337 -67010
rect 59125 -66881 59501 -66847
rect 59125 -66989 59501 -66955
rect 59125 -67097 59501 -67063
rect 54081 -68822 54857 -68788
rect 54081 -68950 54857 -68916
rect 56430 -68275 56464 -67499
rect 56558 -68275 56592 -67499
rect 59044 -67747 59078 -67371
rect 59162 -67747 59196 -67371
rect 60459 -67807 60493 -67773
rect 60527 -67807 60561 -67773
rect 60595 -67807 60629 -67773
rect 60823 -67807 60857 -67773
rect 60891 -67807 60925 -67773
rect 60959 -67807 60993 -67773
rect 60459 -67891 60493 -67857
rect 60527 -67891 60561 -67857
rect 60595 -67891 60629 -67857
rect 60823 -67891 60857 -67857
rect 60891 -67891 60925 -67857
rect 60959 -67891 60993 -67857
rect 59044 -68477 59078 -68101
rect 59162 -68477 59196 -68101
rect 60527 -67975 60561 -67941
rect 60595 -67975 60629 -67941
rect 60823 -67975 60857 -67941
rect 60891 -67975 60925 -67941
rect 60459 -68059 60493 -68025
rect 60527 -68059 60561 -68025
rect 60595 -68059 60629 -68025
rect 60823 -68059 60857 -68025
rect 60891 -68059 60925 -68025
rect 60959 -68059 60993 -68025
rect 60595 -68143 60629 -68109
rect 60823 -68143 60857 -68109
rect 57131 -68791 57165 -68757
rect 57131 -68859 57165 -68825
rect 57217 -68791 57251 -68757
rect 57217 -68859 57251 -68825
rect 57303 -68778 57337 -68744
rect 57303 -68859 57337 -68825
rect 59125 -68788 59501 -68754
rect 59125 -68896 59501 -68862
rect 59125 -69004 59501 -68970
rect 54081 -69178 54857 -69144
rect 54081 -69306 54857 -69272
rect 54091 -71906 54867 -71872
rect 54091 -72034 54867 -72000
rect 54091 -72262 54867 -72228
rect 54091 -72390 54867 -72356
rect 57131 -72363 57165 -72329
rect 57131 -72431 57165 -72397
rect 57217 -72363 57251 -72329
rect 57217 -72431 57251 -72397
rect 57303 -72363 57337 -72329
rect 57303 -72444 57337 -72410
rect 59125 -72281 59501 -72247
rect 59125 -72389 59501 -72355
rect 59125 -72497 59501 -72463
rect 54081 -74222 54857 -74188
rect 54081 -74350 54857 -74316
rect 56430 -73675 56464 -72899
rect 56558 -73675 56592 -72899
rect 59044 -73147 59078 -72771
rect 59162 -73147 59196 -72771
rect 60459 -73207 60493 -73173
rect 60527 -73207 60561 -73173
rect 60595 -73207 60629 -73173
rect 60823 -73207 60857 -73173
rect 60891 -73207 60925 -73173
rect 60959 -73207 60993 -73173
rect 60459 -73291 60493 -73257
rect 60527 -73291 60561 -73257
rect 60595 -73291 60629 -73257
rect 60823 -73291 60857 -73257
rect 60891 -73291 60925 -73257
rect 60959 -73291 60993 -73257
rect 59044 -73877 59078 -73501
rect 59162 -73877 59196 -73501
rect 60527 -73375 60561 -73341
rect 60595 -73375 60629 -73341
rect 60823 -73375 60857 -73341
rect 60891 -73375 60925 -73341
rect 60459 -73459 60493 -73425
rect 60527 -73459 60561 -73425
rect 60595 -73459 60629 -73425
rect 60823 -73459 60857 -73425
rect 60891 -73459 60925 -73425
rect 60959 -73459 60993 -73425
rect 60595 -73543 60629 -73509
rect 60823 -73543 60857 -73509
rect 57131 -74191 57165 -74157
rect 57131 -74259 57165 -74225
rect 57217 -74191 57251 -74157
rect 57217 -74259 57251 -74225
rect 57303 -74178 57337 -74144
rect 57303 -74259 57337 -74225
rect 59125 -74188 59501 -74154
rect 59125 -74296 59501 -74262
rect 59125 -74404 59501 -74370
rect 54081 -74578 54857 -74544
rect 54081 -74706 54857 -74672
rect 54091 -77306 54867 -77272
rect 54091 -77434 54867 -77400
rect 54091 -77662 54867 -77628
rect 54091 -77790 54867 -77756
rect 57131 -77763 57165 -77729
rect 57131 -77831 57165 -77797
rect 57217 -77763 57251 -77729
rect 57217 -77831 57251 -77797
rect 57303 -77763 57337 -77729
rect 57303 -77844 57337 -77810
rect 59125 -77681 59501 -77647
rect 59125 -77789 59501 -77755
rect 59125 -77897 59501 -77863
rect 54081 -79622 54857 -79588
rect 54081 -79750 54857 -79716
rect 56430 -79075 56464 -78299
rect 56558 -79075 56592 -78299
rect 59044 -78547 59078 -78171
rect 59162 -78547 59196 -78171
rect 60459 -78607 60493 -78573
rect 60527 -78607 60561 -78573
rect 60595 -78607 60629 -78573
rect 60823 -78607 60857 -78573
rect 60891 -78607 60925 -78573
rect 60959 -78607 60993 -78573
rect 60459 -78691 60493 -78657
rect 60527 -78691 60561 -78657
rect 60595 -78691 60629 -78657
rect 60823 -78691 60857 -78657
rect 60891 -78691 60925 -78657
rect 60959 -78691 60993 -78657
rect 59044 -79277 59078 -78901
rect 59162 -79277 59196 -78901
rect 60527 -78775 60561 -78741
rect 60595 -78775 60629 -78741
rect 60823 -78775 60857 -78741
rect 60891 -78775 60925 -78741
rect 60459 -78859 60493 -78825
rect 60527 -78859 60561 -78825
rect 60595 -78859 60629 -78825
rect 60823 -78859 60857 -78825
rect 60891 -78859 60925 -78825
rect 60959 -78859 60993 -78825
rect 60595 -78943 60629 -78909
rect 60823 -78943 60857 -78909
rect 57131 -79591 57165 -79557
rect 57131 -79659 57165 -79625
rect 57217 -79591 57251 -79557
rect 57217 -79659 57251 -79625
rect 57303 -79578 57337 -79544
rect 57303 -79659 57337 -79625
rect 59125 -79588 59501 -79554
rect 59125 -79696 59501 -79662
rect 59125 -79804 59501 -79770
rect 54081 -79978 54857 -79944
rect 54081 -80106 54857 -80072
rect 54091 -82706 54867 -82672
rect 54091 -82834 54867 -82800
rect 54091 -83062 54867 -83028
rect 54091 -83190 54867 -83156
rect 57131 -83163 57165 -83129
rect 57131 -83231 57165 -83197
rect 57217 -83163 57251 -83129
rect 57217 -83231 57251 -83197
rect 57303 -83163 57337 -83129
rect 57303 -83244 57337 -83210
rect 59125 -83081 59501 -83047
rect 59125 -83189 59501 -83155
rect 59125 -83297 59501 -83263
rect 54081 -85022 54857 -84988
rect 54081 -85150 54857 -85116
rect 56430 -84475 56464 -83699
rect 56558 -84475 56592 -83699
rect 59044 -83947 59078 -83571
rect 59162 -83947 59196 -83571
rect 60459 -84007 60493 -83973
rect 60527 -84007 60561 -83973
rect 60595 -84007 60629 -83973
rect 60823 -84007 60857 -83973
rect 60891 -84007 60925 -83973
rect 60959 -84007 60993 -83973
rect 60459 -84091 60493 -84057
rect 60527 -84091 60561 -84057
rect 60595 -84091 60629 -84057
rect 60823 -84091 60857 -84057
rect 60891 -84091 60925 -84057
rect 60959 -84091 60993 -84057
rect 59044 -84677 59078 -84301
rect 59162 -84677 59196 -84301
rect 60527 -84175 60561 -84141
rect 60595 -84175 60629 -84141
rect 60823 -84175 60857 -84141
rect 60891 -84175 60925 -84141
rect 60459 -84259 60493 -84225
rect 60527 -84259 60561 -84225
rect 60595 -84259 60629 -84225
rect 60823 -84259 60857 -84225
rect 60891 -84259 60925 -84225
rect 60959 -84259 60993 -84225
rect 60595 -84343 60629 -84309
rect 60823 -84343 60857 -84309
rect 57131 -84991 57165 -84957
rect 57131 -85059 57165 -85025
rect 57217 -84991 57251 -84957
rect 57217 -85059 57251 -85025
rect 57303 -84978 57337 -84944
rect 57303 -85059 57337 -85025
rect 59125 -84988 59501 -84954
rect 59125 -85096 59501 -85062
rect 59125 -85204 59501 -85170
rect 54081 -85378 54857 -85344
rect 54081 -85506 54857 -85472
<< psubdiff >>
rect 53350 -2038 53790 -2004
rect 53350 -2100 53384 -2038
rect 53756 -2664 53790 -2038
rect 55706 -1988 55802 -1954
rect 56050 -1988 56146 -1954
rect 55706 -2050 55740 -1988
rect 55176 -2100 55272 -2066
rect 55430 -2100 55526 -2066
rect 55176 -2162 55210 -2100
rect 55492 -2162 55526 -2100
rect 55176 -2518 55210 -2456
rect 55492 -2518 55526 -2456
rect 54870 -2552 55272 -2518
rect 55430 -2552 55706 -2518
rect 54870 -2558 55706 -2552
rect 54870 -2664 54904 -2558
rect 53756 -2698 53852 -2664
rect 54808 -2698 54904 -2664
rect 53756 -2760 53790 -2698
rect 54870 -2760 54904 -2698
rect 53756 -3070 53790 -3008
rect 54870 -3068 54904 -3008
rect 55700 -3006 55706 -2558
rect 56112 -2050 56146 -1988
rect 55700 -3068 55740 -3006
rect 59772 -2294 59868 -2260
rect 60424 -2294 60520 -2260
rect 59772 -2356 59806 -2294
rect 56112 -3068 56146 -3006
rect 54870 -3070 55160 -3068
rect 53756 -3104 53852 -3070
rect 54808 -3104 55160 -3070
rect 53756 -3166 53790 -3104
rect 54870 -3108 55160 -3104
rect 55600 -3102 55802 -3068
rect 56050 -3102 56146 -3068
rect 55600 -3108 55740 -3102
rect 54870 -3166 54904 -3108
rect 53756 -3476 53790 -3414
rect 55700 -3164 55740 -3108
rect 54870 -3476 54904 -3414
rect 53756 -3510 53852 -3476
rect 54808 -3510 54904 -3476
rect 53350 -4136 53384 -4074
rect 53756 -4136 53790 -3510
rect 54870 -3618 54904 -3510
rect 55700 -3618 55706 -3164
rect 54870 -3624 55706 -3618
rect 54870 -3658 55262 -3624
rect 55420 -3658 55706 -3624
rect 55166 -3720 55200 -3658
rect 53350 -4170 53446 -4136
rect 53694 -4170 53790 -4136
rect 55482 -3720 55516 -3658
rect 55166 -4076 55200 -4014
rect 55482 -4076 55516 -4014
rect 55166 -4110 55262 -4076
rect 55420 -4110 55516 -4076
rect 56112 -3164 56146 -3102
rect 55706 -4182 55740 -4120
rect 57086 -2710 57376 -2680
rect 57086 -2780 57116 -2710
rect 57346 -2780 57376 -2710
rect 57086 -2810 57376 -2780
rect 60486 -2356 60520 -2294
rect 59772 -2596 59806 -2534
rect 60486 -2596 60520 -2534
rect 59388 -2630 59484 -2596
rect 59642 -2630 59800 -2596
rect 59958 -2630 60520 -2596
rect 59388 -2692 59422 -2630
rect 59388 -3109 59422 -3048
rect 59704 -3109 59738 -2630
rect 60020 -2692 60054 -2630
rect 61186 -2800 61286 -2790
rect 61186 -2820 61366 -2800
rect 61186 -2860 61216 -2820
rect 61336 -2860 61366 -2820
rect 61186 -2880 61366 -2860
rect 61186 -2890 61286 -2880
rect 60020 -3109 60054 -3048
rect 57056 -3370 57416 -3340
rect 57056 -3450 57096 -3370
rect 57376 -3450 57416 -3370
rect 57056 -3480 57416 -3450
rect 59387 -3144 60054 -3109
rect 59387 -3205 59421 -3144
rect 59387 -3623 59421 -3561
rect 59703 -3623 59737 -3144
rect 60019 -3205 60053 -3144
rect 60019 -3623 60053 -3561
rect 59387 -3657 59483 -3623
rect 59641 -3657 59799 -3623
rect 59957 -3626 60053 -3623
rect 59957 -3657 60520 -3626
rect 59772 -3660 60520 -3657
rect 59772 -3722 59806 -3660
rect 56112 -4182 56146 -4120
rect 55706 -4216 55802 -4182
rect 56050 -4216 56146 -4182
rect 60486 -3722 60520 -3660
rect 59772 -3962 59806 -3900
rect 60486 -3962 60520 -3900
rect 59772 -3996 59868 -3962
rect 60424 -3996 60520 -3962
rect 55176 -4478 55272 -4444
rect 55566 -4478 55662 -4444
rect 55176 -4540 55210 -4478
rect 55628 -4540 55662 -4478
rect 55176 -4760 55210 -4698
rect 55628 -4760 55662 -4698
rect 55176 -4794 55272 -4760
rect 55566 -4794 55662 -4760
rect 53350 -7438 53790 -7404
rect 53350 -7500 53384 -7438
rect 53756 -8064 53790 -7438
rect 55706 -7388 55802 -7354
rect 56050 -7388 56146 -7354
rect 55706 -7450 55740 -7388
rect 55176 -7500 55272 -7466
rect 55430 -7500 55526 -7466
rect 55176 -7562 55210 -7500
rect 55492 -7562 55526 -7500
rect 55176 -7918 55210 -7856
rect 55492 -7918 55526 -7856
rect 54870 -7952 55272 -7918
rect 55430 -7952 55706 -7918
rect 54870 -7958 55706 -7952
rect 54870 -8064 54904 -7958
rect 53756 -8098 53852 -8064
rect 54808 -8098 54904 -8064
rect 53756 -8160 53790 -8098
rect 54870 -8160 54904 -8098
rect 53756 -8470 53790 -8408
rect 54870 -8468 54904 -8408
rect 55700 -8406 55706 -7958
rect 56112 -7450 56146 -7388
rect 55700 -8468 55740 -8406
rect 59772 -7694 59868 -7660
rect 60424 -7694 60520 -7660
rect 59772 -7756 59806 -7694
rect 56112 -8468 56146 -8406
rect 54870 -8470 55160 -8468
rect 53756 -8504 53852 -8470
rect 54808 -8504 55160 -8470
rect 53756 -8566 53790 -8504
rect 54870 -8508 55160 -8504
rect 55600 -8502 55802 -8468
rect 56050 -8502 56146 -8468
rect 55600 -8508 55740 -8502
rect 54870 -8566 54904 -8508
rect 53756 -8876 53790 -8814
rect 55700 -8564 55740 -8508
rect 54870 -8876 54904 -8814
rect 53756 -8910 53852 -8876
rect 54808 -8910 54904 -8876
rect 53350 -9536 53384 -9474
rect 53756 -9536 53790 -8910
rect 54870 -9018 54904 -8910
rect 55700 -9018 55706 -8564
rect 54870 -9024 55706 -9018
rect 54870 -9058 55262 -9024
rect 55420 -9058 55706 -9024
rect 55166 -9120 55200 -9058
rect 53350 -9570 53446 -9536
rect 53694 -9570 53790 -9536
rect 55482 -9120 55516 -9058
rect 55166 -9476 55200 -9414
rect 55482 -9476 55516 -9414
rect 55166 -9510 55262 -9476
rect 55420 -9510 55516 -9476
rect 56112 -8564 56146 -8502
rect 55706 -9582 55740 -9520
rect 57086 -8110 57376 -8080
rect 57086 -8180 57116 -8110
rect 57346 -8180 57376 -8110
rect 57086 -8210 57376 -8180
rect 60486 -7756 60520 -7694
rect 59772 -7996 59806 -7934
rect 60486 -7996 60520 -7934
rect 59388 -8030 59484 -7996
rect 59642 -8030 59800 -7996
rect 59958 -8030 60520 -7996
rect 59388 -8092 59422 -8030
rect 59388 -8509 59422 -8448
rect 59704 -8509 59738 -8030
rect 60020 -8092 60054 -8030
rect 61186 -8200 61286 -8190
rect 61186 -8220 61366 -8200
rect 61186 -8260 61216 -8220
rect 61336 -8260 61366 -8220
rect 61186 -8280 61366 -8260
rect 61186 -8290 61286 -8280
rect 60020 -8509 60054 -8448
rect 57056 -8770 57416 -8740
rect 57056 -8850 57096 -8770
rect 57376 -8850 57416 -8770
rect 57056 -8880 57416 -8850
rect 59387 -8544 60054 -8509
rect 59387 -8605 59421 -8544
rect 59387 -9023 59421 -8961
rect 59703 -9023 59737 -8544
rect 60019 -8605 60053 -8544
rect 60019 -9023 60053 -8961
rect 59387 -9057 59483 -9023
rect 59641 -9057 59799 -9023
rect 59957 -9026 60053 -9023
rect 59957 -9057 60520 -9026
rect 59772 -9060 60520 -9057
rect 59772 -9122 59806 -9060
rect 56112 -9582 56146 -9520
rect 55706 -9616 55802 -9582
rect 56050 -9616 56146 -9582
rect 60486 -9122 60520 -9060
rect 59772 -9362 59806 -9300
rect 60486 -9362 60520 -9300
rect 59772 -9396 59868 -9362
rect 60424 -9396 60520 -9362
rect 55176 -9878 55272 -9844
rect 55566 -9878 55662 -9844
rect 55176 -9940 55210 -9878
rect 55628 -9940 55662 -9878
rect 55176 -10160 55210 -10098
rect 55628 -10160 55662 -10098
rect 55176 -10194 55272 -10160
rect 55566 -10194 55662 -10160
rect 20156 -11850 20252 -11816
rect 20430 -11850 20526 -11816
rect 20156 -11912 20190 -11850
rect 20492 -11912 20526 -11850
rect 20156 -12132 20190 -12070
rect 20492 -12132 20526 -12070
rect 20156 -12143 20526 -12132
rect 16439 -12177 16535 -12143
rect 16783 -12177 16941 -12143
rect 17189 -12177 17347 -12143
rect 17595 -12177 17753 -12143
rect 18001 -12177 18159 -12143
rect 18407 -12177 18565 -12143
rect 18813 -12177 18971 -12143
rect 19219 -12177 19377 -12143
rect 19625 -12177 19783 -12143
rect 20031 -12177 20189 -12143
rect 20437 -12177 20595 -12143
rect 20843 -12177 21001 -12143
rect 21249 -12177 21407 -12143
rect 21655 -12177 21813 -12143
rect 22061 -12177 22219 -12143
rect 22467 -12177 22625 -12143
rect 22873 -12177 23031 -12143
rect 23279 -12177 23437 -12143
rect 23685 -12177 23843 -12143
rect 24091 -12177 24249 -12143
rect 24497 -12177 24655 -12143
rect 24903 -12177 25061 -12143
rect 25309 -12177 25405 -12143
rect 16439 -12239 16473 -12177
rect 16845 -12239 16879 -12177
rect 16439 -13257 16473 -13195
rect 17251 -12239 17285 -12177
rect 16845 -13257 16879 -13195
rect 17657 -12239 17691 -12177
rect 17251 -13257 17285 -13195
rect 18063 -12239 18097 -12177
rect 17657 -13257 17691 -13195
rect 18469 -12239 18503 -12177
rect 18063 -13257 18097 -13195
rect 18875 -12239 18909 -12177
rect 18469 -13257 18503 -13195
rect 19281 -12239 19315 -12177
rect 18875 -13257 18909 -13195
rect 19687 -12239 19721 -12177
rect 19281 -13257 19315 -13195
rect 20093 -12239 20127 -12177
rect 19687 -13257 19721 -13195
rect 20499 -12239 20533 -12177
rect 20093 -13257 20127 -13195
rect 20905 -12239 20939 -12177
rect 20499 -13257 20533 -13195
rect 21311 -12239 21345 -12177
rect 20905 -13257 20939 -13195
rect 21717 -12239 21751 -12177
rect 21311 -13257 21345 -13195
rect 22123 -12239 22157 -12177
rect 21717 -13257 21751 -13195
rect 22529 -12239 22563 -12177
rect 22123 -13257 22157 -13195
rect 22935 -12239 22969 -12177
rect 22529 -13257 22563 -13195
rect 23341 -12239 23375 -12177
rect 22935 -13257 22969 -13195
rect 23747 -12239 23781 -12177
rect 23341 -13257 23375 -13195
rect 24153 -12239 24187 -12177
rect 23747 -13257 23781 -13195
rect 24559 -12239 24593 -12177
rect 24153 -13257 24187 -13195
rect 24965 -12239 24999 -12177
rect 24559 -13257 24593 -13195
rect 25371 -12239 25405 -12177
rect 24965 -13257 24999 -13195
rect 25371 -13257 25405 -13195
rect 16439 -13291 16535 -13257
rect 16783 -13291 16941 -13257
rect 17189 -13291 17347 -13257
rect 17595 -13291 17753 -13257
rect 18001 -13291 18159 -13257
rect 18407 -13291 18565 -13257
rect 18813 -13291 18971 -13257
rect 19219 -13291 19377 -13257
rect 19625 -13291 19783 -13257
rect 20031 -13291 20189 -13257
rect 20437 -13291 20595 -13257
rect 20843 -13291 21001 -13257
rect 21249 -13291 21407 -13257
rect 21655 -13291 21813 -13257
rect 22061 -13291 22219 -13257
rect 22467 -13291 22625 -13257
rect 22873 -13291 23031 -13257
rect 23279 -13291 23437 -13257
rect 23685 -13291 23843 -13257
rect 24091 -13291 24249 -13257
rect 24497 -13291 24655 -13257
rect 24903 -13291 25061 -13257
rect 25309 -13291 25405 -13257
rect 53350 -12838 53790 -12804
rect 53350 -12900 53384 -12838
rect 16436 -13420 16532 -13386
rect 34620 -13420 34716 -13386
rect 16436 -13482 16470 -13420
rect 34682 -13482 34716 -13420
rect 16436 -14758 16470 -14696
rect 34682 -14758 34716 -14696
rect 16436 -14792 16532 -14758
rect 34620 -14792 34716 -14758
rect 16436 -14854 16470 -14792
rect 34682 -14854 34716 -14792
rect 16436 -16130 16470 -16068
rect 53756 -13464 53790 -12838
rect 55706 -12788 55802 -12754
rect 56050 -12788 56146 -12754
rect 55706 -12850 55740 -12788
rect 55176 -12900 55272 -12866
rect 55430 -12900 55526 -12866
rect 55176 -12962 55210 -12900
rect 55492 -12962 55526 -12900
rect 55176 -13318 55210 -13256
rect 55492 -13318 55526 -13256
rect 54870 -13352 55272 -13318
rect 55430 -13352 55706 -13318
rect 54870 -13358 55706 -13352
rect 54870 -13464 54904 -13358
rect 53756 -13498 53852 -13464
rect 54808 -13498 54904 -13464
rect 53756 -13560 53790 -13498
rect 54870 -13560 54904 -13498
rect 53756 -13870 53790 -13808
rect 54870 -13868 54904 -13808
rect 55700 -13806 55706 -13358
rect 56112 -12850 56146 -12788
rect 55700 -13868 55740 -13806
rect 59772 -13094 59868 -13060
rect 60424 -13094 60520 -13060
rect 59772 -13156 59806 -13094
rect 56112 -13868 56146 -13806
rect 54870 -13870 55160 -13868
rect 53756 -13904 53852 -13870
rect 54808 -13904 55160 -13870
rect 53756 -13966 53790 -13904
rect 54870 -13908 55160 -13904
rect 55600 -13902 55802 -13868
rect 56050 -13902 56146 -13868
rect 55600 -13908 55740 -13902
rect 54870 -13966 54904 -13908
rect 53756 -14276 53790 -14214
rect 55700 -13964 55740 -13908
rect 54870 -14276 54904 -14214
rect 53756 -14310 53852 -14276
rect 54808 -14310 54904 -14276
rect 53350 -14936 53384 -14874
rect 53756 -14936 53790 -14310
rect 54870 -14418 54904 -14310
rect 55700 -14418 55706 -13964
rect 54870 -14424 55706 -14418
rect 54870 -14458 55262 -14424
rect 55420 -14458 55706 -14424
rect 55166 -14520 55200 -14458
rect 53350 -14970 53446 -14936
rect 53694 -14970 53790 -14936
rect 55482 -14520 55516 -14458
rect 55166 -14876 55200 -14814
rect 55482 -14876 55516 -14814
rect 55166 -14910 55262 -14876
rect 55420 -14910 55516 -14876
rect 56112 -13964 56146 -13902
rect 55706 -14982 55740 -14920
rect 57086 -13510 57376 -13480
rect 57086 -13580 57116 -13510
rect 57346 -13580 57376 -13510
rect 57086 -13610 57376 -13580
rect 60486 -13156 60520 -13094
rect 59772 -13396 59806 -13334
rect 60486 -13396 60520 -13334
rect 59388 -13430 59484 -13396
rect 59642 -13430 59800 -13396
rect 59958 -13430 60520 -13396
rect 59388 -13492 59422 -13430
rect 59388 -13909 59422 -13848
rect 59704 -13909 59738 -13430
rect 60020 -13492 60054 -13430
rect 61186 -13600 61286 -13590
rect 61186 -13620 61366 -13600
rect 61186 -13660 61216 -13620
rect 61336 -13660 61366 -13620
rect 61186 -13680 61366 -13660
rect 61186 -13690 61286 -13680
rect 60020 -13909 60054 -13848
rect 57056 -14170 57416 -14140
rect 57056 -14250 57096 -14170
rect 57376 -14250 57416 -14170
rect 57056 -14280 57416 -14250
rect 59387 -13944 60054 -13909
rect 59387 -14005 59421 -13944
rect 59387 -14423 59421 -14361
rect 59703 -14423 59737 -13944
rect 60019 -14005 60053 -13944
rect 60019 -14423 60053 -14361
rect 59387 -14457 59483 -14423
rect 59641 -14457 59799 -14423
rect 59957 -14426 60053 -14423
rect 59957 -14457 60520 -14426
rect 59772 -14460 60520 -14457
rect 59772 -14522 59806 -14460
rect 56112 -14982 56146 -14920
rect 55706 -15016 55802 -14982
rect 56050 -15016 56146 -14982
rect 60486 -14522 60520 -14460
rect 59772 -14762 59806 -14700
rect 60486 -14762 60520 -14700
rect 59772 -14796 59868 -14762
rect 60424 -14796 60520 -14762
rect 55176 -15278 55272 -15244
rect 55566 -15278 55662 -15244
rect 55176 -15340 55210 -15278
rect 55628 -15340 55662 -15278
rect 55176 -15560 55210 -15498
rect 55628 -15560 55662 -15498
rect 55176 -15594 55272 -15560
rect 55566 -15594 55662 -15560
rect 34682 -16130 34716 -16068
rect 16436 -16164 16532 -16130
rect 34620 -16164 34716 -16130
rect 53350 -18238 53790 -18204
rect 53350 -18300 53384 -18238
rect 53756 -18864 53790 -18238
rect 55706 -18188 55802 -18154
rect 56050 -18188 56146 -18154
rect 55706 -18250 55740 -18188
rect 55176 -18300 55272 -18266
rect 55430 -18300 55526 -18266
rect 55176 -18362 55210 -18300
rect 55492 -18362 55526 -18300
rect 55176 -18718 55210 -18656
rect 55492 -18718 55526 -18656
rect 54870 -18752 55272 -18718
rect 55430 -18752 55706 -18718
rect 54870 -18758 55706 -18752
rect 54870 -18864 54904 -18758
rect 53756 -18898 53852 -18864
rect 54808 -18898 54904 -18864
rect 53756 -18960 53790 -18898
rect 54870 -18960 54904 -18898
rect 53756 -19270 53790 -19208
rect 54870 -19268 54904 -19208
rect 55700 -19206 55706 -18758
rect 56112 -18250 56146 -18188
rect 55700 -19268 55740 -19206
rect 59772 -18494 59868 -18460
rect 60424 -18494 60520 -18460
rect 59772 -18556 59806 -18494
rect 56112 -19268 56146 -19206
rect 54870 -19270 55160 -19268
rect 53756 -19304 53852 -19270
rect 54808 -19304 55160 -19270
rect 53756 -19366 53790 -19304
rect 54870 -19308 55160 -19304
rect 55600 -19302 55802 -19268
rect 56050 -19302 56146 -19268
rect 55600 -19308 55740 -19302
rect 54870 -19366 54904 -19308
rect 53756 -19676 53790 -19614
rect 55700 -19364 55740 -19308
rect 54870 -19676 54904 -19614
rect 53756 -19710 53852 -19676
rect 54808 -19710 54904 -19676
rect 53350 -20336 53384 -20274
rect 53756 -20336 53790 -19710
rect 54870 -19818 54904 -19710
rect 55700 -19818 55706 -19364
rect 54870 -19824 55706 -19818
rect 54870 -19858 55262 -19824
rect 55420 -19858 55706 -19824
rect 55166 -19920 55200 -19858
rect 53350 -20370 53446 -20336
rect 53694 -20370 53790 -20336
rect 55482 -19920 55516 -19858
rect 55166 -20276 55200 -20214
rect 55482 -20276 55516 -20214
rect 55166 -20310 55262 -20276
rect 55420 -20310 55516 -20276
rect 56112 -19364 56146 -19302
rect 55706 -20382 55740 -20320
rect 57086 -18910 57376 -18880
rect 57086 -18980 57116 -18910
rect 57346 -18980 57376 -18910
rect 57086 -19010 57376 -18980
rect 60486 -18556 60520 -18494
rect 59772 -18796 59806 -18734
rect 60486 -18796 60520 -18734
rect 59388 -18830 59484 -18796
rect 59642 -18830 59800 -18796
rect 59958 -18830 60520 -18796
rect 59388 -18892 59422 -18830
rect 59388 -19309 59422 -19248
rect 59704 -19309 59738 -18830
rect 60020 -18892 60054 -18830
rect 61186 -19000 61286 -18990
rect 61186 -19020 61366 -19000
rect 61186 -19060 61216 -19020
rect 61336 -19060 61366 -19020
rect 61186 -19080 61366 -19060
rect 61186 -19090 61286 -19080
rect 60020 -19309 60054 -19248
rect 57056 -19570 57416 -19540
rect 57056 -19650 57096 -19570
rect 57376 -19650 57416 -19570
rect 57056 -19680 57416 -19650
rect 59387 -19344 60054 -19309
rect 59387 -19405 59421 -19344
rect 59387 -19823 59421 -19761
rect 59703 -19823 59737 -19344
rect 60019 -19405 60053 -19344
rect 60019 -19823 60053 -19761
rect 59387 -19857 59483 -19823
rect 59641 -19857 59799 -19823
rect 59957 -19826 60053 -19823
rect 59957 -19857 60520 -19826
rect 59772 -19860 60520 -19857
rect 59772 -19922 59806 -19860
rect 56112 -20382 56146 -20320
rect 55706 -20416 55802 -20382
rect 56050 -20416 56146 -20382
rect 60486 -19922 60520 -19860
rect 59772 -20162 59806 -20100
rect 60486 -20162 60520 -20100
rect 59772 -20196 59868 -20162
rect 60424 -20196 60520 -20162
rect 55176 -20678 55272 -20644
rect 55566 -20678 55662 -20644
rect 55176 -20740 55210 -20678
rect 55628 -20740 55662 -20678
rect 55176 -20960 55210 -20898
rect 55628 -20960 55662 -20898
rect 55176 -20994 55272 -20960
rect 55566 -20994 55662 -20960
rect 53350 -23638 53790 -23604
rect 53350 -23700 53384 -23638
rect 53756 -24264 53790 -23638
rect 55706 -23588 55802 -23554
rect 56050 -23588 56146 -23554
rect 55706 -23650 55740 -23588
rect 55176 -23700 55272 -23666
rect 55430 -23700 55526 -23666
rect 55176 -23762 55210 -23700
rect 55492 -23762 55526 -23700
rect 55176 -24118 55210 -24056
rect 55492 -24118 55526 -24056
rect 54870 -24152 55272 -24118
rect 55430 -24152 55706 -24118
rect 54870 -24158 55706 -24152
rect 54870 -24264 54904 -24158
rect 53756 -24298 53852 -24264
rect 54808 -24298 54904 -24264
rect 53756 -24360 53790 -24298
rect 54870 -24360 54904 -24298
rect 53756 -24670 53790 -24608
rect 54870 -24668 54904 -24608
rect 55700 -24606 55706 -24158
rect 56112 -23650 56146 -23588
rect 55700 -24668 55740 -24606
rect 59772 -23894 59868 -23860
rect 60424 -23894 60520 -23860
rect 59772 -23956 59806 -23894
rect 56112 -24668 56146 -24606
rect 54870 -24670 55160 -24668
rect 53756 -24704 53852 -24670
rect 54808 -24704 55160 -24670
rect 53756 -24766 53790 -24704
rect 54870 -24708 55160 -24704
rect 55600 -24702 55802 -24668
rect 56050 -24702 56146 -24668
rect 55600 -24708 55740 -24702
rect 54870 -24766 54904 -24708
rect 53756 -25076 53790 -25014
rect 55700 -24764 55740 -24708
rect 54870 -25076 54904 -25014
rect 53756 -25110 53852 -25076
rect 54808 -25110 54904 -25076
rect 53350 -25736 53384 -25674
rect 53756 -25736 53790 -25110
rect 54870 -25218 54904 -25110
rect 55700 -25218 55706 -24764
rect 54870 -25224 55706 -25218
rect 54870 -25258 55262 -25224
rect 55420 -25258 55706 -25224
rect 55166 -25320 55200 -25258
rect 53350 -25770 53446 -25736
rect 53694 -25770 53790 -25736
rect 55482 -25320 55516 -25258
rect 55166 -25676 55200 -25614
rect 55482 -25676 55516 -25614
rect 55166 -25710 55262 -25676
rect 55420 -25710 55516 -25676
rect 56112 -24764 56146 -24702
rect 55706 -25782 55740 -25720
rect 57086 -24310 57376 -24280
rect 57086 -24380 57116 -24310
rect 57346 -24380 57376 -24310
rect 57086 -24410 57376 -24380
rect 60486 -23956 60520 -23894
rect 59772 -24196 59806 -24134
rect 60486 -24196 60520 -24134
rect 59388 -24230 59484 -24196
rect 59642 -24230 59800 -24196
rect 59958 -24230 60520 -24196
rect 59388 -24292 59422 -24230
rect 59388 -24709 59422 -24648
rect 59704 -24709 59738 -24230
rect 60020 -24292 60054 -24230
rect 61186 -24400 61286 -24390
rect 61186 -24420 61366 -24400
rect 61186 -24460 61216 -24420
rect 61336 -24460 61366 -24420
rect 61186 -24480 61366 -24460
rect 61186 -24490 61286 -24480
rect 60020 -24709 60054 -24648
rect 57056 -24970 57416 -24940
rect 57056 -25050 57096 -24970
rect 57376 -25050 57416 -24970
rect 57056 -25080 57416 -25050
rect 59387 -24744 60054 -24709
rect 59387 -24805 59421 -24744
rect 59387 -25223 59421 -25161
rect 59703 -25223 59737 -24744
rect 60019 -24805 60053 -24744
rect 60019 -25223 60053 -25161
rect 59387 -25257 59483 -25223
rect 59641 -25257 59799 -25223
rect 59957 -25226 60053 -25223
rect 59957 -25257 60520 -25226
rect 59772 -25260 60520 -25257
rect 59772 -25322 59806 -25260
rect 56112 -25782 56146 -25720
rect 55706 -25816 55802 -25782
rect 56050 -25816 56146 -25782
rect 60486 -25322 60520 -25260
rect 59772 -25562 59806 -25500
rect 60486 -25562 60520 -25500
rect 59772 -25596 59868 -25562
rect 60424 -25596 60520 -25562
rect 55176 -26078 55272 -26044
rect 55566 -26078 55662 -26044
rect 55176 -26140 55210 -26078
rect 55628 -26140 55662 -26078
rect 55176 -26360 55210 -26298
rect 55628 -26360 55662 -26298
rect 55176 -26394 55272 -26360
rect 55566 -26394 55662 -26360
rect 53350 -29038 53790 -29004
rect 53350 -29100 53384 -29038
rect 25738 -31032 35838 -30998
rect 25738 -31094 25772 -31032
rect 35804 -31094 35838 -31032
rect 25738 -32592 25772 -32530
rect 53756 -29664 53790 -29038
rect 55706 -28988 55802 -28954
rect 56050 -28988 56146 -28954
rect 55706 -29050 55740 -28988
rect 55176 -29100 55272 -29066
rect 55430 -29100 55526 -29066
rect 55176 -29162 55210 -29100
rect 55492 -29162 55526 -29100
rect 55176 -29518 55210 -29456
rect 55492 -29518 55526 -29456
rect 54870 -29552 55272 -29518
rect 55430 -29552 55706 -29518
rect 54870 -29558 55706 -29552
rect 54870 -29664 54904 -29558
rect 53756 -29698 53852 -29664
rect 54808 -29698 54904 -29664
rect 53756 -29760 53790 -29698
rect 54870 -29760 54904 -29698
rect 53756 -30070 53790 -30008
rect 54870 -30068 54904 -30008
rect 55700 -30006 55706 -29558
rect 56112 -29050 56146 -28988
rect 55700 -30068 55740 -30006
rect 59772 -29294 59868 -29260
rect 60424 -29294 60520 -29260
rect 59772 -29356 59806 -29294
rect 56112 -30068 56146 -30006
rect 54870 -30070 55160 -30068
rect 53756 -30104 53852 -30070
rect 54808 -30104 55160 -30070
rect 53756 -30166 53790 -30104
rect 54870 -30108 55160 -30104
rect 55600 -30102 55802 -30068
rect 56050 -30102 56146 -30068
rect 55600 -30108 55740 -30102
rect 54870 -30166 54904 -30108
rect 53756 -30476 53790 -30414
rect 55700 -30164 55740 -30108
rect 54870 -30476 54904 -30414
rect 53756 -30510 53852 -30476
rect 54808 -30510 54904 -30476
rect 53350 -31136 53384 -31074
rect 53756 -31136 53790 -30510
rect 54870 -30618 54904 -30510
rect 55700 -30618 55706 -30164
rect 54870 -30624 55706 -30618
rect 54870 -30658 55262 -30624
rect 55420 -30658 55706 -30624
rect 55166 -30720 55200 -30658
rect 53350 -31170 53446 -31136
rect 53694 -31170 53790 -31136
rect 55482 -30720 55516 -30658
rect 55166 -31076 55200 -31014
rect 55482 -31076 55516 -31014
rect 55166 -31110 55262 -31076
rect 55420 -31110 55516 -31076
rect 56112 -30164 56146 -30102
rect 55706 -31182 55740 -31120
rect 57086 -29710 57376 -29680
rect 57086 -29780 57116 -29710
rect 57346 -29780 57376 -29710
rect 57086 -29810 57376 -29780
rect 60486 -29356 60520 -29294
rect 59772 -29596 59806 -29534
rect 60486 -29596 60520 -29534
rect 59388 -29630 59484 -29596
rect 59642 -29630 59800 -29596
rect 59958 -29630 60520 -29596
rect 59388 -29692 59422 -29630
rect 59388 -30109 59422 -30048
rect 59704 -30109 59738 -29630
rect 60020 -29692 60054 -29630
rect 61186 -29800 61286 -29790
rect 61186 -29820 61366 -29800
rect 61186 -29860 61216 -29820
rect 61336 -29860 61366 -29820
rect 61186 -29880 61366 -29860
rect 61186 -29890 61286 -29880
rect 60020 -30109 60054 -30048
rect 57056 -30370 57416 -30340
rect 57056 -30450 57096 -30370
rect 57376 -30450 57416 -30370
rect 57056 -30480 57416 -30450
rect 59387 -30144 60054 -30109
rect 59387 -30205 59421 -30144
rect 59387 -30623 59421 -30561
rect 59703 -30623 59737 -30144
rect 60019 -30205 60053 -30144
rect 60019 -30623 60053 -30561
rect 59387 -30657 59483 -30623
rect 59641 -30657 59799 -30623
rect 59957 -30626 60053 -30623
rect 59957 -30657 60520 -30626
rect 59772 -30660 60520 -30657
rect 59772 -30722 59806 -30660
rect 56112 -31182 56146 -31120
rect 55706 -31216 55802 -31182
rect 56050 -31216 56146 -31182
rect 60486 -30722 60520 -30660
rect 59772 -30962 59806 -30900
rect 60486 -30962 60520 -30900
rect 59772 -30996 59868 -30962
rect 60424 -30996 60520 -30962
rect 55176 -31478 55272 -31444
rect 55566 -31478 55662 -31444
rect 55176 -31540 55210 -31478
rect 55628 -31540 55662 -31478
rect 55176 -31760 55210 -31698
rect 55628 -31760 55662 -31698
rect 55176 -31794 55272 -31760
rect 55566 -31794 55662 -31760
rect 35804 -32592 35838 -32530
rect 25738 -32596 35838 -32592
rect 25736 -32626 35838 -32596
rect 25736 -32630 35836 -32626
rect 25736 -32692 25770 -32630
rect 35802 -32692 35836 -32630
rect 25736 -34190 25770 -34128
rect 35802 -34190 35836 -34128
rect 25736 -34228 35836 -34190
rect 25736 -34290 25770 -34228
rect 35802 -34290 35836 -34228
rect 25736 -35788 25770 -35726
rect 35802 -35788 35836 -35726
rect 25736 -35830 35836 -35788
rect 25736 -35892 25770 -35830
rect 35802 -35892 35836 -35830
rect 25736 -37390 25770 -37328
rect 53350 -34438 53790 -34404
rect 53350 -34500 53384 -34438
rect 53756 -35064 53790 -34438
rect 55706 -34388 55802 -34354
rect 56050 -34388 56146 -34354
rect 55706 -34450 55740 -34388
rect 55176 -34500 55272 -34466
rect 55430 -34500 55526 -34466
rect 55176 -34562 55210 -34500
rect 55492 -34562 55526 -34500
rect 55176 -34918 55210 -34856
rect 55492 -34918 55526 -34856
rect 54870 -34952 55272 -34918
rect 55430 -34952 55706 -34918
rect 54870 -34958 55706 -34952
rect 54870 -35064 54904 -34958
rect 53756 -35098 53852 -35064
rect 54808 -35098 54904 -35064
rect 53756 -35160 53790 -35098
rect 54870 -35160 54904 -35098
rect 53756 -35470 53790 -35408
rect 54870 -35468 54904 -35408
rect 55700 -35406 55706 -34958
rect 56112 -34450 56146 -34388
rect 55700 -35468 55740 -35406
rect 59772 -34694 59868 -34660
rect 60424 -34694 60520 -34660
rect 59772 -34756 59806 -34694
rect 56112 -35468 56146 -35406
rect 54870 -35470 55160 -35468
rect 53756 -35504 53852 -35470
rect 54808 -35504 55160 -35470
rect 53756 -35566 53790 -35504
rect 54870 -35508 55160 -35504
rect 55600 -35502 55802 -35468
rect 56050 -35502 56146 -35468
rect 55600 -35508 55740 -35502
rect 54870 -35566 54904 -35508
rect 53756 -35876 53790 -35814
rect 55700 -35564 55740 -35508
rect 54870 -35876 54904 -35814
rect 53756 -35910 53852 -35876
rect 54808 -35910 54904 -35876
rect 53350 -36536 53384 -36474
rect 53756 -36536 53790 -35910
rect 54870 -36018 54904 -35910
rect 55700 -36018 55706 -35564
rect 54870 -36024 55706 -36018
rect 54870 -36058 55262 -36024
rect 55420 -36058 55706 -36024
rect 55166 -36120 55200 -36058
rect 53350 -36570 53446 -36536
rect 53694 -36570 53790 -36536
rect 55482 -36120 55516 -36058
rect 55166 -36476 55200 -36414
rect 55482 -36476 55516 -36414
rect 55166 -36510 55262 -36476
rect 55420 -36510 55516 -36476
rect 56112 -35564 56146 -35502
rect 55706 -36582 55740 -36520
rect 57086 -35110 57376 -35080
rect 57086 -35180 57116 -35110
rect 57346 -35180 57376 -35110
rect 57086 -35210 57376 -35180
rect 60486 -34756 60520 -34694
rect 59772 -34996 59806 -34934
rect 60486 -34996 60520 -34934
rect 59388 -35030 59484 -34996
rect 59642 -35030 59800 -34996
rect 59958 -35030 60520 -34996
rect 59388 -35092 59422 -35030
rect 59388 -35509 59422 -35448
rect 59704 -35509 59738 -35030
rect 60020 -35092 60054 -35030
rect 61186 -35200 61286 -35190
rect 61186 -35220 61366 -35200
rect 61186 -35260 61216 -35220
rect 61336 -35260 61366 -35220
rect 61186 -35280 61366 -35260
rect 61186 -35290 61286 -35280
rect 60020 -35509 60054 -35448
rect 57056 -35770 57416 -35740
rect 57056 -35850 57096 -35770
rect 57376 -35850 57416 -35770
rect 57056 -35880 57416 -35850
rect 59387 -35544 60054 -35509
rect 59387 -35605 59421 -35544
rect 59387 -36023 59421 -35961
rect 59703 -36023 59737 -35544
rect 60019 -35605 60053 -35544
rect 60019 -36023 60053 -35961
rect 59387 -36057 59483 -36023
rect 59641 -36057 59799 -36023
rect 59957 -36026 60053 -36023
rect 59957 -36057 60520 -36026
rect 59772 -36060 60520 -36057
rect 59772 -36122 59806 -36060
rect 56112 -36582 56146 -36520
rect 55706 -36616 55802 -36582
rect 56050 -36616 56146 -36582
rect 60486 -36122 60520 -36060
rect 59772 -36362 59806 -36300
rect 60486 -36362 60520 -36300
rect 59772 -36396 59868 -36362
rect 60424 -36396 60520 -36362
rect 55176 -36878 55272 -36844
rect 55566 -36878 55662 -36844
rect 55176 -36940 55210 -36878
rect 55628 -36940 55662 -36878
rect 55176 -37160 55210 -37098
rect 55628 -37160 55662 -37098
rect 55176 -37194 55272 -37160
rect 55566 -37194 55662 -37160
rect 35802 -37390 35836 -37328
rect 25736 -37430 35836 -37390
rect 25736 -37492 25770 -37430
rect 35802 -37492 35836 -37430
rect 25736 -38990 25770 -38928
rect 77110 -38370 77220 -38350
rect 77110 -38420 77140 -38370
rect 77190 -38420 77220 -38370
rect 77110 -38490 77220 -38420
rect 77110 -38540 77140 -38490
rect 77190 -38540 77220 -38490
rect 77110 -38570 77220 -38540
rect 35802 -38990 35836 -38928
rect 25736 -38998 35836 -38990
rect 25736 -39024 35838 -38998
rect 25738 -39032 35838 -39024
rect 25738 -39094 25772 -39032
rect 35804 -39094 35838 -39032
rect 25738 -40592 25772 -40530
rect 77420 -39490 77540 -39460
rect 77420 -39550 77450 -39490
rect 77510 -39550 77540 -39490
rect 77420 -39580 77540 -39550
rect 35804 -40592 35838 -40530
rect 25738 -40596 35838 -40592
rect 25736 -40626 35838 -40596
rect 53350 -39838 53790 -39804
rect 53350 -39900 53384 -39838
rect 25736 -40630 35836 -40626
rect 25736 -40692 25770 -40630
rect 35802 -40692 35836 -40630
rect 25736 -42190 25770 -42128
rect 53756 -40464 53790 -39838
rect 55706 -39788 55802 -39754
rect 56050 -39788 56146 -39754
rect 55706 -39850 55740 -39788
rect 55176 -39900 55272 -39866
rect 55430 -39900 55526 -39866
rect 55176 -39962 55210 -39900
rect 55492 -39962 55526 -39900
rect 55176 -40318 55210 -40256
rect 55492 -40318 55526 -40256
rect 54870 -40352 55272 -40318
rect 55430 -40352 55706 -40318
rect 54870 -40358 55706 -40352
rect 54870 -40464 54904 -40358
rect 53756 -40498 53852 -40464
rect 54808 -40498 54904 -40464
rect 53756 -40560 53790 -40498
rect 54870 -40560 54904 -40498
rect 53756 -40870 53790 -40808
rect 54870 -40868 54904 -40808
rect 55700 -40806 55706 -40358
rect 56112 -39850 56146 -39788
rect 77420 -39690 77540 -39660
rect 55700 -40868 55740 -40806
rect 77420 -39750 77450 -39690
rect 77510 -39750 77540 -39690
rect 77420 -39780 77540 -39750
rect 82490 -39770 82660 -39740
rect 81590 -39800 81760 -39770
rect 81590 -39910 81620 -39800
rect 81730 -39910 81760 -39800
rect 82490 -39880 82520 -39770
rect 82630 -39880 82660 -39770
rect 82490 -39910 82660 -39880
rect 83750 -39780 83920 -39750
rect 83750 -39890 83780 -39780
rect 83890 -39890 83920 -39780
rect 81590 -39940 81760 -39910
rect 83750 -39920 83920 -39890
rect 85160 -39770 85330 -39740
rect 85160 -39880 85190 -39770
rect 85300 -39880 85330 -39770
rect 85160 -39910 85330 -39880
rect 86320 -39780 86490 -39750
rect 86320 -39890 86350 -39780
rect 86460 -39890 86490 -39780
rect 86320 -39920 86490 -39890
rect 87390 -39770 87560 -39740
rect 87390 -39880 87420 -39770
rect 87530 -39880 87560 -39770
rect 87390 -39910 87560 -39880
rect 88500 -39760 88670 -39730
rect 88500 -39870 88530 -39760
rect 88640 -39870 88670 -39760
rect 88500 -39900 88670 -39870
rect 59772 -40094 59868 -40060
rect 60424 -40094 60520 -40060
rect 59772 -40156 59806 -40094
rect 56112 -40868 56146 -40806
rect 54870 -40870 55160 -40868
rect 53756 -40904 53852 -40870
rect 54808 -40904 55160 -40870
rect 53756 -40966 53790 -40904
rect 54870 -40908 55160 -40904
rect 55600 -40902 55802 -40868
rect 56050 -40902 56146 -40868
rect 55600 -40908 55740 -40902
rect 54870 -40966 54904 -40908
rect 53756 -41276 53790 -41214
rect 55700 -40964 55740 -40908
rect 54870 -41276 54904 -41214
rect 53756 -41310 53852 -41276
rect 54808 -41310 54904 -41276
rect 53350 -41936 53384 -41874
rect 53756 -41936 53790 -41310
rect 54870 -41418 54904 -41310
rect 55700 -41418 55706 -40964
rect 54870 -41424 55706 -41418
rect 54870 -41458 55262 -41424
rect 55420 -41458 55706 -41424
rect 55166 -41520 55200 -41458
rect 53350 -41970 53446 -41936
rect 53694 -41970 53790 -41936
rect 35802 -42190 35836 -42128
rect 25736 -42228 35836 -42190
rect 25736 -42290 25770 -42228
rect 35802 -42290 35836 -42228
rect 25736 -43788 25770 -43726
rect 55482 -41520 55516 -41458
rect 55166 -41876 55200 -41814
rect 55482 -41876 55516 -41814
rect 55166 -41910 55262 -41876
rect 55420 -41910 55516 -41876
rect 56112 -40964 56146 -40902
rect 55706 -41982 55740 -41920
rect 57086 -40510 57376 -40480
rect 57086 -40580 57116 -40510
rect 57346 -40580 57376 -40510
rect 57086 -40610 57376 -40580
rect 60486 -40156 60520 -40094
rect 59772 -40396 59806 -40334
rect 60486 -40396 60520 -40334
rect 59388 -40430 59484 -40396
rect 59642 -40430 59800 -40396
rect 59958 -40430 60520 -40396
rect 59388 -40492 59422 -40430
rect 59388 -40909 59422 -40848
rect 59704 -40909 59738 -40430
rect 60020 -40492 60054 -40430
rect 61186 -40600 61286 -40590
rect 61186 -40620 61366 -40600
rect 61186 -40660 61216 -40620
rect 61336 -40660 61366 -40620
rect 61186 -40680 61366 -40660
rect 61186 -40690 61286 -40680
rect 77400 -40730 77520 -40700
rect 77400 -40790 77430 -40730
rect 77490 -40790 77520 -40730
rect 77400 -40820 77520 -40790
rect 60020 -40909 60054 -40848
rect 57056 -41170 57416 -41140
rect 57056 -41250 57096 -41170
rect 57376 -41250 57416 -41170
rect 57056 -41280 57416 -41250
rect 59387 -40944 60054 -40909
rect 59387 -41005 59421 -40944
rect 59387 -41423 59421 -41361
rect 59703 -41423 59737 -40944
rect 60019 -41005 60053 -40944
rect 77400 -40980 77520 -40950
rect 77400 -41040 77430 -40980
rect 77490 -41040 77520 -40980
rect 77400 -41070 77520 -41040
rect 60019 -41423 60053 -41361
rect 59387 -41457 59483 -41423
rect 59641 -41457 59799 -41423
rect 59957 -41426 60053 -41423
rect 59957 -41457 60520 -41426
rect 59772 -41460 60520 -41457
rect 59772 -41522 59806 -41460
rect 56112 -41982 56146 -41920
rect 55706 -42016 55802 -41982
rect 56050 -42016 56146 -41982
rect 60486 -41522 60520 -41460
rect 59772 -41762 59806 -41700
rect 60486 -41762 60520 -41700
rect 59772 -41796 59868 -41762
rect 60424 -41796 60520 -41762
rect 77420 -41990 77540 -41960
rect 77420 -42050 77450 -41990
rect 77510 -42050 77540 -41990
rect 77420 -42160 77540 -42050
rect 77420 -42220 77450 -42160
rect 77510 -42220 77540 -42160
rect 55176 -42278 55272 -42244
rect 55566 -42278 55662 -42244
rect 77420 -42250 77540 -42220
rect 55176 -42340 55210 -42278
rect 55628 -42340 55662 -42278
rect 55176 -42560 55210 -42498
rect 55628 -42560 55662 -42498
rect 55176 -42594 55272 -42560
rect 55566 -42594 55662 -42560
rect 77410 -43240 77530 -43210
rect 77410 -43300 77440 -43240
rect 77500 -43300 77530 -43240
rect 77410 -43330 77530 -43300
rect 77410 -43420 77530 -43390
rect 77410 -43480 77440 -43420
rect 77500 -43480 77530 -43420
rect 77410 -43510 77530 -43480
rect 35802 -43788 35836 -43726
rect 25736 -43830 35836 -43788
rect 25736 -43892 25770 -43830
rect 35802 -43892 35836 -43830
rect 25736 -45390 25770 -45328
rect 83480 -44240 83650 -44210
rect 77400 -44410 77520 -44380
rect 77400 -44470 77430 -44410
rect 77490 -44470 77520 -44410
rect 83480 -44350 83510 -44240
rect 83620 -44350 83650 -44240
rect 83480 -44380 83650 -44350
rect 85120 -44250 85290 -44220
rect 85120 -44360 85150 -44250
rect 85260 -44360 85290 -44250
rect 85120 -44390 85290 -44360
rect 86530 -44240 86700 -44210
rect 86530 -44350 86560 -44240
rect 86670 -44350 86700 -44240
rect 86530 -44380 86700 -44350
rect 87910 -44240 88080 -44210
rect 87910 -44350 87940 -44240
rect 88050 -44350 88080 -44240
rect 87910 -44380 88080 -44350
rect 89450 -44250 89620 -44220
rect 89450 -44360 89480 -44250
rect 89590 -44360 89620 -44250
rect 89450 -44390 89620 -44360
rect 90730 -44250 90900 -44220
rect 90730 -44360 90760 -44250
rect 90870 -44360 90900 -44250
rect 90730 -44390 90900 -44360
rect 77400 -44500 77520 -44470
rect 77400 -44660 77520 -44630
rect 77400 -44720 77430 -44660
rect 77490 -44720 77520 -44660
rect 77400 -44750 77520 -44720
rect 35802 -45390 35836 -45328
rect 25736 -45428 35836 -45390
rect 25736 -45490 25770 -45428
rect 35802 -45490 35836 -45428
rect 25736 -46988 25770 -46926
rect 35802 -46988 35836 -46926
rect 25736 -47022 35836 -46988
rect 25736 -47084 25770 -47022
rect 35802 -47084 35836 -47022
rect 25736 -48582 25770 -48520
rect 53350 -45238 53790 -45204
rect 53350 -45300 53384 -45238
rect 53756 -45864 53790 -45238
rect 55706 -45188 55802 -45154
rect 56050 -45188 56146 -45154
rect 55706 -45250 55740 -45188
rect 55176 -45300 55272 -45266
rect 55430 -45300 55526 -45266
rect 55176 -45362 55210 -45300
rect 55492 -45362 55526 -45300
rect 55176 -45718 55210 -45656
rect 55492 -45718 55526 -45656
rect 54870 -45752 55272 -45718
rect 55430 -45752 55706 -45718
rect 54870 -45758 55706 -45752
rect 54870 -45864 54904 -45758
rect 53756 -45898 53852 -45864
rect 54808 -45898 54904 -45864
rect 53756 -45960 53790 -45898
rect 54870 -45960 54904 -45898
rect 53756 -46270 53790 -46208
rect 54870 -46268 54904 -46208
rect 55700 -46206 55706 -45758
rect 56112 -45250 56146 -45188
rect 55700 -46268 55740 -46206
rect 59772 -45494 59868 -45460
rect 60424 -45494 60520 -45460
rect 59772 -45556 59806 -45494
rect 56112 -46268 56146 -46206
rect 54870 -46270 55160 -46268
rect 53756 -46304 53852 -46270
rect 54808 -46304 55160 -46270
rect 53756 -46366 53790 -46304
rect 54870 -46308 55160 -46304
rect 55600 -46302 55802 -46268
rect 56050 -46302 56146 -46268
rect 55600 -46308 55740 -46302
rect 54870 -46366 54904 -46308
rect 53756 -46676 53790 -46614
rect 55700 -46364 55740 -46308
rect 54870 -46676 54904 -46614
rect 53756 -46710 53852 -46676
rect 54808 -46710 54904 -46676
rect 53350 -47336 53384 -47274
rect 53756 -47336 53790 -46710
rect 54870 -46818 54904 -46710
rect 55700 -46818 55706 -46364
rect 54870 -46824 55706 -46818
rect 54870 -46858 55262 -46824
rect 55420 -46858 55706 -46824
rect 55166 -46920 55200 -46858
rect 53350 -47370 53446 -47336
rect 53694 -47370 53790 -47336
rect 55482 -46920 55516 -46858
rect 55166 -47276 55200 -47214
rect 55482 -47276 55516 -47214
rect 55166 -47310 55262 -47276
rect 55420 -47310 55516 -47276
rect 56112 -46364 56146 -46302
rect 55706 -47382 55740 -47320
rect 57086 -45910 57376 -45880
rect 57086 -45980 57116 -45910
rect 57346 -45980 57376 -45910
rect 57086 -46010 57376 -45980
rect 60486 -45556 60520 -45494
rect 59772 -45796 59806 -45734
rect 60486 -45796 60520 -45734
rect 77390 -45660 77510 -45630
rect 77390 -45720 77420 -45660
rect 77480 -45720 77510 -45660
rect 77390 -45750 77510 -45720
rect 59388 -45830 59484 -45796
rect 59642 -45830 59800 -45796
rect 59958 -45830 60520 -45796
rect 59388 -45892 59422 -45830
rect 59388 -46309 59422 -46248
rect 59704 -46309 59738 -45830
rect 60020 -45892 60054 -45830
rect 61186 -46000 61286 -45990
rect 61186 -46020 61366 -46000
rect 61186 -46060 61216 -46020
rect 61336 -46060 61366 -46020
rect 61186 -46080 61366 -46060
rect 61186 -46090 61286 -46080
rect 60020 -46309 60054 -46248
rect 57056 -46570 57416 -46540
rect 57056 -46650 57096 -46570
rect 57376 -46650 57416 -46570
rect 57056 -46680 57416 -46650
rect 59387 -46344 60054 -46309
rect 59387 -46405 59421 -46344
rect 59387 -46823 59421 -46761
rect 59703 -46823 59737 -46344
rect 60019 -46405 60053 -46344
rect 77110 -46410 77220 -46390
rect 77110 -46460 77140 -46410
rect 77190 -46460 77220 -46410
rect 77110 -46530 77220 -46460
rect 77110 -46580 77140 -46530
rect 77190 -46580 77220 -46530
rect 77110 -46610 77220 -46580
rect 60019 -46823 60053 -46761
rect 59387 -46857 59483 -46823
rect 59641 -46857 59799 -46823
rect 59957 -46826 60053 -46823
rect 59957 -46857 60520 -46826
rect 59772 -46860 60520 -46857
rect 59772 -46922 59806 -46860
rect 56112 -47382 56146 -47320
rect 55706 -47416 55802 -47382
rect 56050 -47416 56146 -47382
rect 60486 -46922 60520 -46860
rect 59772 -47162 59806 -47100
rect 60486 -47162 60520 -47100
rect 59772 -47196 59868 -47162
rect 60424 -47196 60520 -47162
rect 77420 -47530 77540 -47500
rect 77420 -47590 77450 -47530
rect 77510 -47590 77540 -47530
rect 77420 -47620 77540 -47590
rect 55176 -47678 55272 -47644
rect 55566 -47678 55662 -47644
rect 55176 -47740 55210 -47678
rect 55628 -47740 55662 -47678
rect 55176 -47960 55210 -47898
rect 77420 -47730 77540 -47700
rect 77420 -47790 77450 -47730
rect 77510 -47790 77540 -47730
rect 77420 -47820 77540 -47790
rect 55628 -47960 55662 -47898
rect 55176 -47994 55272 -47960
rect 55566 -47994 55662 -47960
rect 83484 -48378 83654 -48348
rect 35802 -48582 35836 -48520
rect 25736 -48586 35836 -48582
rect 25736 -48620 25832 -48586
rect 35740 -48620 35836 -48586
rect 25736 -48682 25770 -48620
rect 35802 -48682 35836 -48620
rect 25736 -50180 25770 -50118
rect 83484 -48488 83514 -48378
rect 83624 -48488 83654 -48378
rect 83484 -48518 83654 -48488
rect 85124 -48388 85294 -48358
rect 85124 -48498 85154 -48388
rect 85264 -48498 85294 -48388
rect 85124 -48528 85294 -48498
rect 86534 -48378 86704 -48348
rect 86534 -48488 86564 -48378
rect 86674 -48488 86704 -48378
rect 86534 -48518 86704 -48488
rect 87914 -48378 88084 -48348
rect 87914 -48488 87944 -48378
rect 88054 -48488 88084 -48378
rect 87914 -48518 88084 -48488
rect 89454 -48388 89624 -48358
rect 89454 -48498 89484 -48388
rect 89594 -48498 89624 -48388
rect 89454 -48528 89624 -48498
rect 90734 -48388 90904 -48358
rect 90734 -48498 90764 -48388
rect 90874 -48498 90904 -48388
rect 90734 -48528 90904 -48498
rect 77400 -48770 77520 -48740
rect 77400 -48830 77430 -48770
rect 77490 -48830 77520 -48770
rect 77400 -48860 77520 -48830
rect 77400 -49020 77520 -48990
rect 77400 -49080 77430 -49020
rect 77490 -49080 77520 -49020
rect 77400 -49110 77520 -49080
rect 35802 -50180 35836 -50118
rect 77420 -50030 77540 -50000
rect 77420 -50090 77450 -50030
rect 77510 -50090 77540 -50030
rect 25736 -50214 25832 -50180
rect 35740 -50214 35836 -50180
rect 25736 -50222 35836 -50214
rect 25736 -50284 25770 -50222
rect 35802 -50284 35836 -50222
rect 25736 -51782 25770 -51720
rect 77420 -50200 77540 -50090
rect 77420 -50260 77450 -50200
rect 77510 -50260 77540 -50200
rect 77420 -50290 77540 -50260
rect 35802 -51782 35836 -51720
rect 25736 -51820 35836 -51782
rect 25736 -51882 25770 -51820
rect 35802 -51882 35836 -51820
rect 25736 -53380 25770 -53318
rect 53350 -50638 53790 -50604
rect 53350 -50700 53384 -50638
rect 53756 -51264 53790 -50638
rect 55706 -50588 55802 -50554
rect 56050 -50588 56146 -50554
rect 55706 -50650 55740 -50588
rect 55176 -50700 55272 -50666
rect 55430 -50700 55526 -50666
rect 55176 -50762 55210 -50700
rect 55492 -50762 55526 -50700
rect 55176 -51118 55210 -51056
rect 55492 -51118 55526 -51056
rect 54870 -51152 55272 -51118
rect 55430 -51152 55706 -51118
rect 54870 -51158 55706 -51152
rect 54870 -51264 54904 -51158
rect 53756 -51298 53852 -51264
rect 54808 -51298 54904 -51264
rect 53756 -51360 53790 -51298
rect 54870 -51360 54904 -51298
rect 53756 -51670 53790 -51608
rect 54870 -51668 54904 -51608
rect 55700 -51606 55706 -51158
rect 56112 -50650 56146 -50588
rect 55700 -51668 55740 -51606
rect 59772 -50894 59868 -50860
rect 60424 -50894 60520 -50860
rect 59772 -50956 59806 -50894
rect 56112 -51668 56146 -51606
rect 54870 -51670 55160 -51668
rect 53756 -51704 53852 -51670
rect 54808 -51704 55160 -51670
rect 53756 -51766 53790 -51704
rect 54870 -51708 55160 -51704
rect 55600 -51702 55802 -51668
rect 56050 -51702 56146 -51668
rect 55600 -51708 55740 -51702
rect 54870 -51766 54904 -51708
rect 53756 -52076 53790 -52014
rect 55700 -51764 55740 -51708
rect 54870 -52076 54904 -52014
rect 53756 -52110 53852 -52076
rect 54808 -52110 54904 -52076
rect 53350 -52736 53384 -52674
rect 53756 -52736 53790 -52110
rect 54870 -52218 54904 -52110
rect 55700 -52218 55706 -51764
rect 54870 -52224 55706 -52218
rect 54870 -52258 55262 -52224
rect 55420 -52258 55706 -52224
rect 55166 -52320 55200 -52258
rect 53350 -52770 53446 -52736
rect 53694 -52770 53790 -52736
rect 55482 -52320 55516 -52258
rect 55166 -52676 55200 -52614
rect 55482 -52676 55516 -52614
rect 55166 -52710 55262 -52676
rect 55420 -52710 55516 -52676
rect 56112 -51764 56146 -51702
rect 55706 -52782 55740 -52720
rect 57086 -51310 57376 -51280
rect 57086 -51380 57116 -51310
rect 57346 -51380 57376 -51310
rect 57086 -51410 57376 -51380
rect 60486 -50956 60520 -50894
rect 59772 -51196 59806 -51134
rect 60486 -51196 60520 -51134
rect 59388 -51230 59484 -51196
rect 59642 -51230 59800 -51196
rect 59958 -51230 60520 -51196
rect 59388 -51292 59422 -51230
rect 59388 -51709 59422 -51648
rect 59704 -51709 59738 -51230
rect 60020 -51292 60054 -51230
rect 77410 -51280 77530 -51250
rect 77410 -51340 77440 -51280
rect 77500 -51340 77530 -51280
rect 77410 -51370 77530 -51340
rect 61186 -51400 61286 -51390
rect 61186 -51420 61366 -51400
rect 61186 -51460 61216 -51420
rect 61336 -51460 61366 -51420
rect 61186 -51480 61366 -51460
rect 77410 -51460 77530 -51430
rect 61186 -51490 61286 -51480
rect 77410 -51520 77440 -51460
rect 77500 -51520 77530 -51460
rect 77410 -51550 77530 -51520
rect 60020 -51709 60054 -51648
rect 57056 -51970 57416 -51940
rect 57056 -52050 57096 -51970
rect 57376 -52050 57416 -51970
rect 57056 -52080 57416 -52050
rect 59387 -51744 60054 -51709
rect 59387 -51805 59421 -51744
rect 59387 -52223 59421 -52161
rect 59703 -52223 59737 -51744
rect 60019 -51805 60053 -51744
rect 83480 -52030 83650 -52000
rect 60019 -52223 60053 -52161
rect 59387 -52257 59483 -52223
rect 59641 -52257 59799 -52223
rect 59957 -52226 60053 -52223
rect 59957 -52257 60520 -52226
rect 59772 -52260 60520 -52257
rect 59772 -52322 59806 -52260
rect 56112 -52782 56146 -52720
rect 55706 -52816 55802 -52782
rect 56050 -52816 56146 -52782
rect 60486 -52322 60520 -52260
rect 59772 -52562 59806 -52500
rect 83480 -52140 83510 -52030
rect 83620 -52140 83650 -52030
rect 83480 -52170 83650 -52140
rect 85120 -52040 85290 -52010
rect 85120 -52150 85150 -52040
rect 85260 -52150 85290 -52040
rect 85120 -52180 85290 -52150
rect 86530 -52030 86700 -52000
rect 86530 -52140 86560 -52030
rect 86670 -52140 86700 -52030
rect 86530 -52170 86700 -52140
rect 87910 -52030 88080 -52000
rect 87910 -52140 87940 -52030
rect 88050 -52140 88080 -52030
rect 87910 -52170 88080 -52140
rect 89450 -52040 89620 -52010
rect 89450 -52150 89480 -52040
rect 89590 -52150 89620 -52040
rect 89450 -52180 89620 -52150
rect 90730 -52040 90900 -52010
rect 90730 -52150 90760 -52040
rect 90870 -52150 90900 -52040
rect 90730 -52180 90900 -52150
rect 60486 -52562 60520 -52500
rect 77400 -52450 77520 -52420
rect 77400 -52510 77430 -52450
rect 77490 -52510 77520 -52450
rect 77400 -52540 77520 -52510
rect 59772 -52596 59868 -52562
rect 60424 -52596 60520 -52562
rect 77400 -52700 77520 -52670
rect 77400 -52760 77430 -52700
rect 77490 -52760 77520 -52700
rect 77400 -52790 77520 -52760
rect 55176 -53078 55272 -53044
rect 55566 -53078 55662 -53044
rect 55176 -53140 55210 -53078
rect 35802 -53380 35836 -53318
rect 25736 -53388 35836 -53380
rect 55628 -53140 55662 -53078
rect 55176 -53360 55210 -53298
rect 55628 -53360 55662 -53298
rect 25736 -53414 35838 -53388
rect 55176 -53394 55272 -53360
rect 55566 -53394 55662 -53360
rect 25738 -53422 35838 -53414
rect 25738 -53484 25772 -53422
rect 35804 -53484 35838 -53422
rect 25738 -54982 25772 -54920
rect 77390 -53700 77510 -53670
rect 77390 -53760 77420 -53700
rect 77480 -53760 77510 -53700
rect 77390 -53790 77510 -53760
rect 35804 -54982 35838 -54920
rect 25738 -54986 35838 -54982
rect 25736 -55016 35838 -54986
rect 25736 -55020 35836 -55016
rect 25736 -55082 25770 -55020
rect 35802 -55082 35836 -55020
rect 25736 -56580 25770 -56518
rect 35802 -56580 35836 -56518
rect 25736 -56620 35836 -56580
rect 25736 -56682 25770 -56620
rect 35802 -56682 35836 -56620
rect 25736 -58180 25770 -58118
rect 35802 -58180 35836 -58118
rect 53350 -56038 53790 -56004
rect 53350 -56100 53384 -56038
rect 53756 -56664 53790 -56038
rect 55706 -55988 55802 -55954
rect 56050 -55988 56146 -55954
rect 55706 -56050 55740 -55988
rect 55176 -56100 55272 -56066
rect 55430 -56100 55526 -56066
rect 55176 -56162 55210 -56100
rect 55492 -56162 55526 -56100
rect 55176 -56518 55210 -56456
rect 55492 -56518 55526 -56456
rect 54870 -56552 55272 -56518
rect 55430 -56552 55706 -56518
rect 54870 -56558 55706 -56552
rect 54870 -56664 54904 -56558
rect 53756 -56698 53852 -56664
rect 54808 -56698 54904 -56664
rect 53756 -56760 53790 -56698
rect 54870 -56760 54904 -56698
rect 53756 -57070 53790 -57008
rect 54870 -57068 54904 -57008
rect 55700 -57006 55706 -56558
rect 56112 -56050 56146 -55988
rect 55700 -57068 55740 -57006
rect 59772 -56294 59868 -56260
rect 60424 -56294 60520 -56260
rect 59772 -56356 59806 -56294
rect 56112 -57068 56146 -57006
rect 54870 -57070 55160 -57068
rect 53756 -57104 53852 -57070
rect 54808 -57104 55160 -57070
rect 53756 -57166 53790 -57104
rect 54870 -57108 55160 -57104
rect 55600 -57102 55802 -57068
rect 56050 -57102 56146 -57068
rect 55600 -57108 55740 -57102
rect 54870 -57166 54904 -57108
rect 53756 -57476 53790 -57414
rect 55700 -57164 55740 -57108
rect 54870 -57476 54904 -57414
rect 53756 -57510 53852 -57476
rect 54808 -57510 54904 -57476
rect 53350 -58136 53384 -58074
rect 53756 -58136 53790 -57510
rect 54870 -57618 54904 -57510
rect 55700 -57618 55706 -57164
rect 54870 -57624 55706 -57618
rect 54870 -57658 55262 -57624
rect 55420 -57658 55706 -57624
rect 55166 -57720 55200 -57658
rect 53350 -58170 53446 -58136
rect 53694 -58170 53790 -58136
rect 25736 -58214 25832 -58180
rect 35740 -58214 35836 -58180
rect 55482 -57720 55516 -57658
rect 55166 -58076 55200 -58014
rect 55482 -58076 55516 -58014
rect 55166 -58110 55262 -58076
rect 55420 -58110 55516 -58076
rect 56112 -57164 56146 -57102
rect 55706 -58182 55740 -58120
rect 57086 -56710 57376 -56680
rect 57086 -56780 57116 -56710
rect 57346 -56780 57376 -56710
rect 57086 -56810 57376 -56780
rect 60486 -56356 60520 -56294
rect 59772 -56596 59806 -56534
rect 60486 -56596 60520 -56534
rect 59388 -56630 59484 -56596
rect 59642 -56630 59800 -56596
rect 59958 -56630 60520 -56596
rect 59388 -56692 59422 -56630
rect 59388 -57109 59422 -57048
rect 59704 -57109 59738 -56630
rect 60020 -56692 60054 -56630
rect 61186 -56800 61286 -56790
rect 61186 -56820 61366 -56800
rect 61186 -56860 61216 -56820
rect 61336 -56860 61366 -56820
rect 61186 -56880 61366 -56860
rect 61186 -56890 61286 -56880
rect 60020 -57109 60054 -57048
rect 57056 -57370 57416 -57340
rect 57056 -57450 57096 -57370
rect 57376 -57450 57416 -57370
rect 57056 -57480 57416 -57450
rect 59387 -57144 60054 -57109
rect 59387 -57205 59421 -57144
rect 59387 -57623 59421 -57561
rect 59703 -57623 59737 -57144
rect 60019 -57205 60053 -57144
rect 60019 -57623 60053 -57561
rect 59387 -57657 59483 -57623
rect 59641 -57657 59799 -57623
rect 59957 -57626 60053 -57623
rect 59957 -57657 60520 -57626
rect 59772 -57660 60520 -57657
rect 59772 -57722 59806 -57660
rect 56112 -58182 56146 -58120
rect 55706 -58216 55802 -58182
rect 56050 -58216 56146 -58182
rect 60486 -57722 60520 -57660
rect 59772 -57962 59806 -57900
rect 60486 -57962 60520 -57900
rect 59772 -57996 59868 -57962
rect 60424 -57996 60520 -57962
rect 55176 -58478 55272 -58444
rect 55566 -58478 55662 -58444
rect 55176 -58540 55210 -58478
rect 55628 -58540 55662 -58478
rect 55176 -58760 55210 -58698
rect 55628 -58760 55662 -58698
rect 55176 -58794 55272 -58760
rect 55566 -58794 55662 -58760
rect 53350 -61438 53790 -61404
rect 53350 -61500 53384 -61438
rect 53756 -62064 53790 -61438
rect 55706 -61388 55802 -61354
rect 56050 -61388 56146 -61354
rect 55706 -61450 55740 -61388
rect 55176 -61500 55272 -61466
rect 55430 -61500 55526 -61466
rect 55176 -61562 55210 -61500
rect 55492 -61562 55526 -61500
rect 55176 -61918 55210 -61856
rect 55492 -61918 55526 -61856
rect 54870 -61952 55272 -61918
rect 55430 -61952 55706 -61918
rect 54870 -61958 55706 -61952
rect 54870 -62064 54904 -61958
rect 53756 -62098 53852 -62064
rect 54808 -62098 54904 -62064
rect 53756 -62160 53790 -62098
rect 54870 -62160 54904 -62098
rect 53756 -62470 53790 -62408
rect 54870 -62468 54904 -62408
rect 55700 -62406 55706 -61958
rect 56112 -61450 56146 -61388
rect 55700 -62468 55740 -62406
rect 59772 -61694 59868 -61660
rect 60424 -61694 60520 -61660
rect 59772 -61756 59806 -61694
rect 56112 -62468 56146 -62406
rect 54870 -62470 55160 -62468
rect 53756 -62504 53852 -62470
rect 54808 -62504 55160 -62470
rect 53756 -62566 53790 -62504
rect 54870 -62508 55160 -62504
rect 55600 -62502 55802 -62468
rect 56050 -62502 56146 -62468
rect 55600 -62508 55740 -62502
rect 54870 -62566 54904 -62508
rect 53756 -62876 53790 -62814
rect 55700 -62564 55740 -62508
rect 54870 -62876 54904 -62814
rect 53756 -62910 53852 -62876
rect 54808 -62910 54904 -62876
rect 53350 -63536 53384 -63474
rect 53756 -63536 53790 -62910
rect 54870 -63018 54904 -62910
rect 55700 -63018 55706 -62564
rect 54870 -63024 55706 -63018
rect 54870 -63058 55262 -63024
rect 55420 -63058 55706 -63024
rect 55166 -63120 55200 -63058
rect 53350 -63570 53446 -63536
rect 53694 -63570 53790 -63536
rect 55482 -63120 55516 -63058
rect 55166 -63476 55200 -63414
rect 55482 -63476 55516 -63414
rect 55166 -63510 55262 -63476
rect 55420 -63510 55516 -63476
rect 56112 -62564 56146 -62502
rect 55706 -63582 55740 -63520
rect 57086 -62110 57376 -62080
rect 57086 -62180 57116 -62110
rect 57346 -62180 57376 -62110
rect 57086 -62210 57376 -62180
rect 60486 -61756 60520 -61694
rect 59772 -61996 59806 -61934
rect 60486 -61996 60520 -61934
rect 59388 -62030 59484 -61996
rect 59642 -62030 59800 -61996
rect 59958 -62030 60520 -61996
rect 59388 -62092 59422 -62030
rect 59388 -62509 59422 -62448
rect 59704 -62509 59738 -62030
rect 60020 -62092 60054 -62030
rect 61186 -62200 61286 -62190
rect 61186 -62220 61366 -62200
rect 61186 -62260 61216 -62220
rect 61336 -62260 61366 -62220
rect 61186 -62280 61366 -62260
rect 61186 -62290 61286 -62280
rect 60020 -62509 60054 -62448
rect 57056 -62770 57416 -62740
rect 57056 -62850 57096 -62770
rect 57376 -62850 57416 -62770
rect 57056 -62880 57416 -62850
rect 59387 -62544 60054 -62509
rect 59387 -62605 59421 -62544
rect 59387 -63023 59421 -62961
rect 59703 -63023 59737 -62544
rect 60019 -62605 60053 -62544
rect 60019 -63023 60053 -62961
rect 59387 -63057 59483 -63023
rect 59641 -63057 59799 -63023
rect 59957 -63026 60053 -63023
rect 59957 -63057 60520 -63026
rect 59772 -63060 60520 -63057
rect 59772 -63122 59806 -63060
rect 56112 -63582 56146 -63520
rect 55706 -63616 55802 -63582
rect 56050 -63616 56146 -63582
rect 60486 -63122 60520 -63060
rect 59772 -63362 59806 -63300
rect 60486 -63362 60520 -63300
rect 59772 -63396 59868 -63362
rect 60424 -63396 60520 -63362
rect 55176 -63878 55272 -63844
rect 55566 -63878 55662 -63844
rect 55176 -63940 55210 -63878
rect 55628 -63940 55662 -63878
rect 55176 -64160 55210 -64098
rect 55628 -64160 55662 -64098
rect 55176 -64194 55272 -64160
rect 55566 -64194 55662 -64160
rect 53350 -66838 53790 -66804
rect 53350 -66900 53384 -66838
rect 53756 -67464 53790 -66838
rect 55706 -66788 55802 -66754
rect 56050 -66788 56146 -66754
rect 55706 -66850 55740 -66788
rect 55176 -66900 55272 -66866
rect 55430 -66900 55526 -66866
rect 55176 -66962 55210 -66900
rect 55492 -66962 55526 -66900
rect 55176 -67318 55210 -67256
rect 55492 -67318 55526 -67256
rect 54870 -67352 55272 -67318
rect 55430 -67352 55706 -67318
rect 54870 -67358 55706 -67352
rect 54870 -67464 54904 -67358
rect 53756 -67498 53852 -67464
rect 54808 -67498 54904 -67464
rect 53756 -67560 53790 -67498
rect 54870 -67560 54904 -67498
rect 53756 -67870 53790 -67808
rect 54870 -67868 54904 -67808
rect 55700 -67806 55706 -67358
rect 56112 -66850 56146 -66788
rect 55700 -67868 55740 -67806
rect 59772 -67094 59868 -67060
rect 60424 -67094 60520 -67060
rect 59772 -67156 59806 -67094
rect 56112 -67868 56146 -67806
rect 54870 -67870 55160 -67868
rect 53756 -67904 53852 -67870
rect 54808 -67904 55160 -67870
rect 53756 -67966 53790 -67904
rect 54870 -67908 55160 -67904
rect 55600 -67902 55802 -67868
rect 56050 -67902 56146 -67868
rect 55600 -67908 55740 -67902
rect 54870 -67966 54904 -67908
rect 53756 -68276 53790 -68214
rect 55700 -67964 55740 -67908
rect 54870 -68276 54904 -68214
rect 53756 -68310 53852 -68276
rect 54808 -68310 54904 -68276
rect 53350 -68936 53384 -68874
rect 53756 -68936 53790 -68310
rect 54870 -68418 54904 -68310
rect 55700 -68418 55706 -67964
rect 54870 -68424 55706 -68418
rect 54870 -68458 55262 -68424
rect 55420 -68458 55706 -68424
rect 55166 -68520 55200 -68458
rect 53350 -68970 53446 -68936
rect 53694 -68970 53790 -68936
rect 55482 -68520 55516 -68458
rect 55166 -68876 55200 -68814
rect 55482 -68876 55516 -68814
rect 55166 -68910 55262 -68876
rect 55420 -68910 55516 -68876
rect 56112 -67964 56146 -67902
rect 55706 -68982 55740 -68920
rect 57086 -67510 57376 -67480
rect 57086 -67580 57116 -67510
rect 57346 -67580 57376 -67510
rect 57086 -67610 57376 -67580
rect 60486 -67156 60520 -67094
rect 59772 -67396 59806 -67334
rect 60486 -67396 60520 -67334
rect 59388 -67430 59484 -67396
rect 59642 -67430 59800 -67396
rect 59958 -67430 60520 -67396
rect 59388 -67492 59422 -67430
rect 59388 -67909 59422 -67848
rect 59704 -67909 59738 -67430
rect 60020 -67492 60054 -67430
rect 61186 -67600 61286 -67590
rect 61186 -67620 61366 -67600
rect 61186 -67660 61216 -67620
rect 61336 -67660 61366 -67620
rect 61186 -67680 61366 -67660
rect 61186 -67690 61286 -67680
rect 60020 -67909 60054 -67848
rect 57056 -68170 57416 -68140
rect 57056 -68250 57096 -68170
rect 57376 -68250 57416 -68170
rect 57056 -68280 57416 -68250
rect 59387 -67944 60054 -67909
rect 59387 -68005 59421 -67944
rect 59387 -68423 59421 -68361
rect 59703 -68423 59737 -67944
rect 60019 -68005 60053 -67944
rect 60019 -68423 60053 -68361
rect 59387 -68457 59483 -68423
rect 59641 -68457 59799 -68423
rect 59957 -68426 60053 -68423
rect 59957 -68457 60520 -68426
rect 59772 -68460 60520 -68457
rect 59772 -68522 59806 -68460
rect 56112 -68982 56146 -68920
rect 55706 -69016 55802 -68982
rect 56050 -69016 56146 -68982
rect 60486 -68522 60520 -68460
rect 59772 -68762 59806 -68700
rect 60486 -68762 60520 -68700
rect 59772 -68796 59868 -68762
rect 60424 -68796 60520 -68762
rect 55176 -69278 55272 -69244
rect 55566 -69278 55662 -69244
rect 55176 -69340 55210 -69278
rect 55628 -69340 55662 -69278
rect 55176 -69560 55210 -69498
rect 55628 -69560 55662 -69498
rect 55176 -69594 55272 -69560
rect 55566 -69594 55662 -69560
rect 53350 -72238 53790 -72204
rect 53350 -72300 53384 -72238
rect 53756 -72864 53790 -72238
rect 55706 -72188 55802 -72154
rect 56050 -72188 56146 -72154
rect 55706 -72250 55740 -72188
rect 55176 -72300 55272 -72266
rect 55430 -72300 55526 -72266
rect 55176 -72362 55210 -72300
rect 55492 -72362 55526 -72300
rect 55176 -72718 55210 -72656
rect 55492 -72718 55526 -72656
rect 54870 -72752 55272 -72718
rect 55430 -72752 55706 -72718
rect 54870 -72758 55706 -72752
rect 54870 -72864 54904 -72758
rect 53756 -72898 53852 -72864
rect 54808 -72898 54904 -72864
rect 53756 -72960 53790 -72898
rect 54870 -72960 54904 -72898
rect 53756 -73270 53790 -73208
rect 54870 -73268 54904 -73208
rect 55700 -73206 55706 -72758
rect 56112 -72250 56146 -72188
rect 55700 -73268 55740 -73206
rect 59772 -72494 59868 -72460
rect 60424 -72494 60520 -72460
rect 59772 -72556 59806 -72494
rect 56112 -73268 56146 -73206
rect 54870 -73270 55160 -73268
rect 53756 -73304 53852 -73270
rect 54808 -73304 55160 -73270
rect 53756 -73366 53790 -73304
rect 54870 -73308 55160 -73304
rect 55600 -73302 55802 -73268
rect 56050 -73302 56146 -73268
rect 55600 -73308 55740 -73302
rect 54870 -73366 54904 -73308
rect 53756 -73676 53790 -73614
rect 55700 -73364 55740 -73308
rect 54870 -73676 54904 -73614
rect 53756 -73710 53852 -73676
rect 54808 -73710 54904 -73676
rect 53350 -74336 53384 -74274
rect 53756 -74336 53790 -73710
rect 54870 -73818 54904 -73710
rect 55700 -73818 55706 -73364
rect 54870 -73824 55706 -73818
rect 54870 -73858 55262 -73824
rect 55420 -73858 55706 -73824
rect 55166 -73920 55200 -73858
rect 53350 -74370 53446 -74336
rect 53694 -74370 53790 -74336
rect 55482 -73920 55516 -73858
rect 55166 -74276 55200 -74214
rect 55482 -74276 55516 -74214
rect 55166 -74310 55262 -74276
rect 55420 -74310 55516 -74276
rect 56112 -73364 56146 -73302
rect 55706 -74382 55740 -74320
rect 57086 -72910 57376 -72880
rect 57086 -72980 57116 -72910
rect 57346 -72980 57376 -72910
rect 57086 -73010 57376 -72980
rect 60486 -72556 60520 -72494
rect 59772 -72796 59806 -72734
rect 60486 -72796 60520 -72734
rect 59388 -72830 59484 -72796
rect 59642 -72830 59800 -72796
rect 59958 -72830 60520 -72796
rect 59388 -72892 59422 -72830
rect 59388 -73309 59422 -73248
rect 59704 -73309 59738 -72830
rect 60020 -72892 60054 -72830
rect 61186 -73000 61286 -72990
rect 61186 -73020 61366 -73000
rect 61186 -73060 61216 -73020
rect 61336 -73060 61366 -73020
rect 61186 -73080 61366 -73060
rect 61186 -73090 61286 -73080
rect 60020 -73309 60054 -73248
rect 57056 -73570 57416 -73540
rect 57056 -73650 57096 -73570
rect 57376 -73650 57416 -73570
rect 57056 -73680 57416 -73650
rect 59387 -73344 60054 -73309
rect 59387 -73405 59421 -73344
rect 59387 -73823 59421 -73761
rect 59703 -73823 59737 -73344
rect 60019 -73405 60053 -73344
rect 60019 -73823 60053 -73761
rect 59387 -73857 59483 -73823
rect 59641 -73857 59799 -73823
rect 59957 -73826 60053 -73823
rect 59957 -73857 60520 -73826
rect 59772 -73860 60520 -73857
rect 59772 -73922 59806 -73860
rect 56112 -74382 56146 -74320
rect 55706 -74416 55802 -74382
rect 56050 -74416 56146 -74382
rect 60486 -73922 60520 -73860
rect 59772 -74162 59806 -74100
rect 60486 -74162 60520 -74100
rect 59772 -74196 59868 -74162
rect 60424 -74196 60520 -74162
rect 55176 -74678 55272 -74644
rect 55566 -74678 55662 -74644
rect 55176 -74740 55210 -74678
rect 55628 -74740 55662 -74678
rect 55176 -74960 55210 -74898
rect 55628 -74960 55662 -74898
rect 55176 -74994 55272 -74960
rect 55566 -74994 55662 -74960
rect 53350 -77638 53790 -77604
rect 53350 -77700 53384 -77638
rect 53756 -78264 53790 -77638
rect 55706 -77588 55802 -77554
rect 56050 -77588 56146 -77554
rect 55706 -77650 55740 -77588
rect 55176 -77700 55272 -77666
rect 55430 -77700 55526 -77666
rect 55176 -77762 55210 -77700
rect 55492 -77762 55526 -77700
rect 55176 -78118 55210 -78056
rect 55492 -78118 55526 -78056
rect 54870 -78152 55272 -78118
rect 55430 -78152 55706 -78118
rect 54870 -78158 55706 -78152
rect 54870 -78264 54904 -78158
rect 53756 -78298 53852 -78264
rect 54808 -78298 54904 -78264
rect 53756 -78360 53790 -78298
rect 54870 -78360 54904 -78298
rect 53756 -78670 53790 -78608
rect 54870 -78668 54904 -78608
rect 55700 -78606 55706 -78158
rect 56112 -77650 56146 -77588
rect 55700 -78668 55740 -78606
rect 59772 -77894 59868 -77860
rect 60424 -77894 60520 -77860
rect 59772 -77956 59806 -77894
rect 56112 -78668 56146 -78606
rect 54870 -78670 55160 -78668
rect 53756 -78704 53852 -78670
rect 54808 -78704 55160 -78670
rect 53756 -78766 53790 -78704
rect 54870 -78708 55160 -78704
rect 55600 -78702 55802 -78668
rect 56050 -78702 56146 -78668
rect 55600 -78708 55740 -78702
rect 54870 -78766 54904 -78708
rect 53756 -79076 53790 -79014
rect 55700 -78764 55740 -78708
rect 54870 -79076 54904 -79014
rect 53756 -79110 53852 -79076
rect 54808 -79110 54904 -79076
rect 53350 -79736 53384 -79674
rect 53756 -79736 53790 -79110
rect 54870 -79218 54904 -79110
rect 55700 -79218 55706 -78764
rect 54870 -79224 55706 -79218
rect 54870 -79258 55262 -79224
rect 55420 -79258 55706 -79224
rect 55166 -79320 55200 -79258
rect 53350 -79770 53446 -79736
rect 53694 -79770 53790 -79736
rect 55482 -79320 55516 -79258
rect 55166 -79676 55200 -79614
rect 55482 -79676 55516 -79614
rect 55166 -79710 55262 -79676
rect 55420 -79710 55516 -79676
rect 56112 -78764 56146 -78702
rect 55706 -79782 55740 -79720
rect 57086 -78310 57376 -78280
rect 57086 -78380 57116 -78310
rect 57346 -78380 57376 -78310
rect 57086 -78410 57376 -78380
rect 60486 -77956 60520 -77894
rect 59772 -78196 59806 -78134
rect 60486 -78196 60520 -78134
rect 59388 -78230 59484 -78196
rect 59642 -78230 59800 -78196
rect 59958 -78230 60520 -78196
rect 59388 -78292 59422 -78230
rect 59388 -78709 59422 -78648
rect 59704 -78709 59738 -78230
rect 60020 -78292 60054 -78230
rect 61186 -78400 61286 -78390
rect 61186 -78420 61366 -78400
rect 61186 -78460 61216 -78420
rect 61336 -78460 61366 -78420
rect 61186 -78480 61366 -78460
rect 61186 -78490 61286 -78480
rect 60020 -78709 60054 -78648
rect 57056 -78970 57416 -78940
rect 57056 -79050 57096 -78970
rect 57376 -79050 57416 -78970
rect 57056 -79080 57416 -79050
rect 59387 -78744 60054 -78709
rect 59387 -78805 59421 -78744
rect 59387 -79223 59421 -79161
rect 59703 -79223 59737 -78744
rect 60019 -78805 60053 -78744
rect 60019 -79223 60053 -79161
rect 59387 -79257 59483 -79223
rect 59641 -79257 59799 -79223
rect 59957 -79226 60053 -79223
rect 59957 -79257 60520 -79226
rect 59772 -79260 60520 -79257
rect 59772 -79322 59806 -79260
rect 56112 -79782 56146 -79720
rect 55706 -79816 55802 -79782
rect 56050 -79816 56146 -79782
rect 60486 -79322 60520 -79260
rect 59772 -79562 59806 -79500
rect 60486 -79562 60520 -79500
rect 59772 -79596 59868 -79562
rect 60424 -79596 60520 -79562
rect 55176 -80078 55272 -80044
rect 55566 -80078 55662 -80044
rect 55176 -80140 55210 -80078
rect 55628 -80140 55662 -80078
rect 55176 -80360 55210 -80298
rect 55628 -80360 55662 -80298
rect 55176 -80394 55272 -80360
rect 55566 -80394 55662 -80360
rect 53350 -83038 53790 -83004
rect 53350 -83100 53384 -83038
rect 53756 -83664 53790 -83038
rect 55706 -82988 55802 -82954
rect 56050 -82988 56146 -82954
rect 55706 -83050 55740 -82988
rect 55176 -83100 55272 -83066
rect 55430 -83100 55526 -83066
rect 55176 -83162 55210 -83100
rect 55492 -83162 55526 -83100
rect 55176 -83518 55210 -83456
rect 55492 -83518 55526 -83456
rect 54870 -83552 55272 -83518
rect 55430 -83552 55706 -83518
rect 54870 -83558 55706 -83552
rect 54870 -83664 54904 -83558
rect 53756 -83698 53852 -83664
rect 54808 -83698 54904 -83664
rect 53756 -83760 53790 -83698
rect 54870 -83760 54904 -83698
rect 53756 -84070 53790 -84008
rect 54870 -84068 54904 -84008
rect 55700 -84006 55706 -83558
rect 56112 -83050 56146 -82988
rect 55700 -84068 55740 -84006
rect 59772 -83294 59868 -83260
rect 60424 -83294 60520 -83260
rect 59772 -83356 59806 -83294
rect 56112 -84068 56146 -84006
rect 54870 -84070 55160 -84068
rect 53756 -84104 53852 -84070
rect 54808 -84104 55160 -84070
rect 53756 -84166 53790 -84104
rect 54870 -84108 55160 -84104
rect 55600 -84102 55802 -84068
rect 56050 -84102 56146 -84068
rect 55600 -84108 55740 -84102
rect 54870 -84166 54904 -84108
rect 53756 -84476 53790 -84414
rect 55700 -84164 55740 -84108
rect 54870 -84476 54904 -84414
rect 53756 -84510 53852 -84476
rect 54808 -84510 54904 -84476
rect 53350 -85136 53384 -85074
rect 53756 -85136 53790 -84510
rect 54870 -84618 54904 -84510
rect 55700 -84618 55706 -84164
rect 54870 -84624 55706 -84618
rect 54870 -84658 55262 -84624
rect 55420 -84658 55706 -84624
rect 55166 -84720 55200 -84658
rect 53350 -85170 53446 -85136
rect 53694 -85170 53790 -85136
rect 55482 -84720 55516 -84658
rect 55166 -85076 55200 -85014
rect 55482 -85076 55516 -85014
rect 55166 -85110 55262 -85076
rect 55420 -85110 55516 -85076
rect 56112 -84164 56146 -84102
rect 55706 -85182 55740 -85120
rect 57086 -83710 57376 -83680
rect 57086 -83780 57116 -83710
rect 57346 -83780 57376 -83710
rect 57086 -83810 57376 -83780
rect 60486 -83356 60520 -83294
rect 59772 -83596 59806 -83534
rect 60486 -83596 60520 -83534
rect 59388 -83630 59484 -83596
rect 59642 -83630 59800 -83596
rect 59958 -83630 60520 -83596
rect 59388 -83692 59422 -83630
rect 59388 -84109 59422 -84048
rect 59704 -84109 59738 -83630
rect 60020 -83692 60054 -83630
rect 61186 -83800 61286 -83790
rect 61186 -83820 61366 -83800
rect 61186 -83860 61216 -83820
rect 61336 -83860 61366 -83820
rect 61186 -83880 61366 -83860
rect 61186 -83890 61286 -83880
rect 60020 -84109 60054 -84048
rect 57056 -84370 57416 -84340
rect 57056 -84450 57096 -84370
rect 57376 -84450 57416 -84370
rect 57056 -84480 57416 -84450
rect 59387 -84144 60054 -84109
rect 59387 -84205 59421 -84144
rect 59387 -84623 59421 -84561
rect 59703 -84623 59737 -84144
rect 60019 -84205 60053 -84144
rect 60019 -84623 60053 -84561
rect 59387 -84657 59483 -84623
rect 59641 -84657 59799 -84623
rect 59957 -84626 60053 -84623
rect 59957 -84657 60520 -84626
rect 59772 -84660 60520 -84657
rect 59772 -84722 59806 -84660
rect 56112 -85182 56146 -85120
rect 55706 -85216 55802 -85182
rect 56050 -85216 56146 -85182
rect 60486 -84722 60520 -84660
rect 59772 -84962 59806 -84900
rect 60486 -84962 60520 -84900
rect 59772 -84996 59868 -84962
rect 60424 -84996 60520 -84962
rect 55176 -85478 55272 -85444
rect 55566 -85478 55662 -85444
rect 55176 -85540 55210 -85478
rect 55628 -85540 55662 -85478
rect 55176 -85760 55210 -85698
rect 55628 -85760 55662 -85698
rect 55176 -85794 55272 -85760
rect 55566 -85794 55662 -85760
<< nsubdiff >>
rect 53896 -1592 53992 -1558
rect 54966 -1592 55062 -1558
rect 53896 -1654 53930 -1592
rect 55028 -1654 55062 -1592
rect 53896 -1914 53930 -1852
rect 55028 -1914 55062 -1852
rect 53896 -1948 53992 -1914
rect 54966 -1948 55062 -1914
rect 53896 -2010 53930 -1948
rect 55028 -2010 55062 -1948
rect 57126 -1900 57356 -1870
rect 53896 -2270 53930 -2208
rect 55028 -2270 55062 -2208
rect 53896 -2304 53992 -2270
rect 54966 -2304 55062 -2270
rect 55118 -2674 55518 -2662
rect 55118 -2708 55142 -2674
rect 55494 -2708 55518 -2674
rect 55118 -2759 55518 -2708
rect 55118 -2846 55518 -2795
rect 55118 -2880 55142 -2846
rect 55494 -2880 55518 -2846
rect 55118 -2892 55518 -2880
rect 57126 -1970 57156 -1900
rect 57316 -1970 57356 -1900
rect 57126 -2000 57356 -1970
rect 58930 -1967 59026 -1933
rect 59600 -1967 59696 -1933
rect 58930 -2029 58964 -1967
rect 59662 -2029 59696 -1967
rect 58930 -2376 58964 -2315
rect 58930 -2410 59026 -2376
rect 59214 -2377 59310 -2376
rect 59662 -2377 59696 -2315
rect 59214 -2410 59696 -2377
rect 58930 -2411 59696 -2410
rect 55118 -3296 55518 -3284
rect 55118 -3330 55142 -3296
rect 55494 -3330 55518 -3296
rect 55118 -3381 55518 -3330
rect 55118 -3468 55518 -3417
rect 55118 -3502 55142 -3468
rect 55494 -3502 55518 -3468
rect 55118 -3514 55518 -3502
rect 53886 -3908 53982 -3874
rect 54956 -3908 55052 -3874
rect 53886 -3970 53920 -3908
rect 55018 -3970 55052 -3908
rect 53886 -4230 53920 -4168
rect 55018 -4230 55052 -4168
rect 56316 -2538 56412 -2504
rect 56610 -2538 56706 -2504
rect 56316 -2600 56350 -2538
rect 56672 -2600 56706 -2538
rect 58930 -2472 58964 -2411
rect 56316 -3636 56350 -3574
rect 59276 -2472 59310 -2411
rect 58930 -3106 58964 -3046
rect 59276 -3106 59310 -3046
rect 58930 -3142 59310 -3106
rect 58930 -3202 58964 -3142
rect 56672 -3636 56706 -3574
rect 56316 -3670 56412 -3636
rect 56610 -3670 56706 -3636
rect 59276 -3202 59310 -3142
rect 58930 -3838 58964 -3776
rect 60466 -3460 60546 -3430
rect 60466 -3500 60486 -3460
rect 60526 -3500 60546 -3460
rect 60466 -3530 60546 -3500
rect 60606 -3460 60686 -3430
rect 60606 -3500 60626 -3460
rect 60666 -3500 60686 -3460
rect 60606 -3530 60686 -3500
rect 60746 -3460 60826 -3430
rect 60746 -3500 60766 -3460
rect 60806 -3500 60826 -3460
rect 60746 -3530 60826 -3500
rect 60886 -3460 60966 -3430
rect 60886 -3500 60906 -3460
rect 60946 -3500 60966 -3460
rect 60886 -3530 60966 -3500
rect 59276 -3838 59310 -3776
rect 58930 -3872 59026 -3838
rect 59214 -3840 59310 -3838
rect 59214 -3872 59696 -3840
rect 58930 -3874 59696 -3872
rect 58930 -3936 58964 -3874
rect 53886 -4264 53982 -4230
rect 54956 -4264 55052 -4230
rect 59662 -3936 59696 -3874
rect 53886 -4326 53920 -4264
rect 55018 -4326 55052 -4264
rect 53886 -4586 53920 -4524
rect 57156 -4290 57316 -4260
rect 57156 -4390 57186 -4290
rect 57286 -4390 57316 -4290
rect 58930 -4284 58964 -4222
rect 59662 -4284 59696 -4222
rect 58930 -4318 59026 -4284
rect 59600 -4318 59696 -4284
rect 57156 -4420 57316 -4390
rect 55018 -4586 55052 -4524
rect 53886 -4620 53982 -4586
rect 54956 -4620 55052 -4586
rect 53896 -6992 53992 -6958
rect 54966 -6992 55062 -6958
rect 53896 -7054 53930 -6992
rect 55028 -7054 55062 -6992
rect 53896 -7314 53930 -7252
rect 55028 -7314 55062 -7252
rect 53896 -7348 53992 -7314
rect 54966 -7348 55062 -7314
rect 20732 -7707 20828 -7673
rect 21156 -7707 21314 -7673
rect 21642 -7707 21800 -7673
rect 22128 -7707 22224 -7673
rect 20732 -7769 20766 -7707
rect 21218 -7769 21252 -7707
rect 20732 -11805 20766 -11743
rect 21704 -7769 21738 -7707
rect 21218 -11805 21252 -11743
rect 22190 -7769 22224 -7707
rect 21704 -11805 21738 -11743
rect 53896 -7410 53930 -7348
rect 55028 -7410 55062 -7348
rect 57126 -7300 57356 -7270
rect 53896 -7670 53930 -7608
rect 55028 -7670 55062 -7608
rect 53896 -7704 53992 -7670
rect 54966 -7704 55062 -7670
rect 55118 -8074 55518 -8062
rect 55118 -8108 55142 -8074
rect 55494 -8108 55518 -8074
rect 55118 -8159 55518 -8108
rect 55118 -8246 55518 -8195
rect 55118 -8280 55142 -8246
rect 55494 -8280 55518 -8246
rect 55118 -8292 55518 -8280
rect 57126 -7370 57156 -7300
rect 57316 -7370 57356 -7300
rect 57126 -7400 57356 -7370
rect 58930 -7367 59026 -7333
rect 59600 -7367 59696 -7333
rect 58930 -7429 58964 -7367
rect 59662 -7429 59696 -7367
rect 58930 -7776 58964 -7715
rect 58930 -7810 59026 -7776
rect 59214 -7777 59310 -7776
rect 59662 -7777 59696 -7715
rect 59214 -7810 59696 -7777
rect 58930 -7811 59696 -7810
rect 55118 -8696 55518 -8684
rect 55118 -8730 55142 -8696
rect 55494 -8730 55518 -8696
rect 55118 -8781 55518 -8730
rect 55118 -8868 55518 -8817
rect 55118 -8902 55142 -8868
rect 55494 -8902 55518 -8868
rect 55118 -8914 55518 -8902
rect 53886 -9308 53982 -9274
rect 54956 -9308 55052 -9274
rect 53886 -9370 53920 -9308
rect 55018 -9370 55052 -9308
rect 53886 -9630 53920 -9568
rect 55018 -9630 55052 -9568
rect 56316 -7938 56412 -7904
rect 56610 -7938 56706 -7904
rect 56316 -8000 56350 -7938
rect 56672 -8000 56706 -7938
rect 58930 -7872 58964 -7811
rect 56316 -9036 56350 -8974
rect 59276 -7872 59310 -7811
rect 58930 -8506 58964 -8446
rect 59276 -8506 59310 -8446
rect 58930 -8542 59310 -8506
rect 58930 -8602 58964 -8542
rect 56672 -9036 56706 -8974
rect 56316 -9070 56412 -9036
rect 56610 -9070 56706 -9036
rect 59276 -8602 59310 -8542
rect 58930 -9238 58964 -9176
rect 60466 -8860 60546 -8830
rect 60466 -8900 60486 -8860
rect 60526 -8900 60546 -8860
rect 60466 -8930 60546 -8900
rect 60606 -8860 60686 -8830
rect 60606 -8900 60626 -8860
rect 60666 -8900 60686 -8860
rect 60606 -8930 60686 -8900
rect 60746 -8860 60826 -8830
rect 60746 -8900 60766 -8860
rect 60806 -8900 60826 -8860
rect 60746 -8930 60826 -8900
rect 60886 -8860 60966 -8830
rect 60886 -8900 60906 -8860
rect 60946 -8900 60966 -8860
rect 60886 -8930 60966 -8900
rect 59276 -9238 59310 -9176
rect 58930 -9272 59026 -9238
rect 59214 -9240 59310 -9238
rect 59214 -9272 59696 -9240
rect 58930 -9274 59696 -9272
rect 58930 -9336 58964 -9274
rect 53886 -9664 53982 -9630
rect 54956 -9664 55052 -9630
rect 59662 -9336 59696 -9274
rect 53886 -9726 53920 -9664
rect 55018 -9726 55052 -9664
rect 53886 -9986 53920 -9924
rect 57156 -9690 57316 -9660
rect 57156 -9790 57186 -9690
rect 57286 -9790 57316 -9690
rect 58930 -9684 58964 -9622
rect 59662 -9684 59696 -9622
rect 58930 -9718 59026 -9684
rect 59600 -9718 59696 -9684
rect 57156 -9820 57316 -9790
rect 55018 -9986 55052 -9924
rect 53886 -10020 53982 -9986
rect 54956 -10020 55052 -9986
rect 22190 -11805 22224 -11743
rect 20732 -11839 20828 -11805
rect 21156 -11839 21314 -11805
rect 21642 -11839 21800 -11805
rect 22128 -11839 22224 -11805
rect 53896 -12392 53992 -12358
rect 54966 -12392 55062 -12358
rect 53896 -12454 53930 -12392
rect 55028 -12454 55062 -12392
rect 53896 -12714 53930 -12652
rect 55028 -12714 55062 -12652
rect 53896 -12748 53992 -12714
rect 54966 -12748 55062 -12714
rect 53896 -12810 53930 -12748
rect 55028 -12810 55062 -12748
rect 57126 -12700 57356 -12670
rect 53896 -13070 53930 -13008
rect 55028 -13070 55062 -13008
rect 53896 -13104 53992 -13070
rect 54966 -13104 55062 -13070
rect 55118 -13474 55518 -13462
rect 55118 -13508 55142 -13474
rect 55494 -13508 55518 -13474
rect 55118 -13559 55518 -13508
rect 55118 -13646 55518 -13595
rect 55118 -13680 55142 -13646
rect 55494 -13680 55518 -13646
rect 55118 -13692 55518 -13680
rect 57126 -12770 57156 -12700
rect 57316 -12770 57356 -12700
rect 57126 -12800 57356 -12770
rect 58930 -12767 59026 -12733
rect 59600 -12767 59696 -12733
rect 58930 -12829 58964 -12767
rect 59662 -12829 59696 -12767
rect 58930 -13176 58964 -13115
rect 58930 -13210 59026 -13176
rect 59214 -13177 59310 -13176
rect 59662 -13177 59696 -13115
rect 59214 -13210 59696 -13177
rect 58930 -13211 59696 -13210
rect 55118 -14096 55518 -14084
rect 55118 -14130 55142 -14096
rect 55494 -14130 55518 -14096
rect 55118 -14181 55518 -14130
rect 55118 -14268 55518 -14217
rect 55118 -14302 55142 -14268
rect 55494 -14302 55518 -14268
rect 55118 -14314 55518 -14302
rect 53886 -14708 53982 -14674
rect 54956 -14708 55052 -14674
rect 53886 -14770 53920 -14708
rect 55018 -14770 55052 -14708
rect 53886 -15030 53920 -14968
rect 55018 -15030 55052 -14968
rect 56316 -13338 56412 -13304
rect 56610 -13338 56706 -13304
rect 56316 -13400 56350 -13338
rect 56672 -13400 56706 -13338
rect 58930 -13272 58964 -13211
rect 56316 -14436 56350 -14374
rect 59276 -13272 59310 -13211
rect 58930 -13906 58964 -13846
rect 59276 -13906 59310 -13846
rect 58930 -13942 59310 -13906
rect 58930 -14002 58964 -13942
rect 56672 -14436 56706 -14374
rect 56316 -14470 56412 -14436
rect 56610 -14470 56706 -14436
rect 59276 -14002 59310 -13942
rect 58930 -14638 58964 -14576
rect 60466 -14260 60546 -14230
rect 60466 -14300 60486 -14260
rect 60526 -14300 60546 -14260
rect 60466 -14330 60546 -14300
rect 60606 -14260 60686 -14230
rect 60606 -14300 60626 -14260
rect 60666 -14300 60686 -14260
rect 60606 -14330 60686 -14300
rect 60746 -14260 60826 -14230
rect 60746 -14300 60766 -14260
rect 60806 -14300 60826 -14260
rect 60746 -14330 60826 -14300
rect 60886 -14260 60966 -14230
rect 60886 -14300 60906 -14260
rect 60946 -14300 60966 -14260
rect 60886 -14330 60966 -14300
rect 59276 -14638 59310 -14576
rect 58930 -14672 59026 -14638
rect 59214 -14640 59310 -14638
rect 59214 -14672 59696 -14640
rect 58930 -14674 59696 -14672
rect 58930 -14736 58964 -14674
rect 53886 -15064 53982 -15030
rect 54956 -15064 55052 -15030
rect 59662 -14736 59696 -14674
rect 53886 -15126 53920 -15064
rect 55018 -15126 55052 -15064
rect 53886 -15386 53920 -15324
rect 57156 -15090 57316 -15060
rect 57156 -15190 57186 -15090
rect 57286 -15190 57316 -15090
rect 58930 -15084 58964 -15022
rect 59662 -15084 59696 -15022
rect 58930 -15118 59026 -15084
rect 59600 -15118 59696 -15084
rect 57156 -15220 57316 -15190
rect 55018 -15386 55052 -15324
rect 53886 -15420 53982 -15386
rect 54956 -15420 55052 -15386
rect 53896 -17792 53992 -17758
rect 54966 -17792 55062 -17758
rect 53896 -17854 53930 -17792
rect 55028 -17854 55062 -17792
rect 53896 -18114 53930 -18052
rect 55028 -18114 55062 -18052
rect 53896 -18148 53992 -18114
rect 54966 -18148 55062 -18114
rect 53896 -18210 53930 -18148
rect 55028 -18210 55062 -18148
rect 57126 -18100 57356 -18070
rect 53896 -18470 53930 -18408
rect 55028 -18470 55062 -18408
rect 53896 -18504 53992 -18470
rect 54966 -18504 55062 -18470
rect 55118 -18874 55518 -18862
rect 55118 -18908 55142 -18874
rect 55494 -18908 55518 -18874
rect 55118 -18959 55518 -18908
rect 55118 -19046 55518 -18995
rect 55118 -19080 55142 -19046
rect 55494 -19080 55518 -19046
rect 55118 -19092 55518 -19080
rect 57126 -18170 57156 -18100
rect 57316 -18170 57356 -18100
rect 57126 -18200 57356 -18170
rect 58930 -18167 59026 -18133
rect 59600 -18167 59696 -18133
rect 58930 -18229 58964 -18167
rect 59662 -18229 59696 -18167
rect 58930 -18576 58964 -18515
rect 58930 -18610 59026 -18576
rect 59214 -18577 59310 -18576
rect 59662 -18577 59696 -18515
rect 59214 -18610 59696 -18577
rect 58930 -18611 59696 -18610
rect 55118 -19496 55518 -19484
rect 55118 -19530 55142 -19496
rect 55494 -19530 55518 -19496
rect 55118 -19581 55518 -19530
rect 55118 -19668 55518 -19617
rect 55118 -19702 55142 -19668
rect 55494 -19702 55518 -19668
rect 55118 -19714 55518 -19702
rect 53886 -20108 53982 -20074
rect 54956 -20108 55052 -20074
rect 53886 -20170 53920 -20108
rect 55018 -20170 55052 -20108
rect 53886 -20430 53920 -20368
rect 55018 -20430 55052 -20368
rect 56316 -18738 56412 -18704
rect 56610 -18738 56706 -18704
rect 56316 -18800 56350 -18738
rect 56672 -18800 56706 -18738
rect 58930 -18672 58964 -18611
rect 56316 -19836 56350 -19774
rect 59276 -18672 59310 -18611
rect 58930 -19306 58964 -19246
rect 59276 -19306 59310 -19246
rect 58930 -19342 59310 -19306
rect 58930 -19402 58964 -19342
rect 56672 -19836 56706 -19774
rect 56316 -19870 56412 -19836
rect 56610 -19870 56706 -19836
rect 59276 -19402 59310 -19342
rect 58930 -20038 58964 -19976
rect 60466 -19660 60546 -19630
rect 60466 -19700 60486 -19660
rect 60526 -19700 60546 -19660
rect 60466 -19730 60546 -19700
rect 60606 -19660 60686 -19630
rect 60606 -19700 60626 -19660
rect 60666 -19700 60686 -19660
rect 60606 -19730 60686 -19700
rect 60746 -19660 60826 -19630
rect 60746 -19700 60766 -19660
rect 60806 -19700 60826 -19660
rect 60746 -19730 60826 -19700
rect 60886 -19660 60966 -19630
rect 60886 -19700 60906 -19660
rect 60946 -19700 60966 -19660
rect 60886 -19730 60966 -19700
rect 59276 -20038 59310 -19976
rect 58930 -20072 59026 -20038
rect 59214 -20040 59310 -20038
rect 59214 -20072 59696 -20040
rect 58930 -20074 59696 -20072
rect 58930 -20136 58964 -20074
rect 53886 -20464 53982 -20430
rect 54956 -20464 55052 -20430
rect 59662 -20136 59696 -20074
rect 53886 -20526 53920 -20464
rect 55018 -20526 55052 -20464
rect 53886 -20786 53920 -20724
rect 57156 -20490 57316 -20460
rect 57156 -20590 57186 -20490
rect 57286 -20590 57316 -20490
rect 58930 -20484 58964 -20422
rect 59662 -20484 59696 -20422
rect 58930 -20518 59026 -20484
rect 59600 -20518 59696 -20484
rect 57156 -20620 57316 -20590
rect 55018 -20786 55052 -20724
rect 53886 -20820 53982 -20786
rect 54956 -20820 55052 -20786
rect 53896 -23192 53992 -23158
rect 54966 -23192 55062 -23158
rect 53896 -23254 53930 -23192
rect 55028 -23254 55062 -23192
rect 53896 -23514 53930 -23452
rect 55028 -23514 55062 -23452
rect 53896 -23548 53992 -23514
rect 54966 -23548 55062 -23514
rect 53896 -23610 53930 -23548
rect 55028 -23610 55062 -23548
rect 57126 -23500 57356 -23470
rect 53896 -23870 53930 -23808
rect 55028 -23870 55062 -23808
rect 53896 -23904 53992 -23870
rect 54966 -23904 55062 -23870
rect 55118 -24274 55518 -24262
rect 55118 -24308 55142 -24274
rect 55494 -24308 55518 -24274
rect 55118 -24359 55518 -24308
rect 55118 -24446 55518 -24395
rect 55118 -24480 55142 -24446
rect 55494 -24480 55518 -24446
rect 55118 -24492 55518 -24480
rect 57126 -23570 57156 -23500
rect 57316 -23570 57356 -23500
rect 57126 -23600 57356 -23570
rect 58930 -23567 59026 -23533
rect 59600 -23567 59696 -23533
rect 58930 -23629 58964 -23567
rect 59662 -23629 59696 -23567
rect 58930 -23976 58964 -23915
rect 58930 -24010 59026 -23976
rect 59214 -23977 59310 -23976
rect 59662 -23977 59696 -23915
rect 59214 -24010 59696 -23977
rect 58930 -24011 59696 -24010
rect 55118 -24896 55518 -24884
rect 55118 -24930 55142 -24896
rect 55494 -24930 55518 -24896
rect 55118 -24981 55518 -24930
rect 55118 -25068 55518 -25017
rect 55118 -25102 55142 -25068
rect 55494 -25102 55518 -25068
rect 55118 -25114 55518 -25102
rect 53886 -25508 53982 -25474
rect 54956 -25508 55052 -25474
rect 53886 -25570 53920 -25508
rect 55018 -25570 55052 -25508
rect 53886 -25830 53920 -25768
rect 55018 -25830 55052 -25768
rect 56316 -24138 56412 -24104
rect 56610 -24138 56706 -24104
rect 56316 -24200 56350 -24138
rect 56672 -24200 56706 -24138
rect 58930 -24072 58964 -24011
rect 56316 -25236 56350 -25174
rect 59276 -24072 59310 -24011
rect 58930 -24706 58964 -24646
rect 59276 -24706 59310 -24646
rect 58930 -24742 59310 -24706
rect 58930 -24802 58964 -24742
rect 56672 -25236 56706 -25174
rect 56316 -25270 56412 -25236
rect 56610 -25270 56706 -25236
rect 59276 -24802 59310 -24742
rect 58930 -25438 58964 -25376
rect 60466 -25060 60546 -25030
rect 60466 -25100 60486 -25060
rect 60526 -25100 60546 -25060
rect 60466 -25130 60546 -25100
rect 60606 -25060 60686 -25030
rect 60606 -25100 60626 -25060
rect 60666 -25100 60686 -25060
rect 60606 -25130 60686 -25100
rect 60746 -25060 60826 -25030
rect 60746 -25100 60766 -25060
rect 60806 -25100 60826 -25060
rect 60746 -25130 60826 -25100
rect 60886 -25060 60966 -25030
rect 60886 -25100 60906 -25060
rect 60946 -25100 60966 -25060
rect 60886 -25130 60966 -25100
rect 59276 -25438 59310 -25376
rect 58930 -25472 59026 -25438
rect 59214 -25440 59310 -25438
rect 59214 -25472 59696 -25440
rect 58930 -25474 59696 -25472
rect 58930 -25536 58964 -25474
rect 53886 -25864 53982 -25830
rect 54956 -25864 55052 -25830
rect 59662 -25536 59696 -25474
rect 53886 -25926 53920 -25864
rect 55018 -25926 55052 -25864
rect 53886 -26186 53920 -26124
rect 57156 -25890 57316 -25860
rect 57156 -25990 57186 -25890
rect 57286 -25990 57316 -25890
rect 58930 -25884 58964 -25822
rect 59662 -25884 59696 -25822
rect 58930 -25918 59026 -25884
rect 59600 -25918 59696 -25884
rect 57156 -26020 57316 -25990
rect 55018 -26186 55052 -26124
rect 53886 -26220 53982 -26186
rect 54956 -26220 55052 -26186
rect 53896 -28592 53992 -28558
rect 54966 -28592 55062 -28558
rect 53896 -28654 53930 -28592
rect 55028 -28654 55062 -28592
rect 53896 -28914 53930 -28852
rect 55028 -28914 55062 -28852
rect 53896 -28948 53992 -28914
rect 54966 -28948 55062 -28914
rect 53896 -29010 53930 -28948
rect 55028 -29010 55062 -28948
rect 57126 -28900 57356 -28870
rect 53896 -29270 53930 -29208
rect 55028 -29270 55062 -29208
rect 53896 -29304 53992 -29270
rect 54966 -29304 55062 -29270
rect 55118 -29674 55518 -29662
rect 55118 -29708 55142 -29674
rect 55494 -29708 55518 -29674
rect 55118 -29759 55518 -29708
rect 55118 -29846 55518 -29795
rect 55118 -29880 55142 -29846
rect 55494 -29880 55518 -29846
rect 55118 -29892 55518 -29880
rect 57126 -28970 57156 -28900
rect 57316 -28970 57356 -28900
rect 57126 -29000 57356 -28970
rect 58930 -28967 59026 -28933
rect 59600 -28967 59696 -28933
rect 58930 -29029 58964 -28967
rect 59662 -29029 59696 -28967
rect 58930 -29376 58964 -29315
rect 58930 -29410 59026 -29376
rect 59214 -29377 59310 -29376
rect 59662 -29377 59696 -29315
rect 59214 -29410 59696 -29377
rect 58930 -29411 59696 -29410
rect 55118 -30296 55518 -30284
rect 55118 -30330 55142 -30296
rect 55494 -30330 55518 -30296
rect 55118 -30381 55518 -30330
rect 55118 -30468 55518 -30417
rect 55118 -30502 55142 -30468
rect 55494 -30502 55518 -30468
rect 55118 -30514 55518 -30502
rect 53886 -30908 53982 -30874
rect 54956 -30908 55052 -30874
rect 53886 -30970 53920 -30908
rect 55018 -30970 55052 -30908
rect 53886 -31230 53920 -31168
rect 55018 -31230 55052 -31168
rect 56316 -29538 56412 -29504
rect 56610 -29538 56706 -29504
rect 56316 -29600 56350 -29538
rect 56672 -29600 56706 -29538
rect 58930 -29472 58964 -29411
rect 56316 -30636 56350 -30574
rect 59276 -29472 59310 -29411
rect 58930 -30106 58964 -30046
rect 59276 -30106 59310 -30046
rect 58930 -30142 59310 -30106
rect 58930 -30202 58964 -30142
rect 56672 -30636 56706 -30574
rect 56316 -30670 56412 -30636
rect 56610 -30670 56706 -30636
rect 59276 -30202 59310 -30142
rect 58930 -30838 58964 -30776
rect 60466 -30460 60546 -30430
rect 60466 -30500 60486 -30460
rect 60526 -30500 60546 -30460
rect 60466 -30530 60546 -30500
rect 60606 -30460 60686 -30430
rect 60606 -30500 60626 -30460
rect 60666 -30500 60686 -30460
rect 60606 -30530 60686 -30500
rect 60746 -30460 60826 -30430
rect 60746 -30500 60766 -30460
rect 60806 -30500 60826 -30460
rect 60746 -30530 60826 -30500
rect 60886 -30460 60966 -30430
rect 60886 -30500 60906 -30460
rect 60946 -30500 60966 -30460
rect 60886 -30530 60966 -30500
rect 59276 -30838 59310 -30776
rect 58930 -30872 59026 -30838
rect 59214 -30840 59310 -30838
rect 59214 -30872 59696 -30840
rect 58930 -30874 59696 -30872
rect 58930 -30936 58964 -30874
rect 53886 -31264 53982 -31230
rect 54956 -31264 55052 -31230
rect 59662 -30936 59696 -30874
rect 53886 -31326 53920 -31264
rect 55018 -31326 55052 -31264
rect 53886 -31586 53920 -31524
rect 57156 -31290 57316 -31260
rect 57156 -31390 57186 -31290
rect 57286 -31390 57316 -31290
rect 58930 -31284 58964 -31222
rect 59662 -31284 59696 -31222
rect 58930 -31318 59026 -31284
rect 59600 -31318 59696 -31284
rect 57156 -31420 57316 -31390
rect 55018 -31586 55052 -31524
rect 53886 -31620 53982 -31586
rect 54956 -31620 55052 -31586
rect 53896 -33992 53992 -33958
rect 54966 -33992 55062 -33958
rect 53896 -34054 53930 -33992
rect 55028 -34054 55062 -33992
rect 53896 -34314 53930 -34252
rect 55028 -34314 55062 -34252
rect 53896 -34348 53992 -34314
rect 54966 -34348 55062 -34314
rect 53896 -34410 53930 -34348
rect 55028 -34410 55062 -34348
rect 57126 -34300 57356 -34270
rect 53896 -34670 53930 -34608
rect 55028 -34670 55062 -34608
rect 53896 -34704 53992 -34670
rect 54966 -34704 55062 -34670
rect 55118 -35074 55518 -35062
rect 55118 -35108 55142 -35074
rect 55494 -35108 55518 -35074
rect 55118 -35159 55518 -35108
rect 55118 -35246 55518 -35195
rect 55118 -35280 55142 -35246
rect 55494 -35280 55518 -35246
rect 55118 -35292 55518 -35280
rect 57126 -34370 57156 -34300
rect 57316 -34370 57356 -34300
rect 57126 -34400 57356 -34370
rect 58930 -34367 59026 -34333
rect 59600 -34367 59696 -34333
rect 58930 -34429 58964 -34367
rect 59662 -34429 59696 -34367
rect 58930 -34776 58964 -34715
rect 58930 -34810 59026 -34776
rect 59214 -34777 59310 -34776
rect 59662 -34777 59696 -34715
rect 59214 -34810 59696 -34777
rect 58930 -34811 59696 -34810
rect 55118 -35696 55518 -35684
rect 55118 -35730 55142 -35696
rect 55494 -35730 55518 -35696
rect 55118 -35781 55518 -35730
rect 55118 -35868 55518 -35817
rect 55118 -35902 55142 -35868
rect 55494 -35902 55518 -35868
rect 55118 -35914 55518 -35902
rect 53886 -36308 53982 -36274
rect 54956 -36308 55052 -36274
rect 53886 -36370 53920 -36308
rect 55018 -36370 55052 -36308
rect 53886 -36630 53920 -36568
rect 55018 -36630 55052 -36568
rect 56316 -34938 56412 -34904
rect 56610 -34938 56706 -34904
rect 56316 -35000 56350 -34938
rect 56672 -35000 56706 -34938
rect 58930 -34872 58964 -34811
rect 56316 -36036 56350 -35974
rect 59276 -34872 59310 -34811
rect 58930 -35506 58964 -35446
rect 59276 -35506 59310 -35446
rect 58930 -35542 59310 -35506
rect 58930 -35602 58964 -35542
rect 56672 -36036 56706 -35974
rect 56316 -36070 56412 -36036
rect 56610 -36070 56706 -36036
rect 59276 -35602 59310 -35542
rect 58930 -36238 58964 -36176
rect 60466 -35860 60546 -35830
rect 60466 -35900 60486 -35860
rect 60526 -35900 60546 -35860
rect 60466 -35930 60546 -35900
rect 60606 -35860 60686 -35830
rect 60606 -35900 60626 -35860
rect 60666 -35900 60686 -35860
rect 60606 -35930 60686 -35900
rect 60746 -35860 60826 -35830
rect 60746 -35900 60766 -35860
rect 60806 -35900 60826 -35860
rect 60746 -35930 60826 -35900
rect 60886 -35860 60966 -35830
rect 60886 -35900 60906 -35860
rect 60946 -35900 60966 -35860
rect 60886 -35930 60966 -35900
rect 59276 -36238 59310 -36176
rect 58930 -36272 59026 -36238
rect 59214 -36240 59310 -36238
rect 59214 -36272 59696 -36240
rect 58930 -36274 59696 -36272
rect 58930 -36336 58964 -36274
rect 53886 -36664 53982 -36630
rect 54956 -36664 55052 -36630
rect 59662 -36336 59696 -36274
rect 53886 -36726 53920 -36664
rect 55018 -36726 55052 -36664
rect 53886 -36986 53920 -36924
rect 57156 -36690 57316 -36660
rect 57156 -36790 57186 -36690
rect 57286 -36790 57316 -36690
rect 58930 -36684 58964 -36622
rect 59662 -36684 59696 -36622
rect 58930 -36718 59026 -36684
rect 59600 -36718 59696 -36684
rect 57156 -36820 57316 -36790
rect 55018 -36986 55052 -36924
rect 53886 -37020 53982 -36986
rect 54956 -37020 55052 -36986
rect 76930 -38830 77040 -38800
rect 76930 -38880 76960 -38830
rect 77010 -38880 77040 -38830
rect 76930 -38960 77040 -38880
rect 80890 -38820 81070 -38790
rect 80890 -38930 80920 -38820
rect 81030 -38930 81070 -38820
rect 80890 -38960 81070 -38930
rect 81500 -38820 81680 -38790
rect 81500 -38930 81540 -38820
rect 81650 -38930 81680 -38820
rect 81500 -38960 81680 -38930
rect 82110 -38830 82290 -38800
rect 82110 -38940 82140 -38830
rect 82250 -38940 82290 -38830
rect 76930 -39010 76960 -38960
rect 77010 -39010 77040 -38960
rect 82110 -38970 82290 -38940
rect 82760 -38840 82940 -38810
rect 82760 -38950 82790 -38840
rect 82900 -38950 82940 -38840
rect 82760 -38980 82940 -38950
rect 83470 -38830 83650 -38800
rect 83470 -38940 83510 -38830
rect 83620 -38940 83650 -38830
rect 83470 -38970 83650 -38940
rect 84190 -38830 84370 -38800
rect 84190 -38940 84220 -38830
rect 84330 -38940 84370 -38830
rect 84190 -38970 84370 -38940
rect 85840 -38850 86020 -38820
rect 85840 -38960 85880 -38850
rect 85990 -38960 86020 -38850
rect 85840 -38990 86020 -38960
rect 87280 -38860 87460 -38830
rect 87280 -38970 87320 -38860
rect 87430 -38970 87460 -38860
rect 87280 -39000 87460 -38970
rect 76930 -39040 77040 -39010
rect 53896 -39392 53992 -39358
rect 54966 -39392 55062 -39358
rect 53896 -39454 53930 -39392
rect 55028 -39454 55062 -39392
rect 53896 -39714 53930 -39652
rect 55028 -39714 55062 -39652
rect 53896 -39748 53992 -39714
rect 54966 -39748 55062 -39714
rect 53896 -39810 53930 -39748
rect 55028 -39810 55062 -39748
rect 57126 -39700 57356 -39670
rect 53896 -40070 53930 -40008
rect 55028 -40070 55062 -40008
rect 53896 -40104 53992 -40070
rect 54966 -40104 55062 -40070
rect 55118 -40474 55518 -40462
rect 55118 -40508 55142 -40474
rect 55494 -40508 55518 -40474
rect 55118 -40559 55518 -40508
rect 55118 -40646 55518 -40595
rect 55118 -40680 55142 -40646
rect 55494 -40680 55518 -40646
rect 55118 -40692 55518 -40680
rect 57126 -39770 57156 -39700
rect 57316 -39770 57356 -39700
rect 57126 -39800 57356 -39770
rect 58930 -39767 59026 -39733
rect 59600 -39767 59696 -39733
rect 58930 -39829 58964 -39767
rect 59662 -39829 59696 -39767
rect 58930 -40176 58964 -40115
rect 58930 -40210 59026 -40176
rect 59214 -40177 59310 -40176
rect 59662 -40177 59696 -40115
rect 59214 -40210 59696 -40177
rect 58930 -40211 59696 -40210
rect 55118 -41096 55518 -41084
rect 55118 -41130 55142 -41096
rect 55494 -41130 55518 -41096
rect 55118 -41181 55518 -41130
rect 55118 -41268 55518 -41217
rect 55118 -41302 55142 -41268
rect 55494 -41302 55518 -41268
rect 55118 -41314 55518 -41302
rect 53886 -41708 53982 -41674
rect 54956 -41708 55052 -41674
rect 53886 -41770 53920 -41708
rect 55018 -41770 55052 -41708
rect 53886 -42030 53920 -41968
rect 55018 -42030 55052 -41968
rect 56316 -40338 56412 -40304
rect 56610 -40338 56706 -40304
rect 56316 -40400 56350 -40338
rect 56672 -40400 56706 -40338
rect 58930 -40272 58964 -40211
rect 56316 -41436 56350 -41374
rect 59276 -40272 59310 -40211
rect 58930 -40906 58964 -40846
rect 78250 -40250 78360 -40220
rect 78250 -40300 78280 -40250
rect 78330 -40300 78360 -40250
rect 78250 -40330 78360 -40300
rect 78560 -40250 78670 -40220
rect 78560 -40300 78590 -40250
rect 78640 -40300 78670 -40250
rect 78560 -40330 78670 -40300
rect 78800 -40250 78910 -40220
rect 78800 -40300 78830 -40250
rect 78880 -40300 78910 -40250
rect 78800 -40330 78910 -40300
rect 79060 -40250 79170 -40220
rect 79060 -40300 79090 -40250
rect 79140 -40300 79170 -40250
rect 79060 -40330 79170 -40300
rect 59276 -40906 59310 -40846
rect 58930 -40942 59310 -40906
rect 80850 -40360 81020 -40330
rect 80850 -40470 80880 -40360
rect 80990 -40470 81020 -40360
rect 80850 -40500 81020 -40470
rect 58930 -41002 58964 -40942
rect 56672 -41436 56706 -41374
rect 56316 -41470 56412 -41436
rect 56610 -41470 56706 -41436
rect 59276 -41002 59310 -40942
rect 58930 -41638 58964 -41576
rect 60466 -41260 60546 -41230
rect 60466 -41300 60486 -41260
rect 60526 -41300 60546 -41260
rect 60466 -41330 60546 -41300
rect 60606 -41260 60686 -41230
rect 60606 -41300 60626 -41260
rect 60666 -41300 60686 -41260
rect 60606 -41330 60686 -41300
rect 60746 -41260 60826 -41230
rect 60746 -41300 60766 -41260
rect 60806 -41300 60826 -41260
rect 60746 -41330 60826 -41300
rect 60886 -41260 60966 -41230
rect 60886 -41300 60906 -41260
rect 60946 -41300 60966 -41260
rect 60886 -41330 60966 -41300
rect 59276 -41638 59310 -41576
rect 58930 -41672 59026 -41638
rect 59214 -41640 59310 -41638
rect 59214 -41672 59696 -41640
rect 58930 -41674 59696 -41672
rect 58930 -41736 58964 -41674
rect 53886 -42064 53982 -42030
rect 54956 -42064 55052 -42030
rect 59662 -41736 59696 -41674
rect 53886 -42126 53920 -42064
rect 55018 -42126 55052 -42064
rect 53886 -42386 53920 -42324
rect 57156 -42090 57316 -42060
rect 57156 -42190 57186 -42090
rect 57286 -42190 57316 -42090
rect 58930 -42084 58964 -42022
rect 78630 -41490 78740 -41460
rect 78630 -41540 78660 -41490
rect 78710 -41540 78740 -41490
rect 78630 -41570 78740 -41540
rect 78850 -41490 78960 -41460
rect 78850 -41540 78880 -41490
rect 78930 -41540 78960 -41490
rect 78850 -41570 78960 -41540
rect 79090 -41490 79200 -41460
rect 79090 -41540 79120 -41490
rect 79170 -41540 79200 -41490
rect 79090 -41570 79200 -41540
rect 59662 -42084 59696 -42022
rect 58930 -42118 59026 -42084
rect 59600 -42118 59696 -42084
rect 57156 -42220 57316 -42190
rect 55018 -42386 55052 -42324
rect 53886 -42420 53982 -42386
rect 54956 -42420 55052 -42386
rect 78940 -42740 79050 -42710
rect 78940 -42790 78970 -42740
rect 79020 -42790 79050 -42740
rect 78940 -42820 79050 -42790
rect 79130 -42740 79240 -42710
rect 79130 -42790 79160 -42740
rect 79210 -42790 79240 -42740
rect 79130 -42820 79240 -42790
rect 83450 -43410 83620 -43380
rect 83450 -43520 83480 -43410
rect 83590 -43520 83620 -43410
rect 83450 -43550 83620 -43520
rect 85150 -43410 85320 -43380
rect 85150 -43520 85180 -43410
rect 85290 -43520 85320 -43410
rect 85150 -43550 85320 -43520
rect 86530 -43410 86700 -43380
rect 86530 -43520 86560 -43410
rect 86670 -43520 86700 -43410
rect 86530 -43550 86700 -43520
rect 87820 -43410 87990 -43380
rect 87820 -43520 87850 -43410
rect 87960 -43520 87990 -43410
rect 87820 -43550 87990 -43520
rect 89340 -43410 89510 -43380
rect 89340 -43520 89370 -43410
rect 89480 -43520 89510 -43410
rect 89340 -43550 89510 -43520
rect 90750 -43410 90920 -43380
rect 90750 -43520 90780 -43410
rect 90890 -43520 90920 -43410
rect 90750 -43550 90920 -43520
rect 78280 -43970 78390 -43940
rect 78280 -44020 78310 -43970
rect 78360 -44020 78390 -43970
rect 78280 -44050 78390 -44020
rect 78580 -43970 78690 -43940
rect 78580 -44020 78610 -43970
rect 78660 -44020 78690 -43970
rect 78580 -44050 78690 -44020
rect 78880 -43970 78990 -43940
rect 78880 -44020 78910 -43970
rect 78960 -44020 78990 -43970
rect 78880 -44050 78990 -44020
rect 53896 -44792 53992 -44758
rect 54966 -44792 55062 -44758
rect 53896 -44854 53930 -44792
rect 55028 -44854 55062 -44792
rect 53896 -45114 53930 -45052
rect 55028 -45114 55062 -45052
rect 53896 -45148 53992 -45114
rect 54966 -45148 55062 -45114
rect 53896 -45210 53930 -45148
rect 55028 -45210 55062 -45148
rect 57126 -45100 57356 -45070
rect 53896 -45470 53930 -45408
rect 55028 -45470 55062 -45408
rect 53896 -45504 53992 -45470
rect 54966 -45504 55062 -45470
rect 55118 -45874 55518 -45862
rect 55118 -45908 55142 -45874
rect 55494 -45908 55518 -45874
rect 55118 -45959 55518 -45908
rect 55118 -46046 55518 -45995
rect 55118 -46080 55142 -46046
rect 55494 -46080 55518 -46046
rect 55118 -46092 55518 -46080
rect 57126 -45170 57156 -45100
rect 57316 -45170 57356 -45100
rect 57126 -45200 57356 -45170
rect 58930 -45167 59026 -45133
rect 59600 -45167 59696 -45133
rect 58930 -45229 58964 -45167
rect 59662 -45229 59696 -45167
rect 58930 -45576 58964 -45515
rect 79120 -45210 79230 -45180
rect 79120 -45260 79150 -45210
rect 79200 -45260 79230 -45210
rect 79120 -45290 79230 -45260
rect 58930 -45610 59026 -45576
rect 59214 -45577 59310 -45576
rect 59662 -45577 59696 -45515
rect 59214 -45610 59696 -45577
rect 58930 -45611 59696 -45610
rect 55118 -46496 55518 -46484
rect 55118 -46530 55142 -46496
rect 55494 -46530 55518 -46496
rect 55118 -46581 55518 -46530
rect 55118 -46668 55518 -46617
rect 55118 -46702 55142 -46668
rect 55494 -46702 55518 -46668
rect 55118 -46714 55518 -46702
rect 53886 -47108 53982 -47074
rect 54956 -47108 55052 -47074
rect 53886 -47170 53920 -47108
rect 55018 -47170 55052 -47108
rect 53886 -47430 53920 -47368
rect 55018 -47430 55052 -47368
rect 56316 -45738 56412 -45704
rect 56610 -45738 56706 -45704
rect 56316 -45800 56350 -45738
rect 56672 -45800 56706 -45738
rect 58930 -45672 58964 -45611
rect 56316 -46836 56350 -46774
rect 59276 -45672 59310 -45611
rect 58930 -46306 58964 -46246
rect 59276 -46306 59310 -46246
rect 58930 -46342 59310 -46306
rect 58930 -46402 58964 -46342
rect 56672 -46836 56706 -46774
rect 56316 -46870 56412 -46836
rect 56610 -46870 56706 -46836
rect 59276 -46402 59310 -46342
rect 58930 -47038 58964 -46976
rect 60466 -46660 60546 -46630
rect 60466 -46700 60486 -46660
rect 60526 -46700 60546 -46660
rect 60466 -46730 60546 -46700
rect 60606 -46660 60686 -46630
rect 60606 -46700 60626 -46660
rect 60666 -46700 60686 -46660
rect 60606 -46730 60686 -46700
rect 60746 -46660 60826 -46630
rect 60746 -46700 60766 -46660
rect 60806 -46700 60826 -46660
rect 60746 -46730 60826 -46700
rect 60886 -46660 60966 -46630
rect 60886 -46700 60906 -46660
rect 60946 -46700 60966 -46660
rect 60886 -46730 60966 -46700
rect 59276 -47038 59310 -46976
rect 58930 -47072 59026 -47038
rect 59214 -47040 59310 -47038
rect 59214 -47072 59696 -47040
rect 58930 -47074 59696 -47072
rect 58930 -47136 58964 -47074
rect 53886 -47464 53982 -47430
rect 54956 -47464 55052 -47430
rect 59662 -47136 59696 -47074
rect 53886 -47526 53920 -47464
rect 55018 -47526 55052 -47464
rect 53886 -47786 53920 -47724
rect 57156 -47490 57316 -47460
rect 57156 -47590 57186 -47490
rect 57286 -47590 57316 -47490
rect 58930 -47484 58964 -47422
rect 76930 -46870 77040 -46840
rect 76930 -46920 76960 -46870
rect 77010 -46920 77040 -46870
rect 76930 -47000 77040 -46920
rect 76930 -47050 76960 -47000
rect 77010 -47050 77040 -47000
rect 76930 -47080 77040 -47050
rect 59662 -47484 59696 -47422
rect 58930 -47518 59026 -47484
rect 59600 -47518 59696 -47484
rect 57156 -47620 57316 -47590
rect 83454 -47548 83624 -47518
rect 55018 -47786 55052 -47724
rect 53886 -47820 53982 -47786
rect 54956 -47820 55052 -47786
rect 83454 -47658 83484 -47548
rect 83594 -47658 83624 -47548
rect 83454 -47688 83624 -47658
rect 85154 -47548 85324 -47518
rect 85154 -47658 85184 -47548
rect 85294 -47658 85324 -47548
rect 85154 -47688 85324 -47658
rect 86534 -47548 86704 -47518
rect 86534 -47658 86564 -47548
rect 86674 -47658 86704 -47548
rect 86534 -47688 86704 -47658
rect 87824 -47548 87994 -47518
rect 87824 -47658 87854 -47548
rect 87964 -47658 87994 -47548
rect 87824 -47688 87994 -47658
rect 89344 -47548 89514 -47518
rect 89344 -47658 89374 -47548
rect 89484 -47658 89514 -47548
rect 89344 -47688 89514 -47658
rect 90754 -47548 90924 -47518
rect 90754 -47658 90784 -47548
rect 90894 -47658 90924 -47548
rect 90754 -47688 90924 -47658
rect 78250 -48290 78360 -48260
rect 78250 -48340 78280 -48290
rect 78330 -48340 78360 -48290
rect 78250 -48370 78360 -48340
rect 78560 -48290 78670 -48260
rect 78560 -48340 78590 -48290
rect 78640 -48340 78670 -48290
rect 78560 -48370 78670 -48340
rect 78800 -48290 78910 -48260
rect 78800 -48340 78830 -48290
rect 78880 -48340 78910 -48290
rect 78800 -48370 78910 -48340
rect 79060 -48290 79170 -48260
rect 79060 -48340 79090 -48290
rect 79140 -48340 79170 -48290
rect 79060 -48370 79170 -48340
rect 78630 -49530 78740 -49500
rect 78630 -49580 78660 -49530
rect 78710 -49580 78740 -49530
rect 78630 -49610 78740 -49580
rect 78850 -49530 78960 -49500
rect 78850 -49580 78880 -49530
rect 78930 -49580 78960 -49530
rect 78850 -49610 78960 -49580
rect 79090 -49530 79200 -49500
rect 79090 -49580 79120 -49530
rect 79170 -49580 79200 -49530
rect 79090 -49610 79200 -49580
rect 53896 -50192 53992 -50158
rect 54966 -50192 55062 -50158
rect 53896 -50254 53930 -50192
rect 55028 -50254 55062 -50192
rect 53896 -50514 53930 -50452
rect 55028 -50514 55062 -50452
rect 53896 -50548 53992 -50514
rect 54966 -50548 55062 -50514
rect 53896 -50610 53930 -50548
rect 55028 -50610 55062 -50548
rect 57126 -50500 57356 -50470
rect 53896 -50870 53930 -50808
rect 55028 -50870 55062 -50808
rect 53896 -50904 53992 -50870
rect 54966 -50904 55062 -50870
rect 55118 -51274 55518 -51262
rect 55118 -51308 55142 -51274
rect 55494 -51308 55518 -51274
rect 55118 -51359 55518 -51308
rect 55118 -51446 55518 -51395
rect 55118 -51480 55142 -51446
rect 55494 -51480 55518 -51446
rect 55118 -51492 55518 -51480
rect 57126 -50570 57156 -50500
rect 57316 -50570 57356 -50500
rect 57126 -50600 57356 -50570
rect 58930 -50567 59026 -50533
rect 59600 -50567 59696 -50533
rect 58930 -50629 58964 -50567
rect 59662 -50629 59696 -50567
rect 58930 -50976 58964 -50915
rect 78940 -50780 79050 -50750
rect 78940 -50830 78970 -50780
rect 79020 -50830 79050 -50780
rect 58930 -51010 59026 -50976
rect 59214 -50977 59310 -50976
rect 59662 -50977 59696 -50915
rect 59214 -51010 59696 -50977
rect 58930 -51011 59696 -51010
rect 78940 -50860 79050 -50830
rect 79130 -50780 79240 -50750
rect 79130 -50830 79160 -50780
rect 79210 -50830 79240 -50780
rect 79130 -50860 79240 -50830
rect 55118 -51896 55518 -51884
rect 55118 -51930 55142 -51896
rect 55494 -51930 55518 -51896
rect 55118 -51981 55518 -51930
rect 55118 -52068 55518 -52017
rect 55118 -52102 55142 -52068
rect 55494 -52102 55518 -52068
rect 55118 -52114 55518 -52102
rect 53886 -52508 53982 -52474
rect 54956 -52508 55052 -52474
rect 53886 -52570 53920 -52508
rect 55018 -52570 55052 -52508
rect 53886 -52830 53920 -52768
rect 55018 -52830 55052 -52768
rect 56316 -51138 56412 -51104
rect 56610 -51138 56706 -51104
rect 56316 -51200 56350 -51138
rect 56672 -51200 56706 -51138
rect 58930 -51072 58964 -51011
rect 56316 -52236 56350 -52174
rect 59276 -51072 59310 -51011
rect 58930 -51706 58964 -51646
rect 59276 -51706 59310 -51646
rect 58930 -51742 59310 -51706
rect 83450 -51200 83620 -51170
rect 83450 -51310 83480 -51200
rect 83590 -51310 83620 -51200
rect 83450 -51340 83620 -51310
rect 85150 -51200 85320 -51170
rect 85150 -51310 85180 -51200
rect 85290 -51310 85320 -51200
rect 85150 -51340 85320 -51310
rect 86530 -51200 86700 -51170
rect 86530 -51310 86560 -51200
rect 86670 -51310 86700 -51200
rect 86530 -51340 86700 -51310
rect 87820 -51200 87990 -51170
rect 87820 -51310 87850 -51200
rect 87960 -51310 87990 -51200
rect 87820 -51340 87990 -51310
rect 89340 -51200 89510 -51170
rect 89340 -51310 89370 -51200
rect 89480 -51310 89510 -51200
rect 89340 -51340 89510 -51310
rect 90750 -51200 90920 -51170
rect 90750 -51310 90780 -51200
rect 90890 -51310 90920 -51200
rect 90750 -51340 90920 -51310
rect 58930 -51802 58964 -51742
rect 56672 -52236 56706 -52174
rect 56316 -52270 56412 -52236
rect 56610 -52270 56706 -52236
rect 59276 -51802 59310 -51742
rect 58930 -52438 58964 -52376
rect 78280 -52010 78390 -51980
rect 60466 -52060 60546 -52030
rect 60466 -52100 60486 -52060
rect 60526 -52100 60546 -52060
rect 60466 -52130 60546 -52100
rect 60606 -52060 60686 -52030
rect 60606 -52100 60626 -52060
rect 60666 -52100 60686 -52060
rect 60606 -52130 60686 -52100
rect 60746 -52060 60826 -52030
rect 60746 -52100 60766 -52060
rect 60806 -52100 60826 -52060
rect 60746 -52130 60826 -52100
rect 60886 -52060 60966 -52030
rect 60886 -52100 60906 -52060
rect 60946 -52100 60966 -52060
rect 78280 -52060 78310 -52010
rect 78360 -52060 78390 -52010
rect 78280 -52090 78390 -52060
rect 78580 -52010 78690 -51980
rect 78580 -52060 78610 -52010
rect 78660 -52060 78690 -52010
rect 78580 -52090 78690 -52060
rect 78880 -52010 78990 -51980
rect 78880 -52060 78910 -52010
rect 78960 -52060 78990 -52010
rect 78880 -52090 78990 -52060
rect 60886 -52130 60966 -52100
rect 59276 -52438 59310 -52376
rect 58930 -52472 59026 -52438
rect 59214 -52440 59310 -52438
rect 59214 -52472 59696 -52440
rect 58930 -52474 59696 -52472
rect 58930 -52536 58964 -52474
rect 53886 -52864 53982 -52830
rect 54956 -52864 55052 -52830
rect 59662 -52536 59696 -52474
rect 53886 -52926 53920 -52864
rect 55018 -52926 55052 -52864
rect 53886 -53186 53920 -53124
rect 57156 -52890 57316 -52860
rect 57156 -52990 57186 -52890
rect 57286 -52990 57316 -52890
rect 58930 -52884 58964 -52822
rect 59662 -52884 59696 -52822
rect 58930 -52918 59026 -52884
rect 59600 -52918 59696 -52884
rect 57156 -53020 57316 -52990
rect 55018 -53186 55052 -53124
rect 53886 -53220 53982 -53186
rect 54956 -53220 55052 -53186
rect 79120 -53250 79230 -53220
rect 79120 -53300 79150 -53250
rect 79200 -53300 79230 -53250
rect 79120 -53330 79230 -53300
rect 53896 -55592 53992 -55558
rect 54966 -55592 55062 -55558
rect 53896 -55654 53930 -55592
rect 55028 -55654 55062 -55592
rect 53896 -55914 53930 -55852
rect 55028 -55914 55062 -55852
rect 53896 -55948 53992 -55914
rect 54966 -55948 55062 -55914
rect 53896 -56010 53930 -55948
rect 55028 -56010 55062 -55948
rect 57126 -55900 57356 -55870
rect 53896 -56270 53930 -56208
rect 55028 -56270 55062 -56208
rect 53896 -56304 53992 -56270
rect 54966 -56304 55062 -56270
rect 55118 -56674 55518 -56662
rect 55118 -56708 55142 -56674
rect 55494 -56708 55518 -56674
rect 55118 -56759 55518 -56708
rect 55118 -56846 55518 -56795
rect 55118 -56880 55142 -56846
rect 55494 -56880 55518 -56846
rect 55118 -56892 55518 -56880
rect 57126 -55970 57156 -55900
rect 57316 -55970 57356 -55900
rect 57126 -56000 57356 -55970
rect 58930 -55967 59026 -55933
rect 59600 -55967 59696 -55933
rect 58930 -56029 58964 -55967
rect 59662 -56029 59696 -55967
rect 58930 -56376 58964 -56315
rect 58930 -56410 59026 -56376
rect 59214 -56377 59310 -56376
rect 59662 -56377 59696 -56315
rect 59214 -56410 59696 -56377
rect 58930 -56411 59696 -56410
rect 55118 -57296 55518 -57284
rect 55118 -57330 55142 -57296
rect 55494 -57330 55518 -57296
rect 55118 -57381 55518 -57330
rect 55118 -57468 55518 -57417
rect 55118 -57502 55142 -57468
rect 55494 -57502 55518 -57468
rect 55118 -57514 55518 -57502
rect 53886 -57908 53982 -57874
rect 54956 -57908 55052 -57874
rect 53886 -57970 53920 -57908
rect 55018 -57970 55052 -57908
rect 53886 -58230 53920 -58168
rect 55018 -58230 55052 -58168
rect 56316 -56538 56412 -56504
rect 56610 -56538 56706 -56504
rect 56316 -56600 56350 -56538
rect 56672 -56600 56706 -56538
rect 58930 -56472 58964 -56411
rect 56316 -57636 56350 -57574
rect 59276 -56472 59310 -56411
rect 58930 -57106 58964 -57046
rect 59276 -57106 59310 -57046
rect 58930 -57142 59310 -57106
rect 58930 -57202 58964 -57142
rect 56672 -57636 56706 -57574
rect 56316 -57670 56412 -57636
rect 56610 -57670 56706 -57636
rect 59276 -57202 59310 -57142
rect 58930 -57838 58964 -57776
rect 60466 -57460 60546 -57430
rect 60466 -57500 60486 -57460
rect 60526 -57500 60546 -57460
rect 60466 -57530 60546 -57500
rect 60606 -57460 60686 -57430
rect 60606 -57500 60626 -57460
rect 60666 -57500 60686 -57460
rect 60606 -57530 60686 -57500
rect 60746 -57460 60826 -57430
rect 60746 -57500 60766 -57460
rect 60806 -57500 60826 -57460
rect 60746 -57530 60826 -57500
rect 60886 -57460 60966 -57430
rect 60886 -57500 60906 -57460
rect 60946 -57500 60966 -57460
rect 60886 -57530 60966 -57500
rect 59276 -57838 59310 -57776
rect 58930 -57872 59026 -57838
rect 59214 -57840 59310 -57838
rect 59214 -57872 59696 -57840
rect 58930 -57874 59696 -57872
rect 58930 -57936 58964 -57874
rect 53886 -58264 53982 -58230
rect 54956 -58264 55052 -58230
rect 59662 -57936 59696 -57874
rect 53886 -58326 53920 -58264
rect 55018 -58326 55052 -58264
rect 53886 -58586 53920 -58524
rect 57156 -58290 57316 -58260
rect 57156 -58390 57186 -58290
rect 57286 -58390 57316 -58290
rect 58930 -58284 58964 -58222
rect 59662 -58284 59696 -58222
rect 58930 -58318 59026 -58284
rect 59600 -58318 59696 -58284
rect 57156 -58420 57316 -58390
rect 55018 -58586 55052 -58524
rect 53886 -58620 53982 -58586
rect 54956 -58620 55052 -58586
rect 53896 -60992 53992 -60958
rect 54966 -60992 55062 -60958
rect 53896 -61054 53930 -60992
rect 55028 -61054 55062 -60992
rect 53896 -61314 53930 -61252
rect 55028 -61314 55062 -61252
rect 53896 -61348 53992 -61314
rect 54966 -61348 55062 -61314
rect 53896 -61410 53930 -61348
rect 55028 -61410 55062 -61348
rect 57126 -61300 57356 -61270
rect 53896 -61670 53930 -61608
rect 55028 -61670 55062 -61608
rect 53896 -61704 53992 -61670
rect 54966 -61704 55062 -61670
rect 55118 -62074 55518 -62062
rect 55118 -62108 55142 -62074
rect 55494 -62108 55518 -62074
rect 55118 -62159 55518 -62108
rect 55118 -62246 55518 -62195
rect 55118 -62280 55142 -62246
rect 55494 -62280 55518 -62246
rect 55118 -62292 55518 -62280
rect 57126 -61370 57156 -61300
rect 57316 -61370 57356 -61300
rect 57126 -61400 57356 -61370
rect 58930 -61367 59026 -61333
rect 59600 -61367 59696 -61333
rect 58930 -61429 58964 -61367
rect 59662 -61429 59696 -61367
rect 58930 -61776 58964 -61715
rect 58930 -61810 59026 -61776
rect 59214 -61777 59310 -61776
rect 59662 -61777 59696 -61715
rect 59214 -61810 59696 -61777
rect 58930 -61811 59696 -61810
rect 55118 -62696 55518 -62684
rect 55118 -62730 55142 -62696
rect 55494 -62730 55518 -62696
rect 55118 -62781 55518 -62730
rect 55118 -62868 55518 -62817
rect 55118 -62902 55142 -62868
rect 55494 -62902 55518 -62868
rect 55118 -62914 55518 -62902
rect 53886 -63308 53982 -63274
rect 54956 -63308 55052 -63274
rect 53886 -63370 53920 -63308
rect 55018 -63370 55052 -63308
rect 53886 -63630 53920 -63568
rect 55018 -63630 55052 -63568
rect 56316 -61938 56412 -61904
rect 56610 -61938 56706 -61904
rect 56316 -62000 56350 -61938
rect 56672 -62000 56706 -61938
rect 58930 -61872 58964 -61811
rect 56316 -63036 56350 -62974
rect 59276 -61872 59310 -61811
rect 58930 -62506 58964 -62446
rect 59276 -62506 59310 -62446
rect 58930 -62542 59310 -62506
rect 58930 -62602 58964 -62542
rect 56672 -63036 56706 -62974
rect 56316 -63070 56412 -63036
rect 56610 -63070 56706 -63036
rect 59276 -62602 59310 -62542
rect 58930 -63238 58964 -63176
rect 60466 -62860 60546 -62830
rect 60466 -62900 60486 -62860
rect 60526 -62900 60546 -62860
rect 60466 -62930 60546 -62900
rect 60606 -62860 60686 -62830
rect 60606 -62900 60626 -62860
rect 60666 -62900 60686 -62860
rect 60606 -62930 60686 -62900
rect 60746 -62860 60826 -62830
rect 60746 -62900 60766 -62860
rect 60806 -62900 60826 -62860
rect 60746 -62930 60826 -62900
rect 60886 -62860 60966 -62830
rect 60886 -62900 60906 -62860
rect 60946 -62900 60966 -62860
rect 60886 -62930 60966 -62900
rect 59276 -63238 59310 -63176
rect 58930 -63272 59026 -63238
rect 59214 -63240 59310 -63238
rect 59214 -63272 59696 -63240
rect 58930 -63274 59696 -63272
rect 58930 -63336 58964 -63274
rect 53886 -63664 53982 -63630
rect 54956 -63664 55052 -63630
rect 59662 -63336 59696 -63274
rect 53886 -63726 53920 -63664
rect 55018 -63726 55052 -63664
rect 53886 -63986 53920 -63924
rect 57156 -63690 57316 -63660
rect 57156 -63790 57186 -63690
rect 57286 -63790 57316 -63690
rect 58930 -63684 58964 -63622
rect 59662 -63684 59696 -63622
rect 58930 -63718 59026 -63684
rect 59600 -63718 59696 -63684
rect 57156 -63820 57316 -63790
rect 55018 -63986 55052 -63924
rect 53886 -64020 53982 -63986
rect 54956 -64020 55052 -63986
rect 53896 -66392 53992 -66358
rect 54966 -66392 55062 -66358
rect 53896 -66454 53930 -66392
rect 55028 -66454 55062 -66392
rect 53896 -66714 53930 -66652
rect 55028 -66714 55062 -66652
rect 53896 -66748 53992 -66714
rect 54966 -66748 55062 -66714
rect 53896 -66810 53930 -66748
rect 55028 -66810 55062 -66748
rect 57126 -66700 57356 -66670
rect 53896 -67070 53930 -67008
rect 55028 -67070 55062 -67008
rect 53896 -67104 53992 -67070
rect 54966 -67104 55062 -67070
rect 55118 -67474 55518 -67462
rect 55118 -67508 55142 -67474
rect 55494 -67508 55518 -67474
rect 55118 -67559 55518 -67508
rect 55118 -67646 55518 -67595
rect 55118 -67680 55142 -67646
rect 55494 -67680 55518 -67646
rect 55118 -67692 55518 -67680
rect 57126 -66770 57156 -66700
rect 57316 -66770 57356 -66700
rect 57126 -66800 57356 -66770
rect 58930 -66767 59026 -66733
rect 59600 -66767 59696 -66733
rect 58930 -66829 58964 -66767
rect 59662 -66829 59696 -66767
rect 58930 -67176 58964 -67115
rect 58930 -67210 59026 -67176
rect 59214 -67177 59310 -67176
rect 59662 -67177 59696 -67115
rect 59214 -67210 59696 -67177
rect 58930 -67211 59696 -67210
rect 55118 -68096 55518 -68084
rect 55118 -68130 55142 -68096
rect 55494 -68130 55518 -68096
rect 55118 -68181 55518 -68130
rect 55118 -68268 55518 -68217
rect 55118 -68302 55142 -68268
rect 55494 -68302 55518 -68268
rect 55118 -68314 55518 -68302
rect 53886 -68708 53982 -68674
rect 54956 -68708 55052 -68674
rect 53886 -68770 53920 -68708
rect 55018 -68770 55052 -68708
rect 53886 -69030 53920 -68968
rect 55018 -69030 55052 -68968
rect 56316 -67338 56412 -67304
rect 56610 -67338 56706 -67304
rect 56316 -67400 56350 -67338
rect 56672 -67400 56706 -67338
rect 58930 -67272 58964 -67211
rect 56316 -68436 56350 -68374
rect 59276 -67272 59310 -67211
rect 58930 -67906 58964 -67846
rect 59276 -67906 59310 -67846
rect 58930 -67942 59310 -67906
rect 58930 -68002 58964 -67942
rect 56672 -68436 56706 -68374
rect 56316 -68470 56412 -68436
rect 56610 -68470 56706 -68436
rect 59276 -68002 59310 -67942
rect 58930 -68638 58964 -68576
rect 60466 -68260 60546 -68230
rect 60466 -68300 60486 -68260
rect 60526 -68300 60546 -68260
rect 60466 -68330 60546 -68300
rect 60606 -68260 60686 -68230
rect 60606 -68300 60626 -68260
rect 60666 -68300 60686 -68260
rect 60606 -68330 60686 -68300
rect 60746 -68260 60826 -68230
rect 60746 -68300 60766 -68260
rect 60806 -68300 60826 -68260
rect 60746 -68330 60826 -68300
rect 60886 -68260 60966 -68230
rect 60886 -68300 60906 -68260
rect 60946 -68300 60966 -68260
rect 60886 -68330 60966 -68300
rect 59276 -68638 59310 -68576
rect 58930 -68672 59026 -68638
rect 59214 -68640 59310 -68638
rect 59214 -68672 59696 -68640
rect 58930 -68674 59696 -68672
rect 58930 -68736 58964 -68674
rect 53886 -69064 53982 -69030
rect 54956 -69064 55052 -69030
rect 59662 -68736 59696 -68674
rect 53886 -69126 53920 -69064
rect 55018 -69126 55052 -69064
rect 53886 -69386 53920 -69324
rect 57156 -69090 57316 -69060
rect 57156 -69190 57186 -69090
rect 57286 -69190 57316 -69090
rect 58930 -69084 58964 -69022
rect 59662 -69084 59696 -69022
rect 58930 -69118 59026 -69084
rect 59600 -69118 59696 -69084
rect 57156 -69220 57316 -69190
rect 55018 -69386 55052 -69324
rect 53886 -69420 53982 -69386
rect 54956 -69420 55052 -69386
rect 53896 -71792 53992 -71758
rect 54966 -71792 55062 -71758
rect 53896 -71854 53930 -71792
rect 55028 -71854 55062 -71792
rect 53896 -72114 53930 -72052
rect 55028 -72114 55062 -72052
rect 53896 -72148 53992 -72114
rect 54966 -72148 55062 -72114
rect 53896 -72210 53930 -72148
rect 55028 -72210 55062 -72148
rect 57126 -72100 57356 -72070
rect 53896 -72470 53930 -72408
rect 55028 -72470 55062 -72408
rect 53896 -72504 53992 -72470
rect 54966 -72504 55062 -72470
rect 55118 -72874 55518 -72862
rect 55118 -72908 55142 -72874
rect 55494 -72908 55518 -72874
rect 55118 -72959 55518 -72908
rect 55118 -73046 55518 -72995
rect 55118 -73080 55142 -73046
rect 55494 -73080 55518 -73046
rect 55118 -73092 55518 -73080
rect 57126 -72170 57156 -72100
rect 57316 -72170 57356 -72100
rect 57126 -72200 57356 -72170
rect 58930 -72167 59026 -72133
rect 59600 -72167 59696 -72133
rect 58930 -72229 58964 -72167
rect 59662 -72229 59696 -72167
rect 58930 -72576 58964 -72515
rect 58930 -72610 59026 -72576
rect 59214 -72577 59310 -72576
rect 59662 -72577 59696 -72515
rect 59214 -72610 59696 -72577
rect 58930 -72611 59696 -72610
rect 55118 -73496 55518 -73484
rect 55118 -73530 55142 -73496
rect 55494 -73530 55518 -73496
rect 55118 -73581 55518 -73530
rect 55118 -73668 55518 -73617
rect 55118 -73702 55142 -73668
rect 55494 -73702 55518 -73668
rect 55118 -73714 55518 -73702
rect 53886 -74108 53982 -74074
rect 54956 -74108 55052 -74074
rect 53886 -74170 53920 -74108
rect 55018 -74170 55052 -74108
rect 53886 -74430 53920 -74368
rect 55018 -74430 55052 -74368
rect 56316 -72738 56412 -72704
rect 56610 -72738 56706 -72704
rect 56316 -72800 56350 -72738
rect 56672 -72800 56706 -72738
rect 58930 -72672 58964 -72611
rect 56316 -73836 56350 -73774
rect 59276 -72672 59310 -72611
rect 58930 -73306 58964 -73246
rect 59276 -73306 59310 -73246
rect 58930 -73342 59310 -73306
rect 58930 -73402 58964 -73342
rect 56672 -73836 56706 -73774
rect 56316 -73870 56412 -73836
rect 56610 -73870 56706 -73836
rect 59276 -73402 59310 -73342
rect 58930 -74038 58964 -73976
rect 60466 -73660 60546 -73630
rect 60466 -73700 60486 -73660
rect 60526 -73700 60546 -73660
rect 60466 -73730 60546 -73700
rect 60606 -73660 60686 -73630
rect 60606 -73700 60626 -73660
rect 60666 -73700 60686 -73660
rect 60606 -73730 60686 -73700
rect 60746 -73660 60826 -73630
rect 60746 -73700 60766 -73660
rect 60806 -73700 60826 -73660
rect 60746 -73730 60826 -73700
rect 60886 -73660 60966 -73630
rect 60886 -73700 60906 -73660
rect 60946 -73700 60966 -73660
rect 60886 -73730 60966 -73700
rect 59276 -74038 59310 -73976
rect 58930 -74072 59026 -74038
rect 59214 -74040 59310 -74038
rect 59214 -74072 59696 -74040
rect 58930 -74074 59696 -74072
rect 58930 -74136 58964 -74074
rect 53886 -74464 53982 -74430
rect 54956 -74464 55052 -74430
rect 59662 -74136 59696 -74074
rect 53886 -74526 53920 -74464
rect 55018 -74526 55052 -74464
rect 53886 -74786 53920 -74724
rect 57156 -74490 57316 -74460
rect 57156 -74590 57186 -74490
rect 57286 -74590 57316 -74490
rect 58930 -74484 58964 -74422
rect 59662 -74484 59696 -74422
rect 58930 -74518 59026 -74484
rect 59600 -74518 59696 -74484
rect 57156 -74620 57316 -74590
rect 55018 -74786 55052 -74724
rect 53886 -74820 53982 -74786
rect 54956 -74820 55052 -74786
rect 53896 -77192 53992 -77158
rect 54966 -77192 55062 -77158
rect 53896 -77254 53930 -77192
rect 55028 -77254 55062 -77192
rect 53896 -77514 53930 -77452
rect 55028 -77514 55062 -77452
rect 53896 -77548 53992 -77514
rect 54966 -77548 55062 -77514
rect 53896 -77610 53930 -77548
rect 55028 -77610 55062 -77548
rect 57126 -77500 57356 -77470
rect 53896 -77870 53930 -77808
rect 55028 -77870 55062 -77808
rect 53896 -77904 53992 -77870
rect 54966 -77904 55062 -77870
rect 55118 -78274 55518 -78262
rect 55118 -78308 55142 -78274
rect 55494 -78308 55518 -78274
rect 55118 -78359 55518 -78308
rect 55118 -78446 55518 -78395
rect 55118 -78480 55142 -78446
rect 55494 -78480 55518 -78446
rect 55118 -78492 55518 -78480
rect 57126 -77570 57156 -77500
rect 57316 -77570 57356 -77500
rect 57126 -77600 57356 -77570
rect 58930 -77567 59026 -77533
rect 59600 -77567 59696 -77533
rect 58930 -77629 58964 -77567
rect 59662 -77629 59696 -77567
rect 58930 -77976 58964 -77915
rect 58930 -78010 59026 -77976
rect 59214 -77977 59310 -77976
rect 59662 -77977 59696 -77915
rect 59214 -78010 59696 -77977
rect 58930 -78011 59696 -78010
rect 55118 -78896 55518 -78884
rect 55118 -78930 55142 -78896
rect 55494 -78930 55518 -78896
rect 55118 -78981 55518 -78930
rect 55118 -79068 55518 -79017
rect 55118 -79102 55142 -79068
rect 55494 -79102 55518 -79068
rect 55118 -79114 55518 -79102
rect 53886 -79508 53982 -79474
rect 54956 -79508 55052 -79474
rect 53886 -79570 53920 -79508
rect 55018 -79570 55052 -79508
rect 53886 -79830 53920 -79768
rect 55018 -79830 55052 -79768
rect 56316 -78138 56412 -78104
rect 56610 -78138 56706 -78104
rect 56316 -78200 56350 -78138
rect 56672 -78200 56706 -78138
rect 58930 -78072 58964 -78011
rect 56316 -79236 56350 -79174
rect 59276 -78072 59310 -78011
rect 58930 -78706 58964 -78646
rect 59276 -78706 59310 -78646
rect 58930 -78742 59310 -78706
rect 58930 -78802 58964 -78742
rect 56672 -79236 56706 -79174
rect 56316 -79270 56412 -79236
rect 56610 -79270 56706 -79236
rect 59276 -78802 59310 -78742
rect 58930 -79438 58964 -79376
rect 60466 -79060 60546 -79030
rect 60466 -79100 60486 -79060
rect 60526 -79100 60546 -79060
rect 60466 -79130 60546 -79100
rect 60606 -79060 60686 -79030
rect 60606 -79100 60626 -79060
rect 60666 -79100 60686 -79060
rect 60606 -79130 60686 -79100
rect 60746 -79060 60826 -79030
rect 60746 -79100 60766 -79060
rect 60806 -79100 60826 -79060
rect 60746 -79130 60826 -79100
rect 60886 -79060 60966 -79030
rect 60886 -79100 60906 -79060
rect 60946 -79100 60966 -79060
rect 60886 -79130 60966 -79100
rect 59276 -79438 59310 -79376
rect 58930 -79472 59026 -79438
rect 59214 -79440 59310 -79438
rect 59214 -79472 59696 -79440
rect 58930 -79474 59696 -79472
rect 58930 -79536 58964 -79474
rect 53886 -79864 53982 -79830
rect 54956 -79864 55052 -79830
rect 59662 -79536 59696 -79474
rect 53886 -79926 53920 -79864
rect 55018 -79926 55052 -79864
rect 53886 -80186 53920 -80124
rect 57156 -79890 57316 -79860
rect 57156 -79990 57186 -79890
rect 57286 -79990 57316 -79890
rect 58930 -79884 58964 -79822
rect 59662 -79884 59696 -79822
rect 58930 -79918 59026 -79884
rect 59600 -79918 59696 -79884
rect 57156 -80020 57316 -79990
rect 55018 -80186 55052 -80124
rect 53886 -80220 53982 -80186
rect 54956 -80220 55052 -80186
rect 53896 -82592 53992 -82558
rect 54966 -82592 55062 -82558
rect 53896 -82654 53930 -82592
rect 55028 -82654 55062 -82592
rect 53896 -82914 53930 -82852
rect 55028 -82914 55062 -82852
rect 53896 -82948 53992 -82914
rect 54966 -82948 55062 -82914
rect 53896 -83010 53930 -82948
rect 55028 -83010 55062 -82948
rect 57126 -82900 57356 -82870
rect 53896 -83270 53930 -83208
rect 55028 -83270 55062 -83208
rect 53896 -83304 53992 -83270
rect 54966 -83304 55062 -83270
rect 55118 -83674 55518 -83662
rect 55118 -83708 55142 -83674
rect 55494 -83708 55518 -83674
rect 55118 -83759 55518 -83708
rect 55118 -83846 55518 -83795
rect 55118 -83880 55142 -83846
rect 55494 -83880 55518 -83846
rect 55118 -83892 55518 -83880
rect 57126 -82970 57156 -82900
rect 57316 -82970 57356 -82900
rect 57126 -83000 57356 -82970
rect 58930 -82967 59026 -82933
rect 59600 -82967 59696 -82933
rect 58930 -83029 58964 -82967
rect 59662 -83029 59696 -82967
rect 58930 -83376 58964 -83315
rect 58930 -83410 59026 -83376
rect 59214 -83377 59310 -83376
rect 59662 -83377 59696 -83315
rect 59214 -83410 59696 -83377
rect 58930 -83411 59696 -83410
rect 55118 -84296 55518 -84284
rect 55118 -84330 55142 -84296
rect 55494 -84330 55518 -84296
rect 55118 -84381 55518 -84330
rect 55118 -84468 55518 -84417
rect 55118 -84502 55142 -84468
rect 55494 -84502 55518 -84468
rect 55118 -84514 55518 -84502
rect 53886 -84908 53982 -84874
rect 54956 -84908 55052 -84874
rect 53886 -84970 53920 -84908
rect 55018 -84970 55052 -84908
rect 53886 -85230 53920 -85168
rect 55018 -85230 55052 -85168
rect 56316 -83538 56412 -83504
rect 56610 -83538 56706 -83504
rect 56316 -83600 56350 -83538
rect 56672 -83600 56706 -83538
rect 58930 -83472 58964 -83411
rect 56316 -84636 56350 -84574
rect 59276 -83472 59310 -83411
rect 58930 -84106 58964 -84046
rect 59276 -84106 59310 -84046
rect 58930 -84142 59310 -84106
rect 58930 -84202 58964 -84142
rect 56672 -84636 56706 -84574
rect 56316 -84670 56412 -84636
rect 56610 -84670 56706 -84636
rect 59276 -84202 59310 -84142
rect 58930 -84838 58964 -84776
rect 60466 -84460 60546 -84430
rect 60466 -84500 60486 -84460
rect 60526 -84500 60546 -84460
rect 60466 -84530 60546 -84500
rect 60606 -84460 60686 -84430
rect 60606 -84500 60626 -84460
rect 60666 -84500 60686 -84460
rect 60606 -84530 60686 -84500
rect 60746 -84460 60826 -84430
rect 60746 -84500 60766 -84460
rect 60806 -84500 60826 -84460
rect 60746 -84530 60826 -84500
rect 60886 -84460 60966 -84430
rect 60886 -84500 60906 -84460
rect 60946 -84500 60966 -84460
rect 60886 -84530 60966 -84500
rect 59276 -84838 59310 -84776
rect 58930 -84872 59026 -84838
rect 59214 -84840 59310 -84838
rect 59214 -84872 59696 -84840
rect 58930 -84874 59696 -84872
rect 58930 -84936 58964 -84874
rect 53886 -85264 53982 -85230
rect 54956 -85264 55052 -85230
rect 59662 -84936 59696 -84874
rect 53886 -85326 53920 -85264
rect 55018 -85326 55052 -85264
rect 53886 -85586 53920 -85524
rect 57156 -85290 57316 -85260
rect 57156 -85390 57186 -85290
rect 57286 -85390 57316 -85290
rect 58930 -85284 58964 -85222
rect 59662 -85284 59696 -85222
rect 58930 -85318 59026 -85284
rect 59600 -85318 59696 -85284
rect 57156 -85420 57316 -85390
rect 55018 -85586 55052 -85524
rect 53886 -85620 53982 -85586
rect 54956 -85620 55052 -85586
<< psubdiffcont >>
rect 53350 -4074 53384 -2100
rect 55802 -1988 56050 -1954
rect 55272 -2100 55430 -2066
rect 55176 -2456 55210 -2162
rect 55492 -2456 55526 -2162
rect 55272 -2552 55430 -2518
rect 53852 -2698 54808 -2664
rect 53756 -3008 53790 -2760
rect 54870 -3008 54904 -2760
rect 55706 -3006 55740 -2050
rect 56112 -3006 56146 -2050
rect 59868 -2294 60424 -2260
rect 53852 -3104 54808 -3070
rect 53756 -3414 53790 -3166
rect 55160 -3108 55600 -3068
rect 55802 -3102 56050 -3068
rect 54870 -3414 54904 -3166
rect 53852 -3510 54808 -3476
rect 55262 -3658 55420 -3624
rect 53446 -4170 53694 -4136
rect 55166 -4014 55200 -3720
rect 55482 -4014 55516 -3720
rect 55262 -4110 55420 -4076
rect 55706 -4120 55740 -3164
rect 56112 -4120 56146 -3164
rect 57116 -2780 57346 -2710
rect 59772 -2534 59806 -2356
rect 60486 -2534 60520 -2356
rect 59484 -2630 59642 -2596
rect 59800 -2630 59958 -2596
rect 59388 -3048 59422 -2692
rect 60020 -3048 60054 -2692
rect 61216 -2860 61336 -2820
rect 57096 -3450 57376 -3370
rect 59387 -3561 59421 -3205
rect 60019 -3561 60053 -3205
rect 59483 -3657 59641 -3623
rect 59799 -3657 59957 -3623
rect 55802 -4216 56050 -4182
rect 59772 -3900 59806 -3722
rect 60486 -3900 60520 -3722
rect 59868 -3996 60424 -3962
rect 55272 -4478 55566 -4444
rect 55176 -4698 55210 -4540
rect 55628 -4698 55662 -4540
rect 55272 -4794 55566 -4760
rect 53350 -9474 53384 -7500
rect 55802 -7388 56050 -7354
rect 55272 -7500 55430 -7466
rect 55176 -7856 55210 -7562
rect 55492 -7856 55526 -7562
rect 55272 -7952 55430 -7918
rect 53852 -8098 54808 -8064
rect 53756 -8408 53790 -8160
rect 54870 -8408 54904 -8160
rect 55706 -8406 55740 -7450
rect 56112 -8406 56146 -7450
rect 59868 -7694 60424 -7660
rect 53852 -8504 54808 -8470
rect 53756 -8814 53790 -8566
rect 55160 -8508 55600 -8468
rect 55802 -8502 56050 -8468
rect 54870 -8814 54904 -8566
rect 53852 -8910 54808 -8876
rect 55262 -9058 55420 -9024
rect 53446 -9570 53694 -9536
rect 55166 -9414 55200 -9120
rect 55482 -9414 55516 -9120
rect 55262 -9510 55420 -9476
rect 55706 -9520 55740 -8564
rect 56112 -9520 56146 -8564
rect 57116 -8180 57346 -8110
rect 59772 -7934 59806 -7756
rect 60486 -7934 60520 -7756
rect 59484 -8030 59642 -7996
rect 59800 -8030 59958 -7996
rect 59388 -8448 59422 -8092
rect 60020 -8448 60054 -8092
rect 61216 -8260 61336 -8220
rect 57096 -8850 57376 -8770
rect 59387 -8961 59421 -8605
rect 60019 -8961 60053 -8605
rect 59483 -9057 59641 -9023
rect 59799 -9057 59957 -9023
rect 55802 -9616 56050 -9582
rect 59772 -9300 59806 -9122
rect 60486 -9300 60520 -9122
rect 59868 -9396 60424 -9362
rect 55272 -9878 55566 -9844
rect 55176 -10098 55210 -9940
rect 55628 -10098 55662 -9940
rect 55272 -10194 55566 -10160
rect 20252 -11850 20430 -11816
rect 20156 -12070 20190 -11912
rect 20492 -12070 20526 -11912
rect 16535 -12177 16783 -12143
rect 16941 -12177 17189 -12143
rect 17347 -12177 17595 -12143
rect 17753 -12177 18001 -12143
rect 18159 -12177 18407 -12143
rect 18565 -12177 18813 -12143
rect 18971 -12177 19219 -12143
rect 19377 -12177 19625 -12143
rect 19783 -12177 20031 -12143
rect 20189 -12177 20437 -12143
rect 20595 -12177 20843 -12143
rect 21001 -12177 21249 -12143
rect 21407 -12177 21655 -12143
rect 21813 -12177 22061 -12143
rect 22219 -12177 22467 -12143
rect 22625 -12177 22873 -12143
rect 23031 -12177 23279 -12143
rect 23437 -12177 23685 -12143
rect 23843 -12177 24091 -12143
rect 24249 -12177 24497 -12143
rect 24655 -12177 24903 -12143
rect 25061 -12177 25309 -12143
rect 16439 -13195 16473 -12239
rect 16845 -13195 16879 -12239
rect 17251 -13195 17285 -12239
rect 17657 -13195 17691 -12239
rect 18063 -13195 18097 -12239
rect 18469 -13195 18503 -12239
rect 18875 -13195 18909 -12239
rect 19281 -13195 19315 -12239
rect 19687 -13195 19721 -12239
rect 20093 -13195 20127 -12239
rect 20499 -13195 20533 -12239
rect 20905 -13195 20939 -12239
rect 21311 -13195 21345 -12239
rect 21717 -13195 21751 -12239
rect 22123 -13195 22157 -12239
rect 22529 -13195 22563 -12239
rect 22935 -13195 22969 -12239
rect 23341 -13195 23375 -12239
rect 23747 -13195 23781 -12239
rect 24153 -13195 24187 -12239
rect 24559 -13195 24593 -12239
rect 24965 -13195 24999 -12239
rect 25371 -13195 25405 -12239
rect 16535 -13291 16783 -13257
rect 16941 -13291 17189 -13257
rect 17347 -13291 17595 -13257
rect 17753 -13291 18001 -13257
rect 18159 -13291 18407 -13257
rect 18565 -13291 18813 -13257
rect 18971 -13291 19219 -13257
rect 19377 -13291 19625 -13257
rect 19783 -13291 20031 -13257
rect 20189 -13291 20437 -13257
rect 20595 -13291 20843 -13257
rect 21001 -13291 21249 -13257
rect 21407 -13291 21655 -13257
rect 21813 -13291 22061 -13257
rect 22219 -13291 22467 -13257
rect 22625 -13291 22873 -13257
rect 23031 -13291 23279 -13257
rect 23437 -13291 23685 -13257
rect 23843 -13291 24091 -13257
rect 24249 -13291 24497 -13257
rect 24655 -13291 24903 -13257
rect 25061 -13291 25309 -13257
rect 16532 -13420 34620 -13386
rect 16436 -14696 16470 -13482
rect 34682 -14696 34716 -13482
rect 16532 -14792 34620 -14758
rect 16436 -16068 16470 -14854
rect 34682 -16068 34716 -14854
rect 53350 -14874 53384 -12900
rect 55802 -12788 56050 -12754
rect 55272 -12900 55430 -12866
rect 55176 -13256 55210 -12962
rect 55492 -13256 55526 -12962
rect 55272 -13352 55430 -13318
rect 53852 -13498 54808 -13464
rect 53756 -13808 53790 -13560
rect 54870 -13808 54904 -13560
rect 55706 -13806 55740 -12850
rect 56112 -13806 56146 -12850
rect 59868 -13094 60424 -13060
rect 53852 -13904 54808 -13870
rect 53756 -14214 53790 -13966
rect 55160 -13908 55600 -13868
rect 55802 -13902 56050 -13868
rect 54870 -14214 54904 -13966
rect 53852 -14310 54808 -14276
rect 55262 -14458 55420 -14424
rect 53446 -14970 53694 -14936
rect 55166 -14814 55200 -14520
rect 55482 -14814 55516 -14520
rect 55262 -14910 55420 -14876
rect 55706 -14920 55740 -13964
rect 56112 -14920 56146 -13964
rect 57116 -13580 57346 -13510
rect 59772 -13334 59806 -13156
rect 60486 -13334 60520 -13156
rect 59484 -13430 59642 -13396
rect 59800 -13430 59958 -13396
rect 59388 -13848 59422 -13492
rect 60020 -13848 60054 -13492
rect 61216 -13660 61336 -13620
rect 57096 -14250 57376 -14170
rect 59387 -14361 59421 -14005
rect 60019 -14361 60053 -14005
rect 59483 -14457 59641 -14423
rect 59799 -14457 59957 -14423
rect 55802 -15016 56050 -14982
rect 59772 -14700 59806 -14522
rect 60486 -14700 60520 -14522
rect 59868 -14796 60424 -14762
rect 55272 -15278 55566 -15244
rect 55176 -15498 55210 -15340
rect 55628 -15498 55662 -15340
rect 55272 -15594 55566 -15560
rect 16532 -16164 34620 -16130
rect 53350 -20274 53384 -18300
rect 55802 -18188 56050 -18154
rect 55272 -18300 55430 -18266
rect 55176 -18656 55210 -18362
rect 55492 -18656 55526 -18362
rect 55272 -18752 55430 -18718
rect 53852 -18898 54808 -18864
rect 53756 -19208 53790 -18960
rect 54870 -19208 54904 -18960
rect 55706 -19206 55740 -18250
rect 56112 -19206 56146 -18250
rect 59868 -18494 60424 -18460
rect 53852 -19304 54808 -19270
rect 53756 -19614 53790 -19366
rect 55160 -19308 55600 -19268
rect 55802 -19302 56050 -19268
rect 54870 -19614 54904 -19366
rect 53852 -19710 54808 -19676
rect 55262 -19858 55420 -19824
rect 53446 -20370 53694 -20336
rect 55166 -20214 55200 -19920
rect 55482 -20214 55516 -19920
rect 55262 -20310 55420 -20276
rect 55706 -20320 55740 -19364
rect 56112 -20320 56146 -19364
rect 57116 -18980 57346 -18910
rect 59772 -18734 59806 -18556
rect 60486 -18734 60520 -18556
rect 59484 -18830 59642 -18796
rect 59800 -18830 59958 -18796
rect 59388 -19248 59422 -18892
rect 60020 -19248 60054 -18892
rect 61216 -19060 61336 -19020
rect 57096 -19650 57376 -19570
rect 59387 -19761 59421 -19405
rect 60019 -19761 60053 -19405
rect 59483 -19857 59641 -19823
rect 59799 -19857 59957 -19823
rect 55802 -20416 56050 -20382
rect 59772 -20100 59806 -19922
rect 60486 -20100 60520 -19922
rect 59868 -20196 60424 -20162
rect 55272 -20678 55566 -20644
rect 55176 -20898 55210 -20740
rect 55628 -20898 55662 -20740
rect 55272 -20994 55566 -20960
rect 53350 -25674 53384 -23700
rect 55802 -23588 56050 -23554
rect 55272 -23700 55430 -23666
rect 55176 -24056 55210 -23762
rect 55492 -24056 55526 -23762
rect 55272 -24152 55430 -24118
rect 53852 -24298 54808 -24264
rect 53756 -24608 53790 -24360
rect 54870 -24608 54904 -24360
rect 55706 -24606 55740 -23650
rect 56112 -24606 56146 -23650
rect 59868 -23894 60424 -23860
rect 53852 -24704 54808 -24670
rect 53756 -25014 53790 -24766
rect 55160 -24708 55600 -24668
rect 55802 -24702 56050 -24668
rect 54870 -25014 54904 -24766
rect 53852 -25110 54808 -25076
rect 55262 -25258 55420 -25224
rect 53446 -25770 53694 -25736
rect 55166 -25614 55200 -25320
rect 55482 -25614 55516 -25320
rect 55262 -25710 55420 -25676
rect 55706 -25720 55740 -24764
rect 56112 -25720 56146 -24764
rect 57116 -24380 57346 -24310
rect 59772 -24134 59806 -23956
rect 60486 -24134 60520 -23956
rect 59484 -24230 59642 -24196
rect 59800 -24230 59958 -24196
rect 59388 -24648 59422 -24292
rect 60020 -24648 60054 -24292
rect 61216 -24460 61336 -24420
rect 57096 -25050 57376 -24970
rect 59387 -25161 59421 -24805
rect 60019 -25161 60053 -24805
rect 59483 -25257 59641 -25223
rect 59799 -25257 59957 -25223
rect 55802 -25816 56050 -25782
rect 59772 -25500 59806 -25322
rect 60486 -25500 60520 -25322
rect 59868 -25596 60424 -25562
rect 55272 -26078 55566 -26044
rect 55176 -26298 55210 -26140
rect 55628 -26298 55662 -26140
rect 55272 -26394 55566 -26360
rect 25738 -32530 25772 -31094
rect 35804 -32530 35838 -31094
rect 53350 -31074 53384 -29100
rect 55802 -28988 56050 -28954
rect 55272 -29100 55430 -29066
rect 55176 -29456 55210 -29162
rect 55492 -29456 55526 -29162
rect 55272 -29552 55430 -29518
rect 53852 -29698 54808 -29664
rect 53756 -30008 53790 -29760
rect 54870 -30008 54904 -29760
rect 55706 -30006 55740 -29050
rect 56112 -30006 56146 -29050
rect 59868 -29294 60424 -29260
rect 53852 -30104 54808 -30070
rect 53756 -30414 53790 -30166
rect 55160 -30108 55600 -30068
rect 55802 -30102 56050 -30068
rect 54870 -30414 54904 -30166
rect 53852 -30510 54808 -30476
rect 55262 -30658 55420 -30624
rect 53446 -31170 53694 -31136
rect 55166 -31014 55200 -30720
rect 55482 -31014 55516 -30720
rect 55262 -31110 55420 -31076
rect 55706 -31120 55740 -30164
rect 56112 -31120 56146 -30164
rect 57116 -29780 57346 -29710
rect 59772 -29534 59806 -29356
rect 60486 -29534 60520 -29356
rect 59484 -29630 59642 -29596
rect 59800 -29630 59958 -29596
rect 59388 -30048 59422 -29692
rect 60020 -30048 60054 -29692
rect 61216 -29860 61336 -29820
rect 57096 -30450 57376 -30370
rect 59387 -30561 59421 -30205
rect 60019 -30561 60053 -30205
rect 59483 -30657 59641 -30623
rect 59799 -30657 59957 -30623
rect 55802 -31216 56050 -31182
rect 59772 -30900 59806 -30722
rect 60486 -30900 60520 -30722
rect 59868 -30996 60424 -30962
rect 55272 -31478 55566 -31444
rect 55176 -31698 55210 -31540
rect 55628 -31698 55662 -31540
rect 55272 -31794 55566 -31760
rect 25736 -34128 25770 -32692
rect 35802 -34128 35836 -32692
rect 25736 -35726 25770 -34290
rect 35802 -35726 35836 -34290
rect 25736 -37328 25770 -35892
rect 35802 -37328 35836 -35892
rect 53350 -36474 53384 -34500
rect 55802 -34388 56050 -34354
rect 55272 -34500 55430 -34466
rect 55176 -34856 55210 -34562
rect 55492 -34856 55526 -34562
rect 55272 -34952 55430 -34918
rect 53852 -35098 54808 -35064
rect 53756 -35408 53790 -35160
rect 54870 -35408 54904 -35160
rect 55706 -35406 55740 -34450
rect 56112 -35406 56146 -34450
rect 59868 -34694 60424 -34660
rect 53852 -35504 54808 -35470
rect 53756 -35814 53790 -35566
rect 55160 -35508 55600 -35468
rect 55802 -35502 56050 -35468
rect 54870 -35814 54904 -35566
rect 53852 -35910 54808 -35876
rect 55262 -36058 55420 -36024
rect 53446 -36570 53694 -36536
rect 55166 -36414 55200 -36120
rect 55482 -36414 55516 -36120
rect 55262 -36510 55420 -36476
rect 55706 -36520 55740 -35564
rect 56112 -36520 56146 -35564
rect 57116 -35180 57346 -35110
rect 59772 -34934 59806 -34756
rect 60486 -34934 60520 -34756
rect 59484 -35030 59642 -34996
rect 59800 -35030 59958 -34996
rect 59388 -35448 59422 -35092
rect 60020 -35448 60054 -35092
rect 61216 -35260 61336 -35220
rect 57096 -35850 57376 -35770
rect 59387 -35961 59421 -35605
rect 60019 -35961 60053 -35605
rect 59483 -36057 59641 -36023
rect 59799 -36057 59957 -36023
rect 55802 -36616 56050 -36582
rect 59772 -36300 59806 -36122
rect 60486 -36300 60520 -36122
rect 59868 -36396 60424 -36362
rect 55272 -36878 55566 -36844
rect 55176 -37098 55210 -36940
rect 55628 -37098 55662 -36940
rect 55272 -37194 55566 -37160
rect 25736 -38928 25770 -37492
rect 35802 -38928 35836 -37492
rect 77140 -38420 77190 -38370
rect 77140 -38540 77190 -38490
rect 25738 -40530 25772 -39094
rect 35804 -40530 35838 -39094
rect 77450 -39550 77510 -39490
rect 25736 -42128 25770 -40692
rect 35802 -42128 35836 -40692
rect 53350 -41874 53384 -39900
rect 55802 -39788 56050 -39754
rect 55272 -39900 55430 -39866
rect 55176 -40256 55210 -39962
rect 55492 -40256 55526 -39962
rect 55272 -40352 55430 -40318
rect 53852 -40498 54808 -40464
rect 53756 -40808 53790 -40560
rect 54870 -40808 54904 -40560
rect 55706 -40806 55740 -39850
rect 56112 -40806 56146 -39850
rect 77450 -39750 77510 -39690
rect 81620 -39910 81730 -39800
rect 82520 -39880 82630 -39770
rect 83780 -39890 83890 -39780
rect 85190 -39880 85300 -39770
rect 86350 -39890 86460 -39780
rect 87420 -39880 87530 -39770
rect 88530 -39870 88640 -39760
rect 59868 -40094 60424 -40060
rect 53852 -40904 54808 -40870
rect 53756 -41214 53790 -40966
rect 55160 -40908 55600 -40868
rect 55802 -40902 56050 -40868
rect 54870 -41214 54904 -40966
rect 53852 -41310 54808 -41276
rect 55262 -41458 55420 -41424
rect 53446 -41970 53694 -41936
rect 25736 -43726 25770 -42290
rect 35802 -43726 35836 -42290
rect 55166 -41814 55200 -41520
rect 55482 -41814 55516 -41520
rect 55262 -41910 55420 -41876
rect 55706 -41920 55740 -40964
rect 56112 -41920 56146 -40964
rect 57116 -40580 57346 -40510
rect 59772 -40334 59806 -40156
rect 60486 -40334 60520 -40156
rect 59484 -40430 59642 -40396
rect 59800 -40430 59958 -40396
rect 59388 -40848 59422 -40492
rect 60020 -40848 60054 -40492
rect 61216 -40660 61336 -40620
rect 77430 -40790 77490 -40730
rect 57096 -41250 57376 -41170
rect 59387 -41361 59421 -41005
rect 60019 -41361 60053 -41005
rect 77430 -41040 77490 -40980
rect 59483 -41457 59641 -41423
rect 59799 -41457 59957 -41423
rect 55802 -42016 56050 -41982
rect 59772 -41700 59806 -41522
rect 60486 -41700 60520 -41522
rect 59868 -41796 60424 -41762
rect 77450 -42050 77510 -41990
rect 77450 -42220 77510 -42160
rect 55272 -42278 55566 -42244
rect 55176 -42498 55210 -42340
rect 55628 -42498 55662 -42340
rect 55272 -42594 55566 -42560
rect 77440 -43300 77500 -43240
rect 77440 -43480 77500 -43420
rect 25736 -45328 25770 -43892
rect 35802 -45328 35836 -43892
rect 77430 -44470 77490 -44410
rect 83510 -44350 83620 -44240
rect 85150 -44360 85260 -44250
rect 86560 -44350 86670 -44240
rect 87940 -44350 88050 -44240
rect 89480 -44360 89590 -44250
rect 90760 -44360 90870 -44250
rect 77430 -44720 77490 -44660
rect 25736 -46926 25770 -45490
rect 35802 -46926 35836 -45490
rect 25736 -48520 25770 -47084
rect 35802 -48520 35836 -47084
rect 53350 -47274 53384 -45300
rect 55802 -45188 56050 -45154
rect 55272 -45300 55430 -45266
rect 55176 -45656 55210 -45362
rect 55492 -45656 55526 -45362
rect 55272 -45752 55430 -45718
rect 53852 -45898 54808 -45864
rect 53756 -46208 53790 -45960
rect 54870 -46208 54904 -45960
rect 55706 -46206 55740 -45250
rect 56112 -46206 56146 -45250
rect 59868 -45494 60424 -45460
rect 53852 -46304 54808 -46270
rect 53756 -46614 53790 -46366
rect 55160 -46308 55600 -46268
rect 55802 -46302 56050 -46268
rect 54870 -46614 54904 -46366
rect 53852 -46710 54808 -46676
rect 55262 -46858 55420 -46824
rect 53446 -47370 53694 -47336
rect 55166 -47214 55200 -46920
rect 55482 -47214 55516 -46920
rect 55262 -47310 55420 -47276
rect 55706 -47320 55740 -46364
rect 56112 -47320 56146 -46364
rect 57116 -45980 57346 -45910
rect 59772 -45734 59806 -45556
rect 60486 -45734 60520 -45556
rect 77420 -45720 77480 -45660
rect 59484 -45830 59642 -45796
rect 59800 -45830 59958 -45796
rect 59388 -46248 59422 -45892
rect 60020 -46248 60054 -45892
rect 61216 -46060 61336 -46020
rect 57096 -46650 57376 -46570
rect 59387 -46761 59421 -46405
rect 60019 -46761 60053 -46405
rect 77140 -46460 77190 -46410
rect 77140 -46580 77190 -46530
rect 59483 -46857 59641 -46823
rect 59799 -46857 59957 -46823
rect 55802 -47416 56050 -47382
rect 59772 -47100 59806 -46922
rect 60486 -47100 60520 -46922
rect 59868 -47196 60424 -47162
rect 77450 -47590 77510 -47530
rect 55272 -47678 55566 -47644
rect 55176 -47898 55210 -47740
rect 55628 -47898 55662 -47740
rect 77450 -47790 77510 -47730
rect 55272 -47994 55566 -47960
rect 25832 -48620 35740 -48586
rect 25736 -50118 25770 -48682
rect 35802 -50118 35836 -48682
rect 83514 -48488 83624 -48378
rect 85154 -48498 85264 -48388
rect 86564 -48488 86674 -48378
rect 87944 -48488 88054 -48378
rect 89484 -48498 89594 -48388
rect 90764 -48498 90874 -48388
rect 77430 -48830 77490 -48770
rect 77430 -49080 77490 -49020
rect 77450 -50090 77510 -50030
rect 25832 -50214 35740 -50180
rect 25736 -51720 25770 -50284
rect 35802 -51720 35836 -50284
rect 77450 -50260 77510 -50200
rect 25736 -53318 25770 -51882
rect 35802 -53318 35836 -51882
rect 53350 -52674 53384 -50700
rect 55802 -50588 56050 -50554
rect 55272 -50700 55430 -50666
rect 55176 -51056 55210 -50762
rect 55492 -51056 55526 -50762
rect 55272 -51152 55430 -51118
rect 53852 -51298 54808 -51264
rect 53756 -51608 53790 -51360
rect 54870 -51608 54904 -51360
rect 55706 -51606 55740 -50650
rect 56112 -51606 56146 -50650
rect 59868 -50894 60424 -50860
rect 53852 -51704 54808 -51670
rect 53756 -52014 53790 -51766
rect 55160 -51708 55600 -51668
rect 55802 -51702 56050 -51668
rect 54870 -52014 54904 -51766
rect 53852 -52110 54808 -52076
rect 55262 -52258 55420 -52224
rect 53446 -52770 53694 -52736
rect 55166 -52614 55200 -52320
rect 55482 -52614 55516 -52320
rect 55262 -52710 55420 -52676
rect 55706 -52720 55740 -51764
rect 56112 -52720 56146 -51764
rect 57116 -51380 57346 -51310
rect 59772 -51134 59806 -50956
rect 60486 -51134 60520 -50956
rect 59484 -51230 59642 -51196
rect 59800 -51230 59958 -51196
rect 59388 -51648 59422 -51292
rect 60020 -51648 60054 -51292
rect 77440 -51340 77500 -51280
rect 61216 -51460 61336 -51420
rect 77440 -51520 77500 -51460
rect 57096 -52050 57376 -51970
rect 59387 -52161 59421 -51805
rect 60019 -52161 60053 -51805
rect 59483 -52257 59641 -52223
rect 59799 -52257 59957 -52223
rect 55802 -52816 56050 -52782
rect 59772 -52500 59806 -52322
rect 60486 -52500 60520 -52322
rect 83510 -52140 83620 -52030
rect 85150 -52150 85260 -52040
rect 86560 -52140 86670 -52030
rect 87940 -52140 88050 -52030
rect 89480 -52150 89590 -52040
rect 90760 -52150 90870 -52040
rect 77430 -52510 77490 -52450
rect 59868 -52596 60424 -52562
rect 77430 -52760 77490 -52700
rect 55272 -53078 55566 -53044
rect 55176 -53298 55210 -53140
rect 55628 -53298 55662 -53140
rect 55272 -53394 55566 -53360
rect 25738 -54920 25772 -53484
rect 35804 -54920 35838 -53484
rect 77420 -53760 77480 -53700
rect 25736 -56518 25770 -55082
rect 35802 -56518 35836 -55082
rect 25736 -58118 25770 -56682
rect 35802 -58118 35836 -56682
rect 53350 -58074 53384 -56100
rect 55802 -55988 56050 -55954
rect 55272 -56100 55430 -56066
rect 55176 -56456 55210 -56162
rect 55492 -56456 55526 -56162
rect 55272 -56552 55430 -56518
rect 53852 -56698 54808 -56664
rect 53756 -57008 53790 -56760
rect 54870 -57008 54904 -56760
rect 55706 -57006 55740 -56050
rect 56112 -57006 56146 -56050
rect 59868 -56294 60424 -56260
rect 53852 -57104 54808 -57070
rect 53756 -57414 53790 -57166
rect 55160 -57108 55600 -57068
rect 55802 -57102 56050 -57068
rect 54870 -57414 54904 -57166
rect 53852 -57510 54808 -57476
rect 55262 -57658 55420 -57624
rect 53446 -58170 53694 -58136
rect 25832 -58214 35740 -58180
rect 55166 -58014 55200 -57720
rect 55482 -58014 55516 -57720
rect 55262 -58110 55420 -58076
rect 55706 -58120 55740 -57164
rect 56112 -58120 56146 -57164
rect 57116 -56780 57346 -56710
rect 59772 -56534 59806 -56356
rect 60486 -56534 60520 -56356
rect 59484 -56630 59642 -56596
rect 59800 -56630 59958 -56596
rect 59388 -57048 59422 -56692
rect 60020 -57048 60054 -56692
rect 61216 -56860 61336 -56820
rect 57096 -57450 57376 -57370
rect 59387 -57561 59421 -57205
rect 60019 -57561 60053 -57205
rect 59483 -57657 59641 -57623
rect 59799 -57657 59957 -57623
rect 55802 -58216 56050 -58182
rect 59772 -57900 59806 -57722
rect 60486 -57900 60520 -57722
rect 59868 -57996 60424 -57962
rect 55272 -58478 55566 -58444
rect 55176 -58698 55210 -58540
rect 55628 -58698 55662 -58540
rect 55272 -58794 55566 -58760
rect 53350 -63474 53384 -61500
rect 55802 -61388 56050 -61354
rect 55272 -61500 55430 -61466
rect 55176 -61856 55210 -61562
rect 55492 -61856 55526 -61562
rect 55272 -61952 55430 -61918
rect 53852 -62098 54808 -62064
rect 53756 -62408 53790 -62160
rect 54870 -62408 54904 -62160
rect 55706 -62406 55740 -61450
rect 56112 -62406 56146 -61450
rect 59868 -61694 60424 -61660
rect 53852 -62504 54808 -62470
rect 53756 -62814 53790 -62566
rect 55160 -62508 55600 -62468
rect 55802 -62502 56050 -62468
rect 54870 -62814 54904 -62566
rect 53852 -62910 54808 -62876
rect 55262 -63058 55420 -63024
rect 53446 -63570 53694 -63536
rect 55166 -63414 55200 -63120
rect 55482 -63414 55516 -63120
rect 55262 -63510 55420 -63476
rect 55706 -63520 55740 -62564
rect 56112 -63520 56146 -62564
rect 57116 -62180 57346 -62110
rect 59772 -61934 59806 -61756
rect 60486 -61934 60520 -61756
rect 59484 -62030 59642 -61996
rect 59800 -62030 59958 -61996
rect 59388 -62448 59422 -62092
rect 60020 -62448 60054 -62092
rect 61216 -62260 61336 -62220
rect 57096 -62850 57376 -62770
rect 59387 -62961 59421 -62605
rect 60019 -62961 60053 -62605
rect 59483 -63057 59641 -63023
rect 59799 -63057 59957 -63023
rect 55802 -63616 56050 -63582
rect 59772 -63300 59806 -63122
rect 60486 -63300 60520 -63122
rect 59868 -63396 60424 -63362
rect 55272 -63878 55566 -63844
rect 55176 -64098 55210 -63940
rect 55628 -64098 55662 -63940
rect 55272 -64194 55566 -64160
rect 53350 -68874 53384 -66900
rect 55802 -66788 56050 -66754
rect 55272 -66900 55430 -66866
rect 55176 -67256 55210 -66962
rect 55492 -67256 55526 -66962
rect 55272 -67352 55430 -67318
rect 53852 -67498 54808 -67464
rect 53756 -67808 53790 -67560
rect 54870 -67808 54904 -67560
rect 55706 -67806 55740 -66850
rect 56112 -67806 56146 -66850
rect 59868 -67094 60424 -67060
rect 53852 -67904 54808 -67870
rect 53756 -68214 53790 -67966
rect 55160 -67908 55600 -67868
rect 55802 -67902 56050 -67868
rect 54870 -68214 54904 -67966
rect 53852 -68310 54808 -68276
rect 55262 -68458 55420 -68424
rect 53446 -68970 53694 -68936
rect 55166 -68814 55200 -68520
rect 55482 -68814 55516 -68520
rect 55262 -68910 55420 -68876
rect 55706 -68920 55740 -67964
rect 56112 -68920 56146 -67964
rect 57116 -67580 57346 -67510
rect 59772 -67334 59806 -67156
rect 60486 -67334 60520 -67156
rect 59484 -67430 59642 -67396
rect 59800 -67430 59958 -67396
rect 59388 -67848 59422 -67492
rect 60020 -67848 60054 -67492
rect 61216 -67660 61336 -67620
rect 57096 -68250 57376 -68170
rect 59387 -68361 59421 -68005
rect 60019 -68361 60053 -68005
rect 59483 -68457 59641 -68423
rect 59799 -68457 59957 -68423
rect 55802 -69016 56050 -68982
rect 59772 -68700 59806 -68522
rect 60486 -68700 60520 -68522
rect 59868 -68796 60424 -68762
rect 55272 -69278 55566 -69244
rect 55176 -69498 55210 -69340
rect 55628 -69498 55662 -69340
rect 55272 -69594 55566 -69560
rect 53350 -74274 53384 -72300
rect 55802 -72188 56050 -72154
rect 55272 -72300 55430 -72266
rect 55176 -72656 55210 -72362
rect 55492 -72656 55526 -72362
rect 55272 -72752 55430 -72718
rect 53852 -72898 54808 -72864
rect 53756 -73208 53790 -72960
rect 54870 -73208 54904 -72960
rect 55706 -73206 55740 -72250
rect 56112 -73206 56146 -72250
rect 59868 -72494 60424 -72460
rect 53852 -73304 54808 -73270
rect 53756 -73614 53790 -73366
rect 55160 -73308 55600 -73268
rect 55802 -73302 56050 -73268
rect 54870 -73614 54904 -73366
rect 53852 -73710 54808 -73676
rect 55262 -73858 55420 -73824
rect 53446 -74370 53694 -74336
rect 55166 -74214 55200 -73920
rect 55482 -74214 55516 -73920
rect 55262 -74310 55420 -74276
rect 55706 -74320 55740 -73364
rect 56112 -74320 56146 -73364
rect 57116 -72980 57346 -72910
rect 59772 -72734 59806 -72556
rect 60486 -72734 60520 -72556
rect 59484 -72830 59642 -72796
rect 59800 -72830 59958 -72796
rect 59388 -73248 59422 -72892
rect 60020 -73248 60054 -72892
rect 61216 -73060 61336 -73020
rect 57096 -73650 57376 -73570
rect 59387 -73761 59421 -73405
rect 60019 -73761 60053 -73405
rect 59483 -73857 59641 -73823
rect 59799 -73857 59957 -73823
rect 55802 -74416 56050 -74382
rect 59772 -74100 59806 -73922
rect 60486 -74100 60520 -73922
rect 59868 -74196 60424 -74162
rect 55272 -74678 55566 -74644
rect 55176 -74898 55210 -74740
rect 55628 -74898 55662 -74740
rect 55272 -74994 55566 -74960
rect 53350 -79674 53384 -77700
rect 55802 -77588 56050 -77554
rect 55272 -77700 55430 -77666
rect 55176 -78056 55210 -77762
rect 55492 -78056 55526 -77762
rect 55272 -78152 55430 -78118
rect 53852 -78298 54808 -78264
rect 53756 -78608 53790 -78360
rect 54870 -78608 54904 -78360
rect 55706 -78606 55740 -77650
rect 56112 -78606 56146 -77650
rect 59868 -77894 60424 -77860
rect 53852 -78704 54808 -78670
rect 53756 -79014 53790 -78766
rect 55160 -78708 55600 -78668
rect 55802 -78702 56050 -78668
rect 54870 -79014 54904 -78766
rect 53852 -79110 54808 -79076
rect 55262 -79258 55420 -79224
rect 53446 -79770 53694 -79736
rect 55166 -79614 55200 -79320
rect 55482 -79614 55516 -79320
rect 55262 -79710 55420 -79676
rect 55706 -79720 55740 -78764
rect 56112 -79720 56146 -78764
rect 57116 -78380 57346 -78310
rect 59772 -78134 59806 -77956
rect 60486 -78134 60520 -77956
rect 59484 -78230 59642 -78196
rect 59800 -78230 59958 -78196
rect 59388 -78648 59422 -78292
rect 60020 -78648 60054 -78292
rect 61216 -78460 61336 -78420
rect 57096 -79050 57376 -78970
rect 59387 -79161 59421 -78805
rect 60019 -79161 60053 -78805
rect 59483 -79257 59641 -79223
rect 59799 -79257 59957 -79223
rect 55802 -79816 56050 -79782
rect 59772 -79500 59806 -79322
rect 60486 -79500 60520 -79322
rect 59868 -79596 60424 -79562
rect 55272 -80078 55566 -80044
rect 55176 -80298 55210 -80140
rect 55628 -80298 55662 -80140
rect 55272 -80394 55566 -80360
rect 53350 -85074 53384 -83100
rect 55802 -82988 56050 -82954
rect 55272 -83100 55430 -83066
rect 55176 -83456 55210 -83162
rect 55492 -83456 55526 -83162
rect 55272 -83552 55430 -83518
rect 53852 -83698 54808 -83664
rect 53756 -84008 53790 -83760
rect 54870 -84008 54904 -83760
rect 55706 -84006 55740 -83050
rect 56112 -84006 56146 -83050
rect 59868 -83294 60424 -83260
rect 53852 -84104 54808 -84070
rect 53756 -84414 53790 -84166
rect 55160 -84108 55600 -84068
rect 55802 -84102 56050 -84068
rect 54870 -84414 54904 -84166
rect 53852 -84510 54808 -84476
rect 55262 -84658 55420 -84624
rect 53446 -85170 53694 -85136
rect 55166 -85014 55200 -84720
rect 55482 -85014 55516 -84720
rect 55262 -85110 55420 -85076
rect 55706 -85120 55740 -84164
rect 56112 -85120 56146 -84164
rect 57116 -83780 57346 -83710
rect 59772 -83534 59806 -83356
rect 60486 -83534 60520 -83356
rect 59484 -83630 59642 -83596
rect 59800 -83630 59958 -83596
rect 59388 -84048 59422 -83692
rect 60020 -84048 60054 -83692
rect 61216 -83860 61336 -83820
rect 57096 -84450 57376 -84370
rect 59387 -84561 59421 -84205
rect 60019 -84561 60053 -84205
rect 59483 -84657 59641 -84623
rect 59799 -84657 59957 -84623
rect 55802 -85216 56050 -85182
rect 59772 -84900 59806 -84722
rect 60486 -84900 60520 -84722
rect 59868 -84996 60424 -84962
rect 55272 -85478 55566 -85444
rect 55176 -85698 55210 -85540
rect 55628 -85698 55662 -85540
rect 55272 -85794 55566 -85760
<< nsubdiffcont >>
rect 53992 -1592 54966 -1558
rect 53896 -1852 53930 -1654
rect 55028 -1852 55062 -1654
rect 53992 -1948 54966 -1914
rect 53896 -2208 53930 -2010
rect 55028 -2208 55062 -2010
rect 53992 -2304 54966 -2270
rect 55142 -2708 55494 -2674
rect 55142 -2880 55494 -2846
rect 57156 -1970 57316 -1900
rect 59026 -1967 59600 -1933
rect 58930 -2315 58964 -2029
rect 59662 -2315 59696 -2029
rect 59026 -2410 59214 -2376
rect 55142 -3330 55494 -3296
rect 55142 -3502 55494 -3468
rect 53982 -3908 54956 -3874
rect 53886 -4168 53920 -3970
rect 55018 -4168 55052 -3970
rect 56412 -2538 56610 -2504
rect 56316 -3574 56350 -2600
rect 56672 -3574 56706 -2600
rect 58930 -3046 58964 -2472
rect 59276 -3046 59310 -2472
rect 56412 -3670 56610 -3636
rect 58930 -3776 58964 -3202
rect 59276 -3776 59310 -3202
rect 60486 -3500 60526 -3460
rect 60626 -3500 60666 -3460
rect 60766 -3500 60806 -3460
rect 60906 -3500 60946 -3460
rect 59026 -3872 59214 -3838
rect 53982 -4264 54956 -4230
rect 58930 -4222 58964 -3936
rect 53886 -4524 53920 -4326
rect 55018 -4524 55052 -4326
rect 57186 -4390 57286 -4290
rect 59662 -4222 59696 -3936
rect 59026 -4318 59600 -4284
rect 53982 -4620 54956 -4586
rect 53992 -6992 54966 -6958
rect 53896 -7252 53930 -7054
rect 55028 -7252 55062 -7054
rect 53992 -7348 54966 -7314
rect 20828 -7707 21156 -7673
rect 21314 -7707 21642 -7673
rect 21800 -7707 22128 -7673
rect 20732 -11743 20766 -7769
rect 21218 -11743 21252 -7769
rect 21704 -11743 21738 -7769
rect 22190 -11743 22224 -7769
rect 53896 -7608 53930 -7410
rect 55028 -7608 55062 -7410
rect 53992 -7704 54966 -7670
rect 55142 -8108 55494 -8074
rect 55142 -8280 55494 -8246
rect 57156 -7370 57316 -7300
rect 59026 -7367 59600 -7333
rect 58930 -7715 58964 -7429
rect 59662 -7715 59696 -7429
rect 59026 -7810 59214 -7776
rect 55142 -8730 55494 -8696
rect 55142 -8902 55494 -8868
rect 53982 -9308 54956 -9274
rect 53886 -9568 53920 -9370
rect 55018 -9568 55052 -9370
rect 56412 -7938 56610 -7904
rect 56316 -8974 56350 -8000
rect 56672 -8974 56706 -8000
rect 58930 -8446 58964 -7872
rect 59276 -8446 59310 -7872
rect 56412 -9070 56610 -9036
rect 58930 -9176 58964 -8602
rect 59276 -9176 59310 -8602
rect 60486 -8900 60526 -8860
rect 60626 -8900 60666 -8860
rect 60766 -8900 60806 -8860
rect 60906 -8900 60946 -8860
rect 59026 -9272 59214 -9238
rect 53982 -9664 54956 -9630
rect 58930 -9622 58964 -9336
rect 53886 -9924 53920 -9726
rect 55018 -9924 55052 -9726
rect 57186 -9790 57286 -9690
rect 59662 -9622 59696 -9336
rect 59026 -9718 59600 -9684
rect 53982 -10020 54956 -9986
rect 20828 -11839 21156 -11805
rect 21314 -11839 21642 -11805
rect 21800 -11839 22128 -11805
rect 53992 -12392 54966 -12358
rect 53896 -12652 53930 -12454
rect 55028 -12652 55062 -12454
rect 53992 -12748 54966 -12714
rect 53896 -13008 53930 -12810
rect 55028 -13008 55062 -12810
rect 53992 -13104 54966 -13070
rect 55142 -13508 55494 -13474
rect 55142 -13680 55494 -13646
rect 57156 -12770 57316 -12700
rect 59026 -12767 59600 -12733
rect 58930 -13115 58964 -12829
rect 59662 -13115 59696 -12829
rect 59026 -13210 59214 -13176
rect 55142 -14130 55494 -14096
rect 55142 -14302 55494 -14268
rect 53982 -14708 54956 -14674
rect 53886 -14968 53920 -14770
rect 55018 -14968 55052 -14770
rect 56412 -13338 56610 -13304
rect 56316 -14374 56350 -13400
rect 56672 -14374 56706 -13400
rect 58930 -13846 58964 -13272
rect 59276 -13846 59310 -13272
rect 56412 -14470 56610 -14436
rect 58930 -14576 58964 -14002
rect 59276 -14576 59310 -14002
rect 60486 -14300 60526 -14260
rect 60626 -14300 60666 -14260
rect 60766 -14300 60806 -14260
rect 60906 -14300 60946 -14260
rect 59026 -14672 59214 -14638
rect 53982 -15064 54956 -15030
rect 58930 -15022 58964 -14736
rect 53886 -15324 53920 -15126
rect 55018 -15324 55052 -15126
rect 57186 -15190 57286 -15090
rect 59662 -15022 59696 -14736
rect 59026 -15118 59600 -15084
rect 53982 -15420 54956 -15386
rect 53992 -17792 54966 -17758
rect 53896 -18052 53930 -17854
rect 55028 -18052 55062 -17854
rect 53992 -18148 54966 -18114
rect 53896 -18408 53930 -18210
rect 55028 -18408 55062 -18210
rect 53992 -18504 54966 -18470
rect 55142 -18908 55494 -18874
rect 55142 -19080 55494 -19046
rect 57156 -18170 57316 -18100
rect 59026 -18167 59600 -18133
rect 58930 -18515 58964 -18229
rect 59662 -18515 59696 -18229
rect 59026 -18610 59214 -18576
rect 55142 -19530 55494 -19496
rect 55142 -19702 55494 -19668
rect 53982 -20108 54956 -20074
rect 53886 -20368 53920 -20170
rect 55018 -20368 55052 -20170
rect 56412 -18738 56610 -18704
rect 56316 -19774 56350 -18800
rect 56672 -19774 56706 -18800
rect 58930 -19246 58964 -18672
rect 59276 -19246 59310 -18672
rect 56412 -19870 56610 -19836
rect 58930 -19976 58964 -19402
rect 59276 -19976 59310 -19402
rect 60486 -19700 60526 -19660
rect 60626 -19700 60666 -19660
rect 60766 -19700 60806 -19660
rect 60906 -19700 60946 -19660
rect 59026 -20072 59214 -20038
rect 53982 -20464 54956 -20430
rect 58930 -20422 58964 -20136
rect 53886 -20724 53920 -20526
rect 55018 -20724 55052 -20526
rect 57186 -20590 57286 -20490
rect 59662 -20422 59696 -20136
rect 59026 -20518 59600 -20484
rect 53982 -20820 54956 -20786
rect 53992 -23192 54966 -23158
rect 53896 -23452 53930 -23254
rect 55028 -23452 55062 -23254
rect 53992 -23548 54966 -23514
rect 53896 -23808 53930 -23610
rect 55028 -23808 55062 -23610
rect 53992 -23904 54966 -23870
rect 55142 -24308 55494 -24274
rect 55142 -24480 55494 -24446
rect 57156 -23570 57316 -23500
rect 59026 -23567 59600 -23533
rect 58930 -23915 58964 -23629
rect 59662 -23915 59696 -23629
rect 59026 -24010 59214 -23976
rect 55142 -24930 55494 -24896
rect 55142 -25102 55494 -25068
rect 53982 -25508 54956 -25474
rect 53886 -25768 53920 -25570
rect 55018 -25768 55052 -25570
rect 56412 -24138 56610 -24104
rect 56316 -25174 56350 -24200
rect 56672 -25174 56706 -24200
rect 58930 -24646 58964 -24072
rect 59276 -24646 59310 -24072
rect 56412 -25270 56610 -25236
rect 58930 -25376 58964 -24802
rect 59276 -25376 59310 -24802
rect 60486 -25100 60526 -25060
rect 60626 -25100 60666 -25060
rect 60766 -25100 60806 -25060
rect 60906 -25100 60946 -25060
rect 59026 -25472 59214 -25438
rect 53982 -25864 54956 -25830
rect 58930 -25822 58964 -25536
rect 53886 -26124 53920 -25926
rect 55018 -26124 55052 -25926
rect 57186 -25990 57286 -25890
rect 59662 -25822 59696 -25536
rect 59026 -25918 59600 -25884
rect 53982 -26220 54956 -26186
rect 53992 -28592 54966 -28558
rect 53896 -28852 53930 -28654
rect 55028 -28852 55062 -28654
rect 53992 -28948 54966 -28914
rect 53896 -29208 53930 -29010
rect 55028 -29208 55062 -29010
rect 53992 -29304 54966 -29270
rect 55142 -29708 55494 -29674
rect 55142 -29880 55494 -29846
rect 57156 -28970 57316 -28900
rect 59026 -28967 59600 -28933
rect 58930 -29315 58964 -29029
rect 59662 -29315 59696 -29029
rect 59026 -29410 59214 -29376
rect 55142 -30330 55494 -30296
rect 55142 -30502 55494 -30468
rect 53982 -30908 54956 -30874
rect 53886 -31168 53920 -30970
rect 55018 -31168 55052 -30970
rect 56412 -29538 56610 -29504
rect 56316 -30574 56350 -29600
rect 56672 -30574 56706 -29600
rect 58930 -30046 58964 -29472
rect 59276 -30046 59310 -29472
rect 56412 -30670 56610 -30636
rect 58930 -30776 58964 -30202
rect 59276 -30776 59310 -30202
rect 60486 -30500 60526 -30460
rect 60626 -30500 60666 -30460
rect 60766 -30500 60806 -30460
rect 60906 -30500 60946 -30460
rect 59026 -30872 59214 -30838
rect 53982 -31264 54956 -31230
rect 58930 -31222 58964 -30936
rect 53886 -31524 53920 -31326
rect 55018 -31524 55052 -31326
rect 57186 -31390 57286 -31290
rect 59662 -31222 59696 -30936
rect 59026 -31318 59600 -31284
rect 53982 -31620 54956 -31586
rect 53992 -33992 54966 -33958
rect 53896 -34252 53930 -34054
rect 55028 -34252 55062 -34054
rect 53992 -34348 54966 -34314
rect 53896 -34608 53930 -34410
rect 55028 -34608 55062 -34410
rect 53992 -34704 54966 -34670
rect 55142 -35108 55494 -35074
rect 55142 -35280 55494 -35246
rect 57156 -34370 57316 -34300
rect 59026 -34367 59600 -34333
rect 58930 -34715 58964 -34429
rect 59662 -34715 59696 -34429
rect 59026 -34810 59214 -34776
rect 55142 -35730 55494 -35696
rect 55142 -35902 55494 -35868
rect 53982 -36308 54956 -36274
rect 53886 -36568 53920 -36370
rect 55018 -36568 55052 -36370
rect 56412 -34938 56610 -34904
rect 56316 -35974 56350 -35000
rect 56672 -35974 56706 -35000
rect 58930 -35446 58964 -34872
rect 59276 -35446 59310 -34872
rect 56412 -36070 56610 -36036
rect 58930 -36176 58964 -35602
rect 59276 -36176 59310 -35602
rect 60486 -35900 60526 -35860
rect 60626 -35900 60666 -35860
rect 60766 -35900 60806 -35860
rect 60906 -35900 60946 -35860
rect 59026 -36272 59214 -36238
rect 53982 -36664 54956 -36630
rect 58930 -36622 58964 -36336
rect 53886 -36924 53920 -36726
rect 55018 -36924 55052 -36726
rect 57186 -36790 57286 -36690
rect 59662 -36622 59696 -36336
rect 59026 -36718 59600 -36684
rect 53982 -37020 54956 -36986
rect 76960 -38880 77010 -38830
rect 80920 -38930 81030 -38820
rect 81540 -38930 81650 -38820
rect 82140 -38940 82250 -38830
rect 76960 -39010 77010 -38960
rect 82790 -38950 82900 -38840
rect 83510 -38940 83620 -38830
rect 84220 -38940 84330 -38830
rect 85880 -38960 85990 -38850
rect 87320 -38970 87430 -38860
rect 53992 -39392 54966 -39358
rect 53896 -39652 53930 -39454
rect 55028 -39652 55062 -39454
rect 53992 -39748 54966 -39714
rect 53896 -40008 53930 -39810
rect 55028 -40008 55062 -39810
rect 53992 -40104 54966 -40070
rect 55142 -40508 55494 -40474
rect 55142 -40680 55494 -40646
rect 57156 -39770 57316 -39700
rect 59026 -39767 59600 -39733
rect 58930 -40115 58964 -39829
rect 59662 -40115 59696 -39829
rect 59026 -40210 59214 -40176
rect 55142 -41130 55494 -41096
rect 55142 -41302 55494 -41268
rect 53982 -41708 54956 -41674
rect 53886 -41968 53920 -41770
rect 55018 -41968 55052 -41770
rect 56412 -40338 56610 -40304
rect 56316 -41374 56350 -40400
rect 56672 -41374 56706 -40400
rect 58930 -40846 58964 -40272
rect 59276 -40846 59310 -40272
rect 78280 -40300 78330 -40250
rect 78590 -40300 78640 -40250
rect 78830 -40300 78880 -40250
rect 79090 -40300 79140 -40250
rect 80880 -40470 80990 -40360
rect 56412 -41470 56610 -41436
rect 58930 -41576 58964 -41002
rect 59276 -41576 59310 -41002
rect 60486 -41300 60526 -41260
rect 60626 -41300 60666 -41260
rect 60766 -41300 60806 -41260
rect 60906 -41300 60946 -41260
rect 59026 -41672 59214 -41638
rect 53982 -42064 54956 -42030
rect 58930 -42022 58964 -41736
rect 53886 -42324 53920 -42126
rect 55018 -42324 55052 -42126
rect 57186 -42190 57286 -42090
rect 59662 -42022 59696 -41736
rect 78660 -41540 78710 -41490
rect 78880 -41540 78930 -41490
rect 79120 -41540 79170 -41490
rect 59026 -42118 59600 -42084
rect 53982 -42420 54956 -42386
rect 78970 -42790 79020 -42740
rect 79160 -42790 79210 -42740
rect 83480 -43520 83590 -43410
rect 85180 -43520 85290 -43410
rect 86560 -43520 86670 -43410
rect 87850 -43520 87960 -43410
rect 89370 -43520 89480 -43410
rect 90780 -43520 90890 -43410
rect 78310 -44020 78360 -43970
rect 78610 -44020 78660 -43970
rect 78910 -44020 78960 -43970
rect 53992 -44792 54966 -44758
rect 53896 -45052 53930 -44854
rect 55028 -45052 55062 -44854
rect 53992 -45148 54966 -45114
rect 53896 -45408 53930 -45210
rect 55028 -45408 55062 -45210
rect 53992 -45504 54966 -45470
rect 55142 -45908 55494 -45874
rect 55142 -46080 55494 -46046
rect 57156 -45170 57316 -45100
rect 59026 -45167 59600 -45133
rect 58930 -45515 58964 -45229
rect 59662 -45515 59696 -45229
rect 79150 -45260 79200 -45210
rect 59026 -45610 59214 -45576
rect 55142 -46530 55494 -46496
rect 55142 -46702 55494 -46668
rect 53982 -47108 54956 -47074
rect 53886 -47368 53920 -47170
rect 55018 -47368 55052 -47170
rect 56412 -45738 56610 -45704
rect 56316 -46774 56350 -45800
rect 56672 -46774 56706 -45800
rect 58930 -46246 58964 -45672
rect 59276 -46246 59310 -45672
rect 56412 -46870 56610 -46836
rect 58930 -46976 58964 -46402
rect 59276 -46976 59310 -46402
rect 60486 -46700 60526 -46660
rect 60626 -46700 60666 -46660
rect 60766 -46700 60806 -46660
rect 60906 -46700 60946 -46660
rect 59026 -47072 59214 -47038
rect 53982 -47464 54956 -47430
rect 58930 -47422 58964 -47136
rect 53886 -47724 53920 -47526
rect 55018 -47724 55052 -47526
rect 57186 -47590 57286 -47490
rect 59662 -47422 59696 -47136
rect 76960 -46920 77010 -46870
rect 76960 -47050 77010 -47000
rect 59026 -47518 59600 -47484
rect 53982 -47820 54956 -47786
rect 83484 -47658 83594 -47548
rect 85184 -47658 85294 -47548
rect 86564 -47658 86674 -47548
rect 87854 -47658 87964 -47548
rect 89374 -47658 89484 -47548
rect 90784 -47658 90894 -47548
rect 78280 -48340 78330 -48290
rect 78590 -48340 78640 -48290
rect 78830 -48340 78880 -48290
rect 79090 -48340 79140 -48290
rect 78660 -49580 78710 -49530
rect 78880 -49580 78930 -49530
rect 79120 -49580 79170 -49530
rect 53992 -50192 54966 -50158
rect 53896 -50452 53930 -50254
rect 55028 -50452 55062 -50254
rect 53992 -50548 54966 -50514
rect 53896 -50808 53930 -50610
rect 55028 -50808 55062 -50610
rect 53992 -50904 54966 -50870
rect 55142 -51308 55494 -51274
rect 55142 -51480 55494 -51446
rect 57156 -50570 57316 -50500
rect 59026 -50567 59600 -50533
rect 58930 -50915 58964 -50629
rect 59662 -50915 59696 -50629
rect 78970 -50830 79020 -50780
rect 59026 -51010 59214 -50976
rect 79160 -50830 79210 -50780
rect 55142 -51930 55494 -51896
rect 55142 -52102 55494 -52068
rect 53982 -52508 54956 -52474
rect 53886 -52768 53920 -52570
rect 55018 -52768 55052 -52570
rect 56412 -51138 56610 -51104
rect 56316 -52174 56350 -51200
rect 56672 -52174 56706 -51200
rect 58930 -51646 58964 -51072
rect 59276 -51646 59310 -51072
rect 83480 -51310 83590 -51200
rect 85180 -51310 85290 -51200
rect 86560 -51310 86670 -51200
rect 87850 -51310 87960 -51200
rect 89370 -51310 89480 -51200
rect 90780 -51310 90890 -51200
rect 56412 -52270 56610 -52236
rect 58930 -52376 58964 -51802
rect 59276 -52376 59310 -51802
rect 60486 -52100 60526 -52060
rect 60626 -52100 60666 -52060
rect 60766 -52100 60806 -52060
rect 60906 -52100 60946 -52060
rect 78310 -52060 78360 -52010
rect 78610 -52060 78660 -52010
rect 78910 -52060 78960 -52010
rect 59026 -52472 59214 -52438
rect 53982 -52864 54956 -52830
rect 58930 -52822 58964 -52536
rect 53886 -53124 53920 -52926
rect 55018 -53124 55052 -52926
rect 57186 -52990 57286 -52890
rect 59662 -52822 59696 -52536
rect 59026 -52918 59600 -52884
rect 53982 -53220 54956 -53186
rect 79150 -53300 79200 -53250
rect 53992 -55592 54966 -55558
rect 53896 -55852 53930 -55654
rect 55028 -55852 55062 -55654
rect 53992 -55948 54966 -55914
rect 53896 -56208 53930 -56010
rect 55028 -56208 55062 -56010
rect 53992 -56304 54966 -56270
rect 55142 -56708 55494 -56674
rect 55142 -56880 55494 -56846
rect 57156 -55970 57316 -55900
rect 59026 -55967 59600 -55933
rect 58930 -56315 58964 -56029
rect 59662 -56315 59696 -56029
rect 59026 -56410 59214 -56376
rect 55142 -57330 55494 -57296
rect 55142 -57502 55494 -57468
rect 53982 -57908 54956 -57874
rect 53886 -58168 53920 -57970
rect 55018 -58168 55052 -57970
rect 56412 -56538 56610 -56504
rect 56316 -57574 56350 -56600
rect 56672 -57574 56706 -56600
rect 58930 -57046 58964 -56472
rect 59276 -57046 59310 -56472
rect 56412 -57670 56610 -57636
rect 58930 -57776 58964 -57202
rect 59276 -57776 59310 -57202
rect 60486 -57500 60526 -57460
rect 60626 -57500 60666 -57460
rect 60766 -57500 60806 -57460
rect 60906 -57500 60946 -57460
rect 59026 -57872 59214 -57838
rect 53982 -58264 54956 -58230
rect 58930 -58222 58964 -57936
rect 53886 -58524 53920 -58326
rect 55018 -58524 55052 -58326
rect 57186 -58390 57286 -58290
rect 59662 -58222 59696 -57936
rect 59026 -58318 59600 -58284
rect 53982 -58620 54956 -58586
rect 53992 -60992 54966 -60958
rect 53896 -61252 53930 -61054
rect 55028 -61252 55062 -61054
rect 53992 -61348 54966 -61314
rect 53896 -61608 53930 -61410
rect 55028 -61608 55062 -61410
rect 53992 -61704 54966 -61670
rect 55142 -62108 55494 -62074
rect 55142 -62280 55494 -62246
rect 57156 -61370 57316 -61300
rect 59026 -61367 59600 -61333
rect 58930 -61715 58964 -61429
rect 59662 -61715 59696 -61429
rect 59026 -61810 59214 -61776
rect 55142 -62730 55494 -62696
rect 55142 -62902 55494 -62868
rect 53982 -63308 54956 -63274
rect 53886 -63568 53920 -63370
rect 55018 -63568 55052 -63370
rect 56412 -61938 56610 -61904
rect 56316 -62974 56350 -62000
rect 56672 -62974 56706 -62000
rect 58930 -62446 58964 -61872
rect 59276 -62446 59310 -61872
rect 56412 -63070 56610 -63036
rect 58930 -63176 58964 -62602
rect 59276 -63176 59310 -62602
rect 60486 -62900 60526 -62860
rect 60626 -62900 60666 -62860
rect 60766 -62900 60806 -62860
rect 60906 -62900 60946 -62860
rect 59026 -63272 59214 -63238
rect 53982 -63664 54956 -63630
rect 58930 -63622 58964 -63336
rect 53886 -63924 53920 -63726
rect 55018 -63924 55052 -63726
rect 57186 -63790 57286 -63690
rect 59662 -63622 59696 -63336
rect 59026 -63718 59600 -63684
rect 53982 -64020 54956 -63986
rect 53992 -66392 54966 -66358
rect 53896 -66652 53930 -66454
rect 55028 -66652 55062 -66454
rect 53992 -66748 54966 -66714
rect 53896 -67008 53930 -66810
rect 55028 -67008 55062 -66810
rect 53992 -67104 54966 -67070
rect 55142 -67508 55494 -67474
rect 55142 -67680 55494 -67646
rect 57156 -66770 57316 -66700
rect 59026 -66767 59600 -66733
rect 58930 -67115 58964 -66829
rect 59662 -67115 59696 -66829
rect 59026 -67210 59214 -67176
rect 55142 -68130 55494 -68096
rect 55142 -68302 55494 -68268
rect 53982 -68708 54956 -68674
rect 53886 -68968 53920 -68770
rect 55018 -68968 55052 -68770
rect 56412 -67338 56610 -67304
rect 56316 -68374 56350 -67400
rect 56672 -68374 56706 -67400
rect 58930 -67846 58964 -67272
rect 59276 -67846 59310 -67272
rect 56412 -68470 56610 -68436
rect 58930 -68576 58964 -68002
rect 59276 -68576 59310 -68002
rect 60486 -68300 60526 -68260
rect 60626 -68300 60666 -68260
rect 60766 -68300 60806 -68260
rect 60906 -68300 60946 -68260
rect 59026 -68672 59214 -68638
rect 53982 -69064 54956 -69030
rect 58930 -69022 58964 -68736
rect 53886 -69324 53920 -69126
rect 55018 -69324 55052 -69126
rect 57186 -69190 57286 -69090
rect 59662 -69022 59696 -68736
rect 59026 -69118 59600 -69084
rect 53982 -69420 54956 -69386
rect 53992 -71792 54966 -71758
rect 53896 -72052 53930 -71854
rect 55028 -72052 55062 -71854
rect 53992 -72148 54966 -72114
rect 53896 -72408 53930 -72210
rect 55028 -72408 55062 -72210
rect 53992 -72504 54966 -72470
rect 55142 -72908 55494 -72874
rect 55142 -73080 55494 -73046
rect 57156 -72170 57316 -72100
rect 59026 -72167 59600 -72133
rect 58930 -72515 58964 -72229
rect 59662 -72515 59696 -72229
rect 59026 -72610 59214 -72576
rect 55142 -73530 55494 -73496
rect 55142 -73702 55494 -73668
rect 53982 -74108 54956 -74074
rect 53886 -74368 53920 -74170
rect 55018 -74368 55052 -74170
rect 56412 -72738 56610 -72704
rect 56316 -73774 56350 -72800
rect 56672 -73774 56706 -72800
rect 58930 -73246 58964 -72672
rect 59276 -73246 59310 -72672
rect 56412 -73870 56610 -73836
rect 58930 -73976 58964 -73402
rect 59276 -73976 59310 -73402
rect 60486 -73700 60526 -73660
rect 60626 -73700 60666 -73660
rect 60766 -73700 60806 -73660
rect 60906 -73700 60946 -73660
rect 59026 -74072 59214 -74038
rect 53982 -74464 54956 -74430
rect 58930 -74422 58964 -74136
rect 53886 -74724 53920 -74526
rect 55018 -74724 55052 -74526
rect 57186 -74590 57286 -74490
rect 59662 -74422 59696 -74136
rect 59026 -74518 59600 -74484
rect 53982 -74820 54956 -74786
rect 53992 -77192 54966 -77158
rect 53896 -77452 53930 -77254
rect 55028 -77452 55062 -77254
rect 53992 -77548 54966 -77514
rect 53896 -77808 53930 -77610
rect 55028 -77808 55062 -77610
rect 53992 -77904 54966 -77870
rect 55142 -78308 55494 -78274
rect 55142 -78480 55494 -78446
rect 57156 -77570 57316 -77500
rect 59026 -77567 59600 -77533
rect 58930 -77915 58964 -77629
rect 59662 -77915 59696 -77629
rect 59026 -78010 59214 -77976
rect 55142 -78930 55494 -78896
rect 55142 -79102 55494 -79068
rect 53982 -79508 54956 -79474
rect 53886 -79768 53920 -79570
rect 55018 -79768 55052 -79570
rect 56412 -78138 56610 -78104
rect 56316 -79174 56350 -78200
rect 56672 -79174 56706 -78200
rect 58930 -78646 58964 -78072
rect 59276 -78646 59310 -78072
rect 56412 -79270 56610 -79236
rect 58930 -79376 58964 -78802
rect 59276 -79376 59310 -78802
rect 60486 -79100 60526 -79060
rect 60626 -79100 60666 -79060
rect 60766 -79100 60806 -79060
rect 60906 -79100 60946 -79060
rect 59026 -79472 59214 -79438
rect 53982 -79864 54956 -79830
rect 58930 -79822 58964 -79536
rect 53886 -80124 53920 -79926
rect 55018 -80124 55052 -79926
rect 57186 -79990 57286 -79890
rect 59662 -79822 59696 -79536
rect 59026 -79918 59600 -79884
rect 53982 -80220 54956 -80186
rect 53992 -82592 54966 -82558
rect 53896 -82852 53930 -82654
rect 55028 -82852 55062 -82654
rect 53992 -82948 54966 -82914
rect 53896 -83208 53930 -83010
rect 55028 -83208 55062 -83010
rect 53992 -83304 54966 -83270
rect 55142 -83708 55494 -83674
rect 55142 -83880 55494 -83846
rect 57156 -82970 57316 -82900
rect 59026 -82967 59600 -82933
rect 58930 -83315 58964 -83029
rect 59662 -83315 59696 -83029
rect 59026 -83410 59214 -83376
rect 55142 -84330 55494 -84296
rect 55142 -84502 55494 -84468
rect 53982 -84908 54956 -84874
rect 53886 -85168 53920 -84970
rect 55018 -85168 55052 -84970
rect 56412 -83538 56610 -83504
rect 56316 -84574 56350 -83600
rect 56672 -84574 56706 -83600
rect 58930 -84046 58964 -83472
rect 59276 -84046 59310 -83472
rect 56412 -84670 56610 -84636
rect 58930 -84776 58964 -84202
rect 59276 -84776 59310 -84202
rect 60486 -84500 60526 -84460
rect 60626 -84500 60666 -84460
rect 60766 -84500 60806 -84460
rect 60906 -84500 60946 -84460
rect 59026 -84872 59214 -84838
rect 53982 -85264 54956 -85230
rect 58930 -85222 58964 -84936
rect 53886 -85524 53920 -85326
rect 55018 -85524 55052 -85326
rect 57186 -85390 57286 -85290
rect 59662 -85222 59696 -84936
rect 59026 -85318 59600 -85284
rect 53982 -85620 54956 -85586
<< poly >>
rect 53982 -1734 54079 -1718
rect 53982 -1772 53998 -1734
rect 54032 -1772 54079 -1734
rect 53982 -1788 54079 -1772
rect 54879 -1734 54976 -1718
rect 54879 -1772 54926 -1734
rect 54960 -1772 54976 -1734
rect 54879 -1788 54976 -1772
rect 53510 -2106 53630 -2090
rect 53510 -2140 53526 -2106
rect 53614 -2140 53630 -2106
rect 53510 -2178 53630 -2140
rect 53982 -2090 54079 -2074
rect 53982 -2128 53998 -2090
rect 54032 -2128 54079 -2090
rect 53982 -2144 54079 -2128
rect 54879 -2090 54976 -2074
rect 54879 -2128 54926 -2090
rect 54960 -2128 54976 -2090
rect 54879 -2144 54976 -2128
rect 55318 -2168 55384 -2152
rect 55318 -2202 55334 -2168
rect 55368 -2202 55384 -2168
rect 55318 -2218 55384 -2202
rect 55336 -2240 55366 -2218
rect 55336 -2466 55366 -2440
rect 53510 -3016 53630 -2978
rect 53510 -3050 53526 -3016
rect 53614 -3050 53630 -3016
rect 53510 -3066 53630 -3050
rect 53842 -2840 53930 -2824
rect 53842 -2928 53858 -2840
rect 53892 -2928 53930 -2840
rect 53842 -2944 53930 -2928
rect 54730 -2840 54818 -2824
rect 54730 -2928 54768 -2840
rect 54802 -2928 54818 -2840
rect 54730 -2944 54818 -2928
rect 55030 -2759 55096 -2744
rect 55540 -2759 55606 -2744
rect 55030 -2760 55118 -2759
rect 55030 -2794 55046 -2760
rect 55080 -2794 55118 -2760
rect 55030 -2795 55118 -2794
rect 55518 -2760 55606 -2759
rect 55518 -2794 55556 -2760
rect 55590 -2794 55606 -2760
rect 55518 -2795 55606 -2794
rect 55030 -2810 55096 -2795
rect 55540 -2810 55606 -2795
rect 55866 -2056 55986 -2040
rect 55866 -2090 55882 -2056
rect 55970 -2090 55986 -2056
rect 55866 -2128 55986 -2090
rect 55866 -2966 55986 -2928
rect 55866 -3000 55882 -2966
rect 55970 -3000 55986 -2966
rect 55866 -3016 55986 -3000
rect 57175 -2109 57205 -2083
rect 57263 -2109 57293 -2083
rect 57175 -2282 57205 -2267
rect 57169 -2306 57205 -2282
rect 57169 -2341 57199 -2306
rect 57263 -2328 57293 -2267
rect 59544 -2093 59610 -2085
rect 59087 -2143 59113 -2093
rect 59513 -2101 59610 -2093
rect 59513 -2135 59560 -2101
rect 59594 -2135 59610 -2101
rect 59513 -2143 59610 -2135
rect 59544 -2151 59610 -2143
rect 59016 -2201 59082 -2193
rect 59016 -2209 59113 -2201
rect 59016 -2243 59032 -2209
rect 59066 -2243 59113 -2209
rect 59016 -2251 59113 -2243
rect 59513 -2251 59539 -2201
rect 59016 -2259 59082 -2251
rect 57123 -2357 57199 -2341
rect 57123 -2391 57133 -2357
rect 57167 -2391 57199 -2357
rect 57123 -2407 57199 -2391
rect 57241 -2344 57295 -2328
rect 57241 -2378 57251 -2344
rect 57285 -2378 57295 -2344
rect 57241 -2394 57295 -2378
rect 57169 -2416 57199 -2407
rect 57169 -2440 57205 -2416
rect 57175 -2455 57205 -2440
rect 57263 -2455 57293 -2394
rect 53510 -3124 53630 -3108
rect 53510 -3158 53526 -3124
rect 53614 -3158 53630 -3124
rect 53510 -3196 53630 -3158
rect 53842 -3246 53930 -3230
rect 53842 -3334 53858 -3246
rect 53892 -3334 53930 -3246
rect 53842 -3350 53930 -3334
rect 54730 -3246 54818 -3230
rect 54730 -3334 54768 -3246
rect 54802 -3334 54818 -3246
rect 54730 -3350 54818 -3334
rect 55030 -3381 55096 -3366
rect 55540 -3381 55606 -3366
rect 55030 -3382 55118 -3381
rect 55030 -3416 55046 -3382
rect 55080 -3416 55118 -3382
rect 55030 -3417 55118 -3416
rect 55518 -3382 55606 -3381
rect 55518 -3416 55556 -3382
rect 55590 -3416 55606 -3382
rect 55518 -3417 55606 -3416
rect 55030 -3432 55096 -3417
rect 53510 -4034 53630 -3996
rect 53510 -4068 53526 -4034
rect 53614 -4068 53630 -4034
rect 53510 -4084 53630 -4068
rect 55540 -3432 55606 -3417
rect 53972 -4050 54069 -4034
rect 53972 -4088 53988 -4050
rect 54022 -4088 54069 -4050
rect 53972 -4104 54069 -4088
rect 54869 -4050 54966 -4034
rect 54869 -4088 54916 -4050
rect 54950 -4088 54966 -4050
rect 54869 -4104 54966 -4088
rect 55326 -3736 55356 -3710
rect 55326 -3958 55356 -3936
rect 55308 -3974 55374 -3958
rect 55308 -4008 55324 -3974
rect 55358 -4008 55374 -3974
rect 55308 -4024 55374 -4008
rect 55866 -3170 55986 -3154
rect 55866 -3204 55882 -3170
rect 55970 -3204 55986 -3170
rect 55866 -3242 55986 -3204
rect 55866 -4080 55986 -4042
rect 55866 -4114 55882 -4080
rect 55970 -4114 55986 -4080
rect 55866 -4130 55986 -4114
rect 56476 -2606 56546 -2590
rect 56476 -2640 56492 -2606
rect 56530 -2640 56546 -2606
rect 56476 -2687 56546 -2640
rect 57175 -2585 57205 -2559
rect 57263 -2585 57293 -2559
rect 56476 -3534 56546 -3487
rect 56476 -3568 56492 -3534
rect 56530 -3568 56546 -3534
rect 56476 -3584 56546 -3568
rect 59087 -2478 59153 -2462
rect 59087 -2512 59103 -2478
rect 59137 -2512 59153 -2478
rect 59087 -2528 59153 -2512
rect 59090 -2559 59150 -2528
rect 59090 -2990 59150 -2959
rect 59087 -3006 59153 -2990
rect 59087 -3040 59103 -3006
rect 59137 -3040 59153 -3006
rect 59087 -3056 59153 -3040
rect 59858 -2420 59924 -2412
rect 60368 -2420 60434 -2412
rect 59858 -2428 59946 -2420
rect 59858 -2462 59874 -2428
rect 59908 -2462 59946 -2428
rect 59858 -2470 59946 -2462
rect 60346 -2428 60434 -2420
rect 60346 -2462 60384 -2428
rect 60418 -2462 60434 -2428
rect 60346 -2470 60434 -2462
rect 59858 -2478 59924 -2470
rect 60368 -2478 60434 -2470
rect 59530 -2698 59596 -2682
rect 59530 -2732 59546 -2698
rect 59580 -2732 59596 -2698
rect 59530 -2748 59596 -2732
rect 59548 -2770 59578 -2748
rect 59548 -2992 59578 -2970
rect 59530 -3008 59596 -2992
rect 59530 -3042 59546 -3008
rect 59580 -3042 59596 -3008
rect 59530 -3058 59596 -3042
rect 59846 -2698 59912 -2682
rect 59846 -2732 59862 -2698
rect 59896 -2732 59912 -2698
rect 59846 -2748 59912 -2732
rect 59864 -2770 59894 -2748
rect 59864 -2992 59894 -2970
rect 59846 -3008 59912 -2992
rect 59846 -3042 59862 -3008
rect 59896 -3042 59912 -3008
rect 59846 -3058 59912 -3042
rect 60343 -2965 60409 -2949
rect 61043 -2965 61109 -2949
rect 60343 -2999 60359 -2965
rect 60393 -2999 60409 -2965
rect 60343 -3017 60409 -2999
rect 61043 -2999 61059 -2965
rect 61093 -2999 61109 -2965
rect 61043 -3017 61109 -2999
rect 60165 -3047 60191 -3017
rect 60321 -3047 60441 -3017
rect 60641 -3047 60667 -3017
rect 60785 -3047 60811 -3017
rect 61011 -3047 61131 -3017
rect 61261 -3047 61287 -3017
rect 60343 -3057 60409 -3047
rect 60343 -3091 60359 -3057
rect 60393 -3091 60409 -3057
rect 60343 -3101 60409 -3091
rect 61043 -3057 61109 -3047
rect 61043 -3091 61059 -3057
rect 61093 -3091 61109 -3057
rect 61043 -3101 61109 -3091
rect 57175 -3629 57205 -3603
rect 57263 -3629 57293 -3603
rect 57175 -3748 57205 -3733
rect 57169 -3772 57205 -3748
rect 57169 -3781 57199 -3772
rect 57123 -3797 57199 -3781
rect 57263 -3794 57293 -3733
rect 59087 -3208 59153 -3192
rect 59087 -3242 59103 -3208
rect 59137 -3242 59153 -3208
rect 59087 -3258 59153 -3242
rect 59090 -3289 59150 -3258
rect 59090 -3720 59150 -3689
rect 57123 -3831 57133 -3797
rect 57167 -3831 57199 -3797
rect 57123 -3847 57199 -3831
rect 57169 -3882 57199 -3847
rect 57241 -3810 57295 -3794
rect 57241 -3844 57251 -3810
rect 57285 -3844 57295 -3810
rect 57241 -3860 57295 -3844
rect 59087 -3736 59153 -3720
rect 59087 -3770 59103 -3736
rect 59137 -3770 59153 -3736
rect 59087 -3786 59153 -3770
rect 60165 -3131 60191 -3101
rect 60321 -3131 60441 -3101
rect 60641 -3131 60667 -3101
rect 60785 -3131 60811 -3101
rect 61011 -3131 61131 -3101
rect 61261 -3131 61287 -3101
rect 59526 -3211 59596 -3180
rect 59526 -3230 59545 -3211
rect 59529 -3245 59545 -3230
rect 59579 -3230 59596 -3211
rect 59579 -3245 59595 -3230
rect 59529 -3261 59595 -3245
rect 59547 -3283 59577 -3261
rect 59547 -3505 59577 -3483
rect 59529 -3521 59595 -3505
rect 59529 -3555 59545 -3521
rect 59579 -3555 59595 -3521
rect 59529 -3571 59595 -3555
rect 59845 -3211 59911 -3195
rect 59845 -3245 59861 -3211
rect 59895 -3245 59911 -3211
rect 59845 -3261 59911 -3245
rect 60343 -3141 60409 -3131
rect 60343 -3175 60359 -3141
rect 60393 -3175 60409 -3141
rect 60343 -3185 60409 -3175
rect 61043 -3141 61109 -3131
rect 61043 -3175 61059 -3141
rect 61093 -3175 61109 -3141
rect 61043 -3185 61109 -3175
rect 59863 -3283 59893 -3261
rect 59863 -3505 59893 -3483
rect 59845 -3521 59911 -3505
rect 59845 -3555 59861 -3521
rect 59895 -3555 59911 -3521
rect 59845 -3571 59911 -3555
rect 60165 -3215 60191 -3185
rect 60321 -3215 60441 -3185
rect 60641 -3215 60667 -3185
rect 60785 -3215 60811 -3185
rect 61011 -3215 61131 -3185
rect 61261 -3215 61287 -3185
rect 60343 -3225 60409 -3215
rect 60343 -3259 60359 -3225
rect 60393 -3259 60409 -3225
rect 60343 -3269 60409 -3259
rect 61043 -3225 61109 -3215
rect 61043 -3259 61059 -3225
rect 61093 -3259 61109 -3225
rect 61043 -3269 61109 -3259
rect 60165 -3299 60191 -3269
rect 60321 -3299 60441 -3269
rect 60641 -3299 60667 -3269
rect 60785 -3299 60811 -3269
rect 61011 -3299 61131 -3269
rect 61261 -3299 61287 -3269
rect 57169 -3906 57205 -3882
rect 57175 -3921 57205 -3906
rect 57263 -3921 57293 -3860
rect 57175 -4105 57205 -4079
rect 57263 -4105 57293 -4079
rect 59544 -4000 59610 -3992
rect 59087 -4050 59113 -4000
rect 59513 -4008 59610 -4000
rect 59513 -4042 59560 -4008
rect 59594 -4042 59610 -4008
rect 59513 -4050 59610 -4042
rect 59544 -4058 59610 -4050
rect 59016 -4108 59082 -4100
rect 59016 -4116 59113 -4108
rect 59016 -4150 59032 -4116
rect 59066 -4150 59113 -4116
rect 59016 -4158 59113 -4150
rect 59513 -4158 59539 -4108
rect 59016 -4166 59082 -4158
rect 53972 -4406 54069 -4390
rect 53972 -4444 53988 -4406
rect 54022 -4444 54069 -4406
rect 53972 -4460 54069 -4444
rect 54869 -4406 54966 -4390
rect 54869 -4444 54916 -4406
rect 54950 -4444 54966 -4406
rect 54869 -4460 54966 -4444
rect 59858 -3786 59924 -3778
rect 60368 -3786 60434 -3778
rect 59858 -3794 59946 -3786
rect 59858 -3828 59874 -3794
rect 59908 -3828 59946 -3794
rect 59858 -3836 59946 -3828
rect 60346 -3794 60434 -3786
rect 60346 -3828 60384 -3794
rect 60418 -3828 60434 -3794
rect 60346 -3836 60434 -3828
rect 59858 -3844 59924 -3836
rect 60368 -3844 60434 -3836
rect 55510 -4602 55576 -4586
rect 55510 -4604 55526 -4602
rect 55262 -4634 55288 -4604
rect 55488 -4634 55526 -4604
rect 55510 -4636 55526 -4634
rect 55560 -4636 55576 -4602
rect 55510 -4652 55576 -4636
rect 53982 -7134 54079 -7118
rect 53982 -7172 53998 -7134
rect 54032 -7172 54079 -7134
rect 53982 -7188 54079 -7172
rect 54879 -7134 54976 -7118
rect 54879 -7172 54926 -7134
rect 54960 -7172 54976 -7134
rect 54879 -7188 54976 -7172
rect 20892 -7775 21092 -7759
rect 20892 -7809 20908 -7775
rect 21076 -7809 21092 -7775
rect 20892 -7856 21092 -7809
rect 20892 -11703 21092 -11656
rect 20892 -11737 20908 -11703
rect 21076 -11737 21092 -11703
rect 20892 -11753 21092 -11737
rect 21378 -7775 21578 -7759
rect 21378 -7809 21394 -7775
rect 21562 -7809 21578 -7775
rect 21378 -7856 21578 -7809
rect 21378 -11703 21578 -11656
rect 21378 -11737 21394 -11703
rect 21562 -11737 21578 -11703
rect 21378 -11753 21578 -11737
rect 21864 -7775 22064 -7759
rect 21864 -7809 21880 -7775
rect 22048 -7809 22064 -7775
rect 21864 -7856 22064 -7809
rect 21864 -11703 22064 -11656
rect 21864 -11737 21880 -11703
rect 22048 -11737 22064 -11703
rect 21864 -11753 22064 -11737
rect 53510 -7506 53630 -7490
rect 53510 -7540 53526 -7506
rect 53614 -7540 53630 -7506
rect 53510 -7578 53630 -7540
rect 53982 -7490 54079 -7474
rect 53982 -7528 53998 -7490
rect 54032 -7528 54079 -7490
rect 53982 -7544 54079 -7528
rect 54879 -7490 54976 -7474
rect 54879 -7528 54926 -7490
rect 54960 -7528 54976 -7490
rect 54879 -7544 54976 -7528
rect 55318 -7568 55384 -7552
rect 55318 -7602 55334 -7568
rect 55368 -7602 55384 -7568
rect 55318 -7618 55384 -7602
rect 55336 -7640 55366 -7618
rect 55336 -7866 55366 -7840
rect 53510 -8416 53630 -8378
rect 53510 -8450 53526 -8416
rect 53614 -8450 53630 -8416
rect 53510 -8466 53630 -8450
rect 53842 -8240 53930 -8224
rect 53842 -8328 53858 -8240
rect 53892 -8328 53930 -8240
rect 53842 -8344 53930 -8328
rect 54730 -8240 54818 -8224
rect 54730 -8328 54768 -8240
rect 54802 -8328 54818 -8240
rect 54730 -8344 54818 -8328
rect 55030 -8159 55096 -8144
rect 55540 -8159 55606 -8144
rect 55030 -8160 55118 -8159
rect 55030 -8194 55046 -8160
rect 55080 -8194 55118 -8160
rect 55030 -8195 55118 -8194
rect 55518 -8160 55606 -8159
rect 55518 -8194 55556 -8160
rect 55590 -8194 55606 -8160
rect 55518 -8195 55606 -8194
rect 55030 -8210 55096 -8195
rect 55540 -8210 55606 -8195
rect 55866 -7456 55986 -7440
rect 55866 -7490 55882 -7456
rect 55970 -7490 55986 -7456
rect 55866 -7528 55986 -7490
rect 55866 -8366 55986 -8328
rect 55866 -8400 55882 -8366
rect 55970 -8400 55986 -8366
rect 55866 -8416 55986 -8400
rect 57175 -7509 57205 -7483
rect 57263 -7509 57293 -7483
rect 57175 -7682 57205 -7667
rect 57169 -7706 57205 -7682
rect 57169 -7741 57199 -7706
rect 57263 -7728 57293 -7667
rect 59544 -7493 59610 -7485
rect 59087 -7543 59113 -7493
rect 59513 -7501 59610 -7493
rect 59513 -7535 59560 -7501
rect 59594 -7535 59610 -7501
rect 59513 -7543 59610 -7535
rect 59544 -7551 59610 -7543
rect 59016 -7601 59082 -7593
rect 59016 -7609 59113 -7601
rect 59016 -7643 59032 -7609
rect 59066 -7643 59113 -7609
rect 59016 -7651 59113 -7643
rect 59513 -7651 59539 -7601
rect 59016 -7659 59082 -7651
rect 57123 -7757 57199 -7741
rect 57123 -7791 57133 -7757
rect 57167 -7791 57199 -7757
rect 57123 -7807 57199 -7791
rect 57241 -7744 57295 -7728
rect 57241 -7778 57251 -7744
rect 57285 -7778 57295 -7744
rect 57241 -7794 57295 -7778
rect 57169 -7816 57199 -7807
rect 57169 -7840 57205 -7816
rect 57175 -7855 57205 -7840
rect 57263 -7855 57293 -7794
rect 53510 -8524 53630 -8508
rect 53510 -8558 53526 -8524
rect 53614 -8558 53630 -8524
rect 53510 -8596 53630 -8558
rect 53842 -8646 53930 -8630
rect 53842 -8734 53858 -8646
rect 53892 -8734 53930 -8646
rect 53842 -8750 53930 -8734
rect 54730 -8646 54818 -8630
rect 54730 -8734 54768 -8646
rect 54802 -8734 54818 -8646
rect 54730 -8750 54818 -8734
rect 55030 -8781 55096 -8766
rect 55540 -8781 55606 -8766
rect 55030 -8782 55118 -8781
rect 55030 -8816 55046 -8782
rect 55080 -8816 55118 -8782
rect 55030 -8817 55118 -8816
rect 55518 -8782 55606 -8781
rect 55518 -8816 55556 -8782
rect 55590 -8816 55606 -8782
rect 55518 -8817 55606 -8816
rect 55030 -8832 55096 -8817
rect 53510 -9434 53630 -9396
rect 53510 -9468 53526 -9434
rect 53614 -9468 53630 -9434
rect 53510 -9484 53630 -9468
rect 55540 -8832 55606 -8817
rect 53972 -9450 54069 -9434
rect 53972 -9488 53988 -9450
rect 54022 -9488 54069 -9450
rect 53972 -9504 54069 -9488
rect 54869 -9450 54966 -9434
rect 54869 -9488 54916 -9450
rect 54950 -9488 54966 -9450
rect 54869 -9504 54966 -9488
rect 55326 -9136 55356 -9110
rect 55326 -9358 55356 -9336
rect 55308 -9374 55374 -9358
rect 55308 -9408 55324 -9374
rect 55358 -9408 55374 -9374
rect 55308 -9424 55374 -9408
rect 55866 -8570 55986 -8554
rect 55866 -8604 55882 -8570
rect 55970 -8604 55986 -8570
rect 55866 -8642 55986 -8604
rect 55866 -9480 55986 -9442
rect 55866 -9514 55882 -9480
rect 55970 -9514 55986 -9480
rect 55866 -9530 55986 -9514
rect 56476 -8006 56546 -7990
rect 56476 -8040 56492 -8006
rect 56530 -8040 56546 -8006
rect 56476 -8087 56546 -8040
rect 57175 -7985 57205 -7959
rect 57263 -7985 57293 -7959
rect 56476 -8934 56546 -8887
rect 56476 -8968 56492 -8934
rect 56530 -8968 56546 -8934
rect 56476 -8984 56546 -8968
rect 59087 -7878 59153 -7862
rect 59087 -7912 59103 -7878
rect 59137 -7912 59153 -7878
rect 59087 -7928 59153 -7912
rect 59090 -7959 59150 -7928
rect 59090 -8390 59150 -8359
rect 59087 -8406 59153 -8390
rect 59087 -8440 59103 -8406
rect 59137 -8440 59153 -8406
rect 59087 -8456 59153 -8440
rect 59858 -7820 59924 -7812
rect 60368 -7820 60434 -7812
rect 59858 -7828 59946 -7820
rect 59858 -7862 59874 -7828
rect 59908 -7862 59946 -7828
rect 59858 -7870 59946 -7862
rect 60346 -7828 60434 -7820
rect 60346 -7862 60384 -7828
rect 60418 -7862 60434 -7828
rect 60346 -7870 60434 -7862
rect 59858 -7878 59924 -7870
rect 60368 -7878 60434 -7870
rect 59530 -8098 59596 -8082
rect 59530 -8132 59546 -8098
rect 59580 -8132 59596 -8098
rect 59530 -8148 59596 -8132
rect 59548 -8170 59578 -8148
rect 59548 -8392 59578 -8370
rect 59530 -8408 59596 -8392
rect 59530 -8442 59546 -8408
rect 59580 -8442 59596 -8408
rect 59530 -8458 59596 -8442
rect 59846 -8098 59912 -8082
rect 59846 -8132 59862 -8098
rect 59896 -8132 59912 -8098
rect 59846 -8148 59912 -8132
rect 59864 -8170 59894 -8148
rect 59864 -8392 59894 -8370
rect 59846 -8408 59912 -8392
rect 59846 -8442 59862 -8408
rect 59896 -8442 59912 -8408
rect 59846 -8458 59912 -8442
rect 60343 -8365 60409 -8349
rect 61043 -8365 61109 -8349
rect 60343 -8399 60359 -8365
rect 60393 -8399 60409 -8365
rect 60343 -8417 60409 -8399
rect 61043 -8399 61059 -8365
rect 61093 -8399 61109 -8365
rect 61043 -8417 61109 -8399
rect 60165 -8447 60191 -8417
rect 60321 -8447 60441 -8417
rect 60641 -8447 60667 -8417
rect 60785 -8447 60811 -8417
rect 61011 -8447 61131 -8417
rect 61261 -8447 61287 -8417
rect 60343 -8457 60409 -8447
rect 60343 -8491 60359 -8457
rect 60393 -8491 60409 -8457
rect 60343 -8501 60409 -8491
rect 61043 -8457 61109 -8447
rect 61043 -8491 61059 -8457
rect 61093 -8491 61109 -8457
rect 61043 -8501 61109 -8491
rect 57175 -9029 57205 -9003
rect 57263 -9029 57293 -9003
rect 57175 -9148 57205 -9133
rect 57169 -9172 57205 -9148
rect 57169 -9181 57199 -9172
rect 57123 -9197 57199 -9181
rect 57263 -9194 57293 -9133
rect 59087 -8608 59153 -8592
rect 59087 -8642 59103 -8608
rect 59137 -8642 59153 -8608
rect 59087 -8658 59153 -8642
rect 59090 -8689 59150 -8658
rect 59090 -9120 59150 -9089
rect 57123 -9231 57133 -9197
rect 57167 -9231 57199 -9197
rect 57123 -9247 57199 -9231
rect 57169 -9282 57199 -9247
rect 57241 -9210 57295 -9194
rect 57241 -9244 57251 -9210
rect 57285 -9244 57295 -9210
rect 57241 -9260 57295 -9244
rect 59087 -9136 59153 -9120
rect 59087 -9170 59103 -9136
rect 59137 -9170 59153 -9136
rect 59087 -9186 59153 -9170
rect 60165 -8531 60191 -8501
rect 60321 -8531 60441 -8501
rect 60641 -8531 60667 -8501
rect 60785 -8531 60811 -8501
rect 61011 -8531 61131 -8501
rect 61261 -8531 61287 -8501
rect 59526 -8611 59596 -8580
rect 59526 -8630 59545 -8611
rect 59529 -8645 59545 -8630
rect 59579 -8630 59596 -8611
rect 59579 -8645 59595 -8630
rect 59529 -8661 59595 -8645
rect 59547 -8683 59577 -8661
rect 59547 -8905 59577 -8883
rect 59529 -8921 59595 -8905
rect 59529 -8955 59545 -8921
rect 59579 -8955 59595 -8921
rect 59529 -8971 59595 -8955
rect 59845 -8611 59911 -8595
rect 59845 -8645 59861 -8611
rect 59895 -8645 59911 -8611
rect 59845 -8661 59911 -8645
rect 60343 -8541 60409 -8531
rect 60343 -8575 60359 -8541
rect 60393 -8575 60409 -8541
rect 60343 -8585 60409 -8575
rect 61043 -8541 61109 -8531
rect 61043 -8575 61059 -8541
rect 61093 -8575 61109 -8541
rect 61043 -8585 61109 -8575
rect 59863 -8683 59893 -8661
rect 59863 -8905 59893 -8883
rect 59845 -8921 59911 -8905
rect 59845 -8955 59861 -8921
rect 59895 -8955 59911 -8921
rect 59845 -8971 59911 -8955
rect 60165 -8615 60191 -8585
rect 60321 -8615 60441 -8585
rect 60641 -8615 60667 -8585
rect 60785 -8615 60811 -8585
rect 61011 -8615 61131 -8585
rect 61261 -8615 61287 -8585
rect 60343 -8625 60409 -8615
rect 60343 -8659 60359 -8625
rect 60393 -8659 60409 -8625
rect 60343 -8669 60409 -8659
rect 61043 -8625 61109 -8615
rect 61043 -8659 61059 -8625
rect 61093 -8659 61109 -8625
rect 61043 -8669 61109 -8659
rect 60165 -8699 60191 -8669
rect 60321 -8699 60441 -8669
rect 60641 -8699 60667 -8669
rect 60785 -8699 60811 -8669
rect 61011 -8699 61131 -8669
rect 61261 -8699 61287 -8669
rect 57169 -9306 57205 -9282
rect 57175 -9321 57205 -9306
rect 57263 -9321 57293 -9260
rect 57175 -9505 57205 -9479
rect 57263 -9505 57293 -9479
rect 59544 -9400 59610 -9392
rect 59087 -9450 59113 -9400
rect 59513 -9408 59610 -9400
rect 59513 -9442 59560 -9408
rect 59594 -9442 59610 -9408
rect 59513 -9450 59610 -9442
rect 59544 -9458 59610 -9450
rect 59016 -9508 59082 -9500
rect 59016 -9516 59113 -9508
rect 59016 -9550 59032 -9516
rect 59066 -9550 59113 -9516
rect 59016 -9558 59113 -9550
rect 59513 -9558 59539 -9508
rect 59016 -9566 59082 -9558
rect 53972 -9806 54069 -9790
rect 53972 -9844 53988 -9806
rect 54022 -9844 54069 -9806
rect 53972 -9860 54069 -9844
rect 54869 -9806 54966 -9790
rect 54869 -9844 54916 -9806
rect 54950 -9844 54966 -9806
rect 54869 -9860 54966 -9844
rect 59858 -9186 59924 -9178
rect 60368 -9186 60434 -9178
rect 59858 -9194 59946 -9186
rect 59858 -9228 59874 -9194
rect 59908 -9228 59946 -9194
rect 59858 -9236 59946 -9228
rect 60346 -9194 60434 -9186
rect 60346 -9228 60384 -9194
rect 60418 -9228 60434 -9194
rect 60346 -9236 60434 -9228
rect 59858 -9244 59924 -9236
rect 60368 -9244 60434 -9236
rect 55510 -10002 55576 -9986
rect 55510 -10004 55526 -10002
rect 55262 -10034 55288 -10004
rect 55488 -10034 55526 -10004
rect 55510 -10036 55526 -10034
rect 55560 -10036 55576 -10002
rect 55510 -10052 55576 -10036
rect 20374 -11974 20440 -11958
rect 20374 -11976 20390 -11974
rect 20242 -12006 20268 -11976
rect 20352 -12006 20390 -11976
rect 20374 -12008 20390 -12006
rect 20424 -12008 20440 -11974
rect 20374 -12024 20440 -12008
rect 16599 -12245 16719 -12229
rect 16599 -12279 16615 -12245
rect 16703 -12279 16719 -12245
rect 16599 -12317 16719 -12279
rect 16599 -13155 16719 -13117
rect 16599 -13189 16615 -13155
rect 16703 -13189 16719 -13155
rect 16599 -13205 16719 -13189
rect 17005 -12245 17125 -12229
rect 17005 -12279 17021 -12245
rect 17109 -12279 17125 -12245
rect 17005 -12317 17125 -12279
rect 17005 -13155 17125 -13117
rect 17005 -13189 17021 -13155
rect 17109 -13189 17125 -13155
rect 17005 -13205 17125 -13189
rect 17411 -12245 17531 -12229
rect 17411 -12279 17427 -12245
rect 17515 -12279 17531 -12245
rect 17411 -12317 17531 -12279
rect 17411 -13155 17531 -13117
rect 17411 -13189 17427 -13155
rect 17515 -13189 17531 -13155
rect 17411 -13205 17531 -13189
rect 17817 -12245 17937 -12229
rect 17817 -12279 17833 -12245
rect 17921 -12279 17937 -12245
rect 17817 -12317 17937 -12279
rect 17817 -13155 17937 -13117
rect 17817 -13189 17833 -13155
rect 17921 -13189 17937 -13155
rect 17817 -13205 17937 -13189
rect 18223 -12245 18343 -12229
rect 18223 -12279 18239 -12245
rect 18327 -12279 18343 -12245
rect 18223 -12317 18343 -12279
rect 18223 -13155 18343 -13117
rect 18223 -13189 18239 -13155
rect 18327 -13189 18343 -13155
rect 18223 -13205 18343 -13189
rect 18629 -12245 18749 -12229
rect 18629 -12279 18645 -12245
rect 18733 -12279 18749 -12245
rect 18629 -12317 18749 -12279
rect 18629 -13155 18749 -13117
rect 18629 -13189 18645 -13155
rect 18733 -13189 18749 -13155
rect 18629 -13205 18749 -13189
rect 19035 -12245 19155 -12229
rect 19035 -12279 19051 -12245
rect 19139 -12279 19155 -12245
rect 19035 -12317 19155 -12279
rect 19035 -13155 19155 -13117
rect 19035 -13189 19051 -13155
rect 19139 -13189 19155 -13155
rect 19035 -13205 19155 -13189
rect 19441 -12245 19561 -12229
rect 19441 -12279 19457 -12245
rect 19545 -12279 19561 -12245
rect 19441 -12317 19561 -12279
rect 19441 -13155 19561 -13117
rect 19441 -13189 19457 -13155
rect 19545 -13189 19561 -13155
rect 19441 -13205 19561 -13189
rect 19847 -12245 19967 -12229
rect 19847 -12279 19863 -12245
rect 19951 -12279 19967 -12245
rect 19847 -12317 19967 -12279
rect 19847 -13155 19967 -13117
rect 19847 -13189 19863 -13155
rect 19951 -13189 19967 -13155
rect 19847 -13205 19967 -13189
rect 20253 -12245 20373 -12229
rect 20253 -12279 20269 -12245
rect 20357 -12279 20373 -12245
rect 20253 -12317 20373 -12279
rect 20253 -13155 20373 -13117
rect 20253 -13189 20269 -13155
rect 20357 -13189 20373 -13155
rect 20253 -13205 20373 -13189
rect 20659 -12245 20779 -12229
rect 20659 -12279 20675 -12245
rect 20763 -12279 20779 -12245
rect 20659 -12317 20779 -12279
rect 20659 -13155 20779 -13117
rect 20659 -13189 20675 -13155
rect 20763 -13189 20779 -13155
rect 20659 -13205 20779 -13189
rect 21065 -12245 21185 -12229
rect 21065 -12279 21081 -12245
rect 21169 -12279 21185 -12245
rect 21065 -12317 21185 -12279
rect 21065 -13155 21185 -13117
rect 21065 -13189 21081 -13155
rect 21169 -13189 21185 -13155
rect 21065 -13205 21185 -13189
rect 21471 -12245 21591 -12229
rect 21471 -12279 21487 -12245
rect 21575 -12279 21591 -12245
rect 21471 -12317 21591 -12279
rect 21471 -13155 21591 -13117
rect 21471 -13189 21487 -13155
rect 21575 -13189 21591 -13155
rect 21471 -13205 21591 -13189
rect 21877 -12245 21997 -12229
rect 21877 -12279 21893 -12245
rect 21981 -12279 21997 -12245
rect 21877 -12317 21997 -12279
rect 21877 -13155 21997 -13117
rect 21877 -13189 21893 -13155
rect 21981 -13189 21997 -13155
rect 21877 -13205 21997 -13189
rect 22283 -12245 22403 -12229
rect 22283 -12279 22299 -12245
rect 22387 -12279 22403 -12245
rect 22283 -12317 22403 -12279
rect 22283 -13155 22403 -13117
rect 22283 -13189 22299 -13155
rect 22387 -13189 22403 -13155
rect 22283 -13205 22403 -13189
rect 22689 -12245 22809 -12229
rect 22689 -12279 22705 -12245
rect 22793 -12279 22809 -12245
rect 22689 -12317 22809 -12279
rect 22689 -13155 22809 -13117
rect 22689 -13189 22705 -13155
rect 22793 -13189 22809 -13155
rect 22689 -13205 22809 -13189
rect 23095 -12245 23215 -12229
rect 23095 -12279 23111 -12245
rect 23199 -12279 23215 -12245
rect 23095 -12317 23215 -12279
rect 23095 -13155 23215 -13117
rect 23095 -13189 23111 -13155
rect 23199 -13189 23215 -13155
rect 23095 -13205 23215 -13189
rect 23501 -12245 23621 -12229
rect 23501 -12279 23517 -12245
rect 23605 -12279 23621 -12245
rect 23501 -12317 23621 -12279
rect 23501 -13155 23621 -13117
rect 23501 -13189 23517 -13155
rect 23605 -13189 23621 -13155
rect 23501 -13205 23621 -13189
rect 23907 -12245 24027 -12229
rect 23907 -12279 23923 -12245
rect 24011 -12279 24027 -12245
rect 23907 -12317 24027 -12279
rect 23907 -13155 24027 -13117
rect 23907 -13189 23923 -13155
rect 24011 -13189 24027 -13155
rect 23907 -13205 24027 -13189
rect 24313 -12245 24433 -12229
rect 24313 -12279 24329 -12245
rect 24417 -12279 24433 -12245
rect 24313 -12317 24433 -12279
rect 24313 -13155 24433 -13117
rect 24313 -13189 24329 -13155
rect 24417 -13189 24433 -13155
rect 24313 -13205 24433 -13189
rect 24719 -12245 24839 -12229
rect 24719 -12279 24735 -12245
rect 24823 -12279 24839 -12245
rect 24719 -12317 24839 -12279
rect 24719 -13155 24839 -13117
rect 24719 -13189 24735 -13155
rect 24823 -13189 24839 -13155
rect 24719 -13205 24839 -13189
rect 25125 -12245 25245 -12229
rect 25125 -12279 25141 -12245
rect 25229 -12279 25245 -12245
rect 25125 -12317 25245 -12279
rect 25125 -13155 25245 -13117
rect 25125 -13189 25141 -13155
rect 25229 -13189 25245 -13155
rect 25125 -13205 25245 -13189
rect 53982 -12534 54079 -12518
rect 53982 -12572 53998 -12534
rect 54032 -12572 54079 -12534
rect 53982 -12588 54079 -12572
rect 54879 -12534 54976 -12518
rect 54879 -12572 54926 -12534
rect 54960 -12572 54976 -12534
rect 54879 -12588 54976 -12572
rect 53510 -12906 53630 -12890
rect 53510 -12940 53526 -12906
rect 53614 -12940 53630 -12906
rect 53510 -12978 53630 -12940
rect 53982 -12890 54079 -12874
rect 53982 -12928 53998 -12890
rect 54032 -12928 54079 -12890
rect 53982 -12944 54079 -12928
rect 54879 -12890 54976 -12874
rect 54879 -12928 54926 -12890
rect 54960 -12928 54976 -12890
rect 54879 -12944 54976 -12928
rect 55318 -12968 55384 -12952
rect 55318 -13002 55334 -12968
rect 55368 -13002 55384 -12968
rect 55318 -13018 55384 -13002
rect 55336 -13040 55366 -13018
rect 55336 -13266 55366 -13240
rect 53510 -13816 53630 -13778
rect 53510 -13850 53526 -13816
rect 53614 -13850 53630 -13816
rect 53510 -13866 53630 -13850
rect 53842 -13640 53930 -13624
rect 53842 -13728 53858 -13640
rect 53892 -13728 53930 -13640
rect 53842 -13744 53930 -13728
rect 54730 -13640 54818 -13624
rect 54730 -13728 54768 -13640
rect 54802 -13728 54818 -13640
rect 54730 -13744 54818 -13728
rect 55030 -13559 55096 -13544
rect 55540 -13559 55606 -13544
rect 55030 -13560 55118 -13559
rect 55030 -13594 55046 -13560
rect 55080 -13594 55118 -13560
rect 55030 -13595 55118 -13594
rect 55518 -13560 55606 -13559
rect 55518 -13594 55556 -13560
rect 55590 -13594 55606 -13560
rect 55518 -13595 55606 -13594
rect 55030 -13610 55096 -13595
rect 55540 -13610 55606 -13595
rect 55866 -12856 55986 -12840
rect 55866 -12890 55882 -12856
rect 55970 -12890 55986 -12856
rect 55866 -12928 55986 -12890
rect 55866 -13766 55986 -13728
rect 55866 -13800 55882 -13766
rect 55970 -13800 55986 -13766
rect 55866 -13816 55986 -13800
rect 57175 -12909 57205 -12883
rect 57263 -12909 57293 -12883
rect 57175 -13082 57205 -13067
rect 57169 -13106 57205 -13082
rect 57169 -13141 57199 -13106
rect 57263 -13128 57293 -13067
rect 59544 -12893 59610 -12885
rect 59087 -12943 59113 -12893
rect 59513 -12901 59610 -12893
rect 59513 -12935 59560 -12901
rect 59594 -12935 59610 -12901
rect 59513 -12943 59610 -12935
rect 59544 -12951 59610 -12943
rect 59016 -13001 59082 -12993
rect 59016 -13009 59113 -13001
rect 59016 -13043 59032 -13009
rect 59066 -13043 59113 -13009
rect 59016 -13051 59113 -13043
rect 59513 -13051 59539 -13001
rect 59016 -13059 59082 -13051
rect 57123 -13157 57199 -13141
rect 57123 -13191 57133 -13157
rect 57167 -13191 57199 -13157
rect 57123 -13207 57199 -13191
rect 57241 -13144 57295 -13128
rect 57241 -13178 57251 -13144
rect 57285 -13178 57295 -13144
rect 57241 -13194 57295 -13178
rect 57169 -13216 57199 -13207
rect 57169 -13240 57205 -13216
rect 57175 -13255 57205 -13240
rect 57263 -13255 57293 -13194
rect 53510 -13924 53630 -13908
rect 53510 -13958 53526 -13924
rect 53614 -13958 53630 -13924
rect 53510 -13996 53630 -13958
rect 53842 -14046 53930 -14030
rect 53842 -14134 53858 -14046
rect 53892 -14134 53930 -14046
rect 53842 -14150 53930 -14134
rect 54730 -14046 54818 -14030
rect 54730 -14134 54768 -14046
rect 54802 -14134 54818 -14046
rect 54730 -14150 54818 -14134
rect 55030 -14181 55096 -14166
rect 55540 -14181 55606 -14166
rect 55030 -14182 55118 -14181
rect 55030 -14216 55046 -14182
rect 55080 -14216 55118 -14182
rect 55030 -14217 55118 -14216
rect 55518 -14182 55606 -14181
rect 55518 -14216 55556 -14182
rect 55590 -14216 55606 -14182
rect 55518 -14217 55606 -14216
rect 55030 -14232 55096 -14217
rect 53510 -14834 53630 -14796
rect 53510 -14868 53526 -14834
rect 53614 -14868 53630 -14834
rect 53510 -14884 53630 -14868
rect 55540 -14232 55606 -14217
rect 53972 -14850 54069 -14834
rect 53972 -14888 53988 -14850
rect 54022 -14888 54069 -14850
rect 53972 -14904 54069 -14888
rect 54869 -14850 54966 -14834
rect 54869 -14888 54916 -14850
rect 54950 -14888 54966 -14850
rect 54869 -14904 54966 -14888
rect 55326 -14536 55356 -14510
rect 55326 -14758 55356 -14736
rect 55308 -14774 55374 -14758
rect 55308 -14808 55324 -14774
rect 55358 -14808 55374 -14774
rect 55308 -14824 55374 -14808
rect 55866 -13970 55986 -13954
rect 55866 -14004 55882 -13970
rect 55970 -14004 55986 -13970
rect 55866 -14042 55986 -14004
rect 55866 -14880 55986 -14842
rect 55866 -14914 55882 -14880
rect 55970 -14914 55986 -14880
rect 55866 -14930 55986 -14914
rect 56476 -13406 56546 -13390
rect 56476 -13440 56492 -13406
rect 56530 -13440 56546 -13406
rect 56476 -13487 56546 -13440
rect 57175 -13385 57205 -13359
rect 57263 -13385 57293 -13359
rect 56476 -14334 56546 -14287
rect 56476 -14368 56492 -14334
rect 56530 -14368 56546 -14334
rect 56476 -14384 56546 -14368
rect 59087 -13278 59153 -13262
rect 59087 -13312 59103 -13278
rect 59137 -13312 59153 -13278
rect 59087 -13328 59153 -13312
rect 59090 -13359 59150 -13328
rect 59090 -13790 59150 -13759
rect 59087 -13806 59153 -13790
rect 59087 -13840 59103 -13806
rect 59137 -13840 59153 -13806
rect 59087 -13856 59153 -13840
rect 59858 -13220 59924 -13212
rect 60368 -13220 60434 -13212
rect 59858 -13228 59946 -13220
rect 59858 -13262 59874 -13228
rect 59908 -13262 59946 -13228
rect 59858 -13270 59946 -13262
rect 60346 -13228 60434 -13220
rect 60346 -13262 60384 -13228
rect 60418 -13262 60434 -13228
rect 60346 -13270 60434 -13262
rect 59858 -13278 59924 -13270
rect 60368 -13278 60434 -13270
rect 59530 -13498 59596 -13482
rect 59530 -13532 59546 -13498
rect 59580 -13532 59596 -13498
rect 59530 -13548 59596 -13532
rect 59548 -13570 59578 -13548
rect 59548 -13792 59578 -13770
rect 59530 -13808 59596 -13792
rect 59530 -13842 59546 -13808
rect 59580 -13842 59596 -13808
rect 59530 -13858 59596 -13842
rect 59846 -13498 59912 -13482
rect 59846 -13532 59862 -13498
rect 59896 -13532 59912 -13498
rect 59846 -13548 59912 -13532
rect 59864 -13570 59894 -13548
rect 59864 -13792 59894 -13770
rect 59846 -13808 59912 -13792
rect 59846 -13842 59862 -13808
rect 59896 -13842 59912 -13808
rect 59846 -13858 59912 -13842
rect 60343 -13765 60409 -13749
rect 61043 -13765 61109 -13749
rect 60343 -13799 60359 -13765
rect 60393 -13799 60409 -13765
rect 60343 -13817 60409 -13799
rect 61043 -13799 61059 -13765
rect 61093 -13799 61109 -13765
rect 61043 -13817 61109 -13799
rect 60165 -13847 60191 -13817
rect 60321 -13847 60441 -13817
rect 60641 -13847 60667 -13817
rect 60785 -13847 60811 -13817
rect 61011 -13847 61131 -13817
rect 61261 -13847 61287 -13817
rect 60343 -13857 60409 -13847
rect 60343 -13891 60359 -13857
rect 60393 -13891 60409 -13857
rect 60343 -13901 60409 -13891
rect 61043 -13857 61109 -13847
rect 61043 -13891 61059 -13857
rect 61093 -13891 61109 -13857
rect 61043 -13901 61109 -13891
rect 57175 -14429 57205 -14403
rect 57263 -14429 57293 -14403
rect 57175 -14548 57205 -14533
rect 57169 -14572 57205 -14548
rect 57169 -14581 57199 -14572
rect 57123 -14597 57199 -14581
rect 57263 -14594 57293 -14533
rect 59087 -14008 59153 -13992
rect 59087 -14042 59103 -14008
rect 59137 -14042 59153 -14008
rect 59087 -14058 59153 -14042
rect 59090 -14089 59150 -14058
rect 59090 -14520 59150 -14489
rect 57123 -14631 57133 -14597
rect 57167 -14631 57199 -14597
rect 57123 -14647 57199 -14631
rect 57169 -14682 57199 -14647
rect 57241 -14610 57295 -14594
rect 57241 -14644 57251 -14610
rect 57285 -14644 57295 -14610
rect 57241 -14660 57295 -14644
rect 59087 -14536 59153 -14520
rect 59087 -14570 59103 -14536
rect 59137 -14570 59153 -14536
rect 59087 -14586 59153 -14570
rect 60165 -13931 60191 -13901
rect 60321 -13931 60441 -13901
rect 60641 -13931 60667 -13901
rect 60785 -13931 60811 -13901
rect 61011 -13931 61131 -13901
rect 61261 -13931 61287 -13901
rect 59526 -14011 59596 -13980
rect 59526 -14030 59545 -14011
rect 59529 -14045 59545 -14030
rect 59579 -14030 59596 -14011
rect 59579 -14045 59595 -14030
rect 59529 -14061 59595 -14045
rect 59547 -14083 59577 -14061
rect 59547 -14305 59577 -14283
rect 59529 -14321 59595 -14305
rect 59529 -14355 59545 -14321
rect 59579 -14355 59595 -14321
rect 59529 -14371 59595 -14355
rect 59845 -14011 59911 -13995
rect 59845 -14045 59861 -14011
rect 59895 -14045 59911 -14011
rect 59845 -14061 59911 -14045
rect 60343 -13941 60409 -13931
rect 60343 -13975 60359 -13941
rect 60393 -13975 60409 -13941
rect 60343 -13985 60409 -13975
rect 61043 -13941 61109 -13931
rect 61043 -13975 61059 -13941
rect 61093 -13975 61109 -13941
rect 61043 -13985 61109 -13975
rect 59863 -14083 59893 -14061
rect 59863 -14305 59893 -14283
rect 59845 -14321 59911 -14305
rect 59845 -14355 59861 -14321
rect 59895 -14355 59911 -14321
rect 59845 -14371 59911 -14355
rect 60165 -14015 60191 -13985
rect 60321 -14015 60441 -13985
rect 60641 -14015 60667 -13985
rect 60785 -14015 60811 -13985
rect 61011 -14015 61131 -13985
rect 61261 -14015 61287 -13985
rect 60343 -14025 60409 -14015
rect 60343 -14059 60359 -14025
rect 60393 -14059 60409 -14025
rect 60343 -14069 60409 -14059
rect 61043 -14025 61109 -14015
rect 61043 -14059 61059 -14025
rect 61093 -14059 61109 -14025
rect 61043 -14069 61109 -14059
rect 60165 -14099 60191 -14069
rect 60321 -14099 60441 -14069
rect 60641 -14099 60667 -14069
rect 60785 -14099 60811 -14069
rect 61011 -14099 61131 -14069
rect 61261 -14099 61287 -14069
rect 57169 -14706 57205 -14682
rect 57175 -14721 57205 -14706
rect 57263 -14721 57293 -14660
rect 57175 -14905 57205 -14879
rect 57263 -14905 57293 -14879
rect 59544 -14800 59610 -14792
rect 59087 -14850 59113 -14800
rect 59513 -14808 59610 -14800
rect 59513 -14842 59560 -14808
rect 59594 -14842 59610 -14808
rect 59513 -14850 59610 -14842
rect 59544 -14858 59610 -14850
rect 59016 -14908 59082 -14900
rect 59016 -14916 59113 -14908
rect 59016 -14950 59032 -14916
rect 59066 -14950 59113 -14916
rect 59016 -14958 59113 -14950
rect 59513 -14958 59539 -14908
rect 59016 -14966 59082 -14958
rect 53972 -15206 54069 -15190
rect 53972 -15244 53988 -15206
rect 54022 -15244 54069 -15206
rect 53972 -15260 54069 -15244
rect 54869 -15206 54966 -15190
rect 54869 -15244 54916 -15206
rect 54950 -15244 54966 -15206
rect 54869 -15260 54966 -15244
rect 59858 -14586 59924 -14578
rect 60368 -14586 60434 -14578
rect 59858 -14594 59946 -14586
rect 59858 -14628 59874 -14594
rect 59908 -14628 59946 -14594
rect 59858 -14636 59946 -14628
rect 60346 -14594 60434 -14586
rect 60346 -14628 60384 -14594
rect 60418 -14628 60434 -14594
rect 60346 -14636 60434 -14628
rect 59858 -14644 59924 -14636
rect 60368 -14644 60434 -14636
rect 55510 -15402 55576 -15386
rect 55510 -15404 55526 -15402
rect 55262 -15434 55288 -15404
rect 55488 -15434 55526 -15404
rect 55510 -15436 55526 -15434
rect 55560 -15436 55576 -15402
rect 55510 -15452 55576 -15436
rect 53982 -17934 54079 -17918
rect 53982 -17972 53998 -17934
rect 54032 -17972 54079 -17934
rect 53982 -17988 54079 -17972
rect 54879 -17934 54976 -17918
rect 54879 -17972 54926 -17934
rect 54960 -17972 54976 -17934
rect 54879 -17988 54976 -17972
rect 53510 -18306 53630 -18290
rect 53510 -18340 53526 -18306
rect 53614 -18340 53630 -18306
rect 53510 -18378 53630 -18340
rect 53982 -18290 54079 -18274
rect 53982 -18328 53998 -18290
rect 54032 -18328 54079 -18290
rect 53982 -18344 54079 -18328
rect 54879 -18290 54976 -18274
rect 54879 -18328 54926 -18290
rect 54960 -18328 54976 -18290
rect 54879 -18344 54976 -18328
rect 55318 -18368 55384 -18352
rect 55318 -18402 55334 -18368
rect 55368 -18402 55384 -18368
rect 55318 -18418 55384 -18402
rect 55336 -18440 55366 -18418
rect 55336 -18666 55366 -18640
rect 53510 -19216 53630 -19178
rect 53510 -19250 53526 -19216
rect 53614 -19250 53630 -19216
rect 53510 -19266 53630 -19250
rect 53842 -19040 53930 -19024
rect 53842 -19128 53858 -19040
rect 53892 -19128 53930 -19040
rect 53842 -19144 53930 -19128
rect 54730 -19040 54818 -19024
rect 54730 -19128 54768 -19040
rect 54802 -19128 54818 -19040
rect 54730 -19144 54818 -19128
rect 55030 -18959 55096 -18944
rect 55540 -18959 55606 -18944
rect 55030 -18960 55118 -18959
rect 55030 -18994 55046 -18960
rect 55080 -18994 55118 -18960
rect 55030 -18995 55118 -18994
rect 55518 -18960 55606 -18959
rect 55518 -18994 55556 -18960
rect 55590 -18994 55606 -18960
rect 55518 -18995 55606 -18994
rect 55030 -19010 55096 -18995
rect 55540 -19010 55606 -18995
rect 55866 -18256 55986 -18240
rect 55866 -18290 55882 -18256
rect 55970 -18290 55986 -18256
rect 55866 -18328 55986 -18290
rect 55866 -19166 55986 -19128
rect 55866 -19200 55882 -19166
rect 55970 -19200 55986 -19166
rect 55866 -19216 55986 -19200
rect 57175 -18309 57205 -18283
rect 57263 -18309 57293 -18283
rect 57175 -18482 57205 -18467
rect 57169 -18506 57205 -18482
rect 57169 -18541 57199 -18506
rect 57263 -18528 57293 -18467
rect 59544 -18293 59610 -18285
rect 59087 -18343 59113 -18293
rect 59513 -18301 59610 -18293
rect 59513 -18335 59560 -18301
rect 59594 -18335 59610 -18301
rect 59513 -18343 59610 -18335
rect 59544 -18351 59610 -18343
rect 59016 -18401 59082 -18393
rect 59016 -18409 59113 -18401
rect 59016 -18443 59032 -18409
rect 59066 -18443 59113 -18409
rect 59016 -18451 59113 -18443
rect 59513 -18451 59539 -18401
rect 59016 -18459 59082 -18451
rect 57123 -18557 57199 -18541
rect 57123 -18591 57133 -18557
rect 57167 -18591 57199 -18557
rect 57123 -18607 57199 -18591
rect 57241 -18544 57295 -18528
rect 57241 -18578 57251 -18544
rect 57285 -18578 57295 -18544
rect 57241 -18594 57295 -18578
rect 57169 -18616 57199 -18607
rect 57169 -18640 57205 -18616
rect 57175 -18655 57205 -18640
rect 57263 -18655 57293 -18594
rect 53510 -19324 53630 -19308
rect 53510 -19358 53526 -19324
rect 53614 -19358 53630 -19324
rect 53510 -19396 53630 -19358
rect 53842 -19446 53930 -19430
rect 53842 -19534 53858 -19446
rect 53892 -19534 53930 -19446
rect 53842 -19550 53930 -19534
rect 54730 -19446 54818 -19430
rect 54730 -19534 54768 -19446
rect 54802 -19534 54818 -19446
rect 54730 -19550 54818 -19534
rect 55030 -19581 55096 -19566
rect 55540 -19581 55606 -19566
rect 55030 -19582 55118 -19581
rect 55030 -19616 55046 -19582
rect 55080 -19616 55118 -19582
rect 55030 -19617 55118 -19616
rect 55518 -19582 55606 -19581
rect 55518 -19616 55556 -19582
rect 55590 -19616 55606 -19582
rect 55518 -19617 55606 -19616
rect 55030 -19632 55096 -19617
rect 53510 -20234 53630 -20196
rect 53510 -20268 53526 -20234
rect 53614 -20268 53630 -20234
rect 53510 -20284 53630 -20268
rect 55540 -19632 55606 -19617
rect 53972 -20250 54069 -20234
rect 53972 -20288 53988 -20250
rect 54022 -20288 54069 -20250
rect 53972 -20304 54069 -20288
rect 54869 -20250 54966 -20234
rect 54869 -20288 54916 -20250
rect 54950 -20288 54966 -20250
rect 54869 -20304 54966 -20288
rect 55326 -19936 55356 -19910
rect 55326 -20158 55356 -20136
rect 55308 -20174 55374 -20158
rect 55308 -20208 55324 -20174
rect 55358 -20208 55374 -20174
rect 55308 -20224 55374 -20208
rect 55866 -19370 55986 -19354
rect 55866 -19404 55882 -19370
rect 55970 -19404 55986 -19370
rect 55866 -19442 55986 -19404
rect 55866 -20280 55986 -20242
rect 55866 -20314 55882 -20280
rect 55970 -20314 55986 -20280
rect 55866 -20330 55986 -20314
rect 56476 -18806 56546 -18790
rect 56476 -18840 56492 -18806
rect 56530 -18840 56546 -18806
rect 56476 -18887 56546 -18840
rect 57175 -18785 57205 -18759
rect 57263 -18785 57293 -18759
rect 56476 -19734 56546 -19687
rect 56476 -19768 56492 -19734
rect 56530 -19768 56546 -19734
rect 56476 -19784 56546 -19768
rect 59087 -18678 59153 -18662
rect 59087 -18712 59103 -18678
rect 59137 -18712 59153 -18678
rect 59087 -18728 59153 -18712
rect 59090 -18759 59150 -18728
rect 59090 -19190 59150 -19159
rect 59087 -19206 59153 -19190
rect 59087 -19240 59103 -19206
rect 59137 -19240 59153 -19206
rect 59087 -19256 59153 -19240
rect 59858 -18620 59924 -18612
rect 60368 -18620 60434 -18612
rect 59858 -18628 59946 -18620
rect 59858 -18662 59874 -18628
rect 59908 -18662 59946 -18628
rect 59858 -18670 59946 -18662
rect 60346 -18628 60434 -18620
rect 60346 -18662 60384 -18628
rect 60418 -18662 60434 -18628
rect 60346 -18670 60434 -18662
rect 59858 -18678 59924 -18670
rect 60368 -18678 60434 -18670
rect 59530 -18898 59596 -18882
rect 59530 -18932 59546 -18898
rect 59580 -18932 59596 -18898
rect 59530 -18948 59596 -18932
rect 59548 -18970 59578 -18948
rect 59548 -19192 59578 -19170
rect 59530 -19208 59596 -19192
rect 59530 -19242 59546 -19208
rect 59580 -19242 59596 -19208
rect 59530 -19258 59596 -19242
rect 59846 -18898 59912 -18882
rect 59846 -18932 59862 -18898
rect 59896 -18932 59912 -18898
rect 59846 -18948 59912 -18932
rect 59864 -18970 59894 -18948
rect 59864 -19192 59894 -19170
rect 59846 -19208 59912 -19192
rect 59846 -19242 59862 -19208
rect 59896 -19242 59912 -19208
rect 59846 -19258 59912 -19242
rect 60343 -19165 60409 -19149
rect 61043 -19165 61109 -19149
rect 60343 -19199 60359 -19165
rect 60393 -19199 60409 -19165
rect 60343 -19217 60409 -19199
rect 61043 -19199 61059 -19165
rect 61093 -19199 61109 -19165
rect 61043 -19217 61109 -19199
rect 60165 -19247 60191 -19217
rect 60321 -19247 60441 -19217
rect 60641 -19247 60667 -19217
rect 60785 -19247 60811 -19217
rect 61011 -19247 61131 -19217
rect 61261 -19247 61287 -19217
rect 60343 -19257 60409 -19247
rect 60343 -19291 60359 -19257
rect 60393 -19291 60409 -19257
rect 60343 -19301 60409 -19291
rect 61043 -19257 61109 -19247
rect 61043 -19291 61059 -19257
rect 61093 -19291 61109 -19257
rect 61043 -19301 61109 -19291
rect 57175 -19829 57205 -19803
rect 57263 -19829 57293 -19803
rect 57175 -19948 57205 -19933
rect 57169 -19972 57205 -19948
rect 57169 -19981 57199 -19972
rect 57123 -19997 57199 -19981
rect 57263 -19994 57293 -19933
rect 59087 -19408 59153 -19392
rect 59087 -19442 59103 -19408
rect 59137 -19442 59153 -19408
rect 59087 -19458 59153 -19442
rect 59090 -19489 59150 -19458
rect 59090 -19920 59150 -19889
rect 57123 -20031 57133 -19997
rect 57167 -20031 57199 -19997
rect 57123 -20047 57199 -20031
rect 57169 -20082 57199 -20047
rect 57241 -20010 57295 -19994
rect 57241 -20044 57251 -20010
rect 57285 -20044 57295 -20010
rect 57241 -20060 57295 -20044
rect 59087 -19936 59153 -19920
rect 59087 -19970 59103 -19936
rect 59137 -19970 59153 -19936
rect 59087 -19986 59153 -19970
rect 60165 -19331 60191 -19301
rect 60321 -19331 60441 -19301
rect 60641 -19331 60667 -19301
rect 60785 -19331 60811 -19301
rect 61011 -19331 61131 -19301
rect 61261 -19331 61287 -19301
rect 59526 -19411 59596 -19380
rect 59526 -19430 59545 -19411
rect 59529 -19445 59545 -19430
rect 59579 -19430 59596 -19411
rect 59579 -19445 59595 -19430
rect 59529 -19461 59595 -19445
rect 59547 -19483 59577 -19461
rect 59547 -19705 59577 -19683
rect 59529 -19721 59595 -19705
rect 59529 -19755 59545 -19721
rect 59579 -19755 59595 -19721
rect 59529 -19771 59595 -19755
rect 59845 -19411 59911 -19395
rect 59845 -19445 59861 -19411
rect 59895 -19445 59911 -19411
rect 59845 -19461 59911 -19445
rect 60343 -19341 60409 -19331
rect 60343 -19375 60359 -19341
rect 60393 -19375 60409 -19341
rect 60343 -19385 60409 -19375
rect 61043 -19341 61109 -19331
rect 61043 -19375 61059 -19341
rect 61093 -19375 61109 -19341
rect 61043 -19385 61109 -19375
rect 59863 -19483 59893 -19461
rect 59863 -19705 59893 -19683
rect 59845 -19721 59911 -19705
rect 59845 -19755 59861 -19721
rect 59895 -19755 59911 -19721
rect 59845 -19771 59911 -19755
rect 60165 -19415 60191 -19385
rect 60321 -19415 60441 -19385
rect 60641 -19415 60667 -19385
rect 60785 -19415 60811 -19385
rect 61011 -19415 61131 -19385
rect 61261 -19415 61287 -19385
rect 60343 -19425 60409 -19415
rect 60343 -19459 60359 -19425
rect 60393 -19459 60409 -19425
rect 60343 -19469 60409 -19459
rect 61043 -19425 61109 -19415
rect 61043 -19459 61059 -19425
rect 61093 -19459 61109 -19425
rect 61043 -19469 61109 -19459
rect 60165 -19499 60191 -19469
rect 60321 -19499 60441 -19469
rect 60641 -19499 60667 -19469
rect 60785 -19499 60811 -19469
rect 61011 -19499 61131 -19469
rect 61261 -19499 61287 -19469
rect 57169 -20106 57205 -20082
rect 57175 -20121 57205 -20106
rect 57263 -20121 57293 -20060
rect 57175 -20305 57205 -20279
rect 57263 -20305 57293 -20279
rect 59544 -20200 59610 -20192
rect 59087 -20250 59113 -20200
rect 59513 -20208 59610 -20200
rect 59513 -20242 59560 -20208
rect 59594 -20242 59610 -20208
rect 59513 -20250 59610 -20242
rect 59544 -20258 59610 -20250
rect 59016 -20308 59082 -20300
rect 59016 -20316 59113 -20308
rect 59016 -20350 59032 -20316
rect 59066 -20350 59113 -20316
rect 59016 -20358 59113 -20350
rect 59513 -20358 59539 -20308
rect 59016 -20366 59082 -20358
rect 53972 -20606 54069 -20590
rect 53972 -20644 53988 -20606
rect 54022 -20644 54069 -20606
rect 53972 -20660 54069 -20644
rect 54869 -20606 54966 -20590
rect 54869 -20644 54916 -20606
rect 54950 -20644 54966 -20606
rect 54869 -20660 54966 -20644
rect 59858 -19986 59924 -19978
rect 60368 -19986 60434 -19978
rect 59858 -19994 59946 -19986
rect 59858 -20028 59874 -19994
rect 59908 -20028 59946 -19994
rect 59858 -20036 59946 -20028
rect 60346 -19994 60434 -19986
rect 60346 -20028 60384 -19994
rect 60418 -20028 60434 -19994
rect 60346 -20036 60434 -20028
rect 59858 -20044 59924 -20036
rect 60368 -20044 60434 -20036
rect 55510 -20802 55576 -20786
rect 55510 -20804 55526 -20802
rect 55262 -20834 55288 -20804
rect 55488 -20834 55526 -20804
rect 55510 -20836 55526 -20834
rect 55560 -20836 55576 -20802
rect 55510 -20852 55576 -20836
rect 53982 -23334 54079 -23318
rect 53982 -23372 53998 -23334
rect 54032 -23372 54079 -23334
rect 53982 -23388 54079 -23372
rect 54879 -23334 54976 -23318
rect 54879 -23372 54926 -23334
rect 54960 -23372 54976 -23334
rect 54879 -23388 54976 -23372
rect 53510 -23706 53630 -23690
rect 53510 -23740 53526 -23706
rect 53614 -23740 53630 -23706
rect 53510 -23778 53630 -23740
rect 53982 -23690 54079 -23674
rect 53982 -23728 53998 -23690
rect 54032 -23728 54079 -23690
rect 53982 -23744 54079 -23728
rect 54879 -23690 54976 -23674
rect 54879 -23728 54926 -23690
rect 54960 -23728 54976 -23690
rect 54879 -23744 54976 -23728
rect 55318 -23768 55384 -23752
rect 55318 -23802 55334 -23768
rect 55368 -23802 55384 -23768
rect 55318 -23818 55384 -23802
rect 55336 -23840 55366 -23818
rect 55336 -24066 55366 -24040
rect 53510 -24616 53630 -24578
rect 53510 -24650 53526 -24616
rect 53614 -24650 53630 -24616
rect 53510 -24666 53630 -24650
rect 53842 -24440 53930 -24424
rect 53842 -24528 53858 -24440
rect 53892 -24528 53930 -24440
rect 53842 -24544 53930 -24528
rect 54730 -24440 54818 -24424
rect 54730 -24528 54768 -24440
rect 54802 -24528 54818 -24440
rect 54730 -24544 54818 -24528
rect 55030 -24359 55096 -24344
rect 55540 -24359 55606 -24344
rect 55030 -24360 55118 -24359
rect 55030 -24394 55046 -24360
rect 55080 -24394 55118 -24360
rect 55030 -24395 55118 -24394
rect 55518 -24360 55606 -24359
rect 55518 -24394 55556 -24360
rect 55590 -24394 55606 -24360
rect 55518 -24395 55606 -24394
rect 55030 -24410 55096 -24395
rect 55540 -24410 55606 -24395
rect 55866 -23656 55986 -23640
rect 55866 -23690 55882 -23656
rect 55970 -23690 55986 -23656
rect 55866 -23728 55986 -23690
rect 55866 -24566 55986 -24528
rect 55866 -24600 55882 -24566
rect 55970 -24600 55986 -24566
rect 55866 -24616 55986 -24600
rect 57175 -23709 57205 -23683
rect 57263 -23709 57293 -23683
rect 57175 -23882 57205 -23867
rect 57169 -23906 57205 -23882
rect 57169 -23941 57199 -23906
rect 57263 -23928 57293 -23867
rect 59544 -23693 59610 -23685
rect 59087 -23743 59113 -23693
rect 59513 -23701 59610 -23693
rect 59513 -23735 59560 -23701
rect 59594 -23735 59610 -23701
rect 59513 -23743 59610 -23735
rect 59544 -23751 59610 -23743
rect 59016 -23801 59082 -23793
rect 59016 -23809 59113 -23801
rect 59016 -23843 59032 -23809
rect 59066 -23843 59113 -23809
rect 59016 -23851 59113 -23843
rect 59513 -23851 59539 -23801
rect 59016 -23859 59082 -23851
rect 57123 -23957 57199 -23941
rect 57123 -23991 57133 -23957
rect 57167 -23991 57199 -23957
rect 57123 -24007 57199 -23991
rect 57241 -23944 57295 -23928
rect 57241 -23978 57251 -23944
rect 57285 -23978 57295 -23944
rect 57241 -23994 57295 -23978
rect 57169 -24016 57199 -24007
rect 57169 -24040 57205 -24016
rect 57175 -24055 57205 -24040
rect 57263 -24055 57293 -23994
rect 53510 -24724 53630 -24708
rect 53510 -24758 53526 -24724
rect 53614 -24758 53630 -24724
rect 53510 -24796 53630 -24758
rect 53842 -24846 53930 -24830
rect 53842 -24934 53858 -24846
rect 53892 -24934 53930 -24846
rect 53842 -24950 53930 -24934
rect 54730 -24846 54818 -24830
rect 54730 -24934 54768 -24846
rect 54802 -24934 54818 -24846
rect 54730 -24950 54818 -24934
rect 55030 -24981 55096 -24966
rect 55540 -24981 55606 -24966
rect 55030 -24982 55118 -24981
rect 55030 -25016 55046 -24982
rect 55080 -25016 55118 -24982
rect 55030 -25017 55118 -25016
rect 55518 -24982 55606 -24981
rect 55518 -25016 55556 -24982
rect 55590 -25016 55606 -24982
rect 55518 -25017 55606 -25016
rect 55030 -25032 55096 -25017
rect 53510 -25634 53630 -25596
rect 53510 -25668 53526 -25634
rect 53614 -25668 53630 -25634
rect 53510 -25684 53630 -25668
rect 55540 -25032 55606 -25017
rect 53972 -25650 54069 -25634
rect 53972 -25688 53988 -25650
rect 54022 -25688 54069 -25650
rect 53972 -25704 54069 -25688
rect 54869 -25650 54966 -25634
rect 54869 -25688 54916 -25650
rect 54950 -25688 54966 -25650
rect 54869 -25704 54966 -25688
rect 55326 -25336 55356 -25310
rect 55326 -25558 55356 -25536
rect 55308 -25574 55374 -25558
rect 55308 -25608 55324 -25574
rect 55358 -25608 55374 -25574
rect 55308 -25624 55374 -25608
rect 55866 -24770 55986 -24754
rect 55866 -24804 55882 -24770
rect 55970 -24804 55986 -24770
rect 55866 -24842 55986 -24804
rect 55866 -25680 55986 -25642
rect 55866 -25714 55882 -25680
rect 55970 -25714 55986 -25680
rect 55866 -25730 55986 -25714
rect 56476 -24206 56546 -24190
rect 56476 -24240 56492 -24206
rect 56530 -24240 56546 -24206
rect 56476 -24287 56546 -24240
rect 57175 -24185 57205 -24159
rect 57263 -24185 57293 -24159
rect 56476 -25134 56546 -25087
rect 56476 -25168 56492 -25134
rect 56530 -25168 56546 -25134
rect 56476 -25184 56546 -25168
rect 59087 -24078 59153 -24062
rect 59087 -24112 59103 -24078
rect 59137 -24112 59153 -24078
rect 59087 -24128 59153 -24112
rect 59090 -24159 59150 -24128
rect 59090 -24590 59150 -24559
rect 59087 -24606 59153 -24590
rect 59087 -24640 59103 -24606
rect 59137 -24640 59153 -24606
rect 59087 -24656 59153 -24640
rect 59858 -24020 59924 -24012
rect 60368 -24020 60434 -24012
rect 59858 -24028 59946 -24020
rect 59858 -24062 59874 -24028
rect 59908 -24062 59946 -24028
rect 59858 -24070 59946 -24062
rect 60346 -24028 60434 -24020
rect 60346 -24062 60384 -24028
rect 60418 -24062 60434 -24028
rect 60346 -24070 60434 -24062
rect 59858 -24078 59924 -24070
rect 60368 -24078 60434 -24070
rect 59530 -24298 59596 -24282
rect 59530 -24332 59546 -24298
rect 59580 -24332 59596 -24298
rect 59530 -24348 59596 -24332
rect 59548 -24370 59578 -24348
rect 59548 -24592 59578 -24570
rect 59530 -24608 59596 -24592
rect 59530 -24642 59546 -24608
rect 59580 -24642 59596 -24608
rect 59530 -24658 59596 -24642
rect 59846 -24298 59912 -24282
rect 59846 -24332 59862 -24298
rect 59896 -24332 59912 -24298
rect 59846 -24348 59912 -24332
rect 59864 -24370 59894 -24348
rect 59864 -24592 59894 -24570
rect 59846 -24608 59912 -24592
rect 59846 -24642 59862 -24608
rect 59896 -24642 59912 -24608
rect 59846 -24658 59912 -24642
rect 60343 -24565 60409 -24549
rect 61043 -24565 61109 -24549
rect 60343 -24599 60359 -24565
rect 60393 -24599 60409 -24565
rect 60343 -24617 60409 -24599
rect 61043 -24599 61059 -24565
rect 61093 -24599 61109 -24565
rect 61043 -24617 61109 -24599
rect 60165 -24647 60191 -24617
rect 60321 -24647 60441 -24617
rect 60641 -24647 60667 -24617
rect 60785 -24647 60811 -24617
rect 61011 -24647 61131 -24617
rect 61261 -24647 61287 -24617
rect 60343 -24657 60409 -24647
rect 60343 -24691 60359 -24657
rect 60393 -24691 60409 -24657
rect 60343 -24701 60409 -24691
rect 61043 -24657 61109 -24647
rect 61043 -24691 61059 -24657
rect 61093 -24691 61109 -24657
rect 61043 -24701 61109 -24691
rect 57175 -25229 57205 -25203
rect 57263 -25229 57293 -25203
rect 57175 -25348 57205 -25333
rect 57169 -25372 57205 -25348
rect 57169 -25381 57199 -25372
rect 57123 -25397 57199 -25381
rect 57263 -25394 57293 -25333
rect 59087 -24808 59153 -24792
rect 59087 -24842 59103 -24808
rect 59137 -24842 59153 -24808
rect 59087 -24858 59153 -24842
rect 59090 -24889 59150 -24858
rect 59090 -25320 59150 -25289
rect 57123 -25431 57133 -25397
rect 57167 -25431 57199 -25397
rect 57123 -25447 57199 -25431
rect 57169 -25482 57199 -25447
rect 57241 -25410 57295 -25394
rect 57241 -25444 57251 -25410
rect 57285 -25444 57295 -25410
rect 57241 -25460 57295 -25444
rect 59087 -25336 59153 -25320
rect 59087 -25370 59103 -25336
rect 59137 -25370 59153 -25336
rect 59087 -25386 59153 -25370
rect 60165 -24731 60191 -24701
rect 60321 -24731 60441 -24701
rect 60641 -24731 60667 -24701
rect 60785 -24731 60811 -24701
rect 61011 -24731 61131 -24701
rect 61261 -24731 61287 -24701
rect 59526 -24811 59596 -24780
rect 59526 -24830 59545 -24811
rect 59529 -24845 59545 -24830
rect 59579 -24830 59596 -24811
rect 59579 -24845 59595 -24830
rect 59529 -24861 59595 -24845
rect 59547 -24883 59577 -24861
rect 59547 -25105 59577 -25083
rect 59529 -25121 59595 -25105
rect 59529 -25155 59545 -25121
rect 59579 -25155 59595 -25121
rect 59529 -25171 59595 -25155
rect 59845 -24811 59911 -24795
rect 59845 -24845 59861 -24811
rect 59895 -24845 59911 -24811
rect 59845 -24861 59911 -24845
rect 60343 -24741 60409 -24731
rect 60343 -24775 60359 -24741
rect 60393 -24775 60409 -24741
rect 60343 -24785 60409 -24775
rect 61043 -24741 61109 -24731
rect 61043 -24775 61059 -24741
rect 61093 -24775 61109 -24741
rect 61043 -24785 61109 -24775
rect 59863 -24883 59893 -24861
rect 59863 -25105 59893 -25083
rect 59845 -25121 59911 -25105
rect 59845 -25155 59861 -25121
rect 59895 -25155 59911 -25121
rect 59845 -25171 59911 -25155
rect 60165 -24815 60191 -24785
rect 60321 -24815 60441 -24785
rect 60641 -24815 60667 -24785
rect 60785 -24815 60811 -24785
rect 61011 -24815 61131 -24785
rect 61261 -24815 61287 -24785
rect 60343 -24825 60409 -24815
rect 60343 -24859 60359 -24825
rect 60393 -24859 60409 -24825
rect 60343 -24869 60409 -24859
rect 61043 -24825 61109 -24815
rect 61043 -24859 61059 -24825
rect 61093 -24859 61109 -24825
rect 61043 -24869 61109 -24859
rect 60165 -24899 60191 -24869
rect 60321 -24899 60441 -24869
rect 60641 -24899 60667 -24869
rect 60785 -24899 60811 -24869
rect 61011 -24899 61131 -24869
rect 61261 -24899 61287 -24869
rect 57169 -25506 57205 -25482
rect 57175 -25521 57205 -25506
rect 57263 -25521 57293 -25460
rect 57175 -25705 57205 -25679
rect 57263 -25705 57293 -25679
rect 59544 -25600 59610 -25592
rect 59087 -25650 59113 -25600
rect 59513 -25608 59610 -25600
rect 59513 -25642 59560 -25608
rect 59594 -25642 59610 -25608
rect 59513 -25650 59610 -25642
rect 59544 -25658 59610 -25650
rect 59016 -25708 59082 -25700
rect 59016 -25716 59113 -25708
rect 59016 -25750 59032 -25716
rect 59066 -25750 59113 -25716
rect 59016 -25758 59113 -25750
rect 59513 -25758 59539 -25708
rect 59016 -25766 59082 -25758
rect 53972 -26006 54069 -25990
rect 53972 -26044 53988 -26006
rect 54022 -26044 54069 -26006
rect 53972 -26060 54069 -26044
rect 54869 -26006 54966 -25990
rect 54869 -26044 54916 -26006
rect 54950 -26044 54966 -26006
rect 54869 -26060 54966 -26044
rect 59858 -25386 59924 -25378
rect 60368 -25386 60434 -25378
rect 59858 -25394 59946 -25386
rect 59858 -25428 59874 -25394
rect 59908 -25428 59946 -25394
rect 59858 -25436 59946 -25428
rect 60346 -25394 60434 -25386
rect 60346 -25428 60384 -25394
rect 60418 -25428 60434 -25394
rect 60346 -25436 60434 -25428
rect 59858 -25444 59924 -25436
rect 60368 -25444 60434 -25436
rect 55510 -26202 55576 -26186
rect 55510 -26204 55526 -26202
rect 55262 -26234 55288 -26204
rect 55488 -26234 55526 -26204
rect 55510 -26236 55526 -26234
rect 55560 -26236 55576 -26202
rect 55510 -26252 55576 -26236
rect 53982 -28734 54079 -28718
rect 53982 -28772 53998 -28734
rect 54032 -28772 54079 -28734
rect 53982 -28788 54079 -28772
rect 54879 -28734 54976 -28718
rect 54879 -28772 54926 -28734
rect 54960 -28772 54976 -28734
rect 54879 -28788 54976 -28772
rect 53510 -29106 53630 -29090
rect 53510 -29140 53526 -29106
rect 53614 -29140 53630 -29106
rect 53510 -29178 53630 -29140
rect 53982 -29090 54079 -29074
rect 53982 -29128 53998 -29090
rect 54032 -29128 54079 -29090
rect 53982 -29144 54079 -29128
rect 54879 -29090 54976 -29074
rect 54879 -29128 54926 -29090
rect 54960 -29128 54976 -29090
rect 54879 -29144 54976 -29128
rect 55318 -29168 55384 -29152
rect 55318 -29202 55334 -29168
rect 55368 -29202 55384 -29168
rect 55318 -29218 55384 -29202
rect 55336 -29240 55366 -29218
rect 55336 -29466 55366 -29440
rect 53510 -30016 53630 -29978
rect 53510 -30050 53526 -30016
rect 53614 -30050 53630 -30016
rect 53510 -30066 53630 -30050
rect 53842 -29840 53930 -29824
rect 53842 -29928 53858 -29840
rect 53892 -29928 53930 -29840
rect 53842 -29944 53930 -29928
rect 54730 -29840 54818 -29824
rect 54730 -29928 54768 -29840
rect 54802 -29928 54818 -29840
rect 54730 -29944 54818 -29928
rect 55030 -29759 55096 -29744
rect 55540 -29759 55606 -29744
rect 55030 -29760 55118 -29759
rect 55030 -29794 55046 -29760
rect 55080 -29794 55118 -29760
rect 55030 -29795 55118 -29794
rect 55518 -29760 55606 -29759
rect 55518 -29794 55556 -29760
rect 55590 -29794 55606 -29760
rect 55518 -29795 55606 -29794
rect 55030 -29810 55096 -29795
rect 55540 -29810 55606 -29795
rect 55866 -29056 55986 -29040
rect 55866 -29090 55882 -29056
rect 55970 -29090 55986 -29056
rect 55866 -29128 55986 -29090
rect 55866 -29966 55986 -29928
rect 55866 -30000 55882 -29966
rect 55970 -30000 55986 -29966
rect 55866 -30016 55986 -30000
rect 57175 -29109 57205 -29083
rect 57263 -29109 57293 -29083
rect 57175 -29282 57205 -29267
rect 57169 -29306 57205 -29282
rect 57169 -29341 57199 -29306
rect 57263 -29328 57293 -29267
rect 59544 -29093 59610 -29085
rect 59087 -29143 59113 -29093
rect 59513 -29101 59610 -29093
rect 59513 -29135 59560 -29101
rect 59594 -29135 59610 -29101
rect 59513 -29143 59610 -29135
rect 59544 -29151 59610 -29143
rect 59016 -29201 59082 -29193
rect 59016 -29209 59113 -29201
rect 59016 -29243 59032 -29209
rect 59066 -29243 59113 -29209
rect 59016 -29251 59113 -29243
rect 59513 -29251 59539 -29201
rect 59016 -29259 59082 -29251
rect 57123 -29357 57199 -29341
rect 57123 -29391 57133 -29357
rect 57167 -29391 57199 -29357
rect 57123 -29407 57199 -29391
rect 57241 -29344 57295 -29328
rect 57241 -29378 57251 -29344
rect 57285 -29378 57295 -29344
rect 57241 -29394 57295 -29378
rect 57169 -29416 57199 -29407
rect 57169 -29440 57205 -29416
rect 57175 -29455 57205 -29440
rect 57263 -29455 57293 -29394
rect 53510 -30124 53630 -30108
rect 53510 -30158 53526 -30124
rect 53614 -30158 53630 -30124
rect 53510 -30196 53630 -30158
rect 53842 -30246 53930 -30230
rect 53842 -30334 53858 -30246
rect 53892 -30334 53930 -30246
rect 53842 -30350 53930 -30334
rect 54730 -30246 54818 -30230
rect 54730 -30334 54768 -30246
rect 54802 -30334 54818 -30246
rect 54730 -30350 54818 -30334
rect 55030 -30381 55096 -30366
rect 55540 -30381 55606 -30366
rect 55030 -30382 55118 -30381
rect 55030 -30416 55046 -30382
rect 55080 -30416 55118 -30382
rect 55030 -30417 55118 -30416
rect 55518 -30382 55606 -30381
rect 55518 -30416 55556 -30382
rect 55590 -30416 55606 -30382
rect 55518 -30417 55606 -30416
rect 55030 -30432 55096 -30417
rect 53510 -31034 53630 -30996
rect 53510 -31068 53526 -31034
rect 53614 -31068 53630 -31034
rect 53510 -31084 53630 -31068
rect 55540 -30432 55606 -30417
rect 53972 -31050 54069 -31034
rect 53972 -31088 53988 -31050
rect 54022 -31088 54069 -31050
rect 53972 -31104 54069 -31088
rect 54869 -31050 54966 -31034
rect 54869 -31088 54916 -31050
rect 54950 -31088 54966 -31050
rect 54869 -31104 54966 -31088
rect 55326 -30736 55356 -30710
rect 55326 -30958 55356 -30936
rect 55308 -30974 55374 -30958
rect 55308 -31008 55324 -30974
rect 55358 -31008 55374 -30974
rect 55308 -31024 55374 -31008
rect 55866 -30170 55986 -30154
rect 55866 -30204 55882 -30170
rect 55970 -30204 55986 -30170
rect 55866 -30242 55986 -30204
rect 55866 -31080 55986 -31042
rect 55866 -31114 55882 -31080
rect 55970 -31114 55986 -31080
rect 55866 -31130 55986 -31114
rect 56476 -29606 56546 -29590
rect 56476 -29640 56492 -29606
rect 56530 -29640 56546 -29606
rect 56476 -29687 56546 -29640
rect 57175 -29585 57205 -29559
rect 57263 -29585 57293 -29559
rect 56476 -30534 56546 -30487
rect 56476 -30568 56492 -30534
rect 56530 -30568 56546 -30534
rect 56476 -30584 56546 -30568
rect 59087 -29478 59153 -29462
rect 59087 -29512 59103 -29478
rect 59137 -29512 59153 -29478
rect 59087 -29528 59153 -29512
rect 59090 -29559 59150 -29528
rect 59090 -29990 59150 -29959
rect 59087 -30006 59153 -29990
rect 59087 -30040 59103 -30006
rect 59137 -30040 59153 -30006
rect 59087 -30056 59153 -30040
rect 59858 -29420 59924 -29412
rect 60368 -29420 60434 -29412
rect 59858 -29428 59946 -29420
rect 59858 -29462 59874 -29428
rect 59908 -29462 59946 -29428
rect 59858 -29470 59946 -29462
rect 60346 -29428 60434 -29420
rect 60346 -29462 60384 -29428
rect 60418 -29462 60434 -29428
rect 60346 -29470 60434 -29462
rect 59858 -29478 59924 -29470
rect 60368 -29478 60434 -29470
rect 59530 -29698 59596 -29682
rect 59530 -29732 59546 -29698
rect 59580 -29732 59596 -29698
rect 59530 -29748 59596 -29732
rect 59548 -29770 59578 -29748
rect 59548 -29992 59578 -29970
rect 59530 -30008 59596 -29992
rect 59530 -30042 59546 -30008
rect 59580 -30042 59596 -30008
rect 59530 -30058 59596 -30042
rect 59846 -29698 59912 -29682
rect 59846 -29732 59862 -29698
rect 59896 -29732 59912 -29698
rect 59846 -29748 59912 -29732
rect 59864 -29770 59894 -29748
rect 59864 -29992 59894 -29970
rect 59846 -30008 59912 -29992
rect 59846 -30042 59862 -30008
rect 59896 -30042 59912 -30008
rect 59846 -30058 59912 -30042
rect 60343 -29965 60409 -29949
rect 61043 -29965 61109 -29949
rect 60343 -29999 60359 -29965
rect 60393 -29999 60409 -29965
rect 60343 -30017 60409 -29999
rect 61043 -29999 61059 -29965
rect 61093 -29999 61109 -29965
rect 61043 -30017 61109 -29999
rect 60165 -30047 60191 -30017
rect 60321 -30047 60441 -30017
rect 60641 -30047 60667 -30017
rect 60785 -30047 60811 -30017
rect 61011 -30047 61131 -30017
rect 61261 -30047 61287 -30017
rect 60343 -30057 60409 -30047
rect 60343 -30091 60359 -30057
rect 60393 -30091 60409 -30057
rect 60343 -30101 60409 -30091
rect 61043 -30057 61109 -30047
rect 61043 -30091 61059 -30057
rect 61093 -30091 61109 -30057
rect 61043 -30101 61109 -30091
rect 57175 -30629 57205 -30603
rect 57263 -30629 57293 -30603
rect 57175 -30748 57205 -30733
rect 57169 -30772 57205 -30748
rect 57169 -30781 57199 -30772
rect 57123 -30797 57199 -30781
rect 57263 -30794 57293 -30733
rect 59087 -30208 59153 -30192
rect 59087 -30242 59103 -30208
rect 59137 -30242 59153 -30208
rect 59087 -30258 59153 -30242
rect 59090 -30289 59150 -30258
rect 59090 -30720 59150 -30689
rect 57123 -30831 57133 -30797
rect 57167 -30831 57199 -30797
rect 57123 -30847 57199 -30831
rect 57169 -30882 57199 -30847
rect 57241 -30810 57295 -30794
rect 57241 -30844 57251 -30810
rect 57285 -30844 57295 -30810
rect 57241 -30860 57295 -30844
rect 59087 -30736 59153 -30720
rect 59087 -30770 59103 -30736
rect 59137 -30770 59153 -30736
rect 59087 -30786 59153 -30770
rect 60165 -30131 60191 -30101
rect 60321 -30131 60441 -30101
rect 60641 -30131 60667 -30101
rect 60785 -30131 60811 -30101
rect 61011 -30131 61131 -30101
rect 61261 -30131 61287 -30101
rect 59526 -30211 59596 -30180
rect 59526 -30230 59545 -30211
rect 59529 -30245 59545 -30230
rect 59579 -30230 59596 -30211
rect 59579 -30245 59595 -30230
rect 59529 -30261 59595 -30245
rect 59547 -30283 59577 -30261
rect 59547 -30505 59577 -30483
rect 59529 -30521 59595 -30505
rect 59529 -30555 59545 -30521
rect 59579 -30555 59595 -30521
rect 59529 -30571 59595 -30555
rect 59845 -30211 59911 -30195
rect 59845 -30245 59861 -30211
rect 59895 -30245 59911 -30211
rect 59845 -30261 59911 -30245
rect 60343 -30141 60409 -30131
rect 60343 -30175 60359 -30141
rect 60393 -30175 60409 -30141
rect 60343 -30185 60409 -30175
rect 61043 -30141 61109 -30131
rect 61043 -30175 61059 -30141
rect 61093 -30175 61109 -30141
rect 61043 -30185 61109 -30175
rect 59863 -30283 59893 -30261
rect 59863 -30505 59893 -30483
rect 59845 -30521 59911 -30505
rect 59845 -30555 59861 -30521
rect 59895 -30555 59911 -30521
rect 59845 -30571 59911 -30555
rect 60165 -30215 60191 -30185
rect 60321 -30215 60441 -30185
rect 60641 -30215 60667 -30185
rect 60785 -30215 60811 -30185
rect 61011 -30215 61131 -30185
rect 61261 -30215 61287 -30185
rect 60343 -30225 60409 -30215
rect 60343 -30259 60359 -30225
rect 60393 -30259 60409 -30225
rect 60343 -30269 60409 -30259
rect 61043 -30225 61109 -30215
rect 61043 -30259 61059 -30225
rect 61093 -30259 61109 -30225
rect 61043 -30269 61109 -30259
rect 60165 -30299 60191 -30269
rect 60321 -30299 60441 -30269
rect 60641 -30299 60667 -30269
rect 60785 -30299 60811 -30269
rect 61011 -30299 61131 -30269
rect 61261 -30299 61287 -30269
rect 57169 -30906 57205 -30882
rect 57175 -30921 57205 -30906
rect 57263 -30921 57293 -30860
rect 57175 -31105 57205 -31079
rect 57263 -31105 57293 -31079
rect 59544 -31000 59610 -30992
rect 59087 -31050 59113 -31000
rect 59513 -31008 59610 -31000
rect 59513 -31042 59560 -31008
rect 59594 -31042 59610 -31008
rect 59513 -31050 59610 -31042
rect 59544 -31058 59610 -31050
rect 59016 -31108 59082 -31100
rect 59016 -31116 59113 -31108
rect 59016 -31150 59032 -31116
rect 59066 -31150 59113 -31116
rect 59016 -31158 59113 -31150
rect 59513 -31158 59539 -31108
rect 59016 -31166 59082 -31158
rect 53972 -31406 54069 -31390
rect 53972 -31444 53988 -31406
rect 54022 -31444 54069 -31406
rect 53972 -31460 54069 -31444
rect 54869 -31406 54966 -31390
rect 54869 -31444 54916 -31406
rect 54950 -31444 54966 -31406
rect 54869 -31460 54966 -31444
rect 59858 -30786 59924 -30778
rect 60368 -30786 60434 -30778
rect 59858 -30794 59946 -30786
rect 59858 -30828 59874 -30794
rect 59908 -30828 59946 -30794
rect 59858 -30836 59946 -30828
rect 60346 -30794 60434 -30786
rect 60346 -30828 60384 -30794
rect 60418 -30828 60434 -30794
rect 60346 -30836 60434 -30828
rect 59858 -30844 59924 -30836
rect 60368 -30844 60434 -30836
rect 55510 -31602 55576 -31586
rect 55510 -31604 55526 -31602
rect 55262 -31634 55288 -31604
rect 55488 -31634 55526 -31604
rect 55510 -31636 55526 -31634
rect 55560 -31636 55576 -31602
rect 55510 -31652 55576 -31636
rect 53982 -34134 54079 -34118
rect 53982 -34172 53998 -34134
rect 54032 -34172 54079 -34134
rect 53982 -34188 54079 -34172
rect 54879 -34134 54976 -34118
rect 54879 -34172 54926 -34134
rect 54960 -34172 54976 -34134
rect 54879 -34188 54976 -34172
rect 53510 -34506 53630 -34490
rect 53510 -34540 53526 -34506
rect 53614 -34540 53630 -34506
rect 53510 -34578 53630 -34540
rect 53982 -34490 54079 -34474
rect 53982 -34528 53998 -34490
rect 54032 -34528 54079 -34490
rect 53982 -34544 54079 -34528
rect 54879 -34490 54976 -34474
rect 54879 -34528 54926 -34490
rect 54960 -34528 54976 -34490
rect 54879 -34544 54976 -34528
rect 55318 -34568 55384 -34552
rect 55318 -34602 55334 -34568
rect 55368 -34602 55384 -34568
rect 55318 -34618 55384 -34602
rect 55336 -34640 55366 -34618
rect 55336 -34866 55366 -34840
rect 53510 -35416 53630 -35378
rect 53510 -35450 53526 -35416
rect 53614 -35450 53630 -35416
rect 53510 -35466 53630 -35450
rect 53842 -35240 53930 -35224
rect 53842 -35328 53858 -35240
rect 53892 -35328 53930 -35240
rect 53842 -35344 53930 -35328
rect 54730 -35240 54818 -35224
rect 54730 -35328 54768 -35240
rect 54802 -35328 54818 -35240
rect 54730 -35344 54818 -35328
rect 55030 -35159 55096 -35144
rect 55540 -35159 55606 -35144
rect 55030 -35160 55118 -35159
rect 55030 -35194 55046 -35160
rect 55080 -35194 55118 -35160
rect 55030 -35195 55118 -35194
rect 55518 -35160 55606 -35159
rect 55518 -35194 55556 -35160
rect 55590 -35194 55606 -35160
rect 55518 -35195 55606 -35194
rect 55030 -35210 55096 -35195
rect 55540 -35210 55606 -35195
rect 55866 -34456 55986 -34440
rect 55866 -34490 55882 -34456
rect 55970 -34490 55986 -34456
rect 55866 -34528 55986 -34490
rect 55866 -35366 55986 -35328
rect 55866 -35400 55882 -35366
rect 55970 -35400 55986 -35366
rect 55866 -35416 55986 -35400
rect 57175 -34509 57205 -34483
rect 57263 -34509 57293 -34483
rect 57175 -34682 57205 -34667
rect 57169 -34706 57205 -34682
rect 57169 -34741 57199 -34706
rect 57263 -34728 57293 -34667
rect 59544 -34493 59610 -34485
rect 59087 -34543 59113 -34493
rect 59513 -34501 59610 -34493
rect 59513 -34535 59560 -34501
rect 59594 -34535 59610 -34501
rect 59513 -34543 59610 -34535
rect 59544 -34551 59610 -34543
rect 59016 -34601 59082 -34593
rect 59016 -34609 59113 -34601
rect 59016 -34643 59032 -34609
rect 59066 -34643 59113 -34609
rect 59016 -34651 59113 -34643
rect 59513 -34651 59539 -34601
rect 59016 -34659 59082 -34651
rect 57123 -34757 57199 -34741
rect 57123 -34791 57133 -34757
rect 57167 -34791 57199 -34757
rect 57123 -34807 57199 -34791
rect 57241 -34744 57295 -34728
rect 57241 -34778 57251 -34744
rect 57285 -34778 57295 -34744
rect 57241 -34794 57295 -34778
rect 57169 -34816 57199 -34807
rect 57169 -34840 57205 -34816
rect 57175 -34855 57205 -34840
rect 57263 -34855 57293 -34794
rect 53510 -35524 53630 -35508
rect 53510 -35558 53526 -35524
rect 53614 -35558 53630 -35524
rect 53510 -35596 53630 -35558
rect 53842 -35646 53930 -35630
rect 53842 -35734 53858 -35646
rect 53892 -35734 53930 -35646
rect 53842 -35750 53930 -35734
rect 54730 -35646 54818 -35630
rect 54730 -35734 54768 -35646
rect 54802 -35734 54818 -35646
rect 54730 -35750 54818 -35734
rect 55030 -35781 55096 -35766
rect 55540 -35781 55606 -35766
rect 55030 -35782 55118 -35781
rect 55030 -35816 55046 -35782
rect 55080 -35816 55118 -35782
rect 55030 -35817 55118 -35816
rect 55518 -35782 55606 -35781
rect 55518 -35816 55556 -35782
rect 55590 -35816 55606 -35782
rect 55518 -35817 55606 -35816
rect 55030 -35832 55096 -35817
rect 53510 -36434 53630 -36396
rect 53510 -36468 53526 -36434
rect 53614 -36468 53630 -36434
rect 53510 -36484 53630 -36468
rect 55540 -35832 55606 -35817
rect 53972 -36450 54069 -36434
rect 53972 -36488 53988 -36450
rect 54022 -36488 54069 -36450
rect 53972 -36504 54069 -36488
rect 54869 -36450 54966 -36434
rect 54869 -36488 54916 -36450
rect 54950 -36488 54966 -36450
rect 54869 -36504 54966 -36488
rect 55326 -36136 55356 -36110
rect 55326 -36358 55356 -36336
rect 55308 -36374 55374 -36358
rect 55308 -36408 55324 -36374
rect 55358 -36408 55374 -36374
rect 55308 -36424 55374 -36408
rect 55866 -35570 55986 -35554
rect 55866 -35604 55882 -35570
rect 55970 -35604 55986 -35570
rect 55866 -35642 55986 -35604
rect 55866 -36480 55986 -36442
rect 55866 -36514 55882 -36480
rect 55970 -36514 55986 -36480
rect 55866 -36530 55986 -36514
rect 56476 -35006 56546 -34990
rect 56476 -35040 56492 -35006
rect 56530 -35040 56546 -35006
rect 56476 -35087 56546 -35040
rect 57175 -34985 57205 -34959
rect 57263 -34985 57293 -34959
rect 56476 -35934 56546 -35887
rect 56476 -35968 56492 -35934
rect 56530 -35968 56546 -35934
rect 56476 -35984 56546 -35968
rect 59087 -34878 59153 -34862
rect 59087 -34912 59103 -34878
rect 59137 -34912 59153 -34878
rect 59087 -34928 59153 -34912
rect 59090 -34959 59150 -34928
rect 59090 -35390 59150 -35359
rect 59087 -35406 59153 -35390
rect 59087 -35440 59103 -35406
rect 59137 -35440 59153 -35406
rect 59087 -35456 59153 -35440
rect 59858 -34820 59924 -34812
rect 60368 -34820 60434 -34812
rect 59858 -34828 59946 -34820
rect 59858 -34862 59874 -34828
rect 59908 -34862 59946 -34828
rect 59858 -34870 59946 -34862
rect 60346 -34828 60434 -34820
rect 60346 -34862 60384 -34828
rect 60418 -34862 60434 -34828
rect 60346 -34870 60434 -34862
rect 59858 -34878 59924 -34870
rect 60368 -34878 60434 -34870
rect 59530 -35098 59596 -35082
rect 59530 -35132 59546 -35098
rect 59580 -35132 59596 -35098
rect 59530 -35148 59596 -35132
rect 59548 -35170 59578 -35148
rect 59548 -35392 59578 -35370
rect 59530 -35408 59596 -35392
rect 59530 -35442 59546 -35408
rect 59580 -35442 59596 -35408
rect 59530 -35458 59596 -35442
rect 59846 -35098 59912 -35082
rect 59846 -35132 59862 -35098
rect 59896 -35132 59912 -35098
rect 59846 -35148 59912 -35132
rect 59864 -35170 59894 -35148
rect 59864 -35392 59894 -35370
rect 59846 -35408 59912 -35392
rect 59846 -35442 59862 -35408
rect 59896 -35442 59912 -35408
rect 59846 -35458 59912 -35442
rect 60343 -35365 60409 -35349
rect 61043 -35365 61109 -35349
rect 60343 -35399 60359 -35365
rect 60393 -35399 60409 -35365
rect 60343 -35417 60409 -35399
rect 61043 -35399 61059 -35365
rect 61093 -35399 61109 -35365
rect 61043 -35417 61109 -35399
rect 60165 -35447 60191 -35417
rect 60321 -35447 60441 -35417
rect 60641 -35447 60667 -35417
rect 60785 -35447 60811 -35417
rect 61011 -35447 61131 -35417
rect 61261 -35447 61287 -35417
rect 60343 -35457 60409 -35447
rect 60343 -35491 60359 -35457
rect 60393 -35491 60409 -35457
rect 60343 -35501 60409 -35491
rect 61043 -35457 61109 -35447
rect 61043 -35491 61059 -35457
rect 61093 -35491 61109 -35457
rect 61043 -35501 61109 -35491
rect 57175 -36029 57205 -36003
rect 57263 -36029 57293 -36003
rect 57175 -36148 57205 -36133
rect 57169 -36172 57205 -36148
rect 57169 -36181 57199 -36172
rect 57123 -36197 57199 -36181
rect 57263 -36194 57293 -36133
rect 59087 -35608 59153 -35592
rect 59087 -35642 59103 -35608
rect 59137 -35642 59153 -35608
rect 59087 -35658 59153 -35642
rect 59090 -35689 59150 -35658
rect 59090 -36120 59150 -36089
rect 57123 -36231 57133 -36197
rect 57167 -36231 57199 -36197
rect 57123 -36247 57199 -36231
rect 57169 -36282 57199 -36247
rect 57241 -36210 57295 -36194
rect 57241 -36244 57251 -36210
rect 57285 -36244 57295 -36210
rect 57241 -36260 57295 -36244
rect 59087 -36136 59153 -36120
rect 59087 -36170 59103 -36136
rect 59137 -36170 59153 -36136
rect 59087 -36186 59153 -36170
rect 60165 -35531 60191 -35501
rect 60321 -35531 60441 -35501
rect 60641 -35531 60667 -35501
rect 60785 -35531 60811 -35501
rect 61011 -35531 61131 -35501
rect 61261 -35531 61287 -35501
rect 59526 -35611 59596 -35580
rect 59526 -35630 59545 -35611
rect 59529 -35645 59545 -35630
rect 59579 -35630 59596 -35611
rect 59579 -35645 59595 -35630
rect 59529 -35661 59595 -35645
rect 59547 -35683 59577 -35661
rect 59547 -35905 59577 -35883
rect 59529 -35921 59595 -35905
rect 59529 -35955 59545 -35921
rect 59579 -35955 59595 -35921
rect 59529 -35971 59595 -35955
rect 59845 -35611 59911 -35595
rect 59845 -35645 59861 -35611
rect 59895 -35645 59911 -35611
rect 59845 -35661 59911 -35645
rect 60343 -35541 60409 -35531
rect 60343 -35575 60359 -35541
rect 60393 -35575 60409 -35541
rect 60343 -35585 60409 -35575
rect 61043 -35541 61109 -35531
rect 61043 -35575 61059 -35541
rect 61093 -35575 61109 -35541
rect 61043 -35585 61109 -35575
rect 59863 -35683 59893 -35661
rect 59863 -35905 59893 -35883
rect 59845 -35921 59911 -35905
rect 59845 -35955 59861 -35921
rect 59895 -35955 59911 -35921
rect 59845 -35971 59911 -35955
rect 60165 -35615 60191 -35585
rect 60321 -35615 60441 -35585
rect 60641 -35615 60667 -35585
rect 60785 -35615 60811 -35585
rect 61011 -35615 61131 -35585
rect 61261 -35615 61287 -35585
rect 60343 -35625 60409 -35615
rect 60343 -35659 60359 -35625
rect 60393 -35659 60409 -35625
rect 60343 -35669 60409 -35659
rect 61043 -35625 61109 -35615
rect 61043 -35659 61059 -35625
rect 61093 -35659 61109 -35625
rect 61043 -35669 61109 -35659
rect 60165 -35699 60191 -35669
rect 60321 -35699 60441 -35669
rect 60641 -35699 60667 -35669
rect 60785 -35699 60811 -35669
rect 61011 -35699 61131 -35669
rect 61261 -35699 61287 -35669
rect 57169 -36306 57205 -36282
rect 57175 -36321 57205 -36306
rect 57263 -36321 57293 -36260
rect 57175 -36505 57205 -36479
rect 57263 -36505 57293 -36479
rect 59544 -36400 59610 -36392
rect 59087 -36450 59113 -36400
rect 59513 -36408 59610 -36400
rect 59513 -36442 59560 -36408
rect 59594 -36442 59610 -36408
rect 59513 -36450 59610 -36442
rect 59544 -36458 59610 -36450
rect 59016 -36508 59082 -36500
rect 59016 -36516 59113 -36508
rect 59016 -36550 59032 -36516
rect 59066 -36550 59113 -36516
rect 59016 -36558 59113 -36550
rect 59513 -36558 59539 -36508
rect 59016 -36566 59082 -36558
rect 53972 -36806 54069 -36790
rect 53972 -36844 53988 -36806
rect 54022 -36844 54069 -36806
rect 53972 -36860 54069 -36844
rect 54869 -36806 54966 -36790
rect 54869 -36844 54916 -36806
rect 54950 -36844 54966 -36806
rect 54869 -36860 54966 -36844
rect 59858 -36186 59924 -36178
rect 60368 -36186 60434 -36178
rect 59858 -36194 59946 -36186
rect 59858 -36228 59874 -36194
rect 59908 -36228 59946 -36194
rect 59858 -36236 59946 -36228
rect 60346 -36194 60434 -36186
rect 60346 -36228 60384 -36194
rect 60418 -36228 60434 -36194
rect 60346 -36236 60434 -36228
rect 59858 -36244 59924 -36236
rect 60368 -36244 60434 -36236
rect 55510 -37002 55576 -36986
rect 55510 -37004 55526 -37002
rect 55262 -37034 55288 -37004
rect 55488 -37034 55526 -37004
rect 55510 -37036 55526 -37034
rect 55560 -37036 55576 -37002
rect 55510 -37052 55576 -37036
rect 75626 -38435 75656 -38409
rect 75902 -38435 75932 -38409
rect 76176 -38435 76206 -38409
rect 76452 -38435 76482 -38409
rect 76728 -38435 76758 -38409
rect 75626 -38587 75656 -38565
rect 75902 -38587 75932 -38565
rect 76176 -38587 76206 -38565
rect 76452 -38587 76482 -38565
rect 76728 -38587 76758 -38565
rect 75570 -38603 75656 -38587
rect 75570 -38637 75586 -38603
rect 75620 -38637 75656 -38603
rect 75570 -38653 75656 -38637
rect 75846 -38603 75932 -38587
rect 75846 -38637 75862 -38603
rect 75896 -38637 75932 -38603
rect 75846 -38653 75932 -38637
rect 76120 -38603 76206 -38587
rect 76120 -38637 76136 -38603
rect 76170 -38637 76206 -38603
rect 76120 -38653 76206 -38637
rect 76396 -38603 76482 -38587
rect 76396 -38637 76412 -38603
rect 76446 -38637 76482 -38603
rect 76396 -38653 76482 -38637
rect 76672 -38603 76758 -38587
rect 76672 -38637 76688 -38603
rect 76722 -38637 76758 -38603
rect 76672 -38653 76758 -38637
rect 75626 -38685 75656 -38653
rect 75902 -38685 75932 -38653
rect 76176 -38685 76206 -38653
rect 76452 -38685 76482 -38653
rect 76728 -38685 76758 -38653
rect 75626 -38911 75656 -38885
rect 75902 -38911 75932 -38885
rect 76176 -38911 76206 -38885
rect 76452 -38911 76482 -38885
rect 76728 -38911 76758 -38885
rect 78019 -39105 78049 -39079
rect 78477 -39105 78507 -39079
rect 78897 -39105 78927 -39079
rect 77819 -39129 77885 -39119
rect 77819 -39163 77835 -39129
rect 77869 -39163 77885 -39129
rect 77819 -39173 77885 -39163
rect 77657 -39221 77687 -39195
rect 77753 -39221 77783 -39195
rect 77825 -39221 77855 -39173
rect 77921 -39221 77951 -39195
rect 78277 -39129 78343 -39119
rect 78277 -39163 78293 -39129
rect 78327 -39163 78343 -39129
rect 78277 -39173 78343 -39163
rect 78211 -39221 78241 -39195
rect 78283 -39221 78313 -39173
rect 78379 -39221 78409 -39195
rect 78705 -39147 78735 -39121
rect 78789 -39147 78819 -39121
rect 77657 -39337 77687 -39305
rect 77753 -39337 77783 -39305
rect 77603 -39353 77687 -39337
rect 77603 -39387 77613 -39353
rect 77647 -39387 77687 -39353
rect 77603 -39403 77687 -39387
rect 77729 -39353 77783 -39337
rect 77729 -39387 77739 -39353
rect 77773 -39387 77783 -39353
rect 77729 -39403 77783 -39387
rect 53982 -39534 54079 -39518
rect 53982 -39572 53998 -39534
rect 54032 -39572 54079 -39534
rect 53982 -39588 54079 -39572
rect 54879 -39534 54976 -39518
rect 54879 -39572 54926 -39534
rect 54960 -39572 54976 -39534
rect 54879 -39588 54976 -39572
rect 77657 -39465 77687 -39403
rect 77753 -39465 77783 -39403
rect 77825 -39420 77855 -39305
rect 77921 -39337 77951 -39305
rect 78019 -39337 78049 -39305
rect 78211 -39337 78241 -39305
rect 77905 -39353 77959 -39337
rect 77905 -39387 77915 -39353
rect 77949 -39387 77959 -39353
rect 77905 -39403 77959 -39387
rect 78001 -39353 78056 -39337
rect 78001 -39387 78011 -39353
rect 78045 -39387 78056 -39353
rect 78001 -39403 78056 -39387
rect 78154 -39353 78241 -39337
rect 78154 -39387 78164 -39353
rect 78198 -39387 78241 -39353
rect 78154 -39403 78241 -39387
rect 77825 -39421 77866 -39420
rect 77825 -39450 77867 -39421
rect 77837 -39465 77867 -39450
rect 77921 -39465 77951 -39403
rect 78019 -39425 78049 -39403
rect 77657 -39575 77687 -39549
rect 77753 -39575 77783 -39549
rect 77837 -39575 77867 -39549
rect 77921 -39575 77951 -39549
rect 78211 -39465 78241 -39403
rect 78283 -39420 78313 -39305
rect 78379 -39337 78409 -39305
rect 78477 -39337 78507 -39305
rect 78705 -39337 78735 -39231
rect 78364 -39353 78418 -39337
rect 78364 -39387 78374 -39353
rect 78408 -39387 78418 -39353
rect 78364 -39403 78418 -39387
rect 78460 -39353 78514 -39337
rect 78460 -39387 78470 -39353
rect 78504 -39387 78514 -39353
rect 78460 -39403 78514 -39387
rect 78648 -39353 78735 -39337
rect 78648 -39387 78664 -39353
rect 78698 -39387 78735 -39353
rect 78648 -39403 78735 -39387
rect 78283 -39450 78325 -39420
rect 78295 -39465 78325 -39450
rect 78379 -39465 78409 -39403
rect 78477 -39425 78507 -39403
rect 78019 -39581 78049 -39555
rect 78211 -39575 78241 -39549
rect 78295 -39575 78325 -39549
rect 78379 -39575 78409 -39549
rect 78705 -39443 78735 -39403
rect 78789 -39337 78819 -39231
rect 80858 -39155 80888 -39129
rect 81103 -39155 81133 -39129
rect 81187 -39155 81217 -39129
rect 81271 -39155 81301 -39129
rect 81355 -39155 81385 -39129
rect 81566 -39155 81596 -39129
rect 81650 -39155 81680 -39129
rect 81734 -39155 81764 -39129
rect 81818 -39155 81848 -39129
rect 81902 -39155 81932 -39129
rect 81986 -39155 82016 -39129
rect 82070 -39155 82100 -39129
rect 82154 -39155 82184 -39129
rect 82238 -39155 82268 -39129
rect 82322 -39155 82352 -39129
rect 82406 -39155 82436 -39129
rect 82490 -39155 82520 -39129
rect 82574 -39155 82604 -39129
rect 82658 -39155 82688 -39129
rect 82742 -39155 82772 -39129
rect 82826 -39155 82856 -39129
rect 83038 -39155 83068 -39129
rect 83122 -39155 83152 -39129
rect 83206 -39155 83236 -39129
rect 83290 -39155 83320 -39129
rect 83374 -39155 83404 -39129
rect 83458 -39155 83488 -39129
rect 83542 -39155 83572 -39129
rect 83626 -39155 83656 -39129
rect 83710 -39155 83740 -39129
rect 83794 -39155 83824 -39129
rect 83878 -39155 83908 -39129
rect 83962 -39155 83992 -39129
rect 84046 -39155 84076 -39129
rect 84130 -39155 84160 -39129
rect 84214 -39155 84244 -39129
rect 84298 -39155 84328 -39129
rect 84510 -39155 84540 -39129
rect 84594 -39155 84624 -39129
rect 84678 -39155 84708 -39129
rect 84762 -39155 84792 -39129
rect 84846 -39155 84876 -39129
rect 84930 -39155 84960 -39129
rect 85014 -39155 85044 -39129
rect 85098 -39155 85128 -39129
rect 85182 -39155 85212 -39129
rect 85266 -39155 85296 -39129
rect 85350 -39155 85380 -39129
rect 85434 -39155 85464 -39129
rect 85518 -39155 85548 -39129
rect 85602 -39155 85632 -39129
rect 85686 -39155 85716 -39129
rect 85770 -39155 85800 -39129
rect 85982 -39155 86012 -39129
rect 86066 -39155 86096 -39129
rect 86150 -39155 86180 -39129
rect 86234 -39155 86264 -39129
rect 86318 -39155 86348 -39129
rect 86402 -39155 86432 -39129
rect 86486 -39155 86516 -39129
rect 86570 -39155 86600 -39129
rect 86654 -39155 86684 -39129
rect 86738 -39155 86768 -39129
rect 86822 -39155 86852 -39129
rect 86906 -39155 86936 -39129
rect 86990 -39155 87020 -39129
rect 87074 -39155 87104 -39129
rect 87158 -39155 87188 -39129
rect 87242 -39155 87272 -39129
rect 87454 -39155 87484 -39129
rect 87538 -39155 87568 -39129
rect 87622 -39155 87652 -39129
rect 87706 -39155 87736 -39129
rect 87790 -39155 87820 -39129
rect 87874 -39155 87904 -39129
rect 87958 -39155 87988 -39129
rect 88042 -39155 88072 -39129
rect 88126 -39155 88156 -39129
rect 88210 -39155 88240 -39129
rect 88294 -39155 88324 -39129
rect 88378 -39155 88408 -39129
rect 88462 -39155 88492 -39129
rect 88546 -39155 88576 -39129
rect 88630 -39155 88660 -39129
rect 88714 -39155 88744 -39129
rect 78897 -39337 78927 -39305
rect 78789 -39353 78855 -39337
rect 78789 -39387 78805 -39353
rect 78839 -39387 78855 -39353
rect 78789 -39403 78855 -39387
rect 78897 -39353 78963 -39337
rect 78897 -39387 78913 -39353
rect 78947 -39387 78963 -39353
rect 80858 -39387 80888 -39355
rect 81103 -39387 81133 -39355
rect 81187 -39387 81217 -39355
rect 81271 -39387 81301 -39355
rect 81355 -39387 81385 -39355
rect 81566 -39387 81596 -39355
rect 81650 -39387 81680 -39355
rect 81734 -39387 81764 -39355
rect 81818 -39387 81848 -39355
rect 81902 -39387 81932 -39355
rect 81986 -39387 82016 -39355
rect 82070 -39387 82100 -39355
rect 82154 -39387 82184 -39355
rect 82238 -39387 82268 -39355
rect 82322 -39387 82352 -39355
rect 82406 -39387 82436 -39355
rect 82490 -39387 82520 -39355
rect 82574 -39387 82604 -39355
rect 82658 -39387 82688 -39355
rect 82742 -39387 82772 -39355
rect 82826 -39387 82856 -39355
rect 83038 -39387 83068 -39355
rect 83122 -39387 83152 -39355
rect 83206 -39387 83236 -39355
rect 83290 -39387 83320 -39355
rect 83374 -39387 83404 -39355
rect 83458 -39387 83488 -39355
rect 83542 -39387 83572 -39355
rect 83626 -39387 83656 -39355
rect 83710 -39387 83740 -39355
rect 83794 -39387 83824 -39355
rect 83878 -39387 83908 -39355
rect 83962 -39387 83992 -39355
rect 84046 -39387 84076 -39355
rect 84130 -39387 84160 -39355
rect 84214 -39387 84244 -39355
rect 84298 -39387 84328 -39355
rect 84510 -39387 84540 -39355
rect 84594 -39387 84624 -39355
rect 84678 -39387 84708 -39355
rect 84762 -39387 84792 -39355
rect 84846 -39387 84876 -39355
rect 84930 -39387 84960 -39355
rect 85014 -39387 85044 -39355
rect 85098 -39387 85128 -39355
rect 85182 -39387 85212 -39355
rect 85266 -39387 85296 -39355
rect 85350 -39387 85380 -39355
rect 85434 -39387 85464 -39355
rect 85518 -39387 85548 -39355
rect 85602 -39387 85632 -39355
rect 85686 -39387 85716 -39355
rect 85770 -39387 85800 -39355
rect 85982 -39387 86012 -39355
rect 86066 -39387 86096 -39355
rect 86150 -39387 86180 -39355
rect 86234 -39387 86264 -39355
rect 86318 -39387 86348 -39355
rect 86402 -39387 86432 -39355
rect 86486 -39387 86516 -39355
rect 86570 -39387 86600 -39355
rect 86654 -39387 86684 -39355
rect 86738 -39387 86768 -39355
rect 86822 -39387 86852 -39355
rect 86906 -39387 86936 -39355
rect 86990 -39387 87020 -39355
rect 87074 -39387 87104 -39355
rect 87158 -39387 87188 -39355
rect 87242 -39387 87272 -39355
rect 87454 -39387 87484 -39355
rect 87538 -39387 87568 -39355
rect 87622 -39387 87652 -39355
rect 87706 -39387 87736 -39355
rect 87790 -39387 87820 -39355
rect 87874 -39387 87904 -39355
rect 87958 -39387 87988 -39355
rect 88042 -39387 88072 -39355
rect 88126 -39387 88156 -39355
rect 88210 -39387 88240 -39355
rect 88294 -39387 88324 -39355
rect 88378 -39387 88408 -39355
rect 88462 -39387 88492 -39355
rect 88546 -39387 88576 -39355
rect 88630 -39387 88660 -39355
rect 88714 -39387 88744 -39355
rect 78897 -39403 78963 -39387
rect 80802 -39403 80888 -39387
rect 78789 -39443 78819 -39403
rect 78897 -39425 78927 -39403
rect 78705 -39553 78735 -39527
rect 78789 -39553 78819 -39527
rect 80802 -39437 80818 -39403
rect 80852 -39437 80888 -39403
rect 80802 -39453 80888 -39437
rect 81035 -39403 81385 -39387
rect 81035 -39437 81051 -39403
rect 81085 -39437 81143 -39403
rect 81177 -39437 81227 -39403
rect 81261 -39437 81311 -39403
rect 81345 -39437 81385 -39403
rect 81035 -39453 81385 -39437
rect 81500 -39403 82856 -39387
rect 81500 -39437 81516 -39403
rect 81550 -39437 81690 -39403
rect 81724 -39437 81858 -39403
rect 81892 -39437 82027 -39403
rect 82061 -39437 82194 -39403
rect 82228 -39437 82362 -39403
rect 82396 -39437 82529 -39403
rect 82563 -39437 82856 -39403
rect 81500 -39453 82856 -39437
rect 82972 -39403 84328 -39387
rect 82972 -39437 82988 -39403
rect 83022 -39437 83162 -39403
rect 83196 -39437 83330 -39403
rect 83364 -39437 83499 -39403
rect 83533 -39437 83666 -39403
rect 83700 -39437 83834 -39403
rect 83868 -39437 84001 -39403
rect 84035 -39437 84328 -39403
rect 82972 -39453 84328 -39437
rect 84444 -39403 85800 -39387
rect 84444 -39437 84460 -39403
rect 84494 -39437 84634 -39403
rect 84668 -39437 84802 -39403
rect 84836 -39437 84971 -39403
rect 85005 -39437 85138 -39403
rect 85172 -39437 85306 -39403
rect 85340 -39437 85473 -39403
rect 85507 -39437 85800 -39403
rect 84444 -39453 85800 -39437
rect 85916 -39403 87272 -39387
rect 85916 -39437 85932 -39403
rect 85966 -39437 86106 -39403
rect 86140 -39437 86274 -39403
rect 86308 -39437 86443 -39403
rect 86477 -39437 86610 -39403
rect 86644 -39437 86778 -39403
rect 86812 -39437 86945 -39403
rect 86979 -39437 87272 -39403
rect 85916 -39453 87272 -39437
rect 87388 -39403 88744 -39387
rect 87388 -39437 87404 -39403
rect 87438 -39437 87578 -39403
rect 87612 -39437 87746 -39403
rect 87780 -39437 87915 -39403
rect 87949 -39437 88082 -39403
rect 88116 -39437 88250 -39403
rect 88284 -39437 88417 -39403
rect 88451 -39437 88744 -39403
rect 87388 -39453 88744 -39437
rect 80858 -39475 80888 -39453
rect 81103 -39475 81133 -39453
rect 81187 -39475 81217 -39453
rect 81271 -39475 81301 -39453
rect 81355 -39475 81385 -39453
rect 81566 -39475 81596 -39453
rect 81650 -39475 81680 -39453
rect 81734 -39475 81764 -39453
rect 81818 -39475 81848 -39453
rect 81902 -39475 81932 -39453
rect 81986 -39475 82016 -39453
rect 82070 -39475 82100 -39453
rect 82154 -39475 82184 -39453
rect 82238 -39475 82268 -39453
rect 82322 -39475 82352 -39453
rect 82406 -39475 82436 -39453
rect 82490 -39475 82520 -39453
rect 82574 -39475 82604 -39453
rect 82658 -39475 82688 -39453
rect 82742 -39475 82772 -39453
rect 82826 -39475 82856 -39453
rect 83038 -39475 83068 -39453
rect 83122 -39475 83152 -39453
rect 83206 -39475 83236 -39453
rect 83290 -39475 83320 -39453
rect 83374 -39475 83404 -39453
rect 83458 -39475 83488 -39453
rect 83542 -39475 83572 -39453
rect 83626 -39475 83656 -39453
rect 83710 -39475 83740 -39453
rect 83794 -39475 83824 -39453
rect 83878 -39475 83908 -39453
rect 83962 -39475 83992 -39453
rect 84046 -39475 84076 -39453
rect 84130 -39475 84160 -39453
rect 84214 -39475 84244 -39453
rect 84298 -39475 84328 -39453
rect 84510 -39475 84540 -39453
rect 84594 -39475 84624 -39453
rect 84678 -39475 84708 -39453
rect 84762 -39475 84792 -39453
rect 84846 -39475 84876 -39453
rect 84930 -39475 84960 -39453
rect 85014 -39475 85044 -39453
rect 85098 -39475 85128 -39453
rect 85182 -39475 85212 -39453
rect 85266 -39475 85296 -39453
rect 85350 -39475 85380 -39453
rect 85434 -39475 85464 -39453
rect 85518 -39475 85548 -39453
rect 85602 -39475 85632 -39453
rect 85686 -39475 85716 -39453
rect 85770 -39475 85800 -39453
rect 85982 -39475 86012 -39453
rect 86066 -39475 86096 -39453
rect 86150 -39475 86180 -39453
rect 86234 -39475 86264 -39453
rect 86318 -39475 86348 -39453
rect 86402 -39475 86432 -39453
rect 86486 -39475 86516 -39453
rect 86570 -39475 86600 -39453
rect 86654 -39475 86684 -39453
rect 86738 -39475 86768 -39453
rect 86822 -39475 86852 -39453
rect 86906 -39475 86936 -39453
rect 86990 -39475 87020 -39453
rect 87074 -39475 87104 -39453
rect 87158 -39475 87188 -39453
rect 87242 -39475 87272 -39453
rect 87454 -39475 87484 -39453
rect 87538 -39475 87568 -39453
rect 87622 -39475 87652 -39453
rect 87706 -39475 87736 -39453
rect 87790 -39475 87820 -39453
rect 87874 -39475 87904 -39453
rect 87958 -39475 87988 -39453
rect 88042 -39475 88072 -39453
rect 88126 -39475 88156 -39453
rect 88210 -39475 88240 -39453
rect 88294 -39475 88324 -39453
rect 88378 -39475 88408 -39453
rect 88462 -39475 88492 -39453
rect 88546 -39475 88576 -39453
rect 88630 -39475 88660 -39453
rect 88714 -39475 88744 -39453
rect 78477 -39581 78507 -39555
rect 78897 -39581 78927 -39555
rect 80858 -39631 80888 -39605
rect 81103 -39631 81133 -39605
rect 81187 -39631 81217 -39605
rect 81271 -39631 81301 -39605
rect 81355 -39631 81385 -39605
rect 81566 -39631 81596 -39605
rect 81650 -39631 81680 -39605
rect 81734 -39631 81764 -39605
rect 81818 -39631 81848 -39605
rect 81902 -39631 81932 -39605
rect 81986 -39631 82016 -39605
rect 82070 -39631 82100 -39605
rect 82154 -39631 82184 -39605
rect 82238 -39631 82268 -39605
rect 82322 -39631 82352 -39605
rect 82406 -39631 82436 -39605
rect 82490 -39631 82520 -39605
rect 82574 -39631 82604 -39605
rect 82658 -39631 82688 -39605
rect 82742 -39631 82772 -39605
rect 82826 -39631 82856 -39605
rect 83038 -39631 83068 -39605
rect 83122 -39631 83152 -39605
rect 83206 -39631 83236 -39605
rect 83290 -39631 83320 -39605
rect 83374 -39631 83404 -39605
rect 83458 -39631 83488 -39605
rect 83542 -39631 83572 -39605
rect 83626 -39631 83656 -39605
rect 83710 -39631 83740 -39605
rect 83794 -39631 83824 -39605
rect 83878 -39631 83908 -39605
rect 83962 -39631 83992 -39605
rect 84046 -39631 84076 -39605
rect 84130 -39631 84160 -39605
rect 84214 -39631 84244 -39605
rect 84298 -39631 84328 -39605
rect 84510 -39631 84540 -39605
rect 84594 -39631 84624 -39605
rect 84678 -39631 84708 -39605
rect 84762 -39631 84792 -39605
rect 84846 -39631 84876 -39605
rect 84930 -39631 84960 -39605
rect 85014 -39631 85044 -39605
rect 85098 -39631 85128 -39605
rect 85182 -39631 85212 -39605
rect 85266 -39631 85296 -39605
rect 85350 -39631 85380 -39605
rect 85434 -39631 85464 -39605
rect 85518 -39631 85548 -39605
rect 85602 -39631 85632 -39605
rect 85686 -39631 85716 -39605
rect 85770 -39631 85800 -39605
rect 85982 -39631 86012 -39605
rect 86066 -39631 86096 -39605
rect 86150 -39631 86180 -39605
rect 86234 -39631 86264 -39605
rect 86318 -39631 86348 -39605
rect 86402 -39631 86432 -39605
rect 86486 -39631 86516 -39605
rect 86570 -39631 86600 -39605
rect 86654 -39631 86684 -39605
rect 86738 -39631 86768 -39605
rect 86822 -39631 86852 -39605
rect 86906 -39631 86936 -39605
rect 86990 -39631 87020 -39605
rect 87074 -39631 87104 -39605
rect 87158 -39631 87188 -39605
rect 87242 -39631 87272 -39605
rect 87454 -39631 87484 -39605
rect 87538 -39631 87568 -39605
rect 87622 -39631 87652 -39605
rect 87706 -39631 87736 -39605
rect 87790 -39631 87820 -39605
rect 87874 -39631 87904 -39605
rect 87958 -39631 87988 -39605
rect 88042 -39631 88072 -39605
rect 88126 -39631 88156 -39605
rect 88210 -39631 88240 -39605
rect 88294 -39631 88324 -39605
rect 88378 -39631 88408 -39605
rect 88462 -39631 88492 -39605
rect 88546 -39631 88576 -39605
rect 88630 -39631 88660 -39605
rect 88714 -39631 88744 -39605
rect 53510 -39906 53630 -39890
rect 53510 -39940 53526 -39906
rect 53614 -39940 53630 -39906
rect 53510 -39978 53630 -39940
rect 53982 -39890 54079 -39874
rect 53982 -39928 53998 -39890
rect 54032 -39928 54079 -39890
rect 53982 -39944 54079 -39928
rect 54879 -39890 54976 -39874
rect 54879 -39928 54926 -39890
rect 54960 -39928 54976 -39890
rect 54879 -39944 54976 -39928
rect 55318 -39968 55384 -39952
rect 55318 -40002 55334 -39968
rect 55368 -40002 55384 -39968
rect 55318 -40018 55384 -40002
rect 55336 -40040 55366 -40018
rect 55336 -40266 55366 -40240
rect 53510 -40816 53630 -40778
rect 53510 -40850 53526 -40816
rect 53614 -40850 53630 -40816
rect 53510 -40866 53630 -40850
rect 53842 -40640 53930 -40624
rect 53842 -40728 53858 -40640
rect 53892 -40728 53930 -40640
rect 53842 -40744 53930 -40728
rect 54730 -40640 54818 -40624
rect 54730 -40728 54768 -40640
rect 54802 -40728 54818 -40640
rect 54730 -40744 54818 -40728
rect 55030 -40559 55096 -40544
rect 55540 -40559 55606 -40544
rect 55030 -40560 55118 -40559
rect 55030 -40594 55046 -40560
rect 55080 -40594 55118 -40560
rect 55030 -40595 55118 -40594
rect 55518 -40560 55606 -40559
rect 55518 -40594 55556 -40560
rect 55590 -40594 55606 -40560
rect 55518 -40595 55606 -40594
rect 55030 -40610 55096 -40595
rect 55540 -40610 55606 -40595
rect 55866 -39856 55986 -39840
rect 55866 -39890 55882 -39856
rect 55970 -39890 55986 -39856
rect 55866 -39928 55986 -39890
rect 55866 -40766 55986 -40728
rect 55866 -40800 55882 -40766
rect 55970 -40800 55986 -40766
rect 55866 -40816 55986 -40800
rect 57175 -39909 57205 -39883
rect 57263 -39909 57293 -39883
rect 57175 -40082 57205 -40067
rect 57169 -40106 57205 -40082
rect 57169 -40141 57199 -40106
rect 57263 -40128 57293 -40067
rect 77657 -39741 77687 -39715
rect 77753 -39741 77783 -39715
rect 77837 -39741 77867 -39715
rect 77921 -39741 77951 -39715
rect 78019 -39735 78049 -39709
rect 59544 -39893 59610 -39885
rect 59087 -39943 59113 -39893
rect 59513 -39901 59610 -39893
rect 59513 -39935 59560 -39901
rect 59594 -39935 59610 -39901
rect 59513 -39943 59610 -39935
rect 59544 -39951 59610 -39943
rect 59016 -40001 59082 -39993
rect 59016 -40009 59113 -40001
rect 59016 -40043 59032 -40009
rect 59066 -40043 59113 -40009
rect 59016 -40051 59113 -40043
rect 59513 -40051 59539 -40001
rect 59016 -40059 59082 -40051
rect 57123 -40157 57199 -40141
rect 57123 -40191 57133 -40157
rect 57167 -40191 57199 -40157
rect 57123 -40207 57199 -40191
rect 57241 -40144 57295 -40128
rect 57241 -40178 57251 -40144
rect 57285 -40178 57295 -40144
rect 57241 -40194 57295 -40178
rect 77657 -39887 77687 -39825
rect 77753 -39887 77783 -39825
rect 77837 -39840 77867 -39825
rect 77603 -39903 77687 -39887
rect 77603 -39937 77613 -39903
rect 77647 -39937 77687 -39903
rect 77603 -39953 77687 -39937
rect 77729 -39903 77783 -39887
rect 77729 -39937 77739 -39903
rect 77773 -39937 77783 -39903
rect 77729 -39953 77783 -39937
rect 77657 -39985 77687 -39953
rect 77753 -39985 77783 -39953
rect 77825 -39869 77867 -39840
rect 77825 -39870 77866 -39869
rect 77825 -39985 77855 -39870
rect 77921 -39887 77951 -39825
rect 80908 -39775 80938 -39749
rect 78019 -39887 78049 -39865
rect 77905 -39903 77959 -39887
rect 77905 -39937 77915 -39903
rect 77949 -39937 77959 -39903
rect 77905 -39953 77959 -39937
rect 78001 -39903 78056 -39887
rect 78001 -39937 78011 -39903
rect 78045 -39937 78056 -39903
rect 80908 -39927 80938 -39905
rect 78001 -39953 78056 -39937
rect 80852 -39943 80938 -39927
rect 77921 -39985 77951 -39953
rect 78019 -39985 78049 -39953
rect 80852 -39977 80868 -39943
rect 80902 -39977 80938 -39943
rect 57169 -40216 57199 -40207
rect 57169 -40240 57205 -40216
rect 57175 -40255 57205 -40240
rect 57263 -40255 57293 -40194
rect 53510 -40924 53630 -40908
rect 53510 -40958 53526 -40924
rect 53614 -40958 53630 -40924
rect 53510 -40996 53630 -40958
rect 53842 -41046 53930 -41030
rect 53842 -41134 53858 -41046
rect 53892 -41134 53930 -41046
rect 53842 -41150 53930 -41134
rect 54730 -41046 54818 -41030
rect 54730 -41134 54768 -41046
rect 54802 -41134 54818 -41046
rect 54730 -41150 54818 -41134
rect 55030 -41181 55096 -41166
rect 55540 -41181 55606 -41166
rect 55030 -41182 55118 -41181
rect 55030 -41216 55046 -41182
rect 55080 -41216 55118 -41182
rect 55030 -41217 55118 -41216
rect 55518 -41182 55606 -41181
rect 55518 -41216 55556 -41182
rect 55590 -41216 55606 -41182
rect 55518 -41217 55606 -41216
rect 55030 -41232 55096 -41217
rect 53510 -41834 53630 -41796
rect 53510 -41868 53526 -41834
rect 53614 -41868 53630 -41834
rect 53510 -41884 53630 -41868
rect 55540 -41232 55606 -41217
rect 53972 -41850 54069 -41834
rect 53972 -41888 53988 -41850
rect 54022 -41888 54069 -41850
rect 53972 -41904 54069 -41888
rect 54869 -41850 54966 -41834
rect 54869 -41888 54916 -41850
rect 54950 -41888 54966 -41850
rect 54869 -41904 54966 -41888
rect 55326 -41536 55356 -41510
rect 55326 -41758 55356 -41736
rect 55308 -41774 55374 -41758
rect 55308 -41808 55324 -41774
rect 55358 -41808 55374 -41774
rect 55308 -41824 55374 -41808
rect 55866 -40970 55986 -40954
rect 55866 -41004 55882 -40970
rect 55970 -41004 55986 -40970
rect 55866 -41042 55986 -41004
rect 55866 -41880 55986 -41842
rect 55866 -41914 55882 -41880
rect 55970 -41914 55986 -41880
rect 55866 -41930 55986 -41914
rect 56476 -40406 56546 -40390
rect 56476 -40440 56492 -40406
rect 56530 -40440 56546 -40406
rect 56476 -40487 56546 -40440
rect 57175 -40385 57205 -40359
rect 57263 -40385 57293 -40359
rect 56476 -41334 56546 -41287
rect 56476 -41368 56492 -41334
rect 56530 -41368 56546 -41334
rect 56476 -41384 56546 -41368
rect 59087 -40278 59153 -40262
rect 59087 -40312 59103 -40278
rect 59137 -40312 59153 -40278
rect 59087 -40328 59153 -40312
rect 59090 -40359 59150 -40328
rect 59090 -40790 59150 -40759
rect 59087 -40806 59153 -40790
rect 59087 -40840 59103 -40806
rect 59137 -40840 59153 -40806
rect 59087 -40856 59153 -40840
rect 77657 -40095 77687 -40069
rect 77753 -40095 77783 -40069
rect 77825 -40117 77855 -40069
rect 77921 -40095 77951 -40069
rect 59858 -40220 59924 -40212
rect 60368 -40220 60434 -40212
rect 59858 -40228 59946 -40220
rect 59858 -40262 59874 -40228
rect 59908 -40262 59946 -40228
rect 59858 -40270 59946 -40262
rect 60346 -40228 60434 -40220
rect 60346 -40262 60384 -40228
rect 60418 -40262 60434 -40228
rect 60346 -40270 60434 -40262
rect 59858 -40278 59924 -40270
rect 60368 -40278 60434 -40270
rect 77819 -40127 77885 -40117
rect 77819 -40161 77835 -40127
rect 77869 -40161 77885 -40127
rect 77819 -40171 77885 -40161
rect 80852 -39993 80938 -39977
rect 80908 -40025 80938 -39993
rect 78019 -40211 78049 -40185
rect 77885 -40355 77915 -40329
rect 80908 -40251 80938 -40225
rect 77693 -40397 77723 -40371
rect 77777 -40397 77807 -40371
rect 59530 -40498 59596 -40482
rect 59530 -40532 59546 -40498
rect 59580 -40532 59596 -40498
rect 59530 -40548 59596 -40532
rect 59548 -40570 59578 -40548
rect 59548 -40792 59578 -40770
rect 59530 -40808 59596 -40792
rect 59530 -40842 59546 -40808
rect 59580 -40842 59596 -40808
rect 59530 -40858 59596 -40842
rect 59846 -40498 59912 -40482
rect 59846 -40532 59862 -40498
rect 59896 -40532 59912 -40498
rect 59846 -40548 59912 -40532
rect 59864 -40570 59894 -40548
rect 59864 -40792 59894 -40770
rect 59846 -40808 59912 -40792
rect 59846 -40842 59862 -40808
rect 59896 -40842 59912 -40808
rect 59846 -40858 59912 -40842
rect 77693 -40587 77723 -40481
rect 77636 -40603 77723 -40587
rect 77636 -40637 77652 -40603
rect 77686 -40637 77723 -40603
rect 77636 -40653 77723 -40637
rect 77693 -40693 77723 -40653
rect 77777 -40587 77807 -40481
rect 77885 -40587 77915 -40555
rect 77777 -40603 77843 -40587
rect 77777 -40637 77793 -40603
rect 77827 -40637 77843 -40603
rect 77777 -40653 77843 -40637
rect 77885 -40603 77951 -40587
rect 77885 -40637 77901 -40603
rect 77935 -40637 77951 -40603
rect 77885 -40653 77951 -40637
rect 77777 -40693 77807 -40653
rect 77885 -40675 77915 -40653
rect 60343 -40765 60409 -40749
rect 61043 -40765 61109 -40749
rect 60343 -40799 60359 -40765
rect 60393 -40799 60409 -40765
rect 60343 -40817 60409 -40799
rect 61043 -40799 61059 -40765
rect 61093 -40799 61109 -40765
rect 61043 -40817 61109 -40799
rect 60165 -40847 60191 -40817
rect 60321 -40847 60441 -40817
rect 60641 -40847 60667 -40817
rect 60785 -40847 60811 -40817
rect 61011 -40847 61131 -40817
rect 61261 -40847 61287 -40817
rect 77693 -40803 77723 -40777
rect 77777 -40803 77807 -40777
rect 77885 -40831 77915 -40805
rect 60343 -40857 60409 -40847
rect 60343 -40891 60359 -40857
rect 60393 -40891 60409 -40857
rect 60343 -40901 60409 -40891
rect 61043 -40857 61109 -40847
rect 61043 -40891 61059 -40857
rect 61093 -40891 61109 -40857
rect 61043 -40901 61109 -40891
rect 57175 -41429 57205 -41403
rect 57263 -41429 57293 -41403
rect 57175 -41548 57205 -41533
rect 57169 -41572 57205 -41548
rect 57169 -41581 57199 -41572
rect 57123 -41597 57199 -41581
rect 57263 -41594 57293 -41533
rect 59087 -41008 59153 -40992
rect 59087 -41042 59103 -41008
rect 59137 -41042 59153 -41008
rect 59087 -41058 59153 -41042
rect 59090 -41089 59150 -41058
rect 59090 -41520 59150 -41489
rect 57123 -41631 57133 -41597
rect 57167 -41631 57199 -41597
rect 57123 -41647 57199 -41631
rect 57169 -41682 57199 -41647
rect 57241 -41610 57295 -41594
rect 57241 -41644 57251 -41610
rect 57285 -41644 57295 -41610
rect 57241 -41660 57295 -41644
rect 59087 -41536 59153 -41520
rect 59087 -41570 59103 -41536
rect 59137 -41570 59153 -41536
rect 59087 -41586 59153 -41570
rect 60165 -40931 60191 -40901
rect 60321 -40931 60441 -40901
rect 60641 -40931 60667 -40901
rect 60785 -40931 60811 -40901
rect 61011 -40931 61131 -40901
rect 61261 -40931 61287 -40901
rect 59526 -41011 59596 -40980
rect 59526 -41030 59545 -41011
rect 59529 -41045 59545 -41030
rect 59579 -41030 59596 -41011
rect 59579 -41045 59595 -41030
rect 59529 -41061 59595 -41045
rect 59547 -41083 59577 -41061
rect 59547 -41305 59577 -41283
rect 59529 -41321 59595 -41305
rect 59529 -41355 59545 -41321
rect 59579 -41355 59595 -41321
rect 59529 -41371 59595 -41355
rect 59845 -41011 59911 -40995
rect 59845 -41045 59861 -41011
rect 59895 -41045 59911 -41011
rect 59845 -41061 59911 -41045
rect 60343 -40941 60409 -40931
rect 60343 -40975 60359 -40941
rect 60393 -40975 60409 -40941
rect 60343 -40985 60409 -40975
rect 61043 -40941 61109 -40931
rect 61043 -40975 61059 -40941
rect 61093 -40975 61109 -40941
rect 61043 -40985 61109 -40975
rect 77885 -40975 77915 -40949
rect 59863 -41083 59893 -41061
rect 59863 -41305 59893 -41283
rect 59845 -41321 59911 -41305
rect 59845 -41355 59861 -41321
rect 59895 -41355 59911 -41321
rect 59845 -41371 59911 -41355
rect 60165 -41015 60191 -40985
rect 60321 -41015 60441 -40985
rect 60641 -41015 60667 -40985
rect 60785 -41015 60811 -40985
rect 61011 -41015 61131 -40985
rect 61261 -41015 61287 -40985
rect 60343 -41025 60409 -41015
rect 60343 -41059 60359 -41025
rect 60393 -41059 60409 -41025
rect 60343 -41069 60409 -41059
rect 61043 -41025 61109 -41015
rect 61043 -41059 61059 -41025
rect 61093 -41059 61109 -41025
rect 61043 -41069 61109 -41059
rect 77693 -41003 77723 -40977
rect 77777 -41003 77807 -40977
rect 60165 -41099 60191 -41069
rect 60321 -41099 60441 -41069
rect 60641 -41099 60667 -41069
rect 60785 -41099 60811 -41069
rect 61011 -41099 61131 -41069
rect 61261 -41099 61287 -41069
rect 77693 -41127 77723 -41087
rect 77636 -41143 77723 -41127
rect 77636 -41177 77652 -41143
rect 77686 -41177 77723 -41143
rect 77636 -41193 77723 -41177
rect 77693 -41299 77723 -41193
rect 77777 -41127 77807 -41087
rect 78117 -40981 78147 -40955
rect 78213 -40981 78243 -40955
rect 78297 -40981 78327 -40955
rect 78381 -40981 78411 -40955
rect 78479 -40975 78509 -40949
rect 77885 -41127 77915 -41105
rect 78117 -41127 78147 -41065
rect 78213 -41127 78243 -41065
rect 78297 -41080 78327 -41065
rect 77777 -41143 77843 -41127
rect 77777 -41177 77793 -41143
rect 77827 -41177 77843 -41143
rect 77777 -41193 77843 -41177
rect 77885 -41143 77951 -41127
rect 77885 -41177 77901 -41143
rect 77935 -41177 77951 -41143
rect 77885 -41193 77951 -41177
rect 78063 -41143 78147 -41127
rect 78063 -41177 78073 -41143
rect 78107 -41177 78147 -41143
rect 78063 -41193 78147 -41177
rect 78189 -41143 78243 -41127
rect 78189 -41177 78199 -41143
rect 78233 -41177 78243 -41143
rect 78189 -41193 78243 -41177
rect 77777 -41299 77807 -41193
rect 77885 -41225 77915 -41193
rect 78117 -41225 78147 -41193
rect 78213 -41225 78243 -41193
rect 78285 -41109 78327 -41080
rect 78285 -41110 78326 -41109
rect 78285 -41225 78315 -41110
rect 78381 -41127 78411 -41065
rect 78479 -41127 78509 -41105
rect 78365 -41143 78419 -41127
rect 78365 -41177 78375 -41143
rect 78409 -41177 78419 -41143
rect 78365 -41193 78419 -41177
rect 78461 -41143 78516 -41127
rect 78461 -41177 78471 -41143
rect 78505 -41177 78516 -41143
rect 78461 -41193 78516 -41177
rect 78381 -41225 78411 -41193
rect 78479 -41225 78509 -41193
rect 77693 -41409 77723 -41383
rect 77777 -41409 77807 -41383
rect 78117 -41335 78147 -41309
rect 78213 -41335 78243 -41309
rect 78285 -41357 78315 -41309
rect 78381 -41335 78411 -41309
rect 78279 -41367 78345 -41357
rect 78279 -41401 78295 -41367
rect 78329 -41401 78345 -41367
rect 78279 -41411 78345 -41401
rect 77885 -41451 77915 -41425
rect 78479 -41451 78509 -41425
rect 57169 -41706 57205 -41682
rect 57175 -41721 57205 -41706
rect 57263 -41721 57293 -41660
rect 57175 -41905 57205 -41879
rect 57263 -41905 57293 -41879
rect 59544 -41800 59610 -41792
rect 59087 -41850 59113 -41800
rect 59513 -41808 59610 -41800
rect 59513 -41842 59560 -41808
rect 59594 -41842 59610 -41808
rect 59513 -41850 59610 -41842
rect 59544 -41858 59610 -41850
rect 59016 -41908 59082 -41900
rect 59016 -41916 59113 -41908
rect 59016 -41950 59032 -41916
rect 59066 -41950 59113 -41916
rect 59016 -41958 59113 -41950
rect 59513 -41958 59539 -41908
rect 59016 -41966 59082 -41958
rect 53972 -42206 54069 -42190
rect 53972 -42244 53988 -42206
rect 54022 -42244 54069 -42206
rect 53972 -42260 54069 -42244
rect 54869 -42206 54966 -42190
rect 54869 -42244 54916 -42206
rect 54950 -42244 54966 -42206
rect 54869 -42260 54966 -42244
rect 59858 -41586 59924 -41578
rect 60368 -41586 60434 -41578
rect 59858 -41594 59946 -41586
rect 59858 -41628 59874 -41594
rect 59908 -41628 59946 -41594
rect 59858 -41636 59946 -41628
rect 60346 -41594 60434 -41586
rect 60346 -41628 60384 -41594
rect 60418 -41628 60434 -41594
rect 60346 -41636 60434 -41628
rect 59858 -41644 59924 -41636
rect 60368 -41644 60434 -41636
rect 77885 -41595 77915 -41569
rect 77693 -41637 77723 -41611
rect 77777 -41637 77807 -41611
rect 77693 -41827 77723 -41721
rect 77636 -41843 77723 -41827
rect 77636 -41877 77652 -41843
rect 77686 -41877 77723 -41843
rect 77636 -41893 77723 -41877
rect 77693 -41933 77723 -41893
rect 77777 -41827 77807 -41721
rect 77885 -41827 77915 -41795
rect 77777 -41843 77843 -41827
rect 77777 -41877 77793 -41843
rect 77827 -41877 77843 -41843
rect 77777 -41893 77843 -41877
rect 77885 -41843 77951 -41827
rect 77885 -41877 77901 -41843
rect 77935 -41877 77951 -41843
rect 77885 -41893 77951 -41877
rect 77777 -41933 77807 -41893
rect 77885 -41915 77915 -41893
rect 77693 -42043 77723 -42017
rect 77777 -42043 77807 -42017
rect 77885 -42071 77915 -42045
rect 77887 -42229 77917 -42203
rect 77695 -42257 77725 -42231
rect 77779 -42257 77809 -42231
rect 55510 -42402 55576 -42386
rect 55510 -42404 55526 -42402
rect 55262 -42434 55288 -42404
rect 55488 -42434 55526 -42404
rect 55510 -42436 55526 -42434
rect 55560 -42436 55576 -42402
rect 55510 -42452 55576 -42436
rect 77695 -42381 77725 -42341
rect 77638 -42397 77725 -42381
rect 77638 -42431 77654 -42397
rect 77688 -42431 77725 -42397
rect 77638 -42447 77725 -42431
rect 77695 -42553 77725 -42447
rect 77779 -42381 77809 -42341
rect 77887 -42381 77917 -42359
rect 77779 -42397 77845 -42381
rect 77779 -42431 77795 -42397
rect 77829 -42431 77845 -42397
rect 77779 -42447 77845 -42431
rect 77887 -42397 77953 -42381
rect 77887 -42431 77903 -42397
rect 77937 -42431 77953 -42397
rect 77887 -42447 77953 -42431
rect 77779 -42553 77809 -42447
rect 77887 -42479 77917 -42447
rect 77695 -42663 77725 -42637
rect 77779 -42663 77809 -42637
rect 77887 -42705 77917 -42679
rect 77657 -42845 77687 -42819
rect 77757 -42845 77787 -42819
rect 77861 -42845 77891 -42819
rect 77947 -42845 77977 -42819
rect 78113 -42845 78143 -42819
rect 78763 -42845 78793 -42819
rect 77657 -43077 77687 -42929
rect 77757 -43077 77787 -42929
rect 77861 -43077 77891 -42929
rect 77947 -43077 77977 -42929
rect 78563 -42869 78629 -42859
rect 78563 -42903 78579 -42869
rect 78613 -42903 78629 -42869
rect 78563 -42913 78629 -42903
rect 78401 -42961 78431 -42935
rect 78497 -42961 78527 -42935
rect 78569 -42961 78599 -42913
rect 78665 -42961 78695 -42935
rect 78113 -43077 78143 -43045
rect 78401 -43077 78431 -43045
rect 78497 -43077 78527 -43045
rect 77599 -43093 77687 -43077
rect 77599 -43127 77609 -43093
rect 77643 -43127 77687 -43093
rect 77599 -43143 77687 -43127
rect 77657 -43211 77687 -43143
rect 77745 -43093 77799 -43077
rect 77745 -43127 77755 -43093
rect 77789 -43127 77799 -43093
rect 77745 -43143 77799 -43127
rect 77851 -43093 77905 -43077
rect 77851 -43127 77861 -43093
rect 77895 -43127 77905 -43093
rect 77851 -43143 77905 -43127
rect 77947 -43093 78011 -43077
rect 77947 -43127 77957 -43093
rect 77991 -43127 78011 -43093
rect 77947 -43143 78011 -43127
rect 78058 -43093 78143 -43077
rect 78058 -43127 78068 -43093
rect 78102 -43127 78143 -43093
rect 78058 -43143 78143 -43127
rect 78347 -43093 78431 -43077
rect 78347 -43127 78357 -43093
rect 78391 -43127 78431 -43093
rect 78347 -43143 78431 -43127
rect 78473 -43093 78527 -43077
rect 78473 -43127 78483 -43093
rect 78517 -43127 78527 -43093
rect 78473 -43143 78527 -43127
rect 77745 -43211 77775 -43143
rect 77851 -43211 77881 -43143
rect 77947 -43211 77977 -43143
rect 78113 -43165 78143 -43143
rect 78401 -43205 78431 -43143
rect 78497 -43205 78527 -43143
rect 78569 -43160 78599 -43045
rect 78665 -43077 78695 -43045
rect 78763 -43077 78793 -43045
rect 78649 -43093 78703 -43077
rect 78649 -43127 78659 -43093
rect 78693 -43127 78703 -43093
rect 78649 -43143 78703 -43127
rect 78745 -43093 78800 -43077
rect 78745 -43127 78755 -43093
rect 78789 -43127 78800 -43093
rect 78745 -43143 78800 -43127
rect 78569 -43161 78610 -43160
rect 78569 -43190 78611 -43161
rect 78581 -43205 78611 -43190
rect 78665 -43205 78695 -43143
rect 78763 -43165 78793 -43143
rect 77657 -43321 77687 -43295
rect 77745 -43321 77775 -43295
rect 77851 -43321 77881 -43295
rect 77947 -43321 77977 -43295
rect 78113 -43321 78143 -43295
rect 78401 -43315 78431 -43289
rect 78497 -43315 78527 -43289
rect 78581 -43315 78611 -43289
rect 78665 -43315 78695 -43289
rect 78763 -43321 78793 -43295
rect 77657 -43461 77687 -43435
rect 77745 -43461 77775 -43435
rect 77851 -43461 77881 -43435
rect 77947 -43461 77977 -43435
rect 78113 -43461 78143 -43435
rect 77657 -43613 77687 -43545
rect 77599 -43629 77687 -43613
rect 77599 -43663 77609 -43629
rect 77643 -43663 77687 -43629
rect 77599 -43679 77687 -43663
rect 77745 -43613 77775 -43545
rect 77851 -43613 77881 -43545
rect 77947 -43613 77977 -43545
rect 78113 -43613 78143 -43591
rect 77745 -43629 77799 -43613
rect 77745 -43663 77755 -43629
rect 77789 -43663 77799 -43629
rect 77745 -43679 77799 -43663
rect 77851 -43629 77905 -43613
rect 77851 -43663 77861 -43629
rect 77895 -43663 77905 -43629
rect 77851 -43679 77905 -43663
rect 77947 -43629 78011 -43613
rect 77947 -43663 77957 -43629
rect 77991 -43663 78011 -43629
rect 77947 -43679 78011 -43663
rect 78058 -43629 78143 -43613
rect 78058 -43663 78068 -43629
rect 78102 -43663 78143 -43629
rect 83127 -43655 83157 -43629
rect 83418 -43655 83448 -43629
rect 83663 -43655 83693 -43629
rect 83747 -43655 83777 -43629
rect 83831 -43655 83861 -43629
rect 83915 -43655 83945 -43629
rect 84126 -43655 84156 -43629
rect 84210 -43655 84240 -43629
rect 84294 -43655 84324 -43629
rect 84378 -43655 84408 -43629
rect 84462 -43655 84492 -43629
rect 84546 -43655 84576 -43629
rect 84630 -43655 84660 -43629
rect 84714 -43655 84744 -43629
rect 84798 -43655 84828 -43629
rect 84882 -43655 84912 -43629
rect 84966 -43655 84996 -43629
rect 85050 -43655 85080 -43629
rect 85134 -43655 85164 -43629
rect 85218 -43655 85248 -43629
rect 85302 -43655 85332 -43629
rect 85386 -43655 85416 -43629
rect 85598 -43655 85628 -43629
rect 85682 -43655 85712 -43629
rect 85766 -43655 85796 -43629
rect 85850 -43655 85880 -43629
rect 85934 -43655 85964 -43629
rect 86018 -43655 86048 -43629
rect 86102 -43655 86132 -43629
rect 86186 -43655 86216 -43629
rect 86270 -43655 86300 -43629
rect 86354 -43655 86384 -43629
rect 86438 -43655 86468 -43629
rect 86522 -43655 86552 -43629
rect 86606 -43655 86636 -43629
rect 86690 -43655 86720 -43629
rect 86774 -43655 86804 -43629
rect 86858 -43655 86888 -43629
rect 87070 -43655 87100 -43629
rect 87154 -43655 87184 -43629
rect 87238 -43655 87268 -43629
rect 87322 -43655 87352 -43629
rect 87406 -43655 87436 -43629
rect 87490 -43655 87520 -43629
rect 87574 -43655 87604 -43629
rect 87658 -43655 87688 -43629
rect 87742 -43655 87772 -43629
rect 87826 -43655 87856 -43629
rect 87910 -43655 87940 -43629
rect 87994 -43655 88024 -43629
rect 88078 -43655 88108 -43629
rect 88162 -43655 88192 -43629
rect 88246 -43655 88276 -43629
rect 88330 -43655 88360 -43629
rect 88542 -43655 88572 -43629
rect 88626 -43655 88656 -43629
rect 88710 -43655 88740 -43629
rect 88794 -43655 88824 -43629
rect 88878 -43655 88908 -43629
rect 88962 -43655 88992 -43629
rect 89046 -43655 89076 -43629
rect 89130 -43655 89160 -43629
rect 89214 -43655 89244 -43629
rect 89298 -43655 89328 -43629
rect 89382 -43655 89412 -43629
rect 89466 -43655 89496 -43629
rect 89550 -43655 89580 -43629
rect 89634 -43655 89664 -43629
rect 89718 -43655 89748 -43629
rect 89802 -43655 89832 -43629
rect 90014 -43655 90044 -43629
rect 90098 -43655 90128 -43629
rect 90182 -43655 90212 -43629
rect 90266 -43655 90296 -43629
rect 90350 -43655 90380 -43629
rect 90434 -43655 90464 -43629
rect 90518 -43655 90548 -43629
rect 90602 -43655 90632 -43629
rect 90686 -43655 90716 -43629
rect 90770 -43655 90800 -43629
rect 90854 -43655 90884 -43629
rect 90938 -43655 90968 -43629
rect 91022 -43655 91052 -43629
rect 91106 -43655 91136 -43629
rect 91190 -43655 91220 -43629
rect 91274 -43655 91304 -43629
rect 78058 -43679 78143 -43663
rect 77657 -43827 77687 -43679
rect 77757 -43827 77787 -43679
rect 77861 -43827 77891 -43679
rect 77947 -43827 77977 -43679
rect 78113 -43711 78143 -43679
rect 82958 -43771 82988 -43745
rect 83030 -43771 83060 -43745
rect 82958 -43887 82988 -43855
rect 82888 -43903 82988 -43887
rect 77657 -43937 77687 -43911
rect 77757 -43937 77787 -43911
rect 77861 -43937 77891 -43911
rect 77947 -43937 77977 -43911
rect 78113 -43937 78143 -43911
rect 82888 -43937 82904 -43903
rect 82938 -43937 82988 -43903
rect 82888 -43953 82988 -43937
rect 83030 -43887 83060 -43855
rect 83127 -43887 83157 -43855
rect 83418 -43887 83448 -43855
rect 83663 -43887 83693 -43855
rect 83747 -43887 83777 -43855
rect 83831 -43887 83861 -43855
rect 83915 -43887 83945 -43855
rect 84126 -43887 84156 -43855
rect 84210 -43887 84240 -43855
rect 84294 -43887 84324 -43855
rect 84378 -43887 84408 -43855
rect 84462 -43887 84492 -43855
rect 84546 -43887 84576 -43855
rect 84630 -43887 84660 -43855
rect 84714 -43887 84744 -43855
rect 84798 -43887 84828 -43855
rect 84882 -43887 84912 -43855
rect 84966 -43887 84996 -43855
rect 85050 -43887 85080 -43855
rect 85134 -43887 85164 -43855
rect 85218 -43887 85248 -43855
rect 85302 -43887 85332 -43855
rect 85386 -43887 85416 -43855
rect 85598 -43887 85628 -43855
rect 85682 -43887 85712 -43855
rect 85766 -43887 85796 -43855
rect 85850 -43887 85880 -43855
rect 85934 -43887 85964 -43855
rect 86018 -43887 86048 -43855
rect 86102 -43887 86132 -43855
rect 86186 -43887 86216 -43855
rect 86270 -43887 86300 -43855
rect 86354 -43887 86384 -43855
rect 86438 -43887 86468 -43855
rect 86522 -43887 86552 -43855
rect 86606 -43887 86636 -43855
rect 86690 -43887 86720 -43855
rect 86774 -43887 86804 -43855
rect 86858 -43887 86888 -43855
rect 87070 -43887 87100 -43855
rect 87154 -43887 87184 -43855
rect 87238 -43887 87268 -43855
rect 87322 -43887 87352 -43855
rect 87406 -43887 87436 -43855
rect 87490 -43887 87520 -43855
rect 87574 -43887 87604 -43855
rect 87658 -43887 87688 -43855
rect 87742 -43887 87772 -43855
rect 87826 -43887 87856 -43855
rect 87910 -43887 87940 -43855
rect 87994 -43887 88024 -43855
rect 88078 -43887 88108 -43855
rect 88162 -43887 88192 -43855
rect 88246 -43887 88276 -43855
rect 88330 -43887 88360 -43855
rect 88542 -43887 88572 -43855
rect 88626 -43887 88656 -43855
rect 88710 -43887 88740 -43855
rect 88794 -43887 88824 -43855
rect 88878 -43887 88908 -43855
rect 88962 -43887 88992 -43855
rect 89046 -43887 89076 -43855
rect 89130 -43887 89160 -43855
rect 89214 -43887 89244 -43855
rect 89298 -43887 89328 -43855
rect 89382 -43887 89412 -43855
rect 89466 -43887 89496 -43855
rect 89550 -43887 89580 -43855
rect 89634 -43887 89664 -43855
rect 89718 -43887 89748 -43855
rect 89802 -43887 89832 -43855
rect 90014 -43887 90044 -43855
rect 90098 -43887 90128 -43855
rect 90182 -43887 90212 -43855
rect 90266 -43887 90296 -43855
rect 90350 -43887 90380 -43855
rect 90434 -43887 90464 -43855
rect 90518 -43887 90548 -43855
rect 90602 -43887 90632 -43855
rect 90686 -43887 90716 -43855
rect 90770 -43887 90800 -43855
rect 90854 -43887 90884 -43855
rect 90938 -43887 90968 -43855
rect 91022 -43887 91052 -43855
rect 91106 -43887 91136 -43855
rect 91190 -43887 91220 -43855
rect 91274 -43887 91304 -43855
rect 83030 -43903 83084 -43887
rect 83030 -43937 83040 -43903
rect 83074 -43937 83084 -43903
rect 83030 -43953 83084 -43937
rect 83127 -43903 83193 -43887
rect 83127 -43937 83143 -43903
rect 83177 -43937 83193 -43903
rect 83127 -43953 83193 -43937
rect 83362 -43903 83448 -43887
rect 83362 -43937 83378 -43903
rect 83412 -43937 83448 -43903
rect 83362 -43953 83448 -43937
rect 83595 -43903 83945 -43887
rect 83595 -43937 83611 -43903
rect 83645 -43937 83703 -43903
rect 83737 -43937 83787 -43903
rect 83821 -43937 83871 -43903
rect 83905 -43937 83945 -43903
rect 83595 -43953 83945 -43937
rect 84060 -43903 85416 -43887
rect 84060 -43937 84076 -43903
rect 84110 -43937 84250 -43903
rect 84284 -43937 84418 -43903
rect 84452 -43937 84587 -43903
rect 84621 -43937 84754 -43903
rect 84788 -43937 84922 -43903
rect 84956 -43937 85089 -43903
rect 85123 -43937 85416 -43903
rect 84060 -43953 85416 -43937
rect 85532 -43903 86888 -43887
rect 85532 -43937 85548 -43903
rect 85582 -43937 85722 -43903
rect 85756 -43937 85890 -43903
rect 85924 -43937 86059 -43903
rect 86093 -43937 86226 -43903
rect 86260 -43937 86394 -43903
rect 86428 -43937 86561 -43903
rect 86595 -43937 86888 -43903
rect 85532 -43953 86888 -43937
rect 87004 -43903 88360 -43887
rect 87004 -43937 87020 -43903
rect 87054 -43937 87194 -43903
rect 87228 -43937 87362 -43903
rect 87396 -43937 87531 -43903
rect 87565 -43937 87698 -43903
rect 87732 -43937 87866 -43903
rect 87900 -43937 88033 -43903
rect 88067 -43937 88360 -43903
rect 87004 -43953 88360 -43937
rect 88476 -43903 89832 -43887
rect 88476 -43937 88492 -43903
rect 88526 -43937 88666 -43903
rect 88700 -43937 88834 -43903
rect 88868 -43937 89003 -43903
rect 89037 -43937 89170 -43903
rect 89204 -43937 89338 -43903
rect 89372 -43937 89505 -43903
rect 89539 -43937 89832 -43903
rect 88476 -43953 89832 -43937
rect 89948 -43903 91304 -43887
rect 89948 -43937 89964 -43903
rect 89998 -43937 90138 -43903
rect 90172 -43937 90306 -43903
rect 90340 -43937 90475 -43903
rect 90509 -43937 90642 -43903
rect 90676 -43937 90810 -43903
rect 90844 -43937 90977 -43903
rect 91011 -43937 91304 -43903
rect 89948 -43953 91304 -43937
rect 82946 -44021 82976 -43953
rect 83030 -44021 83060 -43953
rect 83127 -43975 83157 -43953
rect 83418 -43975 83448 -43953
rect 83663 -43975 83693 -43953
rect 83747 -43975 83777 -43953
rect 83831 -43975 83861 -43953
rect 83915 -43975 83945 -43953
rect 84126 -43975 84156 -43953
rect 84210 -43975 84240 -43953
rect 84294 -43975 84324 -43953
rect 84378 -43975 84408 -43953
rect 84462 -43975 84492 -43953
rect 84546 -43975 84576 -43953
rect 84630 -43975 84660 -43953
rect 84714 -43975 84744 -43953
rect 84798 -43975 84828 -43953
rect 84882 -43975 84912 -43953
rect 84966 -43975 84996 -43953
rect 85050 -43975 85080 -43953
rect 85134 -43975 85164 -43953
rect 85218 -43975 85248 -43953
rect 85302 -43975 85332 -43953
rect 85386 -43975 85416 -43953
rect 85598 -43975 85628 -43953
rect 85682 -43975 85712 -43953
rect 85766 -43975 85796 -43953
rect 85850 -43975 85880 -43953
rect 85934 -43975 85964 -43953
rect 86018 -43975 86048 -43953
rect 86102 -43975 86132 -43953
rect 86186 -43975 86216 -43953
rect 86270 -43975 86300 -43953
rect 86354 -43975 86384 -43953
rect 86438 -43975 86468 -43953
rect 86522 -43975 86552 -43953
rect 86606 -43975 86636 -43953
rect 86690 -43975 86720 -43953
rect 86774 -43975 86804 -43953
rect 86858 -43975 86888 -43953
rect 87070 -43975 87100 -43953
rect 87154 -43975 87184 -43953
rect 87238 -43975 87268 -43953
rect 87322 -43975 87352 -43953
rect 87406 -43975 87436 -43953
rect 87490 -43975 87520 -43953
rect 87574 -43975 87604 -43953
rect 87658 -43975 87688 -43953
rect 87742 -43975 87772 -43953
rect 87826 -43975 87856 -43953
rect 87910 -43975 87940 -43953
rect 87994 -43975 88024 -43953
rect 88078 -43975 88108 -43953
rect 88162 -43975 88192 -43953
rect 88246 -43975 88276 -43953
rect 88330 -43975 88360 -43953
rect 88542 -43975 88572 -43953
rect 88626 -43975 88656 -43953
rect 88710 -43975 88740 -43953
rect 88794 -43975 88824 -43953
rect 88878 -43975 88908 -43953
rect 88962 -43975 88992 -43953
rect 89046 -43975 89076 -43953
rect 89130 -43975 89160 -43953
rect 89214 -43975 89244 -43953
rect 89298 -43975 89328 -43953
rect 89382 -43975 89412 -43953
rect 89466 -43975 89496 -43953
rect 89550 -43975 89580 -43953
rect 89634 -43975 89664 -43953
rect 89718 -43975 89748 -43953
rect 89802 -43975 89832 -43953
rect 90014 -43975 90044 -43953
rect 90098 -43975 90128 -43953
rect 90182 -43975 90212 -43953
rect 90266 -43975 90296 -43953
rect 90350 -43975 90380 -43953
rect 90434 -43975 90464 -43953
rect 90518 -43975 90548 -43953
rect 90602 -43975 90632 -43953
rect 90686 -43975 90716 -43953
rect 90770 -43975 90800 -43953
rect 90854 -43975 90884 -43953
rect 90938 -43975 90968 -43953
rect 91022 -43975 91052 -43953
rect 91106 -43975 91136 -43953
rect 91190 -43975 91220 -43953
rect 91274 -43975 91304 -43953
rect 77657 -44077 77687 -44051
rect 77757 -44077 77787 -44051
rect 77861 -44077 77891 -44051
rect 77947 -44077 77977 -44051
rect 78113 -44077 78143 -44051
rect 77657 -44309 77687 -44161
rect 77757 -44309 77787 -44161
rect 77861 -44309 77891 -44161
rect 77947 -44309 77977 -44161
rect 82946 -44131 82976 -44105
rect 83030 -44131 83060 -44105
rect 83127 -44131 83157 -44105
rect 83418 -44131 83448 -44105
rect 83663 -44131 83693 -44105
rect 83747 -44131 83777 -44105
rect 83831 -44131 83861 -44105
rect 83915 -44131 83945 -44105
rect 84126 -44131 84156 -44105
rect 84210 -44131 84240 -44105
rect 84294 -44131 84324 -44105
rect 84378 -44131 84408 -44105
rect 84462 -44131 84492 -44105
rect 84546 -44131 84576 -44105
rect 84630 -44131 84660 -44105
rect 84714 -44131 84744 -44105
rect 84798 -44131 84828 -44105
rect 84882 -44131 84912 -44105
rect 84966 -44131 84996 -44105
rect 85050 -44131 85080 -44105
rect 85134 -44131 85164 -44105
rect 85218 -44131 85248 -44105
rect 85302 -44131 85332 -44105
rect 85386 -44131 85416 -44105
rect 85598 -44131 85628 -44105
rect 85682 -44131 85712 -44105
rect 85766 -44131 85796 -44105
rect 85850 -44131 85880 -44105
rect 85934 -44131 85964 -44105
rect 86018 -44131 86048 -44105
rect 86102 -44131 86132 -44105
rect 86186 -44131 86216 -44105
rect 86270 -44131 86300 -44105
rect 86354 -44131 86384 -44105
rect 86438 -44131 86468 -44105
rect 86522 -44131 86552 -44105
rect 86606 -44131 86636 -44105
rect 86690 -44131 86720 -44105
rect 86774 -44131 86804 -44105
rect 86858 -44131 86888 -44105
rect 87070 -44131 87100 -44105
rect 87154 -44131 87184 -44105
rect 87238 -44131 87268 -44105
rect 87322 -44131 87352 -44105
rect 87406 -44131 87436 -44105
rect 87490 -44131 87520 -44105
rect 87574 -44131 87604 -44105
rect 87658 -44131 87688 -44105
rect 87742 -44131 87772 -44105
rect 87826 -44131 87856 -44105
rect 87910 -44131 87940 -44105
rect 87994 -44131 88024 -44105
rect 88078 -44131 88108 -44105
rect 88162 -44131 88192 -44105
rect 88246 -44131 88276 -44105
rect 88330 -44131 88360 -44105
rect 88542 -44131 88572 -44105
rect 88626 -44131 88656 -44105
rect 88710 -44131 88740 -44105
rect 88794 -44131 88824 -44105
rect 88878 -44131 88908 -44105
rect 88962 -44131 88992 -44105
rect 89046 -44131 89076 -44105
rect 89130 -44131 89160 -44105
rect 89214 -44131 89244 -44105
rect 89298 -44131 89328 -44105
rect 89382 -44131 89412 -44105
rect 89466 -44131 89496 -44105
rect 89550 -44131 89580 -44105
rect 89634 -44131 89664 -44105
rect 89718 -44131 89748 -44105
rect 89802 -44131 89832 -44105
rect 90014 -44131 90044 -44105
rect 90098 -44131 90128 -44105
rect 90182 -44131 90212 -44105
rect 90266 -44131 90296 -44105
rect 90350 -44131 90380 -44105
rect 90434 -44131 90464 -44105
rect 90518 -44131 90548 -44105
rect 90602 -44131 90632 -44105
rect 90686 -44131 90716 -44105
rect 90770 -44131 90800 -44105
rect 90854 -44131 90884 -44105
rect 90938 -44131 90968 -44105
rect 91022 -44131 91052 -44105
rect 91106 -44131 91136 -44105
rect 91190 -44131 91220 -44105
rect 91274 -44131 91304 -44105
rect 78113 -44309 78143 -44277
rect 77599 -44325 77687 -44309
rect 77599 -44359 77609 -44325
rect 77643 -44359 77687 -44325
rect 77599 -44375 77687 -44359
rect 77657 -44443 77687 -44375
rect 77745 -44325 77799 -44309
rect 77745 -44359 77755 -44325
rect 77789 -44359 77799 -44325
rect 77745 -44375 77799 -44359
rect 77851 -44325 77905 -44309
rect 77851 -44359 77861 -44325
rect 77895 -44359 77905 -44325
rect 77851 -44375 77905 -44359
rect 77947 -44325 78011 -44309
rect 77947 -44359 77957 -44325
rect 77991 -44359 78011 -44325
rect 77947 -44375 78011 -44359
rect 78058 -44325 78143 -44309
rect 78058 -44359 78068 -44325
rect 78102 -44359 78143 -44325
rect 78058 -44375 78143 -44359
rect 77745 -44443 77775 -44375
rect 77851 -44443 77881 -44375
rect 77947 -44443 77977 -44375
rect 78113 -44397 78143 -44375
rect 77657 -44553 77687 -44527
rect 77745 -44553 77775 -44527
rect 77851 -44553 77881 -44527
rect 77947 -44553 77977 -44527
rect 78113 -44553 78143 -44527
rect 77657 -44695 77687 -44669
rect 77745 -44695 77775 -44669
rect 77851 -44695 77881 -44669
rect 77947 -44695 77977 -44669
rect 78113 -44695 78143 -44669
rect 77657 -44847 77687 -44779
rect 53982 -44934 54079 -44918
rect 53982 -44972 53998 -44934
rect 54032 -44972 54079 -44934
rect 53982 -44988 54079 -44972
rect 54879 -44934 54976 -44918
rect 54879 -44972 54926 -44934
rect 54960 -44972 54976 -44934
rect 54879 -44988 54976 -44972
rect 77599 -44863 77687 -44847
rect 77599 -44897 77609 -44863
rect 77643 -44897 77687 -44863
rect 77599 -44913 77687 -44897
rect 77745 -44847 77775 -44779
rect 77851 -44847 77881 -44779
rect 77947 -44847 77977 -44779
rect 78113 -44847 78143 -44825
rect 77745 -44863 77799 -44847
rect 77745 -44897 77755 -44863
rect 77789 -44897 77799 -44863
rect 77745 -44913 77799 -44897
rect 77851 -44863 77905 -44847
rect 77851 -44897 77861 -44863
rect 77895 -44897 77905 -44863
rect 77851 -44913 77905 -44897
rect 77947 -44863 78011 -44847
rect 77947 -44897 77957 -44863
rect 77991 -44897 78011 -44863
rect 77947 -44913 78011 -44897
rect 78058 -44863 78143 -44847
rect 78058 -44897 78068 -44863
rect 78102 -44897 78143 -44863
rect 78058 -44913 78143 -44897
rect 77657 -45061 77687 -44913
rect 77757 -45061 77787 -44913
rect 77861 -45061 77891 -44913
rect 77947 -45061 77977 -44913
rect 78113 -44945 78143 -44913
rect 53510 -45306 53630 -45290
rect 53510 -45340 53526 -45306
rect 53614 -45340 53630 -45306
rect 53510 -45378 53630 -45340
rect 53982 -45290 54079 -45274
rect 53982 -45328 53998 -45290
rect 54032 -45328 54079 -45290
rect 53982 -45344 54079 -45328
rect 54879 -45290 54976 -45274
rect 54879 -45328 54926 -45290
rect 54960 -45328 54976 -45290
rect 54879 -45344 54976 -45328
rect 55318 -45368 55384 -45352
rect 55318 -45402 55334 -45368
rect 55368 -45402 55384 -45368
rect 55318 -45418 55384 -45402
rect 55336 -45440 55366 -45418
rect 55336 -45666 55366 -45640
rect 53510 -46216 53630 -46178
rect 53510 -46250 53526 -46216
rect 53614 -46250 53630 -46216
rect 53510 -46266 53630 -46250
rect 53842 -46040 53930 -46024
rect 53842 -46128 53858 -46040
rect 53892 -46128 53930 -46040
rect 53842 -46144 53930 -46128
rect 54730 -46040 54818 -46024
rect 54730 -46128 54768 -46040
rect 54802 -46128 54818 -46040
rect 54730 -46144 54818 -46128
rect 55030 -45959 55096 -45944
rect 55540 -45959 55606 -45944
rect 55030 -45960 55118 -45959
rect 55030 -45994 55046 -45960
rect 55080 -45994 55118 -45960
rect 55030 -45995 55118 -45994
rect 55518 -45960 55606 -45959
rect 55518 -45994 55556 -45960
rect 55590 -45994 55606 -45960
rect 55518 -45995 55606 -45994
rect 55030 -46010 55096 -45995
rect 55540 -46010 55606 -45995
rect 55866 -45256 55986 -45240
rect 55866 -45290 55882 -45256
rect 55970 -45290 55986 -45256
rect 55866 -45328 55986 -45290
rect 55866 -46166 55986 -46128
rect 55866 -46200 55882 -46166
rect 55970 -46200 55986 -46166
rect 55866 -46216 55986 -46200
rect 57175 -45309 57205 -45283
rect 57263 -45309 57293 -45283
rect 57175 -45482 57205 -45467
rect 57169 -45506 57205 -45482
rect 57169 -45541 57199 -45506
rect 57263 -45528 57293 -45467
rect 77657 -45171 77687 -45145
rect 77757 -45171 77787 -45145
rect 77861 -45171 77891 -45145
rect 77947 -45171 77977 -45145
rect 78113 -45171 78143 -45145
rect 59544 -45293 59610 -45285
rect 59087 -45343 59113 -45293
rect 59513 -45301 59610 -45293
rect 59513 -45335 59560 -45301
rect 59594 -45335 59610 -45301
rect 59513 -45343 59610 -45335
rect 59544 -45351 59610 -45343
rect 59016 -45401 59082 -45393
rect 59016 -45409 59113 -45401
rect 59016 -45443 59032 -45409
rect 59066 -45443 59113 -45409
rect 59016 -45451 59113 -45443
rect 59513 -45451 59539 -45401
rect 59016 -45459 59082 -45451
rect 57123 -45557 57199 -45541
rect 57123 -45591 57133 -45557
rect 57167 -45591 57199 -45557
rect 57123 -45607 57199 -45591
rect 57241 -45544 57295 -45528
rect 57241 -45578 57251 -45544
rect 57285 -45578 57295 -45544
rect 57241 -45594 57295 -45578
rect 77929 -45315 77959 -45289
rect 78345 -45315 78375 -45289
rect 78939 -45315 78969 -45289
rect 77741 -45336 77795 -45320
rect 77741 -45370 77751 -45336
rect 77785 -45370 77795 -45336
rect 77741 -45386 77795 -45370
rect 77657 -45428 77687 -45387
rect 77741 -45428 77771 -45386
rect 77834 -45428 77864 -45402
rect 57169 -45616 57199 -45607
rect 57169 -45640 57205 -45616
rect 57175 -45655 57205 -45640
rect 57263 -45655 57293 -45594
rect 53510 -46324 53630 -46308
rect 53510 -46358 53526 -46324
rect 53614 -46358 53630 -46324
rect 53510 -46396 53630 -46358
rect 53842 -46446 53930 -46430
rect 53842 -46534 53858 -46446
rect 53892 -46534 53930 -46446
rect 53842 -46550 53930 -46534
rect 54730 -46446 54818 -46430
rect 54730 -46534 54768 -46446
rect 54802 -46534 54818 -46446
rect 54730 -46550 54818 -46534
rect 55030 -46581 55096 -46566
rect 55540 -46581 55606 -46566
rect 55030 -46582 55118 -46581
rect 55030 -46616 55046 -46582
rect 55080 -46616 55118 -46582
rect 55030 -46617 55118 -46616
rect 55518 -46582 55606 -46581
rect 55518 -46616 55556 -46582
rect 55590 -46616 55606 -46582
rect 55518 -46617 55606 -46616
rect 55030 -46632 55096 -46617
rect 53510 -47234 53630 -47196
rect 53510 -47268 53526 -47234
rect 53614 -47268 53630 -47234
rect 53510 -47284 53630 -47268
rect 55540 -46632 55606 -46617
rect 53972 -47250 54069 -47234
rect 53972 -47288 53988 -47250
rect 54022 -47288 54069 -47250
rect 53972 -47304 54069 -47288
rect 54869 -47250 54966 -47234
rect 54869 -47288 54916 -47250
rect 54950 -47288 54966 -47250
rect 54869 -47304 54966 -47288
rect 55326 -46936 55356 -46910
rect 55326 -47158 55356 -47136
rect 55308 -47174 55374 -47158
rect 55308 -47208 55324 -47174
rect 55358 -47208 55374 -47174
rect 55308 -47224 55374 -47208
rect 55866 -46370 55986 -46354
rect 55866 -46404 55882 -46370
rect 55970 -46404 55986 -46370
rect 55866 -46442 55986 -46404
rect 55866 -47280 55986 -47242
rect 55866 -47314 55882 -47280
rect 55970 -47314 55986 -47280
rect 55866 -47330 55986 -47314
rect 56476 -45806 56546 -45790
rect 56476 -45840 56492 -45806
rect 56530 -45840 56546 -45806
rect 56476 -45887 56546 -45840
rect 57175 -45785 57205 -45759
rect 57263 -45785 57293 -45759
rect 56476 -46734 56546 -46687
rect 56476 -46768 56492 -46734
rect 56530 -46768 56546 -46734
rect 56476 -46784 56546 -46768
rect 59087 -45678 59153 -45662
rect 59087 -45712 59103 -45678
rect 59137 -45712 59153 -45678
rect 59087 -45728 59153 -45712
rect 59090 -45759 59150 -45728
rect 59090 -46190 59150 -46159
rect 59087 -46206 59153 -46190
rect 59087 -46240 59103 -46206
rect 59137 -46240 59153 -46206
rect 59087 -46256 59153 -46240
rect 59858 -45620 59924 -45612
rect 60368 -45620 60434 -45612
rect 59858 -45628 59946 -45620
rect 59858 -45662 59874 -45628
rect 59908 -45662 59946 -45628
rect 59858 -45670 59946 -45662
rect 60346 -45628 60434 -45620
rect 60346 -45662 60384 -45628
rect 60418 -45662 60434 -45628
rect 60346 -45670 60434 -45662
rect 59858 -45678 59924 -45670
rect 60368 -45678 60434 -45670
rect 77657 -45561 77687 -45512
rect 77741 -45530 77771 -45512
rect 77603 -45609 77687 -45561
rect 77603 -45643 77613 -45609
rect 77647 -45643 77687 -45609
rect 77603 -45666 77687 -45643
rect 77657 -45681 77687 -45666
rect 77729 -45555 77771 -45530
rect 77834 -45553 77864 -45512
rect 78153 -45357 78183 -45331
rect 78237 -45357 78267 -45331
rect 77929 -45547 77959 -45515
rect 78153 -45547 78183 -45441
rect 77729 -45681 77759 -45555
rect 77813 -45569 77867 -45553
rect 77813 -45586 77823 -45569
rect 77801 -45603 77823 -45586
rect 77857 -45603 77867 -45569
rect 77801 -45619 77867 -45603
rect 77909 -45563 77963 -45547
rect 77909 -45597 77919 -45563
rect 77953 -45597 77963 -45563
rect 77909 -45613 77963 -45597
rect 78096 -45563 78183 -45547
rect 78096 -45597 78112 -45563
rect 78146 -45597 78183 -45563
rect 78096 -45613 78183 -45597
rect 77801 -45642 77843 -45619
rect 77929 -45635 77959 -45613
rect 77801 -45666 77838 -45642
rect 77801 -45681 77831 -45666
rect 78153 -45653 78183 -45613
rect 78237 -45547 78267 -45441
rect 78739 -45339 78805 -45329
rect 78739 -45373 78755 -45339
rect 78789 -45373 78805 -45339
rect 78739 -45383 78805 -45373
rect 78577 -45431 78607 -45405
rect 78673 -45431 78703 -45405
rect 78745 -45431 78775 -45383
rect 78841 -45431 78871 -45405
rect 78345 -45547 78375 -45515
rect 78577 -45547 78607 -45515
rect 78673 -45547 78703 -45515
rect 78237 -45563 78303 -45547
rect 78237 -45597 78253 -45563
rect 78287 -45597 78303 -45563
rect 78237 -45613 78303 -45597
rect 78345 -45563 78411 -45547
rect 78345 -45597 78361 -45563
rect 78395 -45597 78411 -45563
rect 78345 -45613 78411 -45597
rect 78523 -45563 78607 -45547
rect 78523 -45597 78533 -45563
rect 78567 -45597 78607 -45563
rect 78523 -45613 78607 -45597
rect 78649 -45563 78703 -45547
rect 78649 -45597 78659 -45563
rect 78693 -45597 78703 -45563
rect 78649 -45613 78703 -45597
rect 78237 -45653 78267 -45613
rect 78345 -45635 78375 -45613
rect 78153 -45763 78183 -45737
rect 78237 -45763 78267 -45737
rect 78577 -45675 78607 -45613
rect 78673 -45675 78703 -45613
rect 78745 -45630 78775 -45515
rect 78841 -45547 78871 -45515
rect 78939 -45547 78969 -45515
rect 78825 -45563 78879 -45547
rect 78825 -45597 78835 -45563
rect 78869 -45597 78879 -45563
rect 78825 -45613 78879 -45597
rect 78921 -45563 78976 -45547
rect 78921 -45597 78931 -45563
rect 78965 -45597 78976 -45563
rect 78921 -45613 78976 -45597
rect 78745 -45631 78786 -45630
rect 78745 -45660 78787 -45631
rect 78757 -45675 78787 -45660
rect 78841 -45675 78871 -45613
rect 78939 -45635 78969 -45613
rect 77657 -45791 77687 -45765
rect 77729 -45791 77759 -45765
rect 77801 -45791 77831 -45765
rect 77929 -45791 77959 -45765
rect 78345 -45791 78375 -45765
rect 78577 -45785 78607 -45759
rect 78673 -45785 78703 -45759
rect 78757 -45785 78787 -45759
rect 78841 -45785 78871 -45759
rect 78939 -45791 78969 -45765
rect 59530 -45898 59596 -45882
rect 59530 -45932 59546 -45898
rect 59580 -45932 59596 -45898
rect 59530 -45948 59596 -45932
rect 59548 -45970 59578 -45948
rect 59548 -46192 59578 -46170
rect 59530 -46208 59596 -46192
rect 59530 -46242 59546 -46208
rect 59580 -46242 59596 -46208
rect 59530 -46258 59596 -46242
rect 59846 -45898 59912 -45882
rect 59846 -45932 59862 -45898
rect 59896 -45932 59912 -45898
rect 59846 -45948 59912 -45932
rect 59864 -45970 59894 -45948
rect 59864 -46192 59894 -46170
rect 59846 -46208 59912 -46192
rect 59846 -46242 59862 -46208
rect 59896 -46242 59912 -46208
rect 59846 -46258 59912 -46242
rect 60343 -46165 60409 -46149
rect 61043 -46165 61109 -46149
rect 60343 -46199 60359 -46165
rect 60393 -46199 60409 -46165
rect 60343 -46217 60409 -46199
rect 61043 -46199 61059 -46165
rect 61093 -46199 61109 -46165
rect 61043 -46217 61109 -46199
rect 60165 -46247 60191 -46217
rect 60321 -46247 60441 -46217
rect 60641 -46247 60667 -46217
rect 60785 -46247 60811 -46217
rect 61011 -46247 61131 -46217
rect 61261 -46247 61287 -46217
rect 60343 -46257 60409 -46247
rect 60343 -46291 60359 -46257
rect 60393 -46291 60409 -46257
rect 60343 -46301 60409 -46291
rect 61043 -46257 61109 -46247
rect 61043 -46291 61059 -46257
rect 61093 -46291 61109 -46257
rect 61043 -46301 61109 -46291
rect 57175 -46829 57205 -46803
rect 57263 -46829 57293 -46803
rect 57175 -46948 57205 -46933
rect 57169 -46972 57205 -46948
rect 57169 -46981 57199 -46972
rect 57123 -46997 57199 -46981
rect 57263 -46994 57293 -46933
rect 59087 -46408 59153 -46392
rect 59087 -46442 59103 -46408
rect 59137 -46442 59153 -46408
rect 59087 -46458 59153 -46442
rect 59090 -46489 59150 -46458
rect 59090 -46920 59150 -46889
rect 57123 -47031 57133 -46997
rect 57167 -47031 57199 -46997
rect 57123 -47047 57199 -47031
rect 57169 -47082 57199 -47047
rect 57241 -47010 57295 -46994
rect 57241 -47044 57251 -47010
rect 57285 -47044 57295 -47010
rect 57241 -47060 57295 -47044
rect 59087 -46936 59153 -46920
rect 59087 -46970 59103 -46936
rect 59137 -46970 59153 -46936
rect 59087 -46986 59153 -46970
rect 60165 -46331 60191 -46301
rect 60321 -46331 60441 -46301
rect 60641 -46331 60667 -46301
rect 60785 -46331 60811 -46301
rect 61011 -46331 61131 -46301
rect 61261 -46331 61287 -46301
rect 59526 -46411 59596 -46380
rect 59526 -46430 59545 -46411
rect 59529 -46445 59545 -46430
rect 59579 -46430 59596 -46411
rect 59579 -46445 59595 -46430
rect 59529 -46461 59595 -46445
rect 59547 -46483 59577 -46461
rect 59547 -46705 59577 -46683
rect 59529 -46721 59595 -46705
rect 59529 -46755 59545 -46721
rect 59579 -46755 59595 -46721
rect 59529 -46771 59595 -46755
rect 59845 -46411 59911 -46395
rect 59845 -46445 59861 -46411
rect 59895 -46445 59911 -46411
rect 59845 -46461 59911 -46445
rect 60343 -46341 60409 -46331
rect 60343 -46375 60359 -46341
rect 60393 -46375 60409 -46341
rect 60343 -46385 60409 -46375
rect 61043 -46341 61109 -46331
rect 61043 -46375 61059 -46341
rect 61093 -46375 61109 -46341
rect 61043 -46385 61109 -46375
rect 59863 -46483 59893 -46461
rect 59863 -46705 59893 -46683
rect 59845 -46721 59911 -46705
rect 59845 -46755 59861 -46721
rect 59895 -46755 59911 -46721
rect 59845 -46771 59911 -46755
rect 60165 -46415 60191 -46385
rect 60321 -46415 60441 -46385
rect 60641 -46415 60667 -46385
rect 60785 -46415 60811 -46385
rect 61011 -46415 61131 -46385
rect 61261 -46415 61287 -46385
rect 60343 -46425 60409 -46415
rect 60343 -46459 60359 -46425
rect 60393 -46459 60409 -46425
rect 60343 -46469 60409 -46459
rect 61043 -46425 61109 -46415
rect 61043 -46459 61059 -46425
rect 61093 -46459 61109 -46425
rect 61043 -46469 61109 -46459
rect 60165 -46499 60191 -46469
rect 60321 -46499 60441 -46469
rect 60641 -46499 60667 -46469
rect 60785 -46499 60811 -46469
rect 61011 -46499 61131 -46469
rect 61261 -46499 61287 -46469
rect 75626 -46475 75656 -46449
rect 75902 -46475 75932 -46449
rect 76176 -46475 76206 -46449
rect 76452 -46475 76482 -46449
rect 76728 -46475 76758 -46449
rect 75626 -46627 75656 -46605
rect 75902 -46627 75932 -46605
rect 76176 -46627 76206 -46605
rect 76452 -46627 76482 -46605
rect 76728 -46627 76758 -46605
rect 75570 -46643 75656 -46627
rect 75570 -46677 75586 -46643
rect 75620 -46677 75656 -46643
rect 75570 -46693 75656 -46677
rect 75846 -46643 75932 -46627
rect 75846 -46677 75862 -46643
rect 75896 -46677 75932 -46643
rect 75846 -46693 75932 -46677
rect 76120 -46643 76206 -46627
rect 76120 -46677 76136 -46643
rect 76170 -46677 76206 -46643
rect 76120 -46693 76206 -46677
rect 76396 -46643 76482 -46627
rect 76396 -46677 76412 -46643
rect 76446 -46677 76482 -46643
rect 76396 -46693 76482 -46677
rect 76672 -46643 76758 -46627
rect 76672 -46677 76688 -46643
rect 76722 -46677 76758 -46643
rect 76672 -46693 76758 -46677
rect 75626 -46725 75656 -46693
rect 75902 -46725 75932 -46693
rect 76176 -46725 76206 -46693
rect 76452 -46725 76482 -46693
rect 76728 -46725 76758 -46693
rect 57169 -47106 57205 -47082
rect 57175 -47121 57205 -47106
rect 57263 -47121 57293 -47060
rect 57175 -47305 57205 -47279
rect 57263 -47305 57293 -47279
rect 59544 -47200 59610 -47192
rect 59087 -47250 59113 -47200
rect 59513 -47208 59610 -47200
rect 59513 -47242 59560 -47208
rect 59594 -47242 59610 -47208
rect 59513 -47250 59610 -47242
rect 59544 -47258 59610 -47250
rect 59016 -47308 59082 -47300
rect 59016 -47316 59113 -47308
rect 59016 -47350 59032 -47316
rect 59066 -47350 59113 -47316
rect 59016 -47358 59113 -47350
rect 59513 -47358 59539 -47308
rect 59016 -47366 59082 -47358
rect 53972 -47606 54069 -47590
rect 53972 -47644 53988 -47606
rect 54022 -47644 54069 -47606
rect 53972 -47660 54069 -47644
rect 54869 -47606 54966 -47590
rect 54869 -47644 54916 -47606
rect 54950 -47644 54966 -47606
rect 54869 -47660 54966 -47644
rect 59858 -46986 59924 -46978
rect 60368 -46986 60434 -46978
rect 59858 -46994 59946 -46986
rect 59858 -47028 59874 -46994
rect 59908 -47028 59946 -46994
rect 59858 -47036 59946 -47028
rect 60346 -46994 60434 -46986
rect 60346 -47028 60384 -46994
rect 60418 -47028 60434 -46994
rect 60346 -47036 60434 -47028
rect 59858 -47044 59924 -47036
rect 60368 -47044 60434 -47036
rect 75626 -46951 75656 -46925
rect 75902 -46951 75932 -46925
rect 76176 -46951 76206 -46925
rect 76452 -46951 76482 -46925
rect 76728 -46951 76758 -46925
rect 78019 -47145 78049 -47119
rect 78477 -47145 78507 -47119
rect 78897 -47145 78927 -47119
rect 77819 -47169 77885 -47159
rect 77819 -47203 77835 -47169
rect 77869 -47203 77885 -47169
rect 77819 -47213 77885 -47203
rect 77657 -47261 77687 -47235
rect 77753 -47261 77783 -47235
rect 77825 -47261 77855 -47213
rect 77921 -47261 77951 -47235
rect 78277 -47169 78343 -47159
rect 78277 -47203 78293 -47169
rect 78327 -47203 78343 -47169
rect 78277 -47213 78343 -47203
rect 78211 -47261 78241 -47235
rect 78283 -47261 78313 -47213
rect 78379 -47261 78409 -47235
rect 78705 -47187 78735 -47161
rect 78789 -47187 78819 -47161
rect 77657 -47377 77687 -47345
rect 77753 -47377 77783 -47345
rect 77603 -47393 77687 -47377
rect 77603 -47427 77613 -47393
rect 77647 -47427 77687 -47393
rect 77603 -47443 77687 -47427
rect 77729 -47393 77783 -47377
rect 77729 -47427 77739 -47393
rect 77773 -47427 77783 -47393
rect 77729 -47443 77783 -47427
rect 77657 -47505 77687 -47443
rect 77753 -47505 77783 -47443
rect 77825 -47460 77855 -47345
rect 77921 -47377 77951 -47345
rect 78019 -47377 78049 -47345
rect 78211 -47377 78241 -47345
rect 77905 -47393 77959 -47377
rect 77905 -47427 77915 -47393
rect 77949 -47427 77959 -47393
rect 77905 -47443 77959 -47427
rect 78001 -47393 78056 -47377
rect 78001 -47427 78011 -47393
rect 78045 -47427 78056 -47393
rect 78001 -47443 78056 -47427
rect 78154 -47393 78241 -47377
rect 78154 -47427 78164 -47393
rect 78198 -47427 78241 -47393
rect 78154 -47443 78241 -47427
rect 77825 -47461 77866 -47460
rect 77825 -47490 77867 -47461
rect 77837 -47505 77867 -47490
rect 77921 -47505 77951 -47443
rect 78019 -47465 78049 -47443
rect 77657 -47615 77687 -47589
rect 77753 -47615 77783 -47589
rect 77837 -47615 77867 -47589
rect 77921 -47615 77951 -47589
rect 78211 -47505 78241 -47443
rect 78283 -47460 78313 -47345
rect 78379 -47377 78409 -47345
rect 78477 -47377 78507 -47345
rect 78705 -47377 78735 -47271
rect 78364 -47393 78418 -47377
rect 78364 -47427 78374 -47393
rect 78408 -47427 78418 -47393
rect 78364 -47443 78418 -47427
rect 78460 -47393 78514 -47377
rect 78460 -47427 78470 -47393
rect 78504 -47427 78514 -47393
rect 78460 -47443 78514 -47427
rect 78648 -47393 78735 -47377
rect 78648 -47427 78664 -47393
rect 78698 -47427 78735 -47393
rect 78648 -47443 78735 -47427
rect 78283 -47490 78325 -47460
rect 78295 -47505 78325 -47490
rect 78379 -47505 78409 -47443
rect 78477 -47465 78507 -47443
rect 78019 -47621 78049 -47595
rect 78211 -47615 78241 -47589
rect 78295 -47615 78325 -47589
rect 78379 -47615 78409 -47589
rect 78705 -47483 78735 -47443
rect 78789 -47377 78819 -47271
rect 78897 -47377 78927 -47345
rect 78789 -47393 78855 -47377
rect 78789 -47427 78805 -47393
rect 78839 -47427 78855 -47393
rect 78789 -47443 78855 -47427
rect 78897 -47393 78963 -47377
rect 78897 -47427 78913 -47393
rect 78947 -47427 78963 -47393
rect 78897 -47443 78963 -47427
rect 78789 -47483 78819 -47443
rect 78897 -47465 78927 -47443
rect 78705 -47593 78735 -47567
rect 78789 -47593 78819 -47567
rect 78477 -47621 78507 -47595
rect 78897 -47621 78927 -47595
rect 55510 -47802 55576 -47786
rect 55510 -47804 55526 -47802
rect 55262 -47834 55288 -47804
rect 55488 -47834 55526 -47804
rect 55510 -47836 55526 -47834
rect 55560 -47836 55576 -47802
rect 55510 -47852 55576 -47836
rect 77657 -47781 77687 -47755
rect 77753 -47781 77783 -47755
rect 77837 -47781 77867 -47755
rect 77921 -47781 77951 -47755
rect 78019 -47775 78049 -47749
rect 77657 -47927 77687 -47865
rect 77753 -47927 77783 -47865
rect 77837 -47880 77867 -47865
rect 77603 -47943 77687 -47927
rect 77603 -47977 77613 -47943
rect 77647 -47977 77687 -47943
rect 77603 -47993 77687 -47977
rect 77729 -47943 77783 -47927
rect 77729 -47977 77739 -47943
rect 77773 -47977 77783 -47943
rect 77729 -47993 77783 -47977
rect 77657 -48025 77687 -47993
rect 77753 -48025 77783 -47993
rect 77825 -47909 77867 -47880
rect 77825 -47910 77866 -47909
rect 77825 -48025 77855 -47910
rect 77921 -47927 77951 -47865
rect 83127 -47795 83157 -47769
rect 83418 -47795 83448 -47769
rect 83663 -47795 83693 -47769
rect 83747 -47795 83777 -47769
rect 83831 -47795 83861 -47769
rect 83915 -47795 83945 -47769
rect 84126 -47795 84156 -47769
rect 84210 -47795 84240 -47769
rect 84294 -47795 84324 -47769
rect 84378 -47795 84408 -47769
rect 84462 -47795 84492 -47769
rect 84546 -47795 84576 -47769
rect 84630 -47795 84660 -47769
rect 84714 -47795 84744 -47769
rect 84798 -47795 84828 -47769
rect 84882 -47795 84912 -47769
rect 84966 -47795 84996 -47769
rect 85050 -47795 85080 -47769
rect 85134 -47795 85164 -47769
rect 85218 -47795 85248 -47769
rect 85302 -47795 85332 -47769
rect 85386 -47795 85416 -47769
rect 85598 -47795 85628 -47769
rect 85682 -47795 85712 -47769
rect 85766 -47795 85796 -47769
rect 85850 -47795 85880 -47769
rect 85934 -47795 85964 -47769
rect 86018 -47795 86048 -47769
rect 86102 -47795 86132 -47769
rect 86186 -47795 86216 -47769
rect 86270 -47795 86300 -47769
rect 86354 -47795 86384 -47769
rect 86438 -47795 86468 -47769
rect 86522 -47795 86552 -47769
rect 86606 -47795 86636 -47769
rect 86690 -47795 86720 -47769
rect 86774 -47795 86804 -47769
rect 86858 -47795 86888 -47769
rect 87070 -47795 87100 -47769
rect 87154 -47795 87184 -47769
rect 87238 -47795 87268 -47769
rect 87322 -47795 87352 -47769
rect 87406 -47795 87436 -47769
rect 87490 -47795 87520 -47769
rect 87574 -47795 87604 -47769
rect 87658 -47795 87688 -47769
rect 87742 -47795 87772 -47769
rect 87826 -47795 87856 -47769
rect 87910 -47795 87940 -47769
rect 87994 -47795 88024 -47769
rect 88078 -47795 88108 -47769
rect 88162 -47795 88192 -47769
rect 88246 -47795 88276 -47769
rect 88330 -47795 88360 -47769
rect 88542 -47795 88572 -47769
rect 88626 -47795 88656 -47769
rect 88710 -47795 88740 -47769
rect 88794 -47795 88824 -47769
rect 88878 -47795 88908 -47769
rect 88962 -47795 88992 -47769
rect 89046 -47795 89076 -47769
rect 89130 -47795 89160 -47769
rect 89214 -47795 89244 -47769
rect 89298 -47795 89328 -47769
rect 89382 -47795 89412 -47769
rect 89466 -47795 89496 -47769
rect 89550 -47795 89580 -47769
rect 89634 -47795 89664 -47769
rect 89718 -47795 89748 -47769
rect 89802 -47795 89832 -47769
rect 90014 -47795 90044 -47769
rect 90098 -47795 90128 -47769
rect 90182 -47795 90212 -47769
rect 90266 -47795 90296 -47769
rect 90350 -47795 90380 -47769
rect 90434 -47795 90464 -47769
rect 90518 -47795 90548 -47769
rect 90602 -47795 90632 -47769
rect 90686 -47795 90716 -47769
rect 90770 -47795 90800 -47769
rect 90854 -47795 90884 -47769
rect 90938 -47795 90968 -47769
rect 91022 -47795 91052 -47769
rect 91106 -47795 91136 -47769
rect 91190 -47795 91220 -47769
rect 91274 -47795 91304 -47769
rect 78019 -47927 78049 -47905
rect 82958 -47911 82988 -47885
rect 83030 -47911 83060 -47885
rect 77905 -47943 77959 -47927
rect 77905 -47977 77915 -47943
rect 77949 -47977 77959 -47943
rect 77905 -47993 77959 -47977
rect 78001 -47943 78056 -47927
rect 78001 -47977 78011 -47943
rect 78045 -47977 78056 -47943
rect 78001 -47993 78056 -47977
rect 77921 -48025 77951 -47993
rect 78019 -48025 78049 -47993
rect 77657 -48135 77687 -48109
rect 77753 -48135 77783 -48109
rect 77825 -48157 77855 -48109
rect 77921 -48135 77951 -48109
rect 77819 -48167 77885 -48157
rect 77819 -48201 77835 -48167
rect 77869 -48201 77885 -48167
rect 77819 -48211 77885 -48201
rect 82958 -48027 82988 -47995
rect 82888 -48043 82988 -48027
rect 82888 -48077 82904 -48043
rect 82938 -48077 82988 -48043
rect 82888 -48093 82988 -48077
rect 83030 -48027 83060 -47995
rect 83127 -48027 83157 -47995
rect 83418 -48027 83448 -47995
rect 83663 -48027 83693 -47995
rect 83747 -48027 83777 -47995
rect 83831 -48027 83861 -47995
rect 83915 -48027 83945 -47995
rect 84126 -48027 84156 -47995
rect 84210 -48027 84240 -47995
rect 84294 -48027 84324 -47995
rect 84378 -48027 84408 -47995
rect 84462 -48027 84492 -47995
rect 84546 -48027 84576 -47995
rect 84630 -48027 84660 -47995
rect 84714 -48027 84744 -47995
rect 84798 -48027 84828 -47995
rect 84882 -48027 84912 -47995
rect 84966 -48027 84996 -47995
rect 85050 -48027 85080 -47995
rect 85134 -48027 85164 -47995
rect 85218 -48027 85248 -47995
rect 85302 -48027 85332 -47995
rect 85386 -48027 85416 -47995
rect 85598 -48027 85628 -47995
rect 85682 -48027 85712 -47995
rect 85766 -48027 85796 -47995
rect 85850 -48027 85880 -47995
rect 85934 -48027 85964 -47995
rect 86018 -48027 86048 -47995
rect 86102 -48027 86132 -47995
rect 86186 -48027 86216 -47995
rect 86270 -48027 86300 -47995
rect 86354 -48027 86384 -47995
rect 86438 -48027 86468 -47995
rect 86522 -48027 86552 -47995
rect 86606 -48027 86636 -47995
rect 86690 -48027 86720 -47995
rect 86774 -48027 86804 -47995
rect 86858 -48027 86888 -47995
rect 87070 -48027 87100 -47995
rect 87154 -48027 87184 -47995
rect 87238 -48027 87268 -47995
rect 87322 -48027 87352 -47995
rect 87406 -48027 87436 -47995
rect 87490 -48027 87520 -47995
rect 87574 -48027 87604 -47995
rect 87658 -48027 87688 -47995
rect 87742 -48027 87772 -47995
rect 87826 -48027 87856 -47995
rect 87910 -48027 87940 -47995
rect 87994 -48027 88024 -47995
rect 88078 -48027 88108 -47995
rect 88162 -48027 88192 -47995
rect 88246 -48027 88276 -47995
rect 88330 -48027 88360 -47995
rect 88542 -48027 88572 -47995
rect 88626 -48027 88656 -47995
rect 88710 -48027 88740 -47995
rect 88794 -48027 88824 -47995
rect 88878 -48027 88908 -47995
rect 88962 -48027 88992 -47995
rect 89046 -48027 89076 -47995
rect 89130 -48027 89160 -47995
rect 89214 -48027 89244 -47995
rect 89298 -48027 89328 -47995
rect 89382 -48027 89412 -47995
rect 89466 -48027 89496 -47995
rect 89550 -48027 89580 -47995
rect 89634 -48027 89664 -47995
rect 89718 -48027 89748 -47995
rect 89802 -48027 89832 -47995
rect 90014 -48027 90044 -47995
rect 90098 -48027 90128 -47995
rect 90182 -48027 90212 -47995
rect 90266 -48027 90296 -47995
rect 90350 -48027 90380 -47995
rect 90434 -48027 90464 -47995
rect 90518 -48027 90548 -47995
rect 90602 -48027 90632 -47995
rect 90686 -48027 90716 -47995
rect 90770 -48027 90800 -47995
rect 90854 -48027 90884 -47995
rect 90938 -48027 90968 -47995
rect 91022 -48027 91052 -47995
rect 91106 -48027 91136 -47995
rect 91190 -48027 91220 -47995
rect 91274 -48027 91304 -47995
rect 83030 -48043 83084 -48027
rect 83030 -48077 83040 -48043
rect 83074 -48077 83084 -48043
rect 83030 -48093 83084 -48077
rect 83127 -48043 83193 -48027
rect 83127 -48077 83143 -48043
rect 83177 -48077 83193 -48043
rect 83127 -48093 83193 -48077
rect 83362 -48043 83448 -48027
rect 83362 -48077 83378 -48043
rect 83412 -48077 83448 -48043
rect 83362 -48093 83448 -48077
rect 83595 -48043 83945 -48027
rect 83595 -48077 83611 -48043
rect 83645 -48077 83703 -48043
rect 83737 -48077 83787 -48043
rect 83821 -48077 83871 -48043
rect 83905 -48077 83945 -48043
rect 83595 -48093 83945 -48077
rect 84060 -48043 85416 -48027
rect 84060 -48077 84076 -48043
rect 84110 -48077 84250 -48043
rect 84284 -48077 84418 -48043
rect 84452 -48077 84587 -48043
rect 84621 -48077 84754 -48043
rect 84788 -48077 84922 -48043
rect 84956 -48077 85089 -48043
rect 85123 -48077 85416 -48043
rect 84060 -48093 85416 -48077
rect 85532 -48043 86888 -48027
rect 85532 -48077 85548 -48043
rect 85582 -48077 85722 -48043
rect 85756 -48077 85890 -48043
rect 85924 -48077 86059 -48043
rect 86093 -48077 86226 -48043
rect 86260 -48077 86394 -48043
rect 86428 -48077 86561 -48043
rect 86595 -48077 86888 -48043
rect 85532 -48093 86888 -48077
rect 87004 -48043 88360 -48027
rect 87004 -48077 87020 -48043
rect 87054 -48077 87194 -48043
rect 87228 -48077 87362 -48043
rect 87396 -48077 87531 -48043
rect 87565 -48077 87698 -48043
rect 87732 -48077 87866 -48043
rect 87900 -48077 88033 -48043
rect 88067 -48077 88360 -48043
rect 87004 -48093 88360 -48077
rect 88476 -48043 89832 -48027
rect 88476 -48077 88492 -48043
rect 88526 -48077 88666 -48043
rect 88700 -48077 88834 -48043
rect 88868 -48077 89003 -48043
rect 89037 -48077 89170 -48043
rect 89204 -48077 89338 -48043
rect 89372 -48077 89505 -48043
rect 89539 -48077 89832 -48043
rect 88476 -48093 89832 -48077
rect 89948 -48043 91304 -48027
rect 89948 -48077 89964 -48043
rect 89998 -48077 90138 -48043
rect 90172 -48077 90306 -48043
rect 90340 -48077 90475 -48043
rect 90509 -48077 90642 -48043
rect 90676 -48077 90810 -48043
rect 90844 -48077 90977 -48043
rect 91011 -48077 91304 -48043
rect 89948 -48093 91304 -48077
rect 82946 -48161 82976 -48093
rect 83030 -48161 83060 -48093
rect 83127 -48115 83157 -48093
rect 83418 -48115 83448 -48093
rect 83663 -48115 83693 -48093
rect 83747 -48115 83777 -48093
rect 83831 -48115 83861 -48093
rect 83915 -48115 83945 -48093
rect 84126 -48115 84156 -48093
rect 84210 -48115 84240 -48093
rect 84294 -48115 84324 -48093
rect 84378 -48115 84408 -48093
rect 84462 -48115 84492 -48093
rect 84546 -48115 84576 -48093
rect 84630 -48115 84660 -48093
rect 84714 -48115 84744 -48093
rect 84798 -48115 84828 -48093
rect 84882 -48115 84912 -48093
rect 84966 -48115 84996 -48093
rect 85050 -48115 85080 -48093
rect 85134 -48115 85164 -48093
rect 85218 -48115 85248 -48093
rect 85302 -48115 85332 -48093
rect 85386 -48115 85416 -48093
rect 85598 -48115 85628 -48093
rect 85682 -48115 85712 -48093
rect 85766 -48115 85796 -48093
rect 85850 -48115 85880 -48093
rect 85934 -48115 85964 -48093
rect 86018 -48115 86048 -48093
rect 86102 -48115 86132 -48093
rect 86186 -48115 86216 -48093
rect 86270 -48115 86300 -48093
rect 86354 -48115 86384 -48093
rect 86438 -48115 86468 -48093
rect 86522 -48115 86552 -48093
rect 86606 -48115 86636 -48093
rect 86690 -48115 86720 -48093
rect 86774 -48115 86804 -48093
rect 86858 -48115 86888 -48093
rect 87070 -48115 87100 -48093
rect 87154 -48115 87184 -48093
rect 87238 -48115 87268 -48093
rect 87322 -48115 87352 -48093
rect 87406 -48115 87436 -48093
rect 87490 -48115 87520 -48093
rect 87574 -48115 87604 -48093
rect 87658 -48115 87688 -48093
rect 87742 -48115 87772 -48093
rect 87826 -48115 87856 -48093
rect 87910 -48115 87940 -48093
rect 87994 -48115 88024 -48093
rect 88078 -48115 88108 -48093
rect 88162 -48115 88192 -48093
rect 88246 -48115 88276 -48093
rect 88330 -48115 88360 -48093
rect 88542 -48115 88572 -48093
rect 88626 -48115 88656 -48093
rect 88710 -48115 88740 -48093
rect 88794 -48115 88824 -48093
rect 88878 -48115 88908 -48093
rect 88962 -48115 88992 -48093
rect 89046 -48115 89076 -48093
rect 89130 -48115 89160 -48093
rect 89214 -48115 89244 -48093
rect 89298 -48115 89328 -48093
rect 89382 -48115 89412 -48093
rect 89466 -48115 89496 -48093
rect 89550 -48115 89580 -48093
rect 89634 -48115 89664 -48093
rect 89718 -48115 89748 -48093
rect 89802 -48115 89832 -48093
rect 90014 -48115 90044 -48093
rect 90098 -48115 90128 -48093
rect 90182 -48115 90212 -48093
rect 90266 -48115 90296 -48093
rect 90350 -48115 90380 -48093
rect 90434 -48115 90464 -48093
rect 90518 -48115 90548 -48093
rect 90602 -48115 90632 -48093
rect 90686 -48115 90716 -48093
rect 90770 -48115 90800 -48093
rect 90854 -48115 90884 -48093
rect 90938 -48115 90968 -48093
rect 91022 -48115 91052 -48093
rect 91106 -48115 91136 -48093
rect 91190 -48115 91220 -48093
rect 91274 -48115 91304 -48093
rect 78019 -48251 78049 -48225
rect 77885 -48395 77915 -48369
rect 82946 -48271 82976 -48245
rect 83030 -48271 83060 -48245
rect 83127 -48271 83157 -48245
rect 83418 -48271 83448 -48245
rect 83663 -48271 83693 -48245
rect 83747 -48271 83777 -48245
rect 83831 -48271 83861 -48245
rect 83915 -48271 83945 -48245
rect 84126 -48271 84156 -48245
rect 84210 -48271 84240 -48245
rect 84294 -48271 84324 -48245
rect 84378 -48271 84408 -48245
rect 84462 -48271 84492 -48245
rect 84546 -48271 84576 -48245
rect 84630 -48271 84660 -48245
rect 84714 -48271 84744 -48245
rect 84798 -48271 84828 -48245
rect 84882 -48271 84912 -48245
rect 84966 -48271 84996 -48245
rect 85050 -48271 85080 -48245
rect 85134 -48271 85164 -48245
rect 85218 -48271 85248 -48245
rect 85302 -48271 85332 -48245
rect 85386 -48271 85416 -48245
rect 85598 -48271 85628 -48245
rect 85682 -48271 85712 -48245
rect 85766 -48271 85796 -48245
rect 85850 -48271 85880 -48245
rect 85934 -48271 85964 -48245
rect 86018 -48271 86048 -48245
rect 86102 -48271 86132 -48245
rect 86186 -48271 86216 -48245
rect 86270 -48271 86300 -48245
rect 86354 -48271 86384 -48245
rect 86438 -48271 86468 -48245
rect 86522 -48271 86552 -48245
rect 86606 -48271 86636 -48245
rect 86690 -48271 86720 -48245
rect 86774 -48271 86804 -48245
rect 86858 -48271 86888 -48245
rect 87070 -48271 87100 -48245
rect 87154 -48271 87184 -48245
rect 87238 -48271 87268 -48245
rect 87322 -48271 87352 -48245
rect 87406 -48271 87436 -48245
rect 87490 -48271 87520 -48245
rect 87574 -48271 87604 -48245
rect 87658 -48271 87688 -48245
rect 87742 -48271 87772 -48245
rect 87826 -48271 87856 -48245
rect 87910 -48271 87940 -48245
rect 87994 -48271 88024 -48245
rect 88078 -48271 88108 -48245
rect 88162 -48271 88192 -48245
rect 88246 -48271 88276 -48245
rect 88330 -48271 88360 -48245
rect 88542 -48271 88572 -48245
rect 88626 -48271 88656 -48245
rect 88710 -48271 88740 -48245
rect 88794 -48271 88824 -48245
rect 88878 -48271 88908 -48245
rect 88962 -48271 88992 -48245
rect 89046 -48271 89076 -48245
rect 89130 -48271 89160 -48245
rect 89214 -48271 89244 -48245
rect 89298 -48271 89328 -48245
rect 89382 -48271 89412 -48245
rect 89466 -48271 89496 -48245
rect 89550 -48271 89580 -48245
rect 89634 -48271 89664 -48245
rect 89718 -48271 89748 -48245
rect 89802 -48271 89832 -48245
rect 90014 -48271 90044 -48245
rect 90098 -48271 90128 -48245
rect 90182 -48271 90212 -48245
rect 90266 -48271 90296 -48245
rect 90350 -48271 90380 -48245
rect 90434 -48271 90464 -48245
rect 90518 -48271 90548 -48245
rect 90602 -48271 90632 -48245
rect 90686 -48271 90716 -48245
rect 90770 -48271 90800 -48245
rect 90854 -48271 90884 -48245
rect 90938 -48271 90968 -48245
rect 91022 -48271 91052 -48245
rect 91106 -48271 91136 -48245
rect 91190 -48271 91220 -48245
rect 91274 -48271 91304 -48245
rect 77693 -48437 77723 -48411
rect 77777 -48437 77807 -48411
rect 77693 -48627 77723 -48521
rect 77636 -48643 77723 -48627
rect 77636 -48677 77652 -48643
rect 77686 -48677 77723 -48643
rect 77636 -48693 77723 -48677
rect 77693 -48733 77723 -48693
rect 77777 -48627 77807 -48521
rect 77885 -48627 77915 -48595
rect 77777 -48643 77843 -48627
rect 77777 -48677 77793 -48643
rect 77827 -48677 77843 -48643
rect 77777 -48693 77843 -48677
rect 77885 -48643 77951 -48627
rect 77885 -48677 77901 -48643
rect 77935 -48677 77951 -48643
rect 77885 -48693 77951 -48677
rect 77777 -48733 77807 -48693
rect 77885 -48715 77915 -48693
rect 77693 -48843 77723 -48817
rect 77777 -48843 77807 -48817
rect 77885 -48871 77915 -48845
rect 77885 -49015 77915 -48989
rect 77693 -49043 77723 -49017
rect 77777 -49043 77807 -49017
rect 77693 -49167 77723 -49127
rect 77636 -49183 77723 -49167
rect 77636 -49217 77652 -49183
rect 77686 -49217 77723 -49183
rect 77636 -49233 77723 -49217
rect 77693 -49339 77723 -49233
rect 77777 -49167 77807 -49127
rect 78117 -49021 78147 -48995
rect 78213 -49021 78243 -48995
rect 78297 -49021 78327 -48995
rect 78381 -49021 78411 -48995
rect 78479 -49015 78509 -48989
rect 77885 -49167 77915 -49145
rect 78117 -49167 78147 -49105
rect 78213 -49167 78243 -49105
rect 78297 -49120 78327 -49105
rect 77777 -49183 77843 -49167
rect 77777 -49217 77793 -49183
rect 77827 -49217 77843 -49183
rect 77777 -49233 77843 -49217
rect 77885 -49183 77951 -49167
rect 77885 -49217 77901 -49183
rect 77935 -49217 77951 -49183
rect 77885 -49233 77951 -49217
rect 78063 -49183 78147 -49167
rect 78063 -49217 78073 -49183
rect 78107 -49217 78147 -49183
rect 78063 -49233 78147 -49217
rect 78189 -49183 78243 -49167
rect 78189 -49217 78199 -49183
rect 78233 -49217 78243 -49183
rect 78189 -49233 78243 -49217
rect 77777 -49339 77807 -49233
rect 77885 -49265 77915 -49233
rect 78117 -49265 78147 -49233
rect 78213 -49265 78243 -49233
rect 78285 -49149 78327 -49120
rect 78285 -49150 78326 -49149
rect 78285 -49265 78315 -49150
rect 78381 -49167 78411 -49105
rect 78479 -49167 78509 -49145
rect 78365 -49183 78419 -49167
rect 78365 -49217 78375 -49183
rect 78409 -49217 78419 -49183
rect 78365 -49233 78419 -49217
rect 78461 -49183 78516 -49167
rect 78461 -49217 78471 -49183
rect 78505 -49217 78516 -49183
rect 78461 -49233 78516 -49217
rect 78381 -49265 78411 -49233
rect 78479 -49265 78509 -49233
rect 77693 -49449 77723 -49423
rect 77777 -49449 77807 -49423
rect 78117 -49375 78147 -49349
rect 78213 -49375 78243 -49349
rect 78285 -49397 78315 -49349
rect 78381 -49375 78411 -49349
rect 78279 -49407 78345 -49397
rect 78279 -49441 78295 -49407
rect 78329 -49441 78345 -49407
rect 78279 -49451 78345 -49441
rect 77885 -49491 77915 -49465
rect 78479 -49491 78509 -49465
rect 77885 -49635 77915 -49609
rect 77693 -49677 77723 -49651
rect 77777 -49677 77807 -49651
rect 77693 -49867 77723 -49761
rect 77636 -49883 77723 -49867
rect 77636 -49917 77652 -49883
rect 77686 -49917 77723 -49883
rect 77636 -49933 77723 -49917
rect 77693 -49973 77723 -49933
rect 77777 -49867 77807 -49761
rect 77885 -49867 77915 -49835
rect 77777 -49883 77843 -49867
rect 77777 -49917 77793 -49883
rect 77827 -49917 77843 -49883
rect 77777 -49933 77843 -49917
rect 77885 -49883 77951 -49867
rect 77885 -49917 77901 -49883
rect 77935 -49917 77951 -49883
rect 77885 -49933 77951 -49917
rect 77777 -49973 77807 -49933
rect 77885 -49955 77915 -49933
rect 77693 -50083 77723 -50057
rect 77777 -50083 77807 -50057
rect 53982 -50334 54079 -50318
rect 53982 -50372 53998 -50334
rect 54032 -50372 54079 -50334
rect 53982 -50388 54079 -50372
rect 54879 -50334 54976 -50318
rect 54879 -50372 54926 -50334
rect 54960 -50372 54976 -50334
rect 54879 -50388 54976 -50372
rect 77885 -50111 77915 -50085
rect 77887 -50269 77917 -50243
rect 77695 -50297 77725 -50271
rect 77779 -50297 77809 -50271
rect 77695 -50421 77725 -50381
rect 77638 -50437 77725 -50421
rect 53510 -50706 53630 -50690
rect 53510 -50740 53526 -50706
rect 53614 -50740 53630 -50706
rect 53510 -50778 53630 -50740
rect 77638 -50471 77654 -50437
rect 77688 -50471 77725 -50437
rect 77638 -50487 77725 -50471
rect 53982 -50690 54079 -50674
rect 53982 -50728 53998 -50690
rect 54032 -50728 54079 -50690
rect 53982 -50744 54079 -50728
rect 54879 -50690 54976 -50674
rect 54879 -50728 54926 -50690
rect 54960 -50728 54976 -50690
rect 54879 -50744 54976 -50728
rect 55318 -50768 55384 -50752
rect 55318 -50802 55334 -50768
rect 55368 -50802 55384 -50768
rect 55318 -50818 55384 -50802
rect 55336 -50840 55366 -50818
rect 55336 -51066 55366 -51040
rect 53510 -51616 53630 -51578
rect 53510 -51650 53526 -51616
rect 53614 -51650 53630 -51616
rect 53510 -51666 53630 -51650
rect 53842 -51440 53930 -51424
rect 53842 -51528 53858 -51440
rect 53892 -51528 53930 -51440
rect 53842 -51544 53930 -51528
rect 54730 -51440 54818 -51424
rect 54730 -51528 54768 -51440
rect 54802 -51528 54818 -51440
rect 54730 -51544 54818 -51528
rect 55030 -51359 55096 -51344
rect 55540 -51359 55606 -51344
rect 55030 -51360 55118 -51359
rect 55030 -51394 55046 -51360
rect 55080 -51394 55118 -51360
rect 55030 -51395 55118 -51394
rect 55518 -51360 55606 -51359
rect 55518 -51394 55556 -51360
rect 55590 -51394 55606 -51360
rect 55518 -51395 55606 -51394
rect 55030 -51410 55096 -51395
rect 55540 -51410 55606 -51395
rect 55866 -50656 55986 -50640
rect 55866 -50690 55882 -50656
rect 55970 -50690 55986 -50656
rect 55866 -50728 55986 -50690
rect 55866 -51566 55986 -51528
rect 55866 -51600 55882 -51566
rect 55970 -51600 55986 -51566
rect 55866 -51616 55986 -51600
rect 57175 -50709 57205 -50683
rect 57263 -50709 57293 -50683
rect 57175 -50882 57205 -50867
rect 57169 -50906 57205 -50882
rect 57169 -50941 57199 -50906
rect 57263 -50928 57293 -50867
rect 77695 -50593 77725 -50487
rect 77779 -50421 77809 -50381
rect 77887 -50421 77917 -50399
rect 77779 -50437 77845 -50421
rect 77779 -50471 77795 -50437
rect 77829 -50471 77845 -50437
rect 77779 -50487 77845 -50471
rect 77887 -50437 77953 -50421
rect 77887 -50471 77903 -50437
rect 77937 -50471 77953 -50437
rect 77887 -50487 77953 -50471
rect 77779 -50593 77809 -50487
rect 77887 -50519 77917 -50487
rect 59544 -50693 59610 -50685
rect 59087 -50743 59113 -50693
rect 59513 -50701 59610 -50693
rect 59513 -50735 59560 -50701
rect 59594 -50735 59610 -50701
rect 59513 -50743 59610 -50735
rect 59544 -50751 59610 -50743
rect 59016 -50801 59082 -50793
rect 59016 -50809 59113 -50801
rect 59016 -50843 59032 -50809
rect 59066 -50843 59113 -50809
rect 59016 -50851 59113 -50843
rect 59513 -50851 59539 -50801
rect 59016 -50859 59082 -50851
rect 57123 -50957 57199 -50941
rect 57123 -50991 57133 -50957
rect 57167 -50991 57199 -50957
rect 57123 -51007 57199 -50991
rect 57241 -50944 57295 -50928
rect 57241 -50978 57251 -50944
rect 57285 -50978 57295 -50944
rect 57241 -50994 57295 -50978
rect 77695 -50703 77725 -50677
rect 77779 -50703 77809 -50677
rect 77887 -50745 77917 -50719
rect 57169 -51016 57199 -51007
rect 57169 -51040 57205 -51016
rect 57175 -51055 57205 -51040
rect 57263 -51055 57293 -50994
rect 77657 -50885 77687 -50859
rect 77757 -50885 77787 -50859
rect 77861 -50885 77891 -50859
rect 77947 -50885 77977 -50859
rect 78113 -50885 78143 -50859
rect 78763 -50885 78793 -50859
rect 53510 -51724 53630 -51708
rect 53510 -51758 53526 -51724
rect 53614 -51758 53630 -51724
rect 53510 -51796 53630 -51758
rect 53842 -51846 53930 -51830
rect 53842 -51934 53858 -51846
rect 53892 -51934 53930 -51846
rect 53842 -51950 53930 -51934
rect 54730 -51846 54818 -51830
rect 54730 -51934 54768 -51846
rect 54802 -51934 54818 -51846
rect 54730 -51950 54818 -51934
rect 55030 -51981 55096 -51966
rect 55540 -51981 55606 -51966
rect 55030 -51982 55118 -51981
rect 55030 -52016 55046 -51982
rect 55080 -52016 55118 -51982
rect 55030 -52017 55118 -52016
rect 55518 -51982 55606 -51981
rect 55518 -52016 55556 -51982
rect 55590 -52016 55606 -51982
rect 55518 -52017 55606 -52016
rect 55030 -52032 55096 -52017
rect 53510 -52634 53630 -52596
rect 53510 -52668 53526 -52634
rect 53614 -52668 53630 -52634
rect 53510 -52684 53630 -52668
rect 55540 -52032 55606 -52017
rect 53972 -52650 54069 -52634
rect 53972 -52688 53988 -52650
rect 54022 -52688 54069 -52650
rect 53972 -52704 54069 -52688
rect 54869 -52650 54966 -52634
rect 54869 -52688 54916 -52650
rect 54950 -52688 54966 -52650
rect 54869 -52704 54966 -52688
rect 55326 -52336 55356 -52310
rect 55326 -52558 55356 -52536
rect 55308 -52574 55374 -52558
rect 55308 -52608 55324 -52574
rect 55358 -52608 55374 -52574
rect 55308 -52624 55374 -52608
rect 55866 -51770 55986 -51754
rect 55866 -51804 55882 -51770
rect 55970 -51804 55986 -51770
rect 55866 -51842 55986 -51804
rect 55866 -52680 55986 -52642
rect 55866 -52714 55882 -52680
rect 55970 -52714 55986 -52680
rect 55866 -52730 55986 -52714
rect 56476 -51206 56546 -51190
rect 56476 -51240 56492 -51206
rect 56530 -51240 56546 -51206
rect 56476 -51287 56546 -51240
rect 57175 -51185 57205 -51159
rect 57263 -51185 57293 -51159
rect 56476 -52134 56546 -52087
rect 56476 -52168 56492 -52134
rect 56530 -52168 56546 -52134
rect 56476 -52184 56546 -52168
rect 59087 -51078 59153 -51062
rect 59087 -51112 59103 -51078
rect 59137 -51112 59153 -51078
rect 59087 -51128 59153 -51112
rect 59090 -51159 59150 -51128
rect 59090 -51590 59150 -51559
rect 59087 -51606 59153 -51590
rect 59087 -51640 59103 -51606
rect 59137 -51640 59153 -51606
rect 59087 -51656 59153 -51640
rect 59858 -51020 59924 -51012
rect 60368 -51020 60434 -51012
rect 59858 -51028 59946 -51020
rect 59858 -51062 59874 -51028
rect 59908 -51062 59946 -51028
rect 59858 -51070 59946 -51062
rect 60346 -51028 60434 -51020
rect 60346 -51062 60384 -51028
rect 60418 -51062 60434 -51028
rect 60346 -51070 60434 -51062
rect 59858 -51078 59924 -51070
rect 60368 -51078 60434 -51070
rect 77657 -51117 77687 -50969
rect 77757 -51117 77787 -50969
rect 77861 -51117 77891 -50969
rect 77947 -51117 77977 -50969
rect 78563 -50909 78629 -50899
rect 78563 -50943 78579 -50909
rect 78613 -50943 78629 -50909
rect 78563 -50953 78629 -50943
rect 78401 -51001 78431 -50975
rect 78497 -51001 78527 -50975
rect 78569 -51001 78599 -50953
rect 78665 -51001 78695 -50975
rect 78113 -51117 78143 -51085
rect 78401 -51117 78431 -51085
rect 78497 -51117 78527 -51085
rect 77599 -51133 77687 -51117
rect 77599 -51167 77609 -51133
rect 77643 -51167 77687 -51133
rect 77599 -51183 77687 -51167
rect 59530 -51298 59596 -51282
rect 59530 -51332 59546 -51298
rect 59580 -51332 59596 -51298
rect 59530 -51348 59596 -51332
rect 59548 -51370 59578 -51348
rect 59548 -51592 59578 -51570
rect 59530 -51608 59596 -51592
rect 59530 -51642 59546 -51608
rect 59580 -51642 59596 -51608
rect 59530 -51658 59596 -51642
rect 59846 -51298 59912 -51282
rect 59846 -51332 59862 -51298
rect 59896 -51332 59912 -51298
rect 59846 -51348 59912 -51332
rect 59864 -51370 59894 -51348
rect 59864 -51592 59894 -51570
rect 59846 -51608 59912 -51592
rect 59846 -51642 59862 -51608
rect 59896 -51642 59912 -51608
rect 59846 -51658 59912 -51642
rect 77657 -51251 77687 -51183
rect 77745 -51133 77799 -51117
rect 77745 -51167 77755 -51133
rect 77789 -51167 77799 -51133
rect 77745 -51183 77799 -51167
rect 77851 -51133 77905 -51117
rect 77851 -51167 77861 -51133
rect 77895 -51167 77905 -51133
rect 77851 -51183 77905 -51167
rect 77947 -51133 78011 -51117
rect 77947 -51167 77957 -51133
rect 77991 -51167 78011 -51133
rect 77947 -51183 78011 -51167
rect 78058 -51133 78143 -51117
rect 78058 -51167 78068 -51133
rect 78102 -51167 78143 -51133
rect 78058 -51183 78143 -51167
rect 78347 -51133 78431 -51117
rect 78347 -51167 78357 -51133
rect 78391 -51167 78431 -51133
rect 78347 -51183 78431 -51167
rect 78473 -51133 78527 -51117
rect 78473 -51167 78483 -51133
rect 78517 -51167 78527 -51133
rect 78473 -51183 78527 -51167
rect 77745 -51251 77775 -51183
rect 77851 -51251 77881 -51183
rect 77947 -51251 77977 -51183
rect 78113 -51205 78143 -51183
rect 78401 -51245 78431 -51183
rect 78497 -51245 78527 -51183
rect 78569 -51200 78599 -51085
rect 78665 -51117 78695 -51085
rect 78763 -51117 78793 -51085
rect 78649 -51133 78703 -51117
rect 78649 -51167 78659 -51133
rect 78693 -51167 78703 -51133
rect 78649 -51183 78703 -51167
rect 78745 -51133 78800 -51117
rect 78745 -51167 78755 -51133
rect 78789 -51167 78800 -51133
rect 78745 -51183 78800 -51167
rect 78569 -51201 78610 -51200
rect 78569 -51230 78611 -51201
rect 78581 -51245 78611 -51230
rect 78665 -51245 78695 -51183
rect 78763 -51205 78793 -51183
rect 77657 -51361 77687 -51335
rect 77745 -51361 77775 -51335
rect 77851 -51361 77881 -51335
rect 77947 -51361 77977 -51335
rect 78113 -51361 78143 -51335
rect 78401 -51355 78431 -51329
rect 78497 -51355 78527 -51329
rect 78581 -51355 78611 -51329
rect 78665 -51355 78695 -51329
rect 78763 -51361 78793 -51335
rect 83127 -51445 83157 -51419
rect 83418 -51445 83448 -51419
rect 83663 -51445 83693 -51419
rect 83747 -51445 83777 -51419
rect 83831 -51445 83861 -51419
rect 83915 -51445 83945 -51419
rect 84126 -51445 84156 -51419
rect 84210 -51445 84240 -51419
rect 84294 -51445 84324 -51419
rect 84378 -51445 84408 -51419
rect 84462 -51445 84492 -51419
rect 84546 -51445 84576 -51419
rect 84630 -51445 84660 -51419
rect 84714 -51445 84744 -51419
rect 84798 -51445 84828 -51419
rect 84882 -51445 84912 -51419
rect 84966 -51445 84996 -51419
rect 85050 -51445 85080 -51419
rect 85134 -51445 85164 -51419
rect 85218 -51445 85248 -51419
rect 85302 -51445 85332 -51419
rect 85386 -51445 85416 -51419
rect 85598 -51445 85628 -51419
rect 85682 -51445 85712 -51419
rect 85766 -51445 85796 -51419
rect 85850 -51445 85880 -51419
rect 85934 -51445 85964 -51419
rect 86018 -51445 86048 -51419
rect 86102 -51445 86132 -51419
rect 86186 -51445 86216 -51419
rect 86270 -51445 86300 -51419
rect 86354 -51445 86384 -51419
rect 86438 -51445 86468 -51419
rect 86522 -51445 86552 -51419
rect 86606 -51445 86636 -51419
rect 86690 -51445 86720 -51419
rect 86774 -51445 86804 -51419
rect 86858 -51445 86888 -51419
rect 87070 -51445 87100 -51419
rect 87154 -51445 87184 -51419
rect 87238 -51445 87268 -51419
rect 87322 -51445 87352 -51419
rect 87406 -51445 87436 -51419
rect 87490 -51445 87520 -51419
rect 87574 -51445 87604 -51419
rect 87658 -51445 87688 -51419
rect 87742 -51445 87772 -51419
rect 87826 -51445 87856 -51419
rect 87910 -51445 87940 -51419
rect 87994 -51445 88024 -51419
rect 88078 -51445 88108 -51419
rect 88162 -51445 88192 -51419
rect 88246 -51445 88276 -51419
rect 88330 -51445 88360 -51419
rect 88542 -51445 88572 -51419
rect 88626 -51445 88656 -51419
rect 88710 -51445 88740 -51419
rect 88794 -51445 88824 -51419
rect 88878 -51445 88908 -51419
rect 88962 -51445 88992 -51419
rect 89046 -51445 89076 -51419
rect 89130 -51445 89160 -51419
rect 89214 -51445 89244 -51419
rect 89298 -51445 89328 -51419
rect 89382 -51445 89412 -51419
rect 89466 -51445 89496 -51419
rect 89550 -51445 89580 -51419
rect 89634 -51445 89664 -51419
rect 89718 -51445 89748 -51419
rect 89802 -51445 89832 -51419
rect 90014 -51445 90044 -51419
rect 90098 -51445 90128 -51419
rect 90182 -51445 90212 -51419
rect 90266 -51445 90296 -51419
rect 90350 -51445 90380 -51419
rect 90434 -51445 90464 -51419
rect 90518 -51445 90548 -51419
rect 90602 -51445 90632 -51419
rect 90686 -51445 90716 -51419
rect 90770 -51445 90800 -51419
rect 90854 -51445 90884 -51419
rect 90938 -51445 90968 -51419
rect 91022 -51445 91052 -51419
rect 91106 -51445 91136 -51419
rect 91190 -51445 91220 -51419
rect 91274 -51445 91304 -51419
rect 77657 -51501 77687 -51475
rect 77745 -51501 77775 -51475
rect 77851 -51501 77881 -51475
rect 77947 -51501 77977 -51475
rect 78113 -51501 78143 -51475
rect 60343 -51565 60409 -51549
rect 61043 -51565 61109 -51549
rect 60343 -51599 60359 -51565
rect 60393 -51599 60409 -51565
rect 60343 -51617 60409 -51599
rect 61043 -51599 61059 -51565
rect 61093 -51599 61109 -51565
rect 61043 -51617 61109 -51599
rect 60165 -51647 60191 -51617
rect 60321 -51647 60441 -51617
rect 60641 -51647 60667 -51617
rect 60785 -51647 60811 -51617
rect 61011 -51647 61131 -51617
rect 61261 -51647 61287 -51617
rect 60343 -51657 60409 -51647
rect 60343 -51691 60359 -51657
rect 60393 -51691 60409 -51657
rect 60343 -51701 60409 -51691
rect 61043 -51657 61109 -51647
rect 61043 -51691 61059 -51657
rect 61093 -51691 61109 -51657
rect 61043 -51701 61109 -51691
rect 77657 -51653 77687 -51585
rect 77599 -51669 77687 -51653
rect 57175 -52229 57205 -52203
rect 57263 -52229 57293 -52203
rect 57175 -52348 57205 -52333
rect 57169 -52372 57205 -52348
rect 57169 -52381 57199 -52372
rect 57123 -52397 57199 -52381
rect 57263 -52394 57293 -52333
rect 59087 -51808 59153 -51792
rect 59087 -51842 59103 -51808
rect 59137 -51842 59153 -51808
rect 59087 -51858 59153 -51842
rect 59090 -51889 59150 -51858
rect 59090 -52320 59150 -52289
rect 57123 -52431 57133 -52397
rect 57167 -52431 57199 -52397
rect 57123 -52447 57199 -52431
rect 57169 -52482 57199 -52447
rect 57241 -52410 57295 -52394
rect 57241 -52444 57251 -52410
rect 57285 -52444 57295 -52410
rect 57241 -52460 57295 -52444
rect 59087 -52336 59153 -52320
rect 59087 -52370 59103 -52336
rect 59137 -52370 59153 -52336
rect 59087 -52386 59153 -52370
rect 60165 -51731 60191 -51701
rect 60321 -51731 60441 -51701
rect 60641 -51731 60667 -51701
rect 60785 -51731 60811 -51701
rect 61011 -51731 61131 -51701
rect 61261 -51731 61287 -51701
rect 77599 -51703 77609 -51669
rect 77643 -51703 77687 -51669
rect 77599 -51719 77687 -51703
rect 77745 -51653 77775 -51585
rect 77851 -51653 77881 -51585
rect 77947 -51653 77977 -51585
rect 82958 -51561 82988 -51535
rect 83030 -51561 83060 -51535
rect 78113 -51653 78143 -51631
rect 77745 -51669 77799 -51653
rect 77745 -51703 77755 -51669
rect 77789 -51703 77799 -51669
rect 77745 -51719 77799 -51703
rect 77851 -51669 77905 -51653
rect 77851 -51703 77861 -51669
rect 77895 -51703 77905 -51669
rect 77851 -51719 77905 -51703
rect 77947 -51669 78011 -51653
rect 77947 -51703 77957 -51669
rect 77991 -51703 78011 -51669
rect 77947 -51719 78011 -51703
rect 78058 -51669 78143 -51653
rect 78058 -51703 78068 -51669
rect 78102 -51703 78143 -51669
rect 82958 -51677 82988 -51645
rect 78058 -51719 78143 -51703
rect 59526 -51811 59596 -51780
rect 59526 -51830 59545 -51811
rect 59529 -51845 59545 -51830
rect 59579 -51830 59596 -51811
rect 59579 -51845 59595 -51830
rect 59529 -51861 59595 -51845
rect 59547 -51883 59577 -51861
rect 59547 -52105 59577 -52083
rect 59529 -52121 59595 -52105
rect 59529 -52155 59545 -52121
rect 59579 -52155 59595 -52121
rect 59529 -52171 59595 -52155
rect 59845 -51811 59911 -51795
rect 59845 -51845 59861 -51811
rect 59895 -51845 59911 -51811
rect 59845 -51861 59911 -51845
rect 60343 -51741 60409 -51731
rect 60343 -51775 60359 -51741
rect 60393 -51775 60409 -51741
rect 60343 -51785 60409 -51775
rect 61043 -51741 61109 -51731
rect 61043 -51775 61059 -51741
rect 61093 -51775 61109 -51741
rect 61043 -51785 61109 -51775
rect 59863 -51883 59893 -51861
rect 59863 -52105 59893 -52083
rect 59845 -52121 59911 -52105
rect 59845 -52155 59861 -52121
rect 59895 -52155 59911 -52121
rect 59845 -52171 59911 -52155
rect 60165 -51815 60191 -51785
rect 60321 -51815 60441 -51785
rect 60641 -51815 60667 -51785
rect 60785 -51815 60811 -51785
rect 61011 -51815 61131 -51785
rect 61261 -51815 61287 -51785
rect 60343 -51825 60409 -51815
rect 60343 -51859 60359 -51825
rect 60393 -51859 60409 -51825
rect 60343 -51869 60409 -51859
rect 61043 -51825 61109 -51815
rect 61043 -51859 61059 -51825
rect 61093 -51859 61109 -51825
rect 61043 -51869 61109 -51859
rect 77657 -51867 77687 -51719
rect 77757 -51867 77787 -51719
rect 77861 -51867 77891 -51719
rect 77947 -51867 77977 -51719
rect 78113 -51751 78143 -51719
rect 82888 -51693 82988 -51677
rect 82888 -51727 82904 -51693
rect 82938 -51727 82988 -51693
rect 82888 -51743 82988 -51727
rect 83030 -51677 83060 -51645
rect 83127 -51677 83157 -51645
rect 83418 -51677 83448 -51645
rect 83663 -51677 83693 -51645
rect 83747 -51677 83777 -51645
rect 83831 -51677 83861 -51645
rect 83915 -51677 83945 -51645
rect 84126 -51677 84156 -51645
rect 84210 -51677 84240 -51645
rect 84294 -51677 84324 -51645
rect 84378 -51677 84408 -51645
rect 84462 -51677 84492 -51645
rect 84546 -51677 84576 -51645
rect 84630 -51677 84660 -51645
rect 84714 -51677 84744 -51645
rect 84798 -51677 84828 -51645
rect 84882 -51677 84912 -51645
rect 84966 -51677 84996 -51645
rect 85050 -51677 85080 -51645
rect 85134 -51677 85164 -51645
rect 85218 -51677 85248 -51645
rect 85302 -51677 85332 -51645
rect 85386 -51677 85416 -51645
rect 85598 -51677 85628 -51645
rect 85682 -51677 85712 -51645
rect 85766 -51677 85796 -51645
rect 85850 -51677 85880 -51645
rect 85934 -51677 85964 -51645
rect 86018 -51677 86048 -51645
rect 86102 -51677 86132 -51645
rect 86186 -51677 86216 -51645
rect 86270 -51677 86300 -51645
rect 86354 -51677 86384 -51645
rect 86438 -51677 86468 -51645
rect 86522 -51677 86552 -51645
rect 86606 -51677 86636 -51645
rect 86690 -51677 86720 -51645
rect 86774 -51677 86804 -51645
rect 86858 -51677 86888 -51645
rect 87070 -51677 87100 -51645
rect 87154 -51677 87184 -51645
rect 87238 -51677 87268 -51645
rect 87322 -51677 87352 -51645
rect 87406 -51677 87436 -51645
rect 87490 -51677 87520 -51645
rect 87574 -51677 87604 -51645
rect 87658 -51677 87688 -51645
rect 87742 -51677 87772 -51645
rect 87826 -51677 87856 -51645
rect 87910 -51677 87940 -51645
rect 87994 -51677 88024 -51645
rect 88078 -51677 88108 -51645
rect 88162 -51677 88192 -51645
rect 88246 -51677 88276 -51645
rect 88330 -51677 88360 -51645
rect 88542 -51677 88572 -51645
rect 88626 -51677 88656 -51645
rect 88710 -51677 88740 -51645
rect 88794 -51677 88824 -51645
rect 88878 -51677 88908 -51645
rect 88962 -51677 88992 -51645
rect 89046 -51677 89076 -51645
rect 89130 -51677 89160 -51645
rect 89214 -51677 89244 -51645
rect 89298 -51677 89328 -51645
rect 89382 -51677 89412 -51645
rect 89466 -51677 89496 -51645
rect 89550 -51677 89580 -51645
rect 89634 -51677 89664 -51645
rect 89718 -51677 89748 -51645
rect 89802 -51677 89832 -51645
rect 90014 -51677 90044 -51645
rect 90098 -51677 90128 -51645
rect 90182 -51677 90212 -51645
rect 90266 -51677 90296 -51645
rect 90350 -51677 90380 -51645
rect 90434 -51677 90464 -51645
rect 90518 -51677 90548 -51645
rect 90602 -51677 90632 -51645
rect 90686 -51677 90716 -51645
rect 90770 -51677 90800 -51645
rect 90854 -51677 90884 -51645
rect 90938 -51677 90968 -51645
rect 91022 -51677 91052 -51645
rect 91106 -51677 91136 -51645
rect 91190 -51677 91220 -51645
rect 91274 -51677 91304 -51645
rect 83030 -51693 83084 -51677
rect 83030 -51727 83040 -51693
rect 83074 -51727 83084 -51693
rect 83030 -51743 83084 -51727
rect 83127 -51693 83193 -51677
rect 83127 -51727 83143 -51693
rect 83177 -51727 83193 -51693
rect 83127 -51743 83193 -51727
rect 83362 -51693 83448 -51677
rect 83362 -51727 83378 -51693
rect 83412 -51727 83448 -51693
rect 83362 -51743 83448 -51727
rect 83595 -51693 83945 -51677
rect 83595 -51727 83611 -51693
rect 83645 -51727 83703 -51693
rect 83737 -51727 83787 -51693
rect 83821 -51727 83871 -51693
rect 83905 -51727 83945 -51693
rect 83595 -51743 83945 -51727
rect 84060 -51693 85416 -51677
rect 84060 -51727 84076 -51693
rect 84110 -51727 84250 -51693
rect 84284 -51727 84418 -51693
rect 84452 -51727 84587 -51693
rect 84621 -51727 84754 -51693
rect 84788 -51727 84922 -51693
rect 84956 -51727 85089 -51693
rect 85123 -51727 85416 -51693
rect 84060 -51743 85416 -51727
rect 85532 -51693 86888 -51677
rect 85532 -51727 85548 -51693
rect 85582 -51727 85722 -51693
rect 85756 -51727 85890 -51693
rect 85924 -51727 86059 -51693
rect 86093 -51727 86226 -51693
rect 86260 -51727 86394 -51693
rect 86428 -51727 86561 -51693
rect 86595 -51727 86888 -51693
rect 85532 -51743 86888 -51727
rect 87004 -51693 88360 -51677
rect 87004 -51727 87020 -51693
rect 87054 -51727 87194 -51693
rect 87228 -51727 87362 -51693
rect 87396 -51727 87531 -51693
rect 87565 -51727 87698 -51693
rect 87732 -51727 87866 -51693
rect 87900 -51727 88033 -51693
rect 88067 -51727 88360 -51693
rect 87004 -51743 88360 -51727
rect 88476 -51693 89832 -51677
rect 88476 -51727 88492 -51693
rect 88526 -51727 88666 -51693
rect 88700 -51727 88834 -51693
rect 88868 -51727 89003 -51693
rect 89037 -51727 89170 -51693
rect 89204 -51727 89338 -51693
rect 89372 -51727 89505 -51693
rect 89539 -51727 89832 -51693
rect 88476 -51743 89832 -51727
rect 89948 -51693 91304 -51677
rect 89948 -51727 89964 -51693
rect 89998 -51727 90138 -51693
rect 90172 -51727 90306 -51693
rect 90340 -51727 90475 -51693
rect 90509 -51727 90642 -51693
rect 90676 -51727 90810 -51693
rect 90844 -51727 90977 -51693
rect 91011 -51727 91304 -51693
rect 89948 -51743 91304 -51727
rect 60165 -51899 60191 -51869
rect 60321 -51899 60441 -51869
rect 60641 -51899 60667 -51869
rect 60785 -51899 60811 -51869
rect 61011 -51899 61131 -51869
rect 61261 -51899 61287 -51869
rect 82946 -51811 82976 -51743
rect 83030 -51811 83060 -51743
rect 83127 -51765 83157 -51743
rect 83418 -51765 83448 -51743
rect 83663 -51765 83693 -51743
rect 83747 -51765 83777 -51743
rect 83831 -51765 83861 -51743
rect 83915 -51765 83945 -51743
rect 84126 -51765 84156 -51743
rect 84210 -51765 84240 -51743
rect 84294 -51765 84324 -51743
rect 84378 -51765 84408 -51743
rect 84462 -51765 84492 -51743
rect 84546 -51765 84576 -51743
rect 84630 -51765 84660 -51743
rect 84714 -51765 84744 -51743
rect 84798 -51765 84828 -51743
rect 84882 -51765 84912 -51743
rect 84966 -51765 84996 -51743
rect 85050 -51765 85080 -51743
rect 85134 -51765 85164 -51743
rect 85218 -51765 85248 -51743
rect 85302 -51765 85332 -51743
rect 85386 -51765 85416 -51743
rect 85598 -51765 85628 -51743
rect 85682 -51765 85712 -51743
rect 85766 -51765 85796 -51743
rect 85850 -51765 85880 -51743
rect 85934 -51765 85964 -51743
rect 86018 -51765 86048 -51743
rect 86102 -51765 86132 -51743
rect 86186 -51765 86216 -51743
rect 86270 -51765 86300 -51743
rect 86354 -51765 86384 -51743
rect 86438 -51765 86468 -51743
rect 86522 -51765 86552 -51743
rect 86606 -51765 86636 -51743
rect 86690 -51765 86720 -51743
rect 86774 -51765 86804 -51743
rect 86858 -51765 86888 -51743
rect 87070 -51765 87100 -51743
rect 87154 -51765 87184 -51743
rect 87238 -51765 87268 -51743
rect 87322 -51765 87352 -51743
rect 87406 -51765 87436 -51743
rect 87490 -51765 87520 -51743
rect 87574 -51765 87604 -51743
rect 87658 -51765 87688 -51743
rect 87742 -51765 87772 -51743
rect 87826 -51765 87856 -51743
rect 87910 -51765 87940 -51743
rect 87994 -51765 88024 -51743
rect 88078 -51765 88108 -51743
rect 88162 -51765 88192 -51743
rect 88246 -51765 88276 -51743
rect 88330 -51765 88360 -51743
rect 88542 -51765 88572 -51743
rect 88626 -51765 88656 -51743
rect 88710 -51765 88740 -51743
rect 88794 -51765 88824 -51743
rect 88878 -51765 88908 -51743
rect 88962 -51765 88992 -51743
rect 89046 -51765 89076 -51743
rect 89130 -51765 89160 -51743
rect 89214 -51765 89244 -51743
rect 89298 -51765 89328 -51743
rect 89382 -51765 89412 -51743
rect 89466 -51765 89496 -51743
rect 89550 -51765 89580 -51743
rect 89634 -51765 89664 -51743
rect 89718 -51765 89748 -51743
rect 89802 -51765 89832 -51743
rect 90014 -51765 90044 -51743
rect 90098 -51765 90128 -51743
rect 90182 -51765 90212 -51743
rect 90266 -51765 90296 -51743
rect 90350 -51765 90380 -51743
rect 90434 -51765 90464 -51743
rect 90518 -51765 90548 -51743
rect 90602 -51765 90632 -51743
rect 90686 -51765 90716 -51743
rect 90770 -51765 90800 -51743
rect 90854 -51765 90884 -51743
rect 90938 -51765 90968 -51743
rect 91022 -51765 91052 -51743
rect 91106 -51765 91136 -51743
rect 91190 -51765 91220 -51743
rect 91274 -51765 91304 -51743
rect 82946 -51921 82976 -51895
rect 83030 -51921 83060 -51895
rect 83127 -51921 83157 -51895
rect 83418 -51921 83448 -51895
rect 83663 -51921 83693 -51895
rect 83747 -51921 83777 -51895
rect 83831 -51921 83861 -51895
rect 83915 -51921 83945 -51895
rect 84126 -51921 84156 -51895
rect 84210 -51921 84240 -51895
rect 84294 -51921 84324 -51895
rect 84378 -51921 84408 -51895
rect 84462 -51921 84492 -51895
rect 84546 -51921 84576 -51895
rect 84630 -51921 84660 -51895
rect 84714 -51921 84744 -51895
rect 84798 -51921 84828 -51895
rect 84882 -51921 84912 -51895
rect 84966 -51921 84996 -51895
rect 85050 -51921 85080 -51895
rect 85134 -51921 85164 -51895
rect 85218 -51921 85248 -51895
rect 85302 -51921 85332 -51895
rect 85386 -51921 85416 -51895
rect 85598 -51921 85628 -51895
rect 85682 -51921 85712 -51895
rect 85766 -51921 85796 -51895
rect 85850 -51921 85880 -51895
rect 85934 -51921 85964 -51895
rect 86018 -51921 86048 -51895
rect 86102 -51921 86132 -51895
rect 86186 -51921 86216 -51895
rect 86270 -51921 86300 -51895
rect 86354 -51921 86384 -51895
rect 86438 -51921 86468 -51895
rect 86522 -51921 86552 -51895
rect 86606 -51921 86636 -51895
rect 86690 -51921 86720 -51895
rect 86774 -51921 86804 -51895
rect 86858 -51921 86888 -51895
rect 87070 -51921 87100 -51895
rect 87154 -51921 87184 -51895
rect 87238 -51921 87268 -51895
rect 87322 -51921 87352 -51895
rect 87406 -51921 87436 -51895
rect 87490 -51921 87520 -51895
rect 87574 -51921 87604 -51895
rect 87658 -51921 87688 -51895
rect 87742 -51921 87772 -51895
rect 87826 -51921 87856 -51895
rect 87910 -51921 87940 -51895
rect 87994 -51921 88024 -51895
rect 88078 -51921 88108 -51895
rect 88162 -51921 88192 -51895
rect 88246 -51921 88276 -51895
rect 88330 -51921 88360 -51895
rect 88542 -51921 88572 -51895
rect 88626 -51921 88656 -51895
rect 88710 -51921 88740 -51895
rect 88794 -51921 88824 -51895
rect 88878 -51921 88908 -51895
rect 88962 -51921 88992 -51895
rect 89046 -51921 89076 -51895
rect 89130 -51921 89160 -51895
rect 89214 -51921 89244 -51895
rect 89298 -51921 89328 -51895
rect 89382 -51921 89412 -51895
rect 89466 -51921 89496 -51895
rect 89550 -51921 89580 -51895
rect 89634 -51921 89664 -51895
rect 89718 -51921 89748 -51895
rect 89802 -51921 89832 -51895
rect 90014 -51921 90044 -51895
rect 90098 -51921 90128 -51895
rect 90182 -51921 90212 -51895
rect 90266 -51921 90296 -51895
rect 90350 -51921 90380 -51895
rect 90434 -51921 90464 -51895
rect 90518 -51921 90548 -51895
rect 90602 -51921 90632 -51895
rect 90686 -51921 90716 -51895
rect 90770 -51921 90800 -51895
rect 90854 -51921 90884 -51895
rect 90938 -51921 90968 -51895
rect 91022 -51921 91052 -51895
rect 91106 -51921 91136 -51895
rect 91190 -51921 91220 -51895
rect 91274 -51921 91304 -51895
rect 77657 -51977 77687 -51951
rect 77757 -51977 77787 -51951
rect 77861 -51977 77891 -51951
rect 77947 -51977 77977 -51951
rect 78113 -51977 78143 -51951
rect 77657 -52117 77687 -52091
rect 77757 -52117 77787 -52091
rect 77861 -52117 77891 -52091
rect 77947 -52117 77977 -52091
rect 78113 -52117 78143 -52091
rect 57169 -52506 57205 -52482
rect 57175 -52521 57205 -52506
rect 57263 -52521 57293 -52460
rect 57175 -52705 57205 -52679
rect 57263 -52705 57293 -52679
rect 59544 -52600 59610 -52592
rect 59087 -52650 59113 -52600
rect 59513 -52608 59610 -52600
rect 59513 -52642 59560 -52608
rect 59594 -52642 59610 -52608
rect 59513 -52650 59610 -52642
rect 59544 -52658 59610 -52650
rect 59016 -52708 59082 -52700
rect 59016 -52716 59113 -52708
rect 59016 -52750 59032 -52716
rect 59066 -52750 59113 -52716
rect 59016 -52758 59113 -52750
rect 59513 -52758 59539 -52708
rect 59016 -52766 59082 -52758
rect 53972 -53006 54069 -52990
rect 53972 -53044 53988 -53006
rect 54022 -53044 54069 -53006
rect 53972 -53060 54069 -53044
rect 54869 -53006 54966 -52990
rect 54869 -53044 54916 -53006
rect 54950 -53044 54966 -53006
rect 54869 -53060 54966 -53044
rect 59858 -52386 59924 -52378
rect 60368 -52386 60434 -52378
rect 59858 -52394 59946 -52386
rect 59858 -52428 59874 -52394
rect 59908 -52428 59946 -52394
rect 59858 -52436 59946 -52428
rect 60346 -52394 60434 -52386
rect 60346 -52428 60384 -52394
rect 60418 -52428 60434 -52394
rect 60346 -52436 60434 -52428
rect 59858 -52444 59924 -52436
rect 60368 -52444 60434 -52436
rect 77657 -52349 77687 -52201
rect 77757 -52349 77787 -52201
rect 77861 -52349 77891 -52201
rect 77947 -52349 77977 -52201
rect 78113 -52349 78143 -52317
rect 77599 -52365 77687 -52349
rect 77599 -52399 77609 -52365
rect 77643 -52399 77687 -52365
rect 77599 -52415 77687 -52399
rect 77657 -52483 77687 -52415
rect 77745 -52365 77799 -52349
rect 77745 -52399 77755 -52365
rect 77789 -52399 77799 -52365
rect 77745 -52415 77799 -52399
rect 77851 -52365 77905 -52349
rect 77851 -52399 77861 -52365
rect 77895 -52399 77905 -52365
rect 77851 -52415 77905 -52399
rect 77947 -52365 78011 -52349
rect 77947 -52399 77957 -52365
rect 77991 -52399 78011 -52365
rect 77947 -52415 78011 -52399
rect 78058 -52365 78143 -52349
rect 78058 -52399 78068 -52365
rect 78102 -52399 78143 -52365
rect 78058 -52415 78143 -52399
rect 77745 -52483 77775 -52415
rect 77851 -52483 77881 -52415
rect 77947 -52483 77977 -52415
rect 78113 -52437 78143 -52415
rect 77657 -52593 77687 -52567
rect 77745 -52593 77775 -52567
rect 77851 -52593 77881 -52567
rect 77947 -52593 77977 -52567
rect 78113 -52593 78143 -52567
rect 77657 -52735 77687 -52709
rect 77745 -52735 77775 -52709
rect 77851 -52735 77881 -52709
rect 77947 -52735 77977 -52709
rect 78113 -52735 78143 -52709
rect 77657 -52887 77687 -52819
rect 77599 -52903 77687 -52887
rect 77599 -52937 77609 -52903
rect 77643 -52937 77687 -52903
rect 77599 -52953 77687 -52937
rect 77745 -52887 77775 -52819
rect 77851 -52887 77881 -52819
rect 77947 -52887 77977 -52819
rect 78113 -52887 78143 -52865
rect 77745 -52903 77799 -52887
rect 77745 -52937 77755 -52903
rect 77789 -52937 77799 -52903
rect 77745 -52953 77799 -52937
rect 77851 -52903 77905 -52887
rect 77851 -52937 77861 -52903
rect 77895 -52937 77905 -52903
rect 77851 -52953 77905 -52937
rect 77947 -52903 78011 -52887
rect 77947 -52937 77957 -52903
rect 77991 -52937 78011 -52903
rect 77947 -52953 78011 -52937
rect 78058 -52903 78143 -52887
rect 78058 -52937 78068 -52903
rect 78102 -52937 78143 -52903
rect 78058 -52953 78143 -52937
rect 77657 -53101 77687 -52953
rect 77757 -53101 77787 -52953
rect 77861 -53101 77891 -52953
rect 77947 -53101 77977 -52953
rect 78113 -52985 78143 -52953
rect 55510 -53202 55576 -53186
rect 55510 -53204 55526 -53202
rect 55262 -53234 55288 -53204
rect 55488 -53234 55526 -53204
rect 55510 -53236 55526 -53234
rect 55560 -53236 55576 -53202
rect 55510 -53252 55576 -53236
rect 77657 -53211 77687 -53185
rect 77757 -53211 77787 -53185
rect 77861 -53211 77891 -53185
rect 77947 -53211 77977 -53185
rect 78113 -53211 78143 -53185
rect 77929 -53355 77959 -53329
rect 78345 -53355 78375 -53329
rect 78939 -53355 78969 -53329
rect 77741 -53376 77795 -53360
rect 77741 -53410 77751 -53376
rect 77785 -53410 77795 -53376
rect 77741 -53426 77795 -53410
rect 77657 -53468 77687 -53427
rect 77741 -53468 77771 -53426
rect 77834 -53468 77864 -53442
rect 77657 -53601 77687 -53552
rect 77741 -53570 77771 -53552
rect 77603 -53649 77687 -53601
rect 77603 -53683 77613 -53649
rect 77647 -53683 77687 -53649
rect 77603 -53706 77687 -53683
rect 77657 -53721 77687 -53706
rect 77729 -53595 77771 -53570
rect 77834 -53593 77864 -53552
rect 78153 -53397 78183 -53371
rect 78237 -53397 78267 -53371
rect 77929 -53587 77959 -53555
rect 78153 -53587 78183 -53481
rect 77729 -53721 77759 -53595
rect 77813 -53609 77867 -53593
rect 77813 -53626 77823 -53609
rect 77801 -53643 77823 -53626
rect 77857 -53643 77867 -53609
rect 77801 -53659 77867 -53643
rect 77909 -53603 77963 -53587
rect 77909 -53637 77919 -53603
rect 77953 -53637 77963 -53603
rect 77909 -53653 77963 -53637
rect 78096 -53603 78183 -53587
rect 78096 -53637 78112 -53603
rect 78146 -53637 78183 -53603
rect 78096 -53653 78183 -53637
rect 77801 -53682 77843 -53659
rect 77929 -53675 77959 -53653
rect 77801 -53706 77838 -53682
rect 77801 -53721 77831 -53706
rect 78153 -53693 78183 -53653
rect 78237 -53587 78267 -53481
rect 78739 -53379 78805 -53369
rect 78739 -53413 78755 -53379
rect 78789 -53413 78805 -53379
rect 78739 -53423 78805 -53413
rect 78577 -53471 78607 -53445
rect 78673 -53471 78703 -53445
rect 78745 -53471 78775 -53423
rect 78841 -53471 78871 -53445
rect 78345 -53587 78375 -53555
rect 78577 -53587 78607 -53555
rect 78673 -53587 78703 -53555
rect 78237 -53603 78303 -53587
rect 78237 -53637 78253 -53603
rect 78287 -53637 78303 -53603
rect 78237 -53653 78303 -53637
rect 78345 -53603 78411 -53587
rect 78345 -53637 78361 -53603
rect 78395 -53637 78411 -53603
rect 78345 -53653 78411 -53637
rect 78523 -53603 78607 -53587
rect 78523 -53637 78533 -53603
rect 78567 -53637 78607 -53603
rect 78523 -53653 78607 -53637
rect 78649 -53603 78703 -53587
rect 78649 -53637 78659 -53603
rect 78693 -53637 78703 -53603
rect 78649 -53653 78703 -53637
rect 78237 -53693 78267 -53653
rect 78345 -53675 78375 -53653
rect 78153 -53803 78183 -53777
rect 78237 -53803 78267 -53777
rect 78577 -53715 78607 -53653
rect 78673 -53715 78703 -53653
rect 78745 -53670 78775 -53555
rect 78841 -53587 78871 -53555
rect 78939 -53587 78969 -53555
rect 78825 -53603 78879 -53587
rect 78825 -53637 78835 -53603
rect 78869 -53637 78879 -53603
rect 78825 -53653 78879 -53637
rect 78921 -53603 78976 -53587
rect 78921 -53637 78931 -53603
rect 78965 -53637 78976 -53603
rect 78921 -53653 78976 -53637
rect 78745 -53671 78786 -53670
rect 78745 -53700 78787 -53671
rect 78757 -53715 78787 -53700
rect 78841 -53715 78871 -53653
rect 78939 -53675 78969 -53653
rect 77657 -53831 77687 -53805
rect 77729 -53831 77759 -53805
rect 77801 -53831 77831 -53805
rect 77929 -53831 77959 -53805
rect 78345 -53831 78375 -53805
rect 78577 -53825 78607 -53799
rect 78673 -53825 78703 -53799
rect 78757 -53825 78787 -53799
rect 78841 -53825 78871 -53799
rect 78939 -53831 78969 -53805
rect 53982 -55734 54079 -55718
rect 53982 -55772 53998 -55734
rect 54032 -55772 54079 -55734
rect 53982 -55788 54079 -55772
rect 54879 -55734 54976 -55718
rect 54879 -55772 54926 -55734
rect 54960 -55772 54976 -55734
rect 54879 -55788 54976 -55772
rect 53510 -56106 53630 -56090
rect 53510 -56140 53526 -56106
rect 53614 -56140 53630 -56106
rect 53510 -56178 53630 -56140
rect 53982 -56090 54079 -56074
rect 53982 -56128 53998 -56090
rect 54032 -56128 54079 -56090
rect 53982 -56144 54079 -56128
rect 54879 -56090 54976 -56074
rect 54879 -56128 54926 -56090
rect 54960 -56128 54976 -56090
rect 54879 -56144 54976 -56128
rect 55318 -56168 55384 -56152
rect 55318 -56202 55334 -56168
rect 55368 -56202 55384 -56168
rect 55318 -56218 55384 -56202
rect 55336 -56240 55366 -56218
rect 55336 -56466 55366 -56440
rect 53510 -57016 53630 -56978
rect 53510 -57050 53526 -57016
rect 53614 -57050 53630 -57016
rect 53510 -57066 53630 -57050
rect 53842 -56840 53930 -56824
rect 53842 -56928 53858 -56840
rect 53892 -56928 53930 -56840
rect 53842 -56944 53930 -56928
rect 54730 -56840 54818 -56824
rect 54730 -56928 54768 -56840
rect 54802 -56928 54818 -56840
rect 54730 -56944 54818 -56928
rect 55030 -56759 55096 -56744
rect 55540 -56759 55606 -56744
rect 55030 -56760 55118 -56759
rect 55030 -56794 55046 -56760
rect 55080 -56794 55118 -56760
rect 55030 -56795 55118 -56794
rect 55518 -56760 55606 -56759
rect 55518 -56794 55556 -56760
rect 55590 -56794 55606 -56760
rect 55518 -56795 55606 -56794
rect 55030 -56810 55096 -56795
rect 55540 -56810 55606 -56795
rect 55866 -56056 55986 -56040
rect 55866 -56090 55882 -56056
rect 55970 -56090 55986 -56056
rect 55866 -56128 55986 -56090
rect 55866 -56966 55986 -56928
rect 55866 -57000 55882 -56966
rect 55970 -57000 55986 -56966
rect 55866 -57016 55986 -57000
rect 57175 -56109 57205 -56083
rect 57263 -56109 57293 -56083
rect 57175 -56282 57205 -56267
rect 57169 -56306 57205 -56282
rect 57169 -56341 57199 -56306
rect 57263 -56328 57293 -56267
rect 59544 -56093 59610 -56085
rect 59087 -56143 59113 -56093
rect 59513 -56101 59610 -56093
rect 59513 -56135 59560 -56101
rect 59594 -56135 59610 -56101
rect 59513 -56143 59610 -56135
rect 59544 -56151 59610 -56143
rect 59016 -56201 59082 -56193
rect 59016 -56209 59113 -56201
rect 59016 -56243 59032 -56209
rect 59066 -56243 59113 -56209
rect 59016 -56251 59113 -56243
rect 59513 -56251 59539 -56201
rect 59016 -56259 59082 -56251
rect 57123 -56357 57199 -56341
rect 57123 -56391 57133 -56357
rect 57167 -56391 57199 -56357
rect 57123 -56407 57199 -56391
rect 57241 -56344 57295 -56328
rect 57241 -56378 57251 -56344
rect 57285 -56378 57295 -56344
rect 57241 -56394 57295 -56378
rect 57169 -56416 57199 -56407
rect 57169 -56440 57205 -56416
rect 57175 -56455 57205 -56440
rect 57263 -56455 57293 -56394
rect 53510 -57124 53630 -57108
rect 53510 -57158 53526 -57124
rect 53614 -57158 53630 -57124
rect 53510 -57196 53630 -57158
rect 53842 -57246 53930 -57230
rect 53842 -57334 53858 -57246
rect 53892 -57334 53930 -57246
rect 53842 -57350 53930 -57334
rect 54730 -57246 54818 -57230
rect 54730 -57334 54768 -57246
rect 54802 -57334 54818 -57246
rect 54730 -57350 54818 -57334
rect 55030 -57381 55096 -57366
rect 55540 -57381 55606 -57366
rect 55030 -57382 55118 -57381
rect 55030 -57416 55046 -57382
rect 55080 -57416 55118 -57382
rect 55030 -57417 55118 -57416
rect 55518 -57382 55606 -57381
rect 55518 -57416 55556 -57382
rect 55590 -57416 55606 -57382
rect 55518 -57417 55606 -57416
rect 55030 -57432 55096 -57417
rect 53510 -58034 53630 -57996
rect 53510 -58068 53526 -58034
rect 53614 -58068 53630 -58034
rect 53510 -58084 53630 -58068
rect 55540 -57432 55606 -57417
rect 53972 -58050 54069 -58034
rect 53972 -58088 53988 -58050
rect 54022 -58088 54069 -58050
rect 53972 -58104 54069 -58088
rect 54869 -58050 54966 -58034
rect 54869 -58088 54916 -58050
rect 54950 -58088 54966 -58050
rect 54869 -58104 54966 -58088
rect 55326 -57736 55356 -57710
rect 55326 -57958 55356 -57936
rect 55308 -57974 55374 -57958
rect 55308 -58008 55324 -57974
rect 55358 -58008 55374 -57974
rect 55308 -58024 55374 -58008
rect 55866 -57170 55986 -57154
rect 55866 -57204 55882 -57170
rect 55970 -57204 55986 -57170
rect 55866 -57242 55986 -57204
rect 55866 -58080 55986 -58042
rect 55866 -58114 55882 -58080
rect 55970 -58114 55986 -58080
rect 55866 -58130 55986 -58114
rect 56476 -56606 56546 -56590
rect 56476 -56640 56492 -56606
rect 56530 -56640 56546 -56606
rect 56476 -56687 56546 -56640
rect 57175 -56585 57205 -56559
rect 57263 -56585 57293 -56559
rect 56476 -57534 56546 -57487
rect 56476 -57568 56492 -57534
rect 56530 -57568 56546 -57534
rect 56476 -57584 56546 -57568
rect 59087 -56478 59153 -56462
rect 59087 -56512 59103 -56478
rect 59137 -56512 59153 -56478
rect 59087 -56528 59153 -56512
rect 59090 -56559 59150 -56528
rect 59090 -56990 59150 -56959
rect 59087 -57006 59153 -56990
rect 59087 -57040 59103 -57006
rect 59137 -57040 59153 -57006
rect 59087 -57056 59153 -57040
rect 59858 -56420 59924 -56412
rect 60368 -56420 60434 -56412
rect 59858 -56428 59946 -56420
rect 59858 -56462 59874 -56428
rect 59908 -56462 59946 -56428
rect 59858 -56470 59946 -56462
rect 60346 -56428 60434 -56420
rect 60346 -56462 60384 -56428
rect 60418 -56462 60434 -56428
rect 60346 -56470 60434 -56462
rect 59858 -56478 59924 -56470
rect 60368 -56478 60434 -56470
rect 59530 -56698 59596 -56682
rect 59530 -56732 59546 -56698
rect 59580 -56732 59596 -56698
rect 59530 -56748 59596 -56732
rect 59548 -56770 59578 -56748
rect 59548 -56992 59578 -56970
rect 59530 -57008 59596 -56992
rect 59530 -57042 59546 -57008
rect 59580 -57042 59596 -57008
rect 59530 -57058 59596 -57042
rect 59846 -56698 59912 -56682
rect 59846 -56732 59862 -56698
rect 59896 -56732 59912 -56698
rect 59846 -56748 59912 -56732
rect 59864 -56770 59894 -56748
rect 59864 -56992 59894 -56970
rect 59846 -57008 59912 -56992
rect 59846 -57042 59862 -57008
rect 59896 -57042 59912 -57008
rect 59846 -57058 59912 -57042
rect 60343 -56965 60409 -56949
rect 61043 -56965 61109 -56949
rect 60343 -56999 60359 -56965
rect 60393 -56999 60409 -56965
rect 60343 -57017 60409 -56999
rect 61043 -56999 61059 -56965
rect 61093 -56999 61109 -56965
rect 61043 -57017 61109 -56999
rect 60165 -57047 60191 -57017
rect 60321 -57047 60441 -57017
rect 60641 -57047 60667 -57017
rect 60785 -57047 60811 -57017
rect 61011 -57047 61131 -57017
rect 61261 -57047 61287 -57017
rect 60343 -57057 60409 -57047
rect 60343 -57091 60359 -57057
rect 60393 -57091 60409 -57057
rect 60343 -57101 60409 -57091
rect 61043 -57057 61109 -57047
rect 61043 -57091 61059 -57057
rect 61093 -57091 61109 -57057
rect 61043 -57101 61109 -57091
rect 57175 -57629 57205 -57603
rect 57263 -57629 57293 -57603
rect 57175 -57748 57205 -57733
rect 57169 -57772 57205 -57748
rect 57169 -57781 57199 -57772
rect 57123 -57797 57199 -57781
rect 57263 -57794 57293 -57733
rect 59087 -57208 59153 -57192
rect 59087 -57242 59103 -57208
rect 59137 -57242 59153 -57208
rect 59087 -57258 59153 -57242
rect 59090 -57289 59150 -57258
rect 59090 -57720 59150 -57689
rect 57123 -57831 57133 -57797
rect 57167 -57831 57199 -57797
rect 57123 -57847 57199 -57831
rect 57169 -57882 57199 -57847
rect 57241 -57810 57295 -57794
rect 57241 -57844 57251 -57810
rect 57285 -57844 57295 -57810
rect 57241 -57860 57295 -57844
rect 59087 -57736 59153 -57720
rect 59087 -57770 59103 -57736
rect 59137 -57770 59153 -57736
rect 59087 -57786 59153 -57770
rect 60165 -57131 60191 -57101
rect 60321 -57131 60441 -57101
rect 60641 -57131 60667 -57101
rect 60785 -57131 60811 -57101
rect 61011 -57131 61131 -57101
rect 61261 -57131 61287 -57101
rect 59526 -57211 59596 -57180
rect 59526 -57230 59545 -57211
rect 59529 -57245 59545 -57230
rect 59579 -57230 59596 -57211
rect 59579 -57245 59595 -57230
rect 59529 -57261 59595 -57245
rect 59547 -57283 59577 -57261
rect 59547 -57505 59577 -57483
rect 59529 -57521 59595 -57505
rect 59529 -57555 59545 -57521
rect 59579 -57555 59595 -57521
rect 59529 -57571 59595 -57555
rect 59845 -57211 59911 -57195
rect 59845 -57245 59861 -57211
rect 59895 -57245 59911 -57211
rect 59845 -57261 59911 -57245
rect 60343 -57141 60409 -57131
rect 60343 -57175 60359 -57141
rect 60393 -57175 60409 -57141
rect 60343 -57185 60409 -57175
rect 61043 -57141 61109 -57131
rect 61043 -57175 61059 -57141
rect 61093 -57175 61109 -57141
rect 61043 -57185 61109 -57175
rect 59863 -57283 59893 -57261
rect 59863 -57505 59893 -57483
rect 59845 -57521 59911 -57505
rect 59845 -57555 59861 -57521
rect 59895 -57555 59911 -57521
rect 59845 -57571 59911 -57555
rect 60165 -57215 60191 -57185
rect 60321 -57215 60441 -57185
rect 60641 -57215 60667 -57185
rect 60785 -57215 60811 -57185
rect 61011 -57215 61131 -57185
rect 61261 -57215 61287 -57185
rect 60343 -57225 60409 -57215
rect 60343 -57259 60359 -57225
rect 60393 -57259 60409 -57225
rect 60343 -57269 60409 -57259
rect 61043 -57225 61109 -57215
rect 61043 -57259 61059 -57225
rect 61093 -57259 61109 -57225
rect 61043 -57269 61109 -57259
rect 60165 -57299 60191 -57269
rect 60321 -57299 60441 -57269
rect 60641 -57299 60667 -57269
rect 60785 -57299 60811 -57269
rect 61011 -57299 61131 -57269
rect 61261 -57299 61287 -57269
rect 57169 -57906 57205 -57882
rect 57175 -57921 57205 -57906
rect 57263 -57921 57293 -57860
rect 57175 -58105 57205 -58079
rect 57263 -58105 57293 -58079
rect 59544 -58000 59610 -57992
rect 59087 -58050 59113 -58000
rect 59513 -58008 59610 -58000
rect 59513 -58042 59560 -58008
rect 59594 -58042 59610 -58008
rect 59513 -58050 59610 -58042
rect 59544 -58058 59610 -58050
rect 59016 -58108 59082 -58100
rect 59016 -58116 59113 -58108
rect 59016 -58150 59032 -58116
rect 59066 -58150 59113 -58116
rect 59016 -58158 59113 -58150
rect 59513 -58158 59539 -58108
rect 59016 -58166 59082 -58158
rect 53972 -58406 54069 -58390
rect 53972 -58444 53988 -58406
rect 54022 -58444 54069 -58406
rect 53972 -58460 54069 -58444
rect 54869 -58406 54966 -58390
rect 54869 -58444 54916 -58406
rect 54950 -58444 54966 -58406
rect 54869 -58460 54966 -58444
rect 59858 -57786 59924 -57778
rect 60368 -57786 60434 -57778
rect 59858 -57794 59946 -57786
rect 59858 -57828 59874 -57794
rect 59908 -57828 59946 -57794
rect 59858 -57836 59946 -57828
rect 60346 -57794 60434 -57786
rect 60346 -57828 60384 -57794
rect 60418 -57828 60434 -57794
rect 60346 -57836 60434 -57828
rect 59858 -57844 59924 -57836
rect 60368 -57844 60434 -57836
rect 55510 -58602 55576 -58586
rect 55510 -58604 55526 -58602
rect 55262 -58634 55288 -58604
rect 55488 -58634 55526 -58604
rect 55510 -58636 55526 -58634
rect 55560 -58636 55576 -58602
rect 55510 -58652 55576 -58636
rect 53982 -61134 54079 -61118
rect 53982 -61172 53998 -61134
rect 54032 -61172 54079 -61134
rect 53982 -61188 54079 -61172
rect 54879 -61134 54976 -61118
rect 54879 -61172 54926 -61134
rect 54960 -61172 54976 -61134
rect 54879 -61188 54976 -61172
rect 53510 -61506 53630 -61490
rect 53510 -61540 53526 -61506
rect 53614 -61540 53630 -61506
rect 53510 -61578 53630 -61540
rect 53982 -61490 54079 -61474
rect 53982 -61528 53998 -61490
rect 54032 -61528 54079 -61490
rect 53982 -61544 54079 -61528
rect 54879 -61490 54976 -61474
rect 54879 -61528 54926 -61490
rect 54960 -61528 54976 -61490
rect 54879 -61544 54976 -61528
rect 55318 -61568 55384 -61552
rect 55318 -61602 55334 -61568
rect 55368 -61602 55384 -61568
rect 55318 -61618 55384 -61602
rect 55336 -61640 55366 -61618
rect 55336 -61866 55366 -61840
rect 53510 -62416 53630 -62378
rect 53510 -62450 53526 -62416
rect 53614 -62450 53630 -62416
rect 53510 -62466 53630 -62450
rect 53842 -62240 53930 -62224
rect 53842 -62328 53858 -62240
rect 53892 -62328 53930 -62240
rect 53842 -62344 53930 -62328
rect 54730 -62240 54818 -62224
rect 54730 -62328 54768 -62240
rect 54802 -62328 54818 -62240
rect 54730 -62344 54818 -62328
rect 55030 -62159 55096 -62144
rect 55540 -62159 55606 -62144
rect 55030 -62160 55118 -62159
rect 55030 -62194 55046 -62160
rect 55080 -62194 55118 -62160
rect 55030 -62195 55118 -62194
rect 55518 -62160 55606 -62159
rect 55518 -62194 55556 -62160
rect 55590 -62194 55606 -62160
rect 55518 -62195 55606 -62194
rect 55030 -62210 55096 -62195
rect 55540 -62210 55606 -62195
rect 55866 -61456 55986 -61440
rect 55866 -61490 55882 -61456
rect 55970 -61490 55986 -61456
rect 55866 -61528 55986 -61490
rect 55866 -62366 55986 -62328
rect 55866 -62400 55882 -62366
rect 55970 -62400 55986 -62366
rect 55866 -62416 55986 -62400
rect 57175 -61509 57205 -61483
rect 57263 -61509 57293 -61483
rect 57175 -61682 57205 -61667
rect 57169 -61706 57205 -61682
rect 57169 -61741 57199 -61706
rect 57263 -61728 57293 -61667
rect 59544 -61493 59610 -61485
rect 59087 -61543 59113 -61493
rect 59513 -61501 59610 -61493
rect 59513 -61535 59560 -61501
rect 59594 -61535 59610 -61501
rect 59513 -61543 59610 -61535
rect 59544 -61551 59610 -61543
rect 59016 -61601 59082 -61593
rect 59016 -61609 59113 -61601
rect 59016 -61643 59032 -61609
rect 59066 -61643 59113 -61609
rect 59016 -61651 59113 -61643
rect 59513 -61651 59539 -61601
rect 59016 -61659 59082 -61651
rect 57123 -61757 57199 -61741
rect 57123 -61791 57133 -61757
rect 57167 -61791 57199 -61757
rect 57123 -61807 57199 -61791
rect 57241 -61744 57295 -61728
rect 57241 -61778 57251 -61744
rect 57285 -61778 57295 -61744
rect 57241 -61794 57295 -61778
rect 57169 -61816 57199 -61807
rect 57169 -61840 57205 -61816
rect 57175 -61855 57205 -61840
rect 57263 -61855 57293 -61794
rect 53510 -62524 53630 -62508
rect 53510 -62558 53526 -62524
rect 53614 -62558 53630 -62524
rect 53510 -62596 53630 -62558
rect 53842 -62646 53930 -62630
rect 53842 -62734 53858 -62646
rect 53892 -62734 53930 -62646
rect 53842 -62750 53930 -62734
rect 54730 -62646 54818 -62630
rect 54730 -62734 54768 -62646
rect 54802 -62734 54818 -62646
rect 54730 -62750 54818 -62734
rect 55030 -62781 55096 -62766
rect 55540 -62781 55606 -62766
rect 55030 -62782 55118 -62781
rect 55030 -62816 55046 -62782
rect 55080 -62816 55118 -62782
rect 55030 -62817 55118 -62816
rect 55518 -62782 55606 -62781
rect 55518 -62816 55556 -62782
rect 55590 -62816 55606 -62782
rect 55518 -62817 55606 -62816
rect 55030 -62832 55096 -62817
rect 53510 -63434 53630 -63396
rect 53510 -63468 53526 -63434
rect 53614 -63468 53630 -63434
rect 53510 -63484 53630 -63468
rect 55540 -62832 55606 -62817
rect 53972 -63450 54069 -63434
rect 53972 -63488 53988 -63450
rect 54022 -63488 54069 -63450
rect 53972 -63504 54069 -63488
rect 54869 -63450 54966 -63434
rect 54869 -63488 54916 -63450
rect 54950 -63488 54966 -63450
rect 54869 -63504 54966 -63488
rect 55326 -63136 55356 -63110
rect 55326 -63358 55356 -63336
rect 55308 -63374 55374 -63358
rect 55308 -63408 55324 -63374
rect 55358 -63408 55374 -63374
rect 55308 -63424 55374 -63408
rect 55866 -62570 55986 -62554
rect 55866 -62604 55882 -62570
rect 55970 -62604 55986 -62570
rect 55866 -62642 55986 -62604
rect 55866 -63480 55986 -63442
rect 55866 -63514 55882 -63480
rect 55970 -63514 55986 -63480
rect 55866 -63530 55986 -63514
rect 56476 -62006 56546 -61990
rect 56476 -62040 56492 -62006
rect 56530 -62040 56546 -62006
rect 56476 -62087 56546 -62040
rect 57175 -61985 57205 -61959
rect 57263 -61985 57293 -61959
rect 56476 -62934 56546 -62887
rect 56476 -62968 56492 -62934
rect 56530 -62968 56546 -62934
rect 56476 -62984 56546 -62968
rect 59087 -61878 59153 -61862
rect 59087 -61912 59103 -61878
rect 59137 -61912 59153 -61878
rect 59087 -61928 59153 -61912
rect 59090 -61959 59150 -61928
rect 59090 -62390 59150 -62359
rect 59087 -62406 59153 -62390
rect 59087 -62440 59103 -62406
rect 59137 -62440 59153 -62406
rect 59087 -62456 59153 -62440
rect 59858 -61820 59924 -61812
rect 60368 -61820 60434 -61812
rect 59858 -61828 59946 -61820
rect 59858 -61862 59874 -61828
rect 59908 -61862 59946 -61828
rect 59858 -61870 59946 -61862
rect 60346 -61828 60434 -61820
rect 60346 -61862 60384 -61828
rect 60418 -61862 60434 -61828
rect 60346 -61870 60434 -61862
rect 59858 -61878 59924 -61870
rect 60368 -61878 60434 -61870
rect 59530 -62098 59596 -62082
rect 59530 -62132 59546 -62098
rect 59580 -62132 59596 -62098
rect 59530 -62148 59596 -62132
rect 59548 -62170 59578 -62148
rect 59548 -62392 59578 -62370
rect 59530 -62408 59596 -62392
rect 59530 -62442 59546 -62408
rect 59580 -62442 59596 -62408
rect 59530 -62458 59596 -62442
rect 59846 -62098 59912 -62082
rect 59846 -62132 59862 -62098
rect 59896 -62132 59912 -62098
rect 59846 -62148 59912 -62132
rect 59864 -62170 59894 -62148
rect 59864 -62392 59894 -62370
rect 59846 -62408 59912 -62392
rect 59846 -62442 59862 -62408
rect 59896 -62442 59912 -62408
rect 59846 -62458 59912 -62442
rect 60343 -62365 60409 -62349
rect 61043 -62365 61109 -62349
rect 60343 -62399 60359 -62365
rect 60393 -62399 60409 -62365
rect 60343 -62417 60409 -62399
rect 61043 -62399 61059 -62365
rect 61093 -62399 61109 -62365
rect 61043 -62417 61109 -62399
rect 60165 -62447 60191 -62417
rect 60321 -62447 60441 -62417
rect 60641 -62447 60667 -62417
rect 60785 -62447 60811 -62417
rect 61011 -62447 61131 -62417
rect 61261 -62447 61287 -62417
rect 60343 -62457 60409 -62447
rect 60343 -62491 60359 -62457
rect 60393 -62491 60409 -62457
rect 60343 -62501 60409 -62491
rect 61043 -62457 61109 -62447
rect 61043 -62491 61059 -62457
rect 61093 -62491 61109 -62457
rect 61043 -62501 61109 -62491
rect 57175 -63029 57205 -63003
rect 57263 -63029 57293 -63003
rect 57175 -63148 57205 -63133
rect 57169 -63172 57205 -63148
rect 57169 -63181 57199 -63172
rect 57123 -63197 57199 -63181
rect 57263 -63194 57293 -63133
rect 59087 -62608 59153 -62592
rect 59087 -62642 59103 -62608
rect 59137 -62642 59153 -62608
rect 59087 -62658 59153 -62642
rect 59090 -62689 59150 -62658
rect 59090 -63120 59150 -63089
rect 57123 -63231 57133 -63197
rect 57167 -63231 57199 -63197
rect 57123 -63247 57199 -63231
rect 57169 -63282 57199 -63247
rect 57241 -63210 57295 -63194
rect 57241 -63244 57251 -63210
rect 57285 -63244 57295 -63210
rect 57241 -63260 57295 -63244
rect 59087 -63136 59153 -63120
rect 59087 -63170 59103 -63136
rect 59137 -63170 59153 -63136
rect 59087 -63186 59153 -63170
rect 60165 -62531 60191 -62501
rect 60321 -62531 60441 -62501
rect 60641 -62531 60667 -62501
rect 60785 -62531 60811 -62501
rect 61011 -62531 61131 -62501
rect 61261 -62531 61287 -62501
rect 59526 -62611 59596 -62580
rect 59526 -62630 59545 -62611
rect 59529 -62645 59545 -62630
rect 59579 -62630 59596 -62611
rect 59579 -62645 59595 -62630
rect 59529 -62661 59595 -62645
rect 59547 -62683 59577 -62661
rect 59547 -62905 59577 -62883
rect 59529 -62921 59595 -62905
rect 59529 -62955 59545 -62921
rect 59579 -62955 59595 -62921
rect 59529 -62971 59595 -62955
rect 59845 -62611 59911 -62595
rect 59845 -62645 59861 -62611
rect 59895 -62645 59911 -62611
rect 59845 -62661 59911 -62645
rect 60343 -62541 60409 -62531
rect 60343 -62575 60359 -62541
rect 60393 -62575 60409 -62541
rect 60343 -62585 60409 -62575
rect 61043 -62541 61109 -62531
rect 61043 -62575 61059 -62541
rect 61093 -62575 61109 -62541
rect 61043 -62585 61109 -62575
rect 59863 -62683 59893 -62661
rect 59863 -62905 59893 -62883
rect 59845 -62921 59911 -62905
rect 59845 -62955 59861 -62921
rect 59895 -62955 59911 -62921
rect 59845 -62971 59911 -62955
rect 60165 -62615 60191 -62585
rect 60321 -62615 60441 -62585
rect 60641 -62615 60667 -62585
rect 60785 -62615 60811 -62585
rect 61011 -62615 61131 -62585
rect 61261 -62615 61287 -62585
rect 60343 -62625 60409 -62615
rect 60343 -62659 60359 -62625
rect 60393 -62659 60409 -62625
rect 60343 -62669 60409 -62659
rect 61043 -62625 61109 -62615
rect 61043 -62659 61059 -62625
rect 61093 -62659 61109 -62625
rect 61043 -62669 61109 -62659
rect 60165 -62699 60191 -62669
rect 60321 -62699 60441 -62669
rect 60641 -62699 60667 -62669
rect 60785 -62699 60811 -62669
rect 61011 -62699 61131 -62669
rect 61261 -62699 61287 -62669
rect 57169 -63306 57205 -63282
rect 57175 -63321 57205 -63306
rect 57263 -63321 57293 -63260
rect 57175 -63505 57205 -63479
rect 57263 -63505 57293 -63479
rect 59544 -63400 59610 -63392
rect 59087 -63450 59113 -63400
rect 59513 -63408 59610 -63400
rect 59513 -63442 59560 -63408
rect 59594 -63442 59610 -63408
rect 59513 -63450 59610 -63442
rect 59544 -63458 59610 -63450
rect 59016 -63508 59082 -63500
rect 59016 -63516 59113 -63508
rect 59016 -63550 59032 -63516
rect 59066 -63550 59113 -63516
rect 59016 -63558 59113 -63550
rect 59513 -63558 59539 -63508
rect 59016 -63566 59082 -63558
rect 53972 -63806 54069 -63790
rect 53972 -63844 53988 -63806
rect 54022 -63844 54069 -63806
rect 53972 -63860 54069 -63844
rect 54869 -63806 54966 -63790
rect 54869 -63844 54916 -63806
rect 54950 -63844 54966 -63806
rect 54869 -63860 54966 -63844
rect 59858 -63186 59924 -63178
rect 60368 -63186 60434 -63178
rect 59858 -63194 59946 -63186
rect 59858 -63228 59874 -63194
rect 59908 -63228 59946 -63194
rect 59858 -63236 59946 -63228
rect 60346 -63194 60434 -63186
rect 60346 -63228 60384 -63194
rect 60418 -63228 60434 -63194
rect 60346 -63236 60434 -63228
rect 59858 -63244 59924 -63236
rect 60368 -63244 60434 -63236
rect 55510 -64002 55576 -63986
rect 55510 -64004 55526 -64002
rect 55262 -64034 55288 -64004
rect 55488 -64034 55526 -64004
rect 55510 -64036 55526 -64034
rect 55560 -64036 55576 -64002
rect 55510 -64052 55576 -64036
rect 53982 -66534 54079 -66518
rect 53982 -66572 53998 -66534
rect 54032 -66572 54079 -66534
rect 53982 -66588 54079 -66572
rect 54879 -66534 54976 -66518
rect 54879 -66572 54926 -66534
rect 54960 -66572 54976 -66534
rect 54879 -66588 54976 -66572
rect 53510 -66906 53630 -66890
rect 53510 -66940 53526 -66906
rect 53614 -66940 53630 -66906
rect 53510 -66978 53630 -66940
rect 53982 -66890 54079 -66874
rect 53982 -66928 53998 -66890
rect 54032 -66928 54079 -66890
rect 53982 -66944 54079 -66928
rect 54879 -66890 54976 -66874
rect 54879 -66928 54926 -66890
rect 54960 -66928 54976 -66890
rect 54879 -66944 54976 -66928
rect 55318 -66968 55384 -66952
rect 55318 -67002 55334 -66968
rect 55368 -67002 55384 -66968
rect 55318 -67018 55384 -67002
rect 55336 -67040 55366 -67018
rect 55336 -67266 55366 -67240
rect 53510 -67816 53630 -67778
rect 53510 -67850 53526 -67816
rect 53614 -67850 53630 -67816
rect 53510 -67866 53630 -67850
rect 53842 -67640 53930 -67624
rect 53842 -67728 53858 -67640
rect 53892 -67728 53930 -67640
rect 53842 -67744 53930 -67728
rect 54730 -67640 54818 -67624
rect 54730 -67728 54768 -67640
rect 54802 -67728 54818 -67640
rect 54730 -67744 54818 -67728
rect 55030 -67559 55096 -67544
rect 55540 -67559 55606 -67544
rect 55030 -67560 55118 -67559
rect 55030 -67594 55046 -67560
rect 55080 -67594 55118 -67560
rect 55030 -67595 55118 -67594
rect 55518 -67560 55606 -67559
rect 55518 -67594 55556 -67560
rect 55590 -67594 55606 -67560
rect 55518 -67595 55606 -67594
rect 55030 -67610 55096 -67595
rect 55540 -67610 55606 -67595
rect 55866 -66856 55986 -66840
rect 55866 -66890 55882 -66856
rect 55970 -66890 55986 -66856
rect 55866 -66928 55986 -66890
rect 55866 -67766 55986 -67728
rect 55866 -67800 55882 -67766
rect 55970 -67800 55986 -67766
rect 55866 -67816 55986 -67800
rect 57175 -66909 57205 -66883
rect 57263 -66909 57293 -66883
rect 57175 -67082 57205 -67067
rect 57169 -67106 57205 -67082
rect 57169 -67141 57199 -67106
rect 57263 -67128 57293 -67067
rect 59544 -66893 59610 -66885
rect 59087 -66943 59113 -66893
rect 59513 -66901 59610 -66893
rect 59513 -66935 59560 -66901
rect 59594 -66935 59610 -66901
rect 59513 -66943 59610 -66935
rect 59544 -66951 59610 -66943
rect 59016 -67001 59082 -66993
rect 59016 -67009 59113 -67001
rect 59016 -67043 59032 -67009
rect 59066 -67043 59113 -67009
rect 59016 -67051 59113 -67043
rect 59513 -67051 59539 -67001
rect 59016 -67059 59082 -67051
rect 57123 -67157 57199 -67141
rect 57123 -67191 57133 -67157
rect 57167 -67191 57199 -67157
rect 57123 -67207 57199 -67191
rect 57241 -67144 57295 -67128
rect 57241 -67178 57251 -67144
rect 57285 -67178 57295 -67144
rect 57241 -67194 57295 -67178
rect 57169 -67216 57199 -67207
rect 57169 -67240 57205 -67216
rect 57175 -67255 57205 -67240
rect 57263 -67255 57293 -67194
rect 53510 -67924 53630 -67908
rect 53510 -67958 53526 -67924
rect 53614 -67958 53630 -67924
rect 53510 -67996 53630 -67958
rect 53842 -68046 53930 -68030
rect 53842 -68134 53858 -68046
rect 53892 -68134 53930 -68046
rect 53842 -68150 53930 -68134
rect 54730 -68046 54818 -68030
rect 54730 -68134 54768 -68046
rect 54802 -68134 54818 -68046
rect 54730 -68150 54818 -68134
rect 55030 -68181 55096 -68166
rect 55540 -68181 55606 -68166
rect 55030 -68182 55118 -68181
rect 55030 -68216 55046 -68182
rect 55080 -68216 55118 -68182
rect 55030 -68217 55118 -68216
rect 55518 -68182 55606 -68181
rect 55518 -68216 55556 -68182
rect 55590 -68216 55606 -68182
rect 55518 -68217 55606 -68216
rect 55030 -68232 55096 -68217
rect 53510 -68834 53630 -68796
rect 53510 -68868 53526 -68834
rect 53614 -68868 53630 -68834
rect 53510 -68884 53630 -68868
rect 55540 -68232 55606 -68217
rect 53972 -68850 54069 -68834
rect 53972 -68888 53988 -68850
rect 54022 -68888 54069 -68850
rect 53972 -68904 54069 -68888
rect 54869 -68850 54966 -68834
rect 54869 -68888 54916 -68850
rect 54950 -68888 54966 -68850
rect 54869 -68904 54966 -68888
rect 55326 -68536 55356 -68510
rect 55326 -68758 55356 -68736
rect 55308 -68774 55374 -68758
rect 55308 -68808 55324 -68774
rect 55358 -68808 55374 -68774
rect 55308 -68824 55374 -68808
rect 55866 -67970 55986 -67954
rect 55866 -68004 55882 -67970
rect 55970 -68004 55986 -67970
rect 55866 -68042 55986 -68004
rect 55866 -68880 55986 -68842
rect 55866 -68914 55882 -68880
rect 55970 -68914 55986 -68880
rect 55866 -68930 55986 -68914
rect 56476 -67406 56546 -67390
rect 56476 -67440 56492 -67406
rect 56530 -67440 56546 -67406
rect 56476 -67487 56546 -67440
rect 57175 -67385 57205 -67359
rect 57263 -67385 57293 -67359
rect 56476 -68334 56546 -68287
rect 56476 -68368 56492 -68334
rect 56530 -68368 56546 -68334
rect 56476 -68384 56546 -68368
rect 59087 -67278 59153 -67262
rect 59087 -67312 59103 -67278
rect 59137 -67312 59153 -67278
rect 59087 -67328 59153 -67312
rect 59090 -67359 59150 -67328
rect 59090 -67790 59150 -67759
rect 59087 -67806 59153 -67790
rect 59087 -67840 59103 -67806
rect 59137 -67840 59153 -67806
rect 59087 -67856 59153 -67840
rect 59858 -67220 59924 -67212
rect 60368 -67220 60434 -67212
rect 59858 -67228 59946 -67220
rect 59858 -67262 59874 -67228
rect 59908 -67262 59946 -67228
rect 59858 -67270 59946 -67262
rect 60346 -67228 60434 -67220
rect 60346 -67262 60384 -67228
rect 60418 -67262 60434 -67228
rect 60346 -67270 60434 -67262
rect 59858 -67278 59924 -67270
rect 60368 -67278 60434 -67270
rect 59530 -67498 59596 -67482
rect 59530 -67532 59546 -67498
rect 59580 -67532 59596 -67498
rect 59530 -67548 59596 -67532
rect 59548 -67570 59578 -67548
rect 59548 -67792 59578 -67770
rect 59530 -67808 59596 -67792
rect 59530 -67842 59546 -67808
rect 59580 -67842 59596 -67808
rect 59530 -67858 59596 -67842
rect 59846 -67498 59912 -67482
rect 59846 -67532 59862 -67498
rect 59896 -67532 59912 -67498
rect 59846 -67548 59912 -67532
rect 59864 -67570 59894 -67548
rect 59864 -67792 59894 -67770
rect 59846 -67808 59912 -67792
rect 59846 -67842 59862 -67808
rect 59896 -67842 59912 -67808
rect 59846 -67858 59912 -67842
rect 60343 -67765 60409 -67749
rect 61043 -67765 61109 -67749
rect 60343 -67799 60359 -67765
rect 60393 -67799 60409 -67765
rect 60343 -67817 60409 -67799
rect 61043 -67799 61059 -67765
rect 61093 -67799 61109 -67765
rect 61043 -67817 61109 -67799
rect 60165 -67847 60191 -67817
rect 60321 -67847 60441 -67817
rect 60641 -67847 60667 -67817
rect 60785 -67847 60811 -67817
rect 61011 -67847 61131 -67817
rect 61261 -67847 61287 -67817
rect 60343 -67857 60409 -67847
rect 60343 -67891 60359 -67857
rect 60393 -67891 60409 -67857
rect 60343 -67901 60409 -67891
rect 61043 -67857 61109 -67847
rect 61043 -67891 61059 -67857
rect 61093 -67891 61109 -67857
rect 61043 -67901 61109 -67891
rect 57175 -68429 57205 -68403
rect 57263 -68429 57293 -68403
rect 57175 -68548 57205 -68533
rect 57169 -68572 57205 -68548
rect 57169 -68581 57199 -68572
rect 57123 -68597 57199 -68581
rect 57263 -68594 57293 -68533
rect 59087 -68008 59153 -67992
rect 59087 -68042 59103 -68008
rect 59137 -68042 59153 -68008
rect 59087 -68058 59153 -68042
rect 59090 -68089 59150 -68058
rect 59090 -68520 59150 -68489
rect 57123 -68631 57133 -68597
rect 57167 -68631 57199 -68597
rect 57123 -68647 57199 -68631
rect 57169 -68682 57199 -68647
rect 57241 -68610 57295 -68594
rect 57241 -68644 57251 -68610
rect 57285 -68644 57295 -68610
rect 57241 -68660 57295 -68644
rect 59087 -68536 59153 -68520
rect 59087 -68570 59103 -68536
rect 59137 -68570 59153 -68536
rect 59087 -68586 59153 -68570
rect 60165 -67931 60191 -67901
rect 60321 -67931 60441 -67901
rect 60641 -67931 60667 -67901
rect 60785 -67931 60811 -67901
rect 61011 -67931 61131 -67901
rect 61261 -67931 61287 -67901
rect 59526 -68011 59596 -67980
rect 59526 -68030 59545 -68011
rect 59529 -68045 59545 -68030
rect 59579 -68030 59596 -68011
rect 59579 -68045 59595 -68030
rect 59529 -68061 59595 -68045
rect 59547 -68083 59577 -68061
rect 59547 -68305 59577 -68283
rect 59529 -68321 59595 -68305
rect 59529 -68355 59545 -68321
rect 59579 -68355 59595 -68321
rect 59529 -68371 59595 -68355
rect 59845 -68011 59911 -67995
rect 59845 -68045 59861 -68011
rect 59895 -68045 59911 -68011
rect 59845 -68061 59911 -68045
rect 60343 -67941 60409 -67931
rect 60343 -67975 60359 -67941
rect 60393 -67975 60409 -67941
rect 60343 -67985 60409 -67975
rect 61043 -67941 61109 -67931
rect 61043 -67975 61059 -67941
rect 61093 -67975 61109 -67941
rect 61043 -67985 61109 -67975
rect 59863 -68083 59893 -68061
rect 59863 -68305 59893 -68283
rect 59845 -68321 59911 -68305
rect 59845 -68355 59861 -68321
rect 59895 -68355 59911 -68321
rect 59845 -68371 59911 -68355
rect 60165 -68015 60191 -67985
rect 60321 -68015 60441 -67985
rect 60641 -68015 60667 -67985
rect 60785 -68015 60811 -67985
rect 61011 -68015 61131 -67985
rect 61261 -68015 61287 -67985
rect 60343 -68025 60409 -68015
rect 60343 -68059 60359 -68025
rect 60393 -68059 60409 -68025
rect 60343 -68069 60409 -68059
rect 61043 -68025 61109 -68015
rect 61043 -68059 61059 -68025
rect 61093 -68059 61109 -68025
rect 61043 -68069 61109 -68059
rect 60165 -68099 60191 -68069
rect 60321 -68099 60441 -68069
rect 60641 -68099 60667 -68069
rect 60785 -68099 60811 -68069
rect 61011 -68099 61131 -68069
rect 61261 -68099 61287 -68069
rect 57169 -68706 57205 -68682
rect 57175 -68721 57205 -68706
rect 57263 -68721 57293 -68660
rect 57175 -68905 57205 -68879
rect 57263 -68905 57293 -68879
rect 59544 -68800 59610 -68792
rect 59087 -68850 59113 -68800
rect 59513 -68808 59610 -68800
rect 59513 -68842 59560 -68808
rect 59594 -68842 59610 -68808
rect 59513 -68850 59610 -68842
rect 59544 -68858 59610 -68850
rect 59016 -68908 59082 -68900
rect 59016 -68916 59113 -68908
rect 59016 -68950 59032 -68916
rect 59066 -68950 59113 -68916
rect 59016 -68958 59113 -68950
rect 59513 -68958 59539 -68908
rect 59016 -68966 59082 -68958
rect 53972 -69206 54069 -69190
rect 53972 -69244 53988 -69206
rect 54022 -69244 54069 -69206
rect 53972 -69260 54069 -69244
rect 54869 -69206 54966 -69190
rect 54869 -69244 54916 -69206
rect 54950 -69244 54966 -69206
rect 54869 -69260 54966 -69244
rect 59858 -68586 59924 -68578
rect 60368 -68586 60434 -68578
rect 59858 -68594 59946 -68586
rect 59858 -68628 59874 -68594
rect 59908 -68628 59946 -68594
rect 59858 -68636 59946 -68628
rect 60346 -68594 60434 -68586
rect 60346 -68628 60384 -68594
rect 60418 -68628 60434 -68594
rect 60346 -68636 60434 -68628
rect 59858 -68644 59924 -68636
rect 60368 -68644 60434 -68636
rect 55510 -69402 55576 -69386
rect 55510 -69404 55526 -69402
rect 55262 -69434 55288 -69404
rect 55488 -69434 55526 -69404
rect 55510 -69436 55526 -69434
rect 55560 -69436 55576 -69402
rect 55510 -69452 55576 -69436
rect 53982 -71934 54079 -71918
rect 53982 -71972 53998 -71934
rect 54032 -71972 54079 -71934
rect 53982 -71988 54079 -71972
rect 54879 -71934 54976 -71918
rect 54879 -71972 54926 -71934
rect 54960 -71972 54976 -71934
rect 54879 -71988 54976 -71972
rect 53510 -72306 53630 -72290
rect 53510 -72340 53526 -72306
rect 53614 -72340 53630 -72306
rect 53510 -72378 53630 -72340
rect 53982 -72290 54079 -72274
rect 53982 -72328 53998 -72290
rect 54032 -72328 54079 -72290
rect 53982 -72344 54079 -72328
rect 54879 -72290 54976 -72274
rect 54879 -72328 54926 -72290
rect 54960 -72328 54976 -72290
rect 54879 -72344 54976 -72328
rect 55318 -72368 55384 -72352
rect 55318 -72402 55334 -72368
rect 55368 -72402 55384 -72368
rect 55318 -72418 55384 -72402
rect 55336 -72440 55366 -72418
rect 55336 -72666 55366 -72640
rect 53510 -73216 53630 -73178
rect 53510 -73250 53526 -73216
rect 53614 -73250 53630 -73216
rect 53510 -73266 53630 -73250
rect 53842 -73040 53930 -73024
rect 53842 -73128 53858 -73040
rect 53892 -73128 53930 -73040
rect 53842 -73144 53930 -73128
rect 54730 -73040 54818 -73024
rect 54730 -73128 54768 -73040
rect 54802 -73128 54818 -73040
rect 54730 -73144 54818 -73128
rect 55030 -72959 55096 -72944
rect 55540 -72959 55606 -72944
rect 55030 -72960 55118 -72959
rect 55030 -72994 55046 -72960
rect 55080 -72994 55118 -72960
rect 55030 -72995 55118 -72994
rect 55518 -72960 55606 -72959
rect 55518 -72994 55556 -72960
rect 55590 -72994 55606 -72960
rect 55518 -72995 55606 -72994
rect 55030 -73010 55096 -72995
rect 55540 -73010 55606 -72995
rect 55866 -72256 55986 -72240
rect 55866 -72290 55882 -72256
rect 55970 -72290 55986 -72256
rect 55866 -72328 55986 -72290
rect 55866 -73166 55986 -73128
rect 55866 -73200 55882 -73166
rect 55970 -73200 55986 -73166
rect 55866 -73216 55986 -73200
rect 57175 -72309 57205 -72283
rect 57263 -72309 57293 -72283
rect 57175 -72482 57205 -72467
rect 57169 -72506 57205 -72482
rect 57169 -72541 57199 -72506
rect 57263 -72528 57293 -72467
rect 59544 -72293 59610 -72285
rect 59087 -72343 59113 -72293
rect 59513 -72301 59610 -72293
rect 59513 -72335 59560 -72301
rect 59594 -72335 59610 -72301
rect 59513 -72343 59610 -72335
rect 59544 -72351 59610 -72343
rect 59016 -72401 59082 -72393
rect 59016 -72409 59113 -72401
rect 59016 -72443 59032 -72409
rect 59066 -72443 59113 -72409
rect 59016 -72451 59113 -72443
rect 59513 -72451 59539 -72401
rect 59016 -72459 59082 -72451
rect 57123 -72557 57199 -72541
rect 57123 -72591 57133 -72557
rect 57167 -72591 57199 -72557
rect 57123 -72607 57199 -72591
rect 57241 -72544 57295 -72528
rect 57241 -72578 57251 -72544
rect 57285 -72578 57295 -72544
rect 57241 -72594 57295 -72578
rect 57169 -72616 57199 -72607
rect 57169 -72640 57205 -72616
rect 57175 -72655 57205 -72640
rect 57263 -72655 57293 -72594
rect 53510 -73324 53630 -73308
rect 53510 -73358 53526 -73324
rect 53614 -73358 53630 -73324
rect 53510 -73396 53630 -73358
rect 53842 -73446 53930 -73430
rect 53842 -73534 53858 -73446
rect 53892 -73534 53930 -73446
rect 53842 -73550 53930 -73534
rect 54730 -73446 54818 -73430
rect 54730 -73534 54768 -73446
rect 54802 -73534 54818 -73446
rect 54730 -73550 54818 -73534
rect 55030 -73581 55096 -73566
rect 55540 -73581 55606 -73566
rect 55030 -73582 55118 -73581
rect 55030 -73616 55046 -73582
rect 55080 -73616 55118 -73582
rect 55030 -73617 55118 -73616
rect 55518 -73582 55606 -73581
rect 55518 -73616 55556 -73582
rect 55590 -73616 55606 -73582
rect 55518 -73617 55606 -73616
rect 55030 -73632 55096 -73617
rect 53510 -74234 53630 -74196
rect 53510 -74268 53526 -74234
rect 53614 -74268 53630 -74234
rect 53510 -74284 53630 -74268
rect 55540 -73632 55606 -73617
rect 53972 -74250 54069 -74234
rect 53972 -74288 53988 -74250
rect 54022 -74288 54069 -74250
rect 53972 -74304 54069 -74288
rect 54869 -74250 54966 -74234
rect 54869 -74288 54916 -74250
rect 54950 -74288 54966 -74250
rect 54869 -74304 54966 -74288
rect 55326 -73936 55356 -73910
rect 55326 -74158 55356 -74136
rect 55308 -74174 55374 -74158
rect 55308 -74208 55324 -74174
rect 55358 -74208 55374 -74174
rect 55308 -74224 55374 -74208
rect 55866 -73370 55986 -73354
rect 55866 -73404 55882 -73370
rect 55970 -73404 55986 -73370
rect 55866 -73442 55986 -73404
rect 55866 -74280 55986 -74242
rect 55866 -74314 55882 -74280
rect 55970 -74314 55986 -74280
rect 55866 -74330 55986 -74314
rect 56476 -72806 56546 -72790
rect 56476 -72840 56492 -72806
rect 56530 -72840 56546 -72806
rect 56476 -72887 56546 -72840
rect 57175 -72785 57205 -72759
rect 57263 -72785 57293 -72759
rect 56476 -73734 56546 -73687
rect 56476 -73768 56492 -73734
rect 56530 -73768 56546 -73734
rect 56476 -73784 56546 -73768
rect 59087 -72678 59153 -72662
rect 59087 -72712 59103 -72678
rect 59137 -72712 59153 -72678
rect 59087 -72728 59153 -72712
rect 59090 -72759 59150 -72728
rect 59090 -73190 59150 -73159
rect 59087 -73206 59153 -73190
rect 59087 -73240 59103 -73206
rect 59137 -73240 59153 -73206
rect 59087 -73256 59153 -73240
rect 59858 -72620 59924 -72612
rect 60368 -72620 60434 -72612
rect 59858 -72628 59946 -72620
rect 59858 -72662 59874 -72628
rect 59908 -72662 59946 -72628
rect 59858 -72670 59946 -72662
rect 60346 -72628 60434 -72620
rect 60346 -72662 60384 -72628
rect 60418 -72662 60434 -72628
rect 60346 -72670 60434 -72662
rect 59858 -72678 59924 -72670
rect 60368 -72678 60434 -72670
rect 59530 -72898 59596 -72882
rect 59530 -72932 59546 -72898
rect 59580 -72932 59596 -72898
rect 59530 -72948 59596 -72932
rect 59548 -72970 59578 -72948
rect 59548 -73192 59578 -73170
rect 59530 -73208 59596 -73192
rect 59530 -73242 59546 -73208
rect 59580 -73242 59596 -73208
rect 59530 -73258 59596 -73242
rect 59846 -72898 59912 -72882
rect 59846 -72932 59862 -72898
rect 59896 -72932 59912 -72898
rect 59846 -72948 59912 -72932
rect 59864 -72970 59894 -72948
rect 59864 -73192 59894 -73170
rect 59846 -73208 59912 -73192
rect 59846 -73242 59862 -73208
rect 59896 -73242 59912 -73208
rect 59846 -73258 59912 -73242
rect 60343 -73165 60409 -73149
rect 61043 -73165 61109 -73149
rect 60343 -73199 60359 -73165
rect 60393 -73199 60409 -73165
rect 60343 -73217 60409 -73199
rect 61043 -73199 61059 -73165
rect 61093 -73199 61109 -73165
rect 61043 -73217 61109 -73199
rect 60165 -73247 60191 -73217
rect 60321 -73247 60441 -73217
rect 60641 -73247 60667 -73217
rect 60785 -73247 60811 -73217
rect 61011 -73247 61131 -73217
rect 61261 -73247 61287 -73217
rect 60343 -73257 60409 -73247
rect 60343 -73291 60359 -73257
rect 60393 -73291 60409 -73257
rect 60343 -73301 60409 -73291
rect 61043 -73257 61109 -73247
rect 61043 -73291 61059 -73257
rect 61093 -73291 61109 -73257
rect 61043 -73301 61109 -73291
rect 57175 -73829 57205 -73803
rect 57263 -73829 57293 -73803
rect 57175 -73948 57205 -73933
rect 57169 -73972 57205 -73948
rect 57169 -73981 57199 -73972
rect 57123 -73997 57199 -73981
rect 57263 -73994 57293 -73933
rect 59087 -73408 59153 -73392
rect 59087 -73442 59103 -73408
rect 59137 -73442 59153 -73408
rect 59087 -73458 59153 -73442
rect 59090 -73489 59150 -73458
rect 59090 -73920 59150 -73889
rect 57123 -74031 57133 -73997
rect 57167 -74031 57199 -73997
rect 57123 -74047 57199 -74031
rect 57169 -74082 57199 -74047
rect 57241 -74010 57295 -73994
rect 57241 -74044 57251 -74010
rect 57285 -74044 57295 -74010
rect 57241 -74060 57295 -74044
rect 59087 -73936 59153 -73920
rect 59087 -73970 59103 -73936
rect 59137 -73970 59153 -73936
rect 59087 -73986 59153 -73970
rect 60165 -73331 60191 -73301
rect 60321 -73331 60441 -73301
rect 60641 -73331 60667 -73301
rect 60785 -73331 60811 -73301
rect 61011 -73331 61131 -73301
rect 61261 -73331 61287 -73301
rect 59526 -73411 59596 -73380
rect 59526 -73430 59545 -73411
rect 59529 -73445 59545 -73430
rect 59579 -73430 59596 -73411
rect 59579 -73445 59595 -73430
rect 59529 -73461 59595 -73445
rect 59547 -73483 59577 -73461
rect 59547 -73705 59577 -73683
rect 59529 -73721 59595 -73705
rect 59529 -73755 59545 -73721
rect 59579 -73755 59595 -73721
rect 59529 -73771 59595 -73755
rect 59845 -73411 59911 -73395
rect 59845 -73445 59861 -73411
rect 59895 -73445 59911 -73411
rect 59845 -73461 59911 -73445
rect 60343 -73341 60409 -73331
rect 60343 -73375 60359 -73341
rect 60393 -73375 60409 -73341
rect 60343 -73385 60409 -73375
rect 61043 -73341 61109 -73331
rect 61043 -73375 61059 -73341
rect 61093 -73375 61109 -73341
rect 61043 -73385 61109 -73375
rect 59863 -73483 59893 -73461
rect 59863 -73705 59893 -73683
rect 59845 -73721 59911 -73705
rect 59845 -73755 59861 -73721
rect 59895 -73755 59911 -73721
rect 59845 -73771 59911 -73755
rect 60165 -73415 60191 -73385
rect 60321 -73415 60441 -73385
rect 60641 -73415 60667 -73385
rect 60785 -73415 60811 -73385
rect 61011 -73415 61131 -73385
rect 61261 -73415 61287 -73385
rect 60343 -73425 60409 -73415
rect 60343 -73459 60359 -73425
rect 60393 -73459 60409 -73425
rect 60343 -73469 60409 -73459
rect 61043 -73425 61109 -73415
rect 61043 -73459 61059 -73425
rect 61093 -73459 61109 -73425
rect 61043 -73469 61109 -73459
rect 60165 -73499 60191 -73469
rect 60321 -73499 60441 -73469
rect 60641 -73499 60667 -73469
rect 60785 -73499 60811 -73469
rect 61011 -73499 61131 -73469
rect 61261 -73499 61287 -73469
rect 57169 -74106 57205 -74082
rect 57175 -74121 57205 -74106
rect 57263 -74121 57293 -74060
rect 57175 -74305 57205 -74279
rect 57263 -74305 57293 -74279
rect 59544 -74200 59610 -74192
rect 59087 -74250 59113 -74200
rect 59513 -74208 59610 -74200
rect 59513 -74242 59560 -74208
rect 59594 -74242 59610 -74208
rect 59513 -74250 59610 -74242
rect 59544 -74258 59610 -74250
rect 59016 -74308 59082 -74300
rect 59016 -74316 59113 -74308
rect 59016 -74350 59032 -74316
rect 59066 -74350 59113 -74316
rect 59016 -74358 59113 -74350
rect 59513 -74358 59539 -74308
rect 59016 -74366 59082 -74358
rect 53972 -74606 54069 -74590
rect 53972 -74644 53988 -74606
rect 54022 -74644 54069 -74606
rect 53972 -74660 54069 -74644
rect 54869 -74606 54966 -74590
rect 54869 -74644 54916 -74606
rect 54950 -74644 54966 -74606
rect 54869 -74660 54966 -74644
rect 59858 -73986 59924 -73978
rect 60368 -73986 60434 -73978
rect 59858 -73994 59946 -73986
rect 59858 -74028 59874 -73994
rect 59908 -74028 59946 -73994
rect 59858 -74036 59946 -74028
rect 60346 -73994 60434 -73986
rect 60346 -74028 60384 -73994
rect 60418 -74028 60434 -73994
rect 60346 -74036 60434 -74028
rect 59858 -74044 59924 -74036
rect 60368 -74044 60434 -74036
rect 55510 -74802 55576 -74786
rect 55510 -74804 55526 -74802
rect 55262 -74834 55288 -74804
rect 55488 -74834 55526 -74804
rect 55510 -74836 55526 -74834
rect 55560 -74836 55576 -74802
rect 55510 -74852 55576 -74836
rect 53982 -77334 54079 -77318
rect 53982 -77372 53998 -77334
rect 54032 -77372 54079 -77334
rect 53982 -77388 54079 -77372
rect 54879 -77334 54976 -77318
rect 54879 -77372 54926 -77334
rect 54960 -77372 54976 -77334
rect 54879 -77388 54976 -77372
rect 53510 -77706 53630 -77690
rect 53510 -77740 53526 -77706
rect 53614 -77740 53630 -77706
rect 53510 -77778 53630 -77740
rect 53982 -77690 54079 -77674
rect 53982 -77728 53998 -77690
rect 54032 -77728 54079 -77690
rect 53982 -77744 54079 -77728
rect 54879 -77690 54976 -77674
rect 54879 -77728 54926 -77690
rect 54960 -77728 54976 -77690
rect 54879 -77744 54976 -77728
rect 55318 -77768 55384 -77752
rect 55318 -77802 55334 -77768
rect 55368 -77802 55384 -77768
rect 55318 -77818 55384 -77802
rect 55336 -77840 55366 -77818
rect 55336 -78066 55366 -78040
rect 53510 -78616 53630 -78578
rect 53510 -78650 53526 -78616
rect 53614 -78650 53630 -78616
rect 53510 -78666 53630 -78650
rect 53842 -78440 53930 -78424
rect 53842 -78528 53858 -78440
rect 53892 -78528 53930 -78440
rect 53842 -78544 53930 -78528
rect 54730 -78440 54818 -78424
rect 54730 -78528 54768 -78440
rect 54802 -78528 54818 -78440
rect 54730 -78544 54818 -78528
rect 55030 -78359 55096 -78344
rect 55540 -78359 55606 -78344
rect 55030 -78360 55118 -78359
rect 55030 -78394 55046 -78360
rect 55080 -78394 55118 -78360
rect 55030 -78395 55118 -78394
rect 55518 -78360 55606 -78359
rect 55518 -78394 55556 -78360
rect 55590 -78394 55606 -78360
rect 55518 -78395 55606 -78394
rect 55030 -78410 55096 -78395
rect 55540 -78410 55606 -78395
rect 55866 -77656 55986 -77640
rect 55866 -77690 55882 -77656
rect 55970 -77690 55986 -77656
rect 55866 -77728 55986 -77690
rect 55866 -78566 55986 -78528
rect 55866 -78600 55882 -78566
rect 55970 -78600 55986 -78566
rect 55866 -78616 55986 -78600
rect 57175 -77709 57205 -77683
rect 57263 -77709 57293 -77683
rect 57175 -77882 57205 -77867
rect 57169 -77906 57205 -77882
rect 57169 -77941 57199 -77906
rect 57263 -77928 57293 -77867
rect 59544 -77693 59610 -77685
rect 59087 -77743 59113 -77693
rect 59513 -77701 59610 -77693
rect 59513 -77735 59560 -77701
rect 59594 -77735 59610 -77701
rect 59513 -77743 59610 -77735
rect 59544 -77751 59610 -77743
rect 59016 -77801 59082 -77793
rect 59016 -77809 59113 -77801
rect 59016 -77843 59032 -77809
rect 59066 -77843 59113 -77809
rect 59016 -77851 59113 -77843
rect 59513 -77851 59539 -77801
rect 59016 -77859 59082 -77851
rect 57123 -77957 57199 -77941
rect 57123 -77991 57133 -77957
rect 57167 -77991 57199 -77957
rect 57123 -78007 57199 -77991
rect 57241 -77944 57295 -77928
rect 57241 -77978 57251 -77944
rect 57285 -77978 57295 -77944
rect 57241 -77994 57295 -77978
rect 57169 -78016 57199 -78007
rect 57169 -78040 57205 -78016
rect 57175 -78055 57205 -78040
rect 57263 -78055 57293 -77994
rect 53510 -78724 53630 -78708
rect 53510 -78758 53526 -78724
rect 53614 -78758 53630 -78724
rect 53510 -78796 53630 -78758
rect 53842 -78846 53930 -78830
rect 53842 -78934 53858 -78846
rect 53892 -78934 53930 -78846
rect 53842 -78950 53930 -78934
rect 54730 -78846 54818 -78830
rect 54730 -78934 54768 -78846
rect 54802 -78934 54818 -78846
rect 54730 -78950 54818 -78934
rect 55030 -78981 55096 -78966
rect 55540 -78981 55606 -78966
rect 55030 -78982 55118 -78981
rect 55030 -79016 55046 -78982
rect 55080 -79016 55118 -78982
rect 55030 -79017 55118 -79016
rect 55518 -78982 55606 -78981
rect 55518 -79016 55556 -78982
rect 55590 -79016 55606 -78982
rect 55518 -79017 55606 -79016
rect 55030 -79032 55096 -79017
rect 53510 -79634 53630 -79596
rect 53510 -79668 53526 -79634
rect 53614 -79668 53630 -79634
rect 53510 -79684 53630 -79668
rect 55540 -79032 55606 -79017
rect 53972 -79650 54069 -79634
rect 53972 -79688 53988 -79650
rect 54022 -79688 54069 -79650
rect 53972 -79704 54069 -79688
rect 54869 -79650 54966 -79634
rect 54869 -79688 54916 -79650
rect 54950 -79688 54966 -79650
rect 54869 -79704 54966 -79688
rect 55326 -79336 55356 -79310
rect 55326 -79558 55356 -79536
rect 55308 -79574 55374 -79558
rect 55308 -79608 55324 -79574
rect 55358 -79608 55374 -79574
rect 55308 -79624 55374 -79608
rect 55866 -78770 55986 -78754
rect 55866 -78804 55882 -78770
rect 55970 -78804 55986 -78770
rect 55866 -78842 55986 -78804
rect 55866 -79680 55986 -79642
rect 55866 -79714 55882 -79680
rect 55970 -79714 55986 -79680
rect 55866 -79730 55986 -79714
rect 56476 -78206 56546 -78190
rect 56476 -78240 56492 -78206
rect 56530 -78240 56546 -78206
rect 56476 -78287 56546 -78240
rect 57175 -78185 57205 -78159
rect 57263 -78185 57293 -78159
rect 56476 -79134 56546 -79087
rect 56476 -79168 56492 -79134
rect 56530 -79168 56546 -79134
rect 56476 -79184 56546 -79168
rect 59087 -78078 59153 -78062
rect 59087 -78112 59103 -78078
rect 59137 -78112 59153 -78078
rect 59087 -78128 59153 -78112
rect 59090 -78159 59150 -78128
rect 59090 -78590 59150 -78559
rect 59087 -78606 59153 -78590
rect 59087 -78640 59103 -78606
rect 59137 -78640 59153 -78606
rect 59087 -78656 59153 -78640
rect 59858 -78020 59924 -78012
rect 60368 -78020 60434 -78012
rect 59858 -78028 59946 -78020
rect 59858 -78062 59874 -78028
rect 59908 -78062 59946 -78028
rect 59858 -78070 59946 -78062
rect 60346 -78028 60434 -78020
rect 60346 -78062 60384 -78028
rect 60418 -78062 60434 -78028
rect 60346 -78070 60434 -78062
rect 59858 -78078 59924 -78070
rect 60368 -78078 60434 -78070
rect 59530 -78298 59596 -78282
rect 59530 -78332 59546 -78298
rect 59580 -78332 59596 -78298
rect 59530 -78348 59596 -78332
rect 59548 -78370 59578 -78348
rect 59548 -78592 59578 -78570
rect 59530 -78608 59596 -78592
rect 59530 -78642 59546 -78608
rect 59580 -78642 59596 -78608
rect 59530 -78658 59596 -78642
rect 59846 -78298 59912 -78282
rect 59846 -78332 59862 -78298
rect 59896 -78332 59912 -78298
rect 59846 -78348 59912 -78332
rect 59864 -78370 59894 -78348
rect 59864 -78592 59894 -78570
rect 59846 -78608 59912 -78592
rect 59846 -78642 59862 -78608
rect 59896 -78642 59912 -78608
rect 59846 -78658 59912 -78642
rect 60343 -78565 60409 -78549
rect 61043 -78565 61109 -78549
rect 60343 -78599 60359 -78565
rect 60393 -78599 60409 -78565
rect 60343 -78617 60409 -78599
rect 61043 -78599 61059 -78565
rect 61093 -78599 61109 -78565
rect 61043 -78617 61109 -78599
rect 60165 -78647 60191 -78617
rect 60321 -78647 60441 -78617
rect 60641 -78647 60667 -78617
rect 60785 -78647 60811 -78617
rect 61011 -78647 61131 -78617
rect 61261 -78647 61287 -78617
rect 60343 -78657 60409 -78647
rect 60343 -78691 60359 -78657
rect 60393 -78691 60409 -78657
rect 60343 -78701 60409 -78691
rect 61043 -78657 61109 -78647
rect 61043 -78691 61059 -78657
rect 61093 -78691 61109 -78657
rect 61043 -78701 61109 -78691
rect 57175 -79229 57205 -79203
rect 57263 -79229 57293 -79203
rect 57175 -79348 57205 -79333
rect 57169 -79372 57205 -79348
rect 57169 -79381 57199 -79372
rect 57123 -79397 57199 -79381
rect 57263 -79394 57293 -79333
rect 59087 -78808 59153 -78792
rect 59087 -78842 59103 -78808
rect 59137 -78842 59153 -78808
rect 59087 -78858 59153 -78842
rect 59090 -78889 59150 -78858
rect 59090 -79320 59150 -79289
rect 57123 -79431 57133 -79397
rect 57167 -79431 57199 -79397
rect 57123 -79447 57199 -79431
rect 57169 -79482 57199 -79447
rect 57241 -79410 57295 -79394
rect 57241 -79444 57251 -79410
rect 57285 -79444 57295 -79410
rect 57241 -79460 57295 -79444
rect 59087 -79336 59153 -79320
rect 59087 -79370 59103 -79336
rect 59137 -79370 59153 -79336
rect 59087 -79386 59153 -79370
rect 60165 -78731 60191 -78701
rect 60321 -78731 60441 -78701
rect 60641 -78731 60667 -78701
rect 60785 -78731 60811 -78701
rect 61011 -78731 61131 -78701
rect 61261 -78731 61287 -78701
rect 59526 -78811 59596 -78780
rect 59526 -78830 59545 -78811
rect 59529 -78845 59545 -78830
rect 59579 -78830 59596 -78811
rect 59579 -78845 59595 -78830
rect 59529 -78861 59595 -78845
rect 59547 -78883 59577 -78861
rect 59547 -79105 59577 -79083
rect 59529 -79121 59595 -79105
rect 59529 -79155 59545 -79121
rect 59579 -79155 59595 -79121
rect 59529 -79171 59595 -79155
rect 59845 -78811 59911 -78795
rect 59845 -78845 59861 -78811
rect 59895 -78845 59911 -78811
rect 59845 -78861 59911 -78845
rect 60343 -78741 60409 -78731
rect 60343 -78775 60359 -78741
rect 60393 -78775 60409 -78741
rect 60343 -78785 60409 -78775
rect 61043 -78741 61109 -78731
rect 61043 -78775 61059 -78741
rect 61093 -78775 61109 -78741
rect 61043 -78785 61109 -78775
rect 59863 -78883 59893 -78861
rect 59863 -79105 59893 -79083
rect 59845 -79121 59911 -79105
rect 59845 -79155 59861 -79121
rect 59895 -79155 59911 -79121
rect 59845 -79171 59911 -79155
rect 60165 -78815 60191 -78785
rect 60321 -78815 60441 -78785
rect 60641 -78815 60667 -78785
rect 60785 -78815 60811 -78785
rect 61011 -78815 61131 -78785
rect 61261 -78815 61287 -78785
rect 60343 -78825 60409 -78815
rect 60343 -78859 60359 -78825
rect 60393 -78859 60409 -78825
rect 60343 -78869 60409 -78859
rect 61043 -78825 61109 -78815
rect 61043 -78859 61059 -78825
rect 61093 -78859 61109 -78825
rect 61043 -78869 61109 -78859
rect 60165 -78899 60191 -78869
rect 60321 -78899 60441 -78869
rect 60641 -78899 60667 -78869
rect 60785 -78899 60811 -78869
rect 61011 -78899 61131 -78869
rect 61261 -78899 61287 -78869
rect 57169 -79506 57205 -79482
rect 57175 -79521 57205 -79506
rect 57263 -79521 57293 -79460
rect 57175 -79705 57205 -79679
rect 57263 -79705 57293 -79679
rect 59544 -79600 59610 -79592
rect 59087 -79650 59113 -79600
rect 59513 -79608 59610 -79600
rect 59513 -79642 59560 -79608
rect 59594 -79642 59610 -79608
rect 59513 -79650 59610 -79642
rect 59544 -79658 59610 -79650
rect 59016 -79708 59082 -79700
rect 59016 -79716 59113 -79708
rect 59016 -79750 59032 -79716
rect 59066 -79750 59113 -79716
rect 59016 -79758 59113 -79750
rect 59513 -79758 59539 -79708
rect 59016 -79766 59082 -79758
rect 53972 -80006 54069 -79990
rect 53972 -80044 53988 -80006
rect 54022 -80044 54069 -80006
rect 53972 -80060 54069 -80044
rect 54869 -80006 54966 -79990
rect 54869 -80044 54916 -80006
rect 54950 -80044 54966 -80006
rect 54869 -80060 54966 -80044
rect 59858 -79386 59924 -79378
rect 60368 -79386 60434 -79378
rect 59858 -79394 59946 -79386
rect 59858 -79428 59874 -79394
rect 59908 -79428 59946 -79394
rect 59858 -79436 59946 -79428
rect 60346 -79394 60434 -79386
rect 60346 -79428 60384 -79394
rect 60418 -79428 60434 -79394
rect 60346 -79436 60434 -79428
rect 59858 -79444 59924 -79436
rect 60368 -79444 60434 -79436
rect 55510 -80202 55576 -80186
rect 55510 -80204 55526 -80202
rect 55262 -80234 55288 -80204
rect 55488 -80234 55526 -80204
rect 55510 -80236 55526 -80234
rect 55560 -80236 55576 -80202
rect 55510 -80252 55576 -80236
rect 53982 -82734 54079 -82718
rect 53982 -82772 53998 -82734
rect 54032 -82772 54079 -82734
rect 53982 -82788 54079 -82772
rect 54879 -82734 54976 -82718
rect 54879 -82772 54926 -82734
rect 54960 -82772 54976 -82734
rect 54879 -82788 54976 -82772
rect 53510 -83106 53630 -83090
rect 53510 -83140 53526 -83106
rect 53614 -83140 53630 -83106
rect 53510 -83178 53630 -83140
rect 53982 -83090 54079 -83074
rect 53982 -83128 53998 -83090
rect 54032 -83128 54079 -83090
rect 53982 -83144 54079 -83128
rect 54879 -83090 54976 -83074
rect 54879 -83128 54926 -83090
rect 54960 -83128 54976 -83090
rect 54879 -83144 54976 -83128
rect 55318 -83168 55384 -83152
rect 55318 -83202 55334 -83168
rect 55368 -83202 55384 -83168
rect 55318 -83218 55384 -83202
rect 55336 -83240 55366 -83218
rect 55336 -83466 55366 -83440
rect 53510 -84016 53630 -83978
rect 53510 -84050 53526 -84016
rect 53614 -84050 53630 -84016
rect 53510 -84066 53630 -84050
rect 53842 -83840 53930 -83824
rect 53842 -83928 53858 -83840
rect 53892 -83928 53930 -83840
rect 53842 -83944 53930 -83928
rect 54730 -83840 54818 -83824
rect 54730 -83928 54768 -83840
rect 54802 -83928 54818 -83840
rect 54730 -83944 54818 -83928
rect 55030 -83759 55096 -83744
rect 55540 -83759 55606 -83744
rect 55030 -83760 55118 -83759
rect 55030 -83794 55046 -83760
rect 55080 -83794 55118 -83760
rect 55030 -83795 55118 -83794
rect 55518 -83760 55606 -83759
rect 55518 -83794 55556 -83760
rect 55590 -83794 55606 -83760
rect 55518 -83795 55606 -83794
rect 55030 -83810 55096 -83795
rect 55540 -83810 55606 -83795
rect 55866 -83056 55986 -83040
rect 55866 -83090 55882 -83056
rect 55970 -83090 55986 -83056
rect 55866 -83128 55986 -83090
rect 55866 -83966 55986 -83928
rect 55866 -84000 55882 -83966
rect 55970 -84000 55986 -83966
rect 55866 -84016 55986 -84000
rect 57175 -83109 57205 -83083
rect 57263 -83109 57293 -83083
rect 57175 -83282 57205 -83267
rect 57169 -83306 57205 -83282
rect 57169 -83341 57199 -83306
rect 57263 -83328 57293 -83267
rect 59544 -83093 59610 -83085
rect 59087 -83143 59113 -83093
rect 59513 -83101 59610 -83093
rect 59513 -83135 59560 -83101
rect 59594 -83135 59610 -83101
rect 59513 -83143 59610 -83135
rect 59544 -83151 59610 -83143
rect 59016 -83201 59082 -83193
rect 59016 -83209 59113 -83201
rect 59016 -83243 59032 -83209
rect 59066 -83243 59113 -83209
rect 59016 -83251 59113 -83243
rect 59513 -83251 59539 -83201
rect 59016 -83259 59082 -83251
rect 57123 -83357 57199 -83341
rect 57123 -83391 57133 -83357
rect 57167 -83391 57199 -83357
rect 57123 -83407 57199 -83391
rect 57241 -83344 57295 -83328
rect 57241 -83378 57251 -83344
rect 57285 -83378 57295 -83344
rect 57241 -83394 57295 -83378
rect 57169 -83416 57199 -83407
rect 57169 -83440 57205 -83416
rect 57175 -83455 57205 -83440
rect 57263 -83455 57293 -83394
rect 53510 -84124 53630 -84108
rect 53510 -84158 53526 -84124
rect 53614 -84158 53630 -84124
rect 53510 -84196 53630 -84158
rect 53842 -84246 53930 -84230
rect 53842 -84334 53858 -84246
rect 53892 -84334 53930 -84246
rect 53842 -84350 53930 -84334
rect 54730 -84246 54818 -84230
rect 54730 -84334 54768 -84246
rect 54802 -84334 54818 -84246
rect 54730 -84350 54818 -84334
rect 55030 -84381 55096 -84366
rect 55540 -84381 55606 -84366
rect 55030 -84382 55118 -84381
rect 55030 -84416 55046 -84382
rect 55080 -84416 55118 -84382
rect 55030 -84417 55118 -84416
rect 55518 -84382 55606 -84381
rect 55518 -84416 55556 -84382
rect 55590 -84416 55606 -84382
rect 55518 -84417 55606 -84416
rect 55030 -84432 55096 -84417
rect 53510 -85034 53630 -84996
rect 53510 -85068 53526 -85034
rect 53614 -85068 53630 -85034
rect 53510 -85084 53630 -85068
rect 55540 -84432 55606 -84417
rect 53972 -85050 54069 -85034
rect 53972 -85088 53988 -85050
rect 54022 -85088 54069 -85050
rect 53972 -85104 54069 -85088
rect 54869 -85050 54966 -85034
rect 54869 -85088 54916 -85050
rect 54950 -85088 54966 -85050
rect 54869 -85104 54966 -85088
rect 55326 -84736 55356 -84710
rect 55326 -84958 55356 -84936
rect 55308 -84974 55374 -84958
rect 55308 -85008 55324 -84974
rect 55358 -85008 55374 -84974
rect 55308 -85024 55374 -85008
rect 55866 -84170 55986 -84154
rect 55866 -84204 55882 -84170
rect 55970 -84204 55986 -84170
rect 55866 -84242 55986 -84204
rect 55866 -85080 55986 -85042
rect 55866 -85114 55882 -85080
rect 55970 -85114 55986 -85080
rect 55866 -85130 55986 -85114
rect 56476 -83606 56546 -83590
rect 56476 -83640 56492 -83606
rect 56530 -83640 56546 -83606
rect 56476 -83687 56546 -83640
rect 57175 -83585 57205 -83559
rect 57263 -83585 57293 -83559
rect 56476 -84534 56546 -84487
rect 56476 -84568 56492 -84534
rect 56530 -84568 56546 -84534
rect 56476 -84584 56546 -84568
rect 59087 -83478 59153 -83462
rect 59087 -83512 59103 -83478
rect 59137 -83512 59153 -83478
rect 59087 -83528 59153 -83512
rect 59090 -83559 59150 -83528
rect 59090 -83990 59150 -83959
rect 59087 -84006 59153 -83990
rect 59087 -84040 59103 -84006
rect 59137 -84040 59153 -84006
rect 59087 -84056 59153 -84040
rect 59858 -83420 59924 -83412
rect 60368 -83420 60434 -83412
rect 59858 -83428 59946 -83420
rect 59858 -83462 59874 -83428
rect 59908 -83462 59946 -83428
rect 59858 -83470 59946 -83462
rect 60346 -83428 60434 -83420
rect 60346 -83462 60384 -83428
rect 60418 -83462 60434 -83428
rect 60346 -83470 60434 -83462
rect 59858 -83478 59924 -83470
rect 60368 -83478 60434 -83470
rect 59530 -83698 59596 -83682
rect 59530 -83732 59546 -83698
rect 59580 -83732 59596 -83698
rect 59530 -83748 59596 -83732
rect 59548 -83770 59578 -83748
rect 59548 -83992 59578 -83970
rect 59530 -84008 59596 -83992
rect 59530 -84042 59546 -84008
rect 59580 -84042 59596 -84008
rect 59530 -84058 59596 -84042
rect 59846 -83698 59912 -83682
rect 59846 -83732 59862 -83698
rect 59896 -83732 59912 -83698
rect 59846 -83748 59912 -83732
rect 59864 -83770 59894 -83748
rect 59864 -83992 59894 -83970
rect 59846 -84008 59912 -83992
rect 59846 -84042 59862 -84008
rect 59896 -84042 59912 -84008
rect 59846 -84058 59912 -84042
rect 60343 -83965 60409 -83949
rect 61043 -83965 61109 -83949
rect 60343 -83999 60359 -83965
rect 60393 -83999 60409 -83965
rect 60343 -84017 60409 -83999
rect 61043 -83999 61059 -83965
rect 61093 -83999 61109 -83965
rect 61043 -84017 61109 -83999
rect 60165 -84047 60191 -84017
rect 60321 -84047 60441 -84017
rect 60641 -84047 60667 -84017
rect 60785 -84047 60811 -84017
rect 61011 -84047 61131 -84017
rect 61261 -84047 61287 -84017
rect 60343 -84057 60409 -84047
rect 60343 -84091 60359 -84057
rect 60393 -84091 60409 -84057
rect 60343 -84101 60409 -84091
rect 61043 -84057 61109 -84047
rect 61043 -84091 61059 -84057
rect 61093 -84091 61109 -84057
rect 61043 -84101 61109 -84091
rect 57175 -84629 57205 -84603
rect 57263 -84629 57293 -84603
rect 57175 -84748 57205 -84733
rect 57169 -84772 57205 -84748
rect 57169 -84781 57199 -84772
rect 57123 -84797 57199 -84781
rect 57263 -84794 57293 -84733
rect 59087 -84208 59153 -84192
rect 59087 -84242 59103 -84208
rect 59137 -84242 59153 -84208
rect 59087 -84258 59153 -84242
rect 59090 -84289 59150 -84258
rect 59090 -84720 59150 -84689
rect 57123 -84831 57133 -84797
rect 57167 -84831 57199 -84797
rect 57123 -84847 57199 -84831
rect 57169 -84882 57199 -84847
rect 57241 -84810 57295 -84794
rect 57241 -84844 57251 -84810
rect 57285 -84844 57295 -84810
rect 57241 -84860 57295 -84844
rect 59087 -84736 59153 -84720
rect 59087 -84770 59103 -84736
rect 59137 -84770 59153 -84736
rect 59087 -84786 59153 -84770
rect 60165 -84131 60191 -84101
rect 60321 -84131 60441 -84101
rect 60641 -84131 60667 -84101
rect 60785 -84131 60811 -84101
rect 61011 -84131 61131 -84101
rect 61261 -84131 61287 -84101
rect 59526 -84211 59596 -84180
rect 59526 -84230 59545 -84211
rect 59529 -84245 59545 -84230
rect 59579 -84230 59596 -84211
rect 59579 -84245 59595 -84230
rect 59529 -84261 59595 -84245
rect 59547 -84283 59577 -84261
rect 59547 -84505 59577 -84483
rect 59529 -84521 59595 -84505
rect 59529 -84555 59545 -84521
rect 59579 -84555 59595 -84521
rect 59529 -84571 59595 -84555
rect 59845 -84211 59911 -84195
rect 59845 -84245 59861 -84211
rect 59895 -84245 59911 -84211
rect 59845 -84261 59911 -84245
rect 60343 -84141 60409 -84131
rect 60343 -84175 60359 -84141
rect 60393 -84175 60409 -84141
rect 60343 -84185 60409 -84175
rect 61043 -84141 61109 -84131
rect 61043 -84175 61059 -84141
rect 61093 -84175 61109 -84141
rect 61043 -84185 61109 -84175
rect 59863 -84283 59893 -84261
rect 59863 -84505 59893 -84483
rect 59845 -84521 59911 -84505
rect 59845 -84555 59861 -84521
rect 59895 -84555 59911 -84521
rect 59845 -84571 59911 -84555
rect 60165 -84215 60191 -84185
rect 60321 -84215 60441 -84185
rect 60641 -84215 60667 -84185
rect 60785 -84215 60811 -84185
rect 61011 -84215 61131 -84185
rect 61261 -84215 61287 -84185
rect 60343 -84225 60409 -84215
rect 60343 -84259 60359 -84225
rect 60393 -84259 60409 -84225
rect 60343 -84269 60409 -84259
rect 61043 -84225 61109 -84215
rect 61043 -84259 61059 -84225
rect 61093 -84259 61109 -84225
rect 61043 -84269 61109 -84259
rect 60165 -84299 60191 -84269
rect 60321 -84299 60441 -84269
rect 60641 -84299 60667 -84269
rect 60785 -84299 60811 -84269
rect 61011 -84299 61131 -84269
rect 61261 -84299 61287 -84269
rect 57169 -84906 57205 -84882
rect 57175 -84921 57205 -84906
rect 57263 -84921 57293 -84860
rect 57175 -85105 57205 -85079
rect 57263 -85105 57293 -85079
rect 59544 -85000 59610 -84992
rect 59087 -85050 59113 -85000
rect 59513 -85008 59610 -85000
rect 59513 -85042 59560 -85008
rect 59594 -85042 59610 -85008
rect 59513 -85050 59610 -85042
rect 59544 -85058 59610 -85050
rect 59016 -85108 59082 -85100
rect 59016 -85116 59113 -85108
rect 59016 -85150 59032 -85116
rect 59066 -85150 59113 -85116
rect 59016 -85158 59113 -85150
rect 59513 -85158 59539 -85108
rect 59016 -85166 59082 -85158
rect 53972 -85406 54069 -85390
rect 53972 -85444 53988 -85406
rect 54022 -85444 54069 -85406
rect 53972 -85460 54069 -85444
rect 54869 -85406 54966 -85390
rect 54869 -85444 54916 -85406
rect 54950 -85444 54966 -85406
rect 54869 -85460 54966 -85444
rect 59858 -84786 59924 -84778
rect 60368 -84786 60434 -84778
rect 59858 -84794 59946 -84786
rect 59858 -84828 59874 -84794
rect 59908 -84828 59946 -84794
rect 59858 -84836 59946 -84828
rect 60346 -84794 60434 -84786
rect 60346 -84828 60384 -84794
rect 60418 -84828 60434 -84794
rect 60346 -84836 60434 -84828
rect 59858 -84844 59924 -84836
rect 60368 -84844 60434 -84836
rect 55510 -85602 55576 -85586
rect 55510 -85604 55526 -85602
rect 55262 -85634 55288 -85604
rect 55488 -85634 55526 -85604
rect 55510 -85636 55526 -85634
rect 55560 -85636 55576 -85602
rect 55510 -85652 55576 -85636
<< polycont >>
rect 53998 -1772 54032 -1734
rect 54926 -1772 54960 -1734
rect 53526 -2140 53614 -2106
rect 53998 -2128 54032 -2090
rect 54926 -2128 54960 -2090
rect 55334 -2202 55368 -2168
rect 53526 -3050 53614 -3016
rect 53858 -2928 53892 -2840
rect 54768 -2928 54802 -2840
rect 55046 -2794 55080 -2760
rect 55556 -2794 55590 -2760
rect 55882 -2090 55970 -2056
rect 55882 -3000 55970 -2966
rect 59560 -2135 59594 -2101
rect 59032 -2243 59066 -2209
rect 57133 -2391 57167 -2357
rect 57251 -2378 57285 -2344
rect 53526 -3158 53614 -3124
rect 53858 -3334 53892 -3246
rect 54768 -3334 54802 -3246
rect 55046 -3416 55080 -3382
rect 55556 -3416 55590 -3382
rect 53526 -4068 53614 -4034
rect 53988 -4088 54022 -4050
rect 54916 -4088 54950 -4050
rect 55324 -4008 55358 -3974
rect 55882 -3204 55970 -3170
rect 55882 -4114 55970 -4080
rect 56492 -2640 56530 -2606
rect 56492 -3568 56530 -3534
rect 59103 -2512 59137 -2478
rect 59103 -3040 59137 -3006
rect 59874 -2462 59908 -2428
rect 60384 -2462 60418 -2428
rect 59546 -2732 59580 -2698
rect 59546 -3042 59580 -3008
rect 59862 -2732 59896 -2698
rect 59862 -3042 59896 -3008
rect 60359 -2999 60393 -2965
rect 61059 -2999 61093 -2965
rect 60359 -3091 60393 -3057
rect 61059 -3091 61093 -3057
rect 59103 -3242 59137 -3208
rect 57133 -3831 57167 -3797
rect 57251 -3844 57285 -3810
rect 59103 -3770 59137 -3736
rect 59545 -3245 59579 -3211
rect 59545 -3555 59579 -3521
rect 59861 -3245 59895 -3211
rect 60359 -3175 60393 -3141
rect 61059 -3175 61093 -3141
rect 59861 -3555 59895 -3521
rect 60359 -3259 60393 -3225
rect 61059 -3259 61093 -3225
rect 59560 -4042 59594 -4008
rect 59032 -4150 59066 -4116
rect 53988 -4444 54022 -4406
rect 54916 -4444 54950 -4406
rect 59874 -3828 59908 -3794
rect 60384 -3828 60418 -3794
rect 55526 -4636 55560 -4602
rect 53998 -7172 54032 -7134
rect 54926 -7172 54960 -7134
rect 20908 -7809 21076 -7775
rect 20908 -11737 21076 -11703
rect 21394 -7809 21562 -7775
rect 21394 -11737 21562 -11703
rect 21880 -7809 22048 -7775
rect 21880 -11737 22048 -11703
rect 53526 -7540 53614 -7506
rect 53998 -7528 54032 -7490
rect 54926 -7528 54960 -7490
rect 55334 -7602 55368 -7568
rect 53526 -8450 53614 -8416
rect 53858 -8328 53892 -8240
rect 54768 -8328 54802 -8240
rect 55046 -8194 55080 -8160
rect 55556 -8194 55590 -8160
rect 55882 -7490 55970 -7456
rect 55882 -8400 55970 -8366
rect 59560 -7535 59594 -7501
rect 59032 -7643 59066 -7609
rect 57133 -7791 57167 -7757
rect 57251 -7778 57285 -7744
rect 53526 -8558 53614 -8524
rect 53858 -8734 53892 -8646
rect 54768 -8734 54802 -8646
rect 55046 -8816 55080 -8782
rect 55556 -8816 55590 -8782
rect 53526 -9468 53614 -9434
rect 53988 -9488 54022 -9450
rect 54916 -9488 54950 -9450
rect 55324 -9408 55358 -9374
rect 55882 -8604 55970 -8570
rect 55882 -9514 55970 -9480
rect 56492 -8040 56530 -8006
rect 56492 -8968 56530 -8934
rect 59103 -7912 59137 -7878
rect 59103 -8440 59137 -8406
rect 59874 -7862 59908 -7828
rect 60384 -7862 60418 -7828
rect 59546 -8132 59580 -8098
rect 59546 -8442 59580 -8408
rect 59862 -8132 59896 -8098
rect 59862 -8442 59896 -8408
rect 60359 -8399 60393 -8365
rect 61059 -8399 61093 -8365
rect 60359 -8491 60393 -8457
rect 61059 -8491 61093 -8457
rect 59103 -8642 59137 -8608
rect 57133 -9231 57167 -9197
rect 57251 -9244 57285 -9210
rect 59103 -9170 59137 -9136
rect 59545 -8645 59579 -8611
rect 59545 -8955 59579 -8921
rect 59861 -8645 59895 -8611
rect 60359 -8575 60393 -8541
rect 61059 -8575 61093 -8541
rect 59861 -8955 59895 -8921
rect 60359 -8659 60393 -8625
rect 61059 -8659 61093 -8625
rect 59560 -9442 59594 -9408
rect 59032 -9550 59066 -9516
rect 53988 -9844 54022 -9806
rect 54916 -9844 54950 -9806
rect 59874 -9228 59908 -9194
rect 60384 -9228 60418 -9194
rect 55526 -10036 55560 -10002
rect 20390 -12008 20424 -11974
rect 16615 -12279 16703 -12245
rect 16615 -13189 16703 -13155
rect 17021 -12279 17109 -12245
rect 17021 -13189 17109 -13155
rect 17427 -12279 17515 -12245
rect 17427 -13189 17515 -13155
rect 17833 -12279 17921 -12245
rect 17833 -13189 17921 -13155
rect 18239 -12279 18327 -12245
rect 18239 -13189 18327 -13155
rect 18645 -12279 18733 -12245
rect 18645 -13189 18733 -13155
rect 19051 -12279 19139 -12245
rect 19051 -13189 19139 -13155
rect 19457 -12279 19545 -12245
rect 19457 -13189 19545 -13155
rect 19863 -12279 19951 -12245
rect 19863 -13189 19951 -13155
rect 20269 -12279 20357 -12245
rect 20269 -13189 20357 -13155
rect 20675 -12279 20763 -12245
rect 20675 -13189 20763 -13155
rect 21081 -12279 21169 -12245
rect 21081 -13189 21169 -13155
rect 21487 -12279 21575 -12245
rect 21487 -13189 21575 -13155
rect 21893 -12279 21981 -12245
rect 21893 -13189 21981 -13155
rect 22299 -12279 22387 -12245
rect 22299 -13189 22387 -13155
rect 22705 -12279 22793 -12245
rect 22705 -13189 22793 -13155
rect 23111 -12279 23199 -12245
rect 23111 -13189 23199 -13155
rect 23517 -12279 23605 -12245
rect 23517 -13189 23605 -13155
rect 23923 -12279 24011 -12245
rect 23923 -13189 24011 -13155
rect 24329 -12279 24417 -12245
rect 24329 -13189 24417 -13155
rect 24735 -12279 24823 -12245
rect 24735 -13189 24823 -13155
rect 25141 -12279 25229 -12245
rect 25141 -13189 25229 -13155
rect 53998 -12572 54032 -12534
rect 54926 -12572 54960 -12534
rect 53526 -12940 53614 -12906
rect 53998 -12928 54032 -12890
rect 54926 -12928 54960 -12890
rect 55334 -13002 55368 -12968
rect 53526 -13850 53614 -13816
rect 53858 -13728 53892 -13640
rect 54768 -13728 54802 -13640
rect 55046 -13594 55080 -13560
rect 55556 -13594 55590 -13560
rect 55882 -12890 55970 -12856
rect 55882 -13800 55970 -13766
rect 59560 -12935 59594 -12901
rect 59032 -13043 59066 -13009
rect 57133 -13191 57167 -13157
rect 57251 -13178 57285 -13144
rect 53526 -13958 53614 -13924
rect 53858 -14134 53892 -14046
rect 54768 -14134 54802 -14046
rect 55046 -14216 55080 -14182
rect 55556 -14216 55590 -14182
rect 53526 -14868 53614 -14834
rect 53988 -14888 54022 -14850
rect 54916 -14888 54950 -14850
rect 55324 -14808 55358 -14774
rect 55882 -14004 55970 -13970
rect 55882 -14914 55970 -14880
rect 56492 -13440 56530 -13406
rect 56492 -14368 56530 -14334
rect 59103 -13312 59137 -13278
rect 59103 -13840 59137 -13806
rect 59874 -13262 59908 -13228
rect 60384 -13262 60418 -13228
rect 59546 -13532 59580 -13498
rect 59546 -13842 59580 -13808
rect 59862 -13532 59896 -13498
rect 59862 -13842 59896 -13808
rect 60359 -13799 60393 -13765
rect 61059 -13799 61093 -13765
rect 60359 -13891 60393 -13857
rect 61059 -13891 61093 -13857
rect 59103 -14042 59137 -14008
rect 57133 -14631 57167 -14597
rect 57251 -14644 57285 -14610
rect 59103 -14570 59137 -14536
rect 59545 -14045 59579 -14011
rect 59545 -14355 59579 -14321
rect 59861 -14045 59895 -14011
rect 60359 -13975 60393 -13941
rect 61059 -13975 61093 -13941
rect 59861 -14355 59895 -14321
rect 60359 -14059 60393 -14025
rect 61059 -14059 61093 -14025
rect 59560 -14842 59594 -14808
rect 59032 -14950 59066 -14916
rect 53988 -15244 54022 -15206
rect 54916 -15244 54950 -15206
rect 59874 -14628 59908 -14594
rect 60384 -14628 60418 -14594
rect 55526 -15436 55560 -15402
rect 53998 -17972 54032 -17934
rect 54926 -17972 54960 -17934
rect 53526 -18340 53614 -18306
rect 53998 -18328 54032 -18290
rect 54926 -18328 54960 -18290
rect 55334 -18402 55368 -18368
rect 53526 -19250 53614 -19216
rect 53858 -19128 53892 -19040
rect 54768 -19128 54802 -19040
rect 55046 -18994 55080 -18960
rect 55556 -18994 55590 -18960
rect 55882 -18290 55970 -18256
rect 55882 -19200 55970 -19166
rect 59560 -18335 59594 -18301
rect 59032 -18443 59066 -18409
rect 57133 -18591 57167 -18557
rect 57251 -18578 57285 -18544
rect 53526 -19358 53614 -19324
rect 53858 -19534 53892 -19446
rect 54768 -19534 54802 -19446
rect 55046 -19616 55080 -19582
rect 55556 -19616 55590 -19582
rect 53526 -20268 53614 -20234
rect 53988 -20288 54022 -20250
rect 54916 -20288 54950 -20250
rect 55324 -20208 55358 -20174
rect 55882 -19404 55970 -19370
rect 55882 -20314 55970 -20280
rect 56492 -18840 56530 -18806
rect 56492 -19768 56530 -19734
rect 59103 -18712 59137 -18678
rect 59103 -19240 59137 -19206
rect 59874 -18662 59908 -18628
rect 60384 -18662 60418 -18628
rect 59546 -18932 59580 -18898
rect 59546 -19242 59580 -19208
rect 59862 -18932 59896 -18898
rect 59862 -19242 59896 -19208
rect 60359 -19199 60393 -19165
rect 61059 -19199 61093 -19165
rect 60359 -19291 60393 -19257
rect 61059 -19291 61093 -19257
rect 59103 -19442 59137 -19408
rect 57133 -20031 57167 -19997
rect 57251 -20044 57285 -20010
rect 59103 -19970 59137 -19936
rect 59545 -19445 59579 -19411
rect 59545 -19755 59579 -19721
rect 59861 -19445 59895 -19411
rect 60359 -19375 60393 -19341
rect 61059 -19375 61093 -19341
rect 59861 -19755 59895 -19721
rect 60359 -19459 60393 -19425
rect 61059 -19459 61093 -19425
rect 59560 -20242 59594 -20208
rect 59032 -20350 59066 -20316
rect 53988 -20644 54022 -20606
rect 54916 -20644 54950 -20606
rect 59874 -20028 59908 -19994
rect 60384 -20028 60418 -19994
rect 55526 -20836 55560 -20802
rect 53998 -23372 54032 -23334
rect 54926 -23372 54960 -23334
rect 53526 -23740 53614 -23706
rect 53998 -23728 54032 -23690
rect 54926 -23728 54960 -23690
rect 55334 -23802 55368 -23768
rect 53526 -24650 53614 -24616
rect 53858 -24528 53892 -24440
rect 54768 -24528 54802 -24440
rect 55046 -24394 55080 -24360
rect 55556 -24394 55590 -24360
rect 55882 -23690 55970 -23656
rect 55882 -24600 55970 -24566
rect 59560 -23735 59594 -23701
rect 59032 -23843 59066 -23809
rect 57133 -23991 57167 -23957
rect 57251 -23978 57285 -23944
rect 53526 -24758 53614 -24724
rect 53858 -24934 53892 -24846
rect 54768 -24934 54802 -24846
rect 55046 -25016 55080 -24982
rect 55556 -25016 55590 -24982
rect 53526 -25668 53614 -25634
rect 53988 -25688 54022 -25650
rect 54916 -25688 54950 -25650
rect 55324 -25608 55358 -25574
rect 55882 -24804 55970 -24770
rect 55882 -25714 55970 -25680
rect 56492 -24240 56530 -24206
rect 56492 -25168 56530 -25134
rect 59103 -24112 59137 -24078
rect 59103 -24640 59137 -24606
rect 59874 -24062 59908 -24028
rect 60384 -24062 60418 -24028
rect 59546 -24332 59580 -24298
rect 59546 -24642 59580 -24608
rect 59862 -24332 59896 -24298
rect 59862 -24642 59896 -24608
rect 60359 -24599 60393 -24565
rect 61059 -24599 61093 -24565
rect 60359 -24691 60393 -24657
rect 61059 -24691 61093 -24657
rect 59103 -24842 59137 -24808
rect 57133 -25431 57167 -25397
rect 57251 -25444 57285 -25410
rect 59103 -25370 59137 -25336
rect 59545 -24845 59579 -24811
rect 59545 -25155 59579 -25121
rect 59861 -24845 59895 -24811
rect 60359 -24775 60393 -24741
rect 61059 -24775 61093 -24741
rect 59861 -25155 59895 -25121
rect 60359 -24859 60393 -24825
rect 61059 -24859 61093 -24825
rect 59560 -25642 59594 -25608
rect 59032 -25750 59066 -25716
rect 53988 -26044 54022 -26006
rect 54916 -26044 54950 -26006
rect 59874 -25428 59908 -25394
rect 60384 -25428 60418 -25394
rect 55526 -26236 55560 -26202
rect 53998 -28772 54032 -28734
rect 54926 -28772 54960 -28734
rect 53526 -29140 53614 -29106
rect 53998 -29128 54032 -29090
rect 54926 -29128 54960 -29090
rect 55334 -29202 55368 -29168
rect 53526 -30050 53614 -30016
rect 53858 -29928 53892 -29840
rect 54768 -29928 54802 -29840
rect 55046 -29794 55080 -29760
rect 55556 -29794 55590 -29760
rect 55882 -29090 55970 -29056
rect 55882 -30000 55970 -29966
rect 59560 -29135 59594 -29101
rect 59032 -29243 59066 -29209
rect 57133 -29391 57167 -29357
rect 57251 -29378 57285 -29344
rect 53526 -30158 53614 -30124
rect 53858 -30334 53892 -30246
rect 54768 -30334 54802 -30246
rect 55046 -30416 55080 -30382
rect 55556 -30416 55590 -30382
rect 53526 -31068 53614 -31034
rect 53988 -31088 54022 -31050
rect 54916 -31088 54950 -31050
rect 55324 -31008 55358 -30974
rect 55882 -30204 55970 -30170
rect 55882 -31114 55970 -31080
rect 56492 -29640 56530 -29606
rect 56492 -30568 56530 -30534
rect 59103 -29512 59137 -29478
rect 59103 -30040 59137 -30006
rect 59874 -29462 59908 -29428
rect 60384 -29462 60418 -29428
rect 59546 -29732 59580 -29698
rect 59546 -30042 59580 -30008
rect 59862 -29732 59896 -29698
rect 59862 -30042 59896 -30008
rect 60359 -29999 60393 -29965
rect 61059 -29999 61093 -29965
rect 60359 -30091 60393 -30057
rect 61059 -30091 61093 -30057
rect 59103 -30242 59137 -30208
rect 57133 -30831 57167 -30797
rect 57251 -30844 57285 -30810
rect 59103 -30770 59137 -30736
rect 59545 -30245 59579 -30211
rect 59545 -30555 59579 -30521
rect 59861 -30245 59895 -30211
rect 60359 -30175 60393 -30141
rect 61059 -30175 61093 -30141
rect 59861 -30555 59895 -30521
rect 60359 -30259 60393 -30225
rect 61059 -30259 61093 -30225
rect 59560 -31042 59594 -31008
rect 59032 -31150 59066 -31116
rect 53988 -31444 54022 -31406
rect 54916 -31444 54950 -31406
rect 59874 -30828 59908 -30794
rect 60384 -30828 60418 -30794
rect 55526 -31636 55560 -31602
rect 53998 -34172 54032 -34134
rect 54926 -34172 54960 -34134
rect 53526 -34540 53614 -34506
rect 53998 -34528 54032 -34490
rect 54926 -34528 54960 -34490
rect 55334 -34602 55368 -34568
rect 53526 -35450 53614 -35416
rect 53858 -35328 53892 -35240
rect 54768 -35328 54802 -35240
rect 55046 -35194 55080 -35160
rect 55556 -35194 55590 -35160
rect 55882 -34490 55970 -34456
rect 55882 -35400 55970 -35366
rect 59560 -34535 59594 -34501
rect 59032 -34643 59066 -34609
rect 57133 -34791 57167 -34757
rect 57251 -34778 57285 -34744
rect 53526 -35558 53614 -35524
rect 53858 -35734 53892 -35646
rect 54768 -35734 54802 -35646
rect 55046 -35816 55080 -35782
rect 55556 -35816 55590 -35782
rect 53526 -36468 53614 -36434
rect 53988 -36488 54022 -36450
rect 54916 -36488 54950 -36450
rect 55324 -36408 55358 -36374
rect 55882 -35604 55970 -35570
rect 55882 -36514 55970 -36480
rect 56492 -35040 56530 -35006
rect 56492 -35968 56530 -35934
rect 59103 -34912 59137 -34878
rect 59103 -35440 59137 -35406
rect 59874 -34862 59908 -34828
rect 60384 -34862 60418 -34828
rect 59546 -35132 59580 -35098
rect 59546 -35442 59580 -35408
rect 59862 -35132 59896 -35098
rect 59862 -35442 59896 -35408
rect 60359 -35399 60393 -35365
rect 61059 -35399 61093 -35365
rect 60359 -35491 60393 -35457
rect 61059 -35491 61093 -35457
rect 59103 -35642 59137 -35608
rect 57133 -36231 57167 -36197
rect 57251 -36244 57285 -36210
rect 59103 -36170 59137 -36136
rect 59545 -35645 59579 -35611
rect 59545 -35955 59579 -35921
rect 59861 -35645 59895 -35611
rect 60359 -35575 60393 -35541
rect 61059 -35575 61093 -35541
rect 59861 -35955 59895 -35921
rect 60359 -35659 60393 -35625
rect 61059 -35659 61093 -35625
rect 59560 -36442 59594 -36408
rect 59032 -36550 59066 -36516
rect 53988 -36844 54022 -36806
rect 54916 -36844 54950 -36806
rect 59874 -36228 59908 -36194
rect 60384 -36228 60418 -36194
rect 55526 -37036 55560 -37002
rect 75586 -38637 75620 -38603
rect 75862 -38637 75896 -38603
rect 76136 -38637 76170 -38603
rect 76412 -38637 76446 -38603
rect 76688 -38637 76722 -38603
rect 77835 -39163 77869 -39129
rect 78293 -39163 78327 -39129
rect 77613 -39387 77647 -39353
rect 77739 -39387 77773 -39353
rect 53998 -39572 54032 -39534
rect 54926 -39572 54960 -39534
rect 77915 -39387 77949 -39353
rect 78011 -39387 78045 -39353
rect 78164 -39387 78198 -39353
rect 78374 -39387 78408 -39353
rect 78470 -39387 78504 -39353
rect 78664 -39387 78698 -39353
rect 78805 -39387 78839 -39353
rect 78913 -39387 78947 -39353
rect 80818 -39437 80852 -39403
rect 81051 -39437 81085 -39403
rect 81143 -39437 81177 -39403
rect 81227 -39437 81261 -39403
rect 81311 -39437 81345 -39403
rect 81516 -39437 81550 -39403
rect 81690 -39437 81724 -39403
rect 81858 -39437 81892 -39403
rect 82027 -39437 82061 -39403
rect 82194 -39437 82228 -39403
rect 82362 -39437 82396 -39403
rect 82529 -39437 82563 -39403
rect 82988 -39437 83022 -39403
rect 83162 -39437 83196 -39403
rect 83330 -39437 83364 -39403
rect 83499 -39437 83533 -39403
rect 83666 -39437 83700 -39403
rect 83834 -39437 83868 -39403
rect 84001 -39437 84035 -39403
rect 84460 -39437 84494 -39403
rect 84634 -39437 84668 -39403
rect 84802 -39437 84836 -39403
rect 84971 -39437 85005 -39403
rect 85138 -39437 85172 -39403
rect 85306 -39437 85340 -39403
rect 85473 -39437 85507 -39403
rect 85932 -39437 85966 -39403
rect 86106 -39437 86140 -39403
rect 86274 -39437 86308 -39403
rect 86443 -39437 86477 -39403
rect 86610 -39437 86644 -39403
rect 86778 -39437 86812 -39403
rect 86945 -39437 86979 -39403
rect 87404 -39437 87438 -39403
rect 87578 -39437 87612 -39403
rect 87746 -39437 87780 -39403
rect 87915 -39437 87949 -39403
rect 88082 -39437 88116 -39403
rect 88250 -39437 88284 -39403
rect 88417 -39437 88451 -39403
rect 53526 -39940 53614 -39906
rect 53998 -39928 54032 -39890
rect 54926 -39928 54960 -39890
rect 55334 -40002 55368 -39968
rect 53526 -40850 53614 -40816
rect 53858 -40728 53892 -40640
rect 54768 -40728 54802 -40640
rect 55046 -40594 55080 -40560
rect 55556 -40594 55590 -40560
rect 55882 -39890 55970 -39856
rect 55882 -40800 55970 -40766
rect 59560 -39935 59594 -39901
rect 59032 -40043 59066 -40009
rect 57133 -40191 57167 -40157
rect 57251 -40178 57285 -40144
rect 77613 -39937 77647 -39903
rect 77739 -39937 77773 -39903
rect 77915 -39937 77949 -39903
rect 78011 -39937 78045 -39903
rect 80868 -39977 80902 -39943
rect 53526 -40958 53614 -40924
rect 53858 -41134 53892 -41046
rect 54768 -41134 54802 -41046
rect 55046 -41216 55080 -41182
rect 55556 -41216 55590 -41182
rect 53526 -41868 53614 -41834
rect 53988 -41888 54022 -41850
rect 54916 -41888 54950 -41850
rect 55324 -41808 55358 -41774
rect 55882 -41004 55970 -40970
rect 55882 -41914 55970 -41880
rect 56492 -40440 56530 -40406
rect 56492 -41368 56530 -41334
rect 59103 -40312 59137 -40278
rect 59103 -40840 59137 -40806
rect 59874 -40262 59908 -40228
rect 60384 -40262 60418 -40228
rect 77835 -40161 77869 -40127
rect 59546 -40532 59580 -40498
rect 59546 -40842 59580 -40808
rect 59862 -40532 59896 -40498
rect 59862 -40842 59896 -40808
rect 77652 -40637 77686 -40603
rect 77793 -40637 77827 -40603
rect 77901 -40637 77935 -40603
rect 60359 -40799 60393 -40765
rect 61059 -40799 61093 -40765
rect 60359 -40891 60393 -40857
rect 61059 -40891 61093 -40857
rect 59103 -41042 59137 -41008
rect 57133 -41631 57167 -41597
rect 57251 -41644 57285 -41610
rect 59103 -41570 59137 -41536
rect 59545 -41045 59579 -41011
rect 59545 -41355 59579 -41321
rect 59861 -41045 59895 -41011
rect 60359 -40975 60393 -40941
rect 61059 -40975 61093 -40941
rect 59861 -41355 59895 -41321
rect 60359 -41059 60393 -41025
rect 61059 -41059 61093 -41025
rect 77652 -41177 77686 -41143
rect 77793 -41177 77827 -41143
rect 77901 -41177 77935 -41143
rect 78073 -41177 78107 -41143
rect 78199 -41177 78233 -41143
rect 78375 -41177 78409 -41143
rect 78471 -41177 78505 -41143
rect 78295 -41401 78329 -41367
rect 59560 -41842 59594 -41808
rect 59032 -41950 59066 -41916
rect 53988 -42244 54022 -42206
rect 54916 -42244 54950 -42206
rect 59874 -41628 59908 -41594
rect 60384 -41628 60418 -41594
rect 77652 -41877 77686 -41843
rect 77793 -41877 77827 -41843
rect 77901 -41877 77935 -41843
rect 55526 -42436 55560 -42402
rect 77654 -42431 77688 -42397
rect 77795 -42431 77829 -42397
rect 77903 -42431 77937 -42397
rect 78579 -42903 78613 -42869
rect 77609 -43127 77643 -43093
rect 77755 -43127 77789 -43093
rect 77861 -43127 77895 -43093
rect 77957 -43127 77991 -43093
rect 78068 -43127 78102 -43093
rect 78357 -43127 78391 -43093
rect 78483 -43127 78517 -43093
rect 78659 -43127 78693 -43093
rect 78755 -43127 78789 -43093
rect 77609 -43663 77643 -43629
rect 77755 -43663 77789 -43629
rect 77861 -43663 77895 -43629
rect 77957 -43663 77991 -43629
rect 78068 -43663 78102 -43629
rect 82904 -43937 82938 -43903
rect 83040 -43937 83074 -43903
rect 83143 -43937 83177 -43903
rect 83378 -43937 83412 -43903
rect 83611 -43937 83645 -43903
rect 83703 -43937 83737 -43903
rect 83787 -43937 83821 -43903
rect 83871 -43937 83905 -43903
rect 84076 -43937 84110 -43903
rect 84250 -43937 84284 -43903
rect 84418 -43937 84452 -43903
rect 84587 -43937 84621 -43903
rect 84754 -43937 84788 -43903
rect 84922 -43937 84956 -43903
rect 85089 -43937 85123 -43903
rect 85548 -43937 85582 -43903
rect 85722 -43937 85756 -43903
rect 85890 -43937 85924 -43903
rect 86059 -43937 86093 -43903
rect 86226 -43937 86260 -43903
rect 86394 -43937 86428 -43903
rect 86561 -43937 86595 -43903
rect 87020 -43937 87054 -43903
rect 87194 -43937 87228 -43903
rect 87362 -43937 87396 -43903
rect 87531 -43937 87565 -43903
rect 87698 -43937 87732 -43903
rect 87866 -43937 87900 -43903
rect 88033 -43937 88067 -43903
rect 88492 -43937 88526 -43903
rect 88666 -43937 88700 -43903
rect 88834 -43937 88868 -43903
rect 89003 -43937 89037 -43903
rect 89170 -43937 89204 -43903
rect 89338 -43937 89372 -43903
rect 89505 -43937 89539 -43903
rect 89964 -43937 89998 -43903
rect 90138 -43937 90172 -43903
rect 90306 -43937 90340 -43903
rect 90475 -43937 90509 -43903
rect 90642 -43937 90676 -43903
rect 90810 -43937 90844 -43903
rect 90977 -43937 91011 -43903
rect 77609 -44359 77643 -44325
rect 77755 -44359 77789 -44325
rect 77861 -44359 77895 -44325
rect 77957 -44359 77991 -44325
rect 78068 -44359 78102 -44325
rect 53998 -44972 54032 -44934
rect 54926 -44972 54960 -44934
rect 77609 -44897 77643 -44863
rect 77755 -44897 77789 -44863
rect 77861 -44897 77895 -44863
rect 77957 -44897 77991 -44863
rect 78068 -44897 78102 -44863
rect 53526 -45340 53614 -45306
rect 53998 -45328 54032 -45290
rect 54926 -45328 54960 -45290
rect 55334 -45402 55368 -45368
rect 53526 -46250 53614 -46216
rect 53858 -46128 53892 -46040
rect 54768 -46128 54802 -46040
rect 55046 -45994 55080 -45960
rect 55556 -45994 55590 -45960
rect 55882 -45290 55970 -45256
rect 55882 -46200 55970 -46166
rect 59560 -45335 59594 -45301
rect 59032 -45443 59066 -45409
rect 57133 -45591 57167 -45557
rect 57251 -45578 57285 -45544
rect 77751 -45370 77785 -45336
rect 53526 -46358 53614 -46324
rect 53858 -46534 53892 -46446
rect 54768 -46534 54802 -46446
rect 55046 -46616 55080 -46582
rect 55556 -46616 55590 -46582
rect 53526 -47268 53614 -47234
rect 53988 -47288 54022 -47250
rect 54916 -47288 54950 -47250
rect 55324 -47208 55358 -47174
rect 55882 -46404 55970 -46370
rect 55882 -47314 55970 -47280
rect 56492 -45840 56530 -45806
rect 56492 -46768 56530 -46734
rect 59103 -45712 59137 -45678
rect 59103 -46240 59137 -46206
rect 59874 -45662 59908 -45628
rect 60384 -45662 60418 -45628
rect 77613 -45643 77647 -45609
rect 77823 -45603 77857 -45569
rect 77919 -45597 77953 -45563
rect 78112 -45597 78146 -45563
rect 78755 -45373 78789 -45339
rect 78253 -45597 78287 -45563
rect 78361 -45597 78395 -45563
rect 78533 -45597 78567 -45563
rect 78659 -45597 78693 -45563
rect 78835 -45597 78869 -45563
rect 78931 -45597 78965 -45563
rect 59546 -45932 59580 -45898
rect 59546 -46242 59580 -46208
rect 59862 -45932 59896 -45898
rect 59862 -46242 59896 -46208
rect 60359 -46199 60393 -46165
rect 61059 -46199 61093 -46165
rect 60359 -46291 60393 -46257
rect 61059 -46291 61093 -46257
rect 59103 -46442 59137 -46408
rect 57133 -47031 57167 -46997
rect 57251 -47044 57285 -47010
rect 59103 -46970 59137 -46936
rect 59545 -46445 59579 -46411
rect 59545 -46755 59579 -46721
rect 59861 -46445 59895 -46411
rect 60359 -46375 60393 -46341
rect 61059 -46375 61093 -46341
rect 59861 -46755 59895 -46721
rect 60359 -46459 60393 -46425
rect 61059 -46459 61093 -46425
rect 75586 -46677 75620 -46643
rect 75862 -46677 75896 -46643
rect 76136 -46677 76170 -46643
rect 76412 -46677 76446 -46643
rect 76688 -46677 76722 -46643
rect 59560 -47242 59594 -47208
rect 59032 -47350 59066 -47316
rect 53988 -47644 54022 -47606
rect 54916 -47644 54950 -47606
rect 59874 -47028 59908 -46994
rect 60384 -47028 60418 -46994
rect 77835 -47203 77869 -47169
rect 78293 -47203 78327 -47169
rect 77613 -47427 77647 -47393
rect 77739 -47427 77773 -47393
rect 77915 -47427 77949 -47393
rect 78011 -47427 78045 -47393
rect 78164 -47427 78198 -47393
rect 78374 -47427 78408 -47393
rect 78470 -47427 78504 -47393
rect 78664 -47427 78698 -47393
rect 78805 -47427 78839 -47393
rect 78913 -47427 78947 -47393
rect 55526 -47836 55560 -47802
rect 77613 -47977 77647 -47943
rect 77739 -47977 77773 -47943
rect 77915 -47977 77949 -47943
rect 78011 -47977 78045 -47943
rect 77835 -48201 77869 -48167
rect 82904 -48077 82938 -48043
rect 83040 -48077 83074 -48043
rect 83143 -48077 83177 -48043
rect 83378 -48077 83412 -48043
rect 83611 -48077 83645 -48043
rect 83703 -48077 83737 -48043
rect 83787 -48077 83821 -48043
rect 83871 -48077 83905 -48043
rect 84076 -48077 84110 -48043
rect 84250 -48077 84284 -48043
rect 84418 -48077 84452 -48043
rect 84587 -48077 84621 -48043
rect 84754 -48077 84788 -48043
rect 84922 -48077 84956 -48043
rect 85089 -48077 85123 -48043
rect 85548 -48077 85582 -48043
rect 85722 -48077 85756 -48043
rect 85890 -48077 85924 -48043
rect 86059 -48077 86093 -48043
rect 86226 -48077 86260 -48043
rect 86394 -48077 86428 -48043
rect 86561 -48077 86595 -48043
rect 87020 -48077 87054 -48043
rect 87194 -48077 87228 -48043
rect 87362 -48077 87396 -48043
rect 87531 -48077 87565 -48043
rect 87698 -48077 87732 -48043
rect 87866 -48077 87900 -48043
rect 88033 -48077 88067 -48043
rect 88492 -48077 88526 -48043
rect 88666 -48077 88700 -48043
rect 88834 -48077 88868 -48043
rect 89003 -48077 89037 -48043
rect 89170 -48077 89204 -48043
rect 89338 -48077 89372 -48043
rect 89505 -48077 89539 -48043
rect 89964 -48077 89998 -48043
rect 90138 -48077 90172 -48043
rect 90306 -48077 90340 -48043
rect 90475 -48077 90509 -48043
rect 90642 -48077 90676 -48043
rect 90810 -48077 90844 -48043
rect 90977 -48077 91011 -48043
rect 77652 -48677 77686 -48643
rect 77793 -48677 77827 -48643
rect 77901 -48677 77935 -48643
rect 77652 -49217 77686 -49183
rect 77793 -49217 77827 -49183
rect 77901 -49217 77935 -49183
rect 78073 -49217 78107 -49183
rect 78199 -49217 78233 -49183
rect 78375 -49217 78409 -49183
rect 78471 -49217 78505 -49183
rect 78295 -49441 78329 -49407
rect 77652 -49917 77686 -49883
rect 77793 -49917 77827 -49883
rect 77901 -49917 77935 -49883
rect 53998 -50372 54032 -50334
rect 54926 -50372 54960 -50334
rect 53526 -50740 53614 -50706
rect 77654 -50471 77688 -50437
rect 53998 -50728 54032 -50690
rect 54926 -50728 54960 -50690
rect 55334 -50802 55368 -50768
rect 53526 -51650 53614 -51616
rect 53858 -51528 53892 -51440
rect 54768 -51528 54802 -51440
rect 55046 -51394 55080 -51360
rect 55556 -51394 55590 -51360
rect 55882 -50690 55970 -50656
rect 55882 -51600 55970 -51566
rect 77795 -50471 77829 -50437
rect 77903 -50471 77937 -50437
rect 59560 -50735 59594 -50701
rect 59032 -50843 59066 -50809
rect 57133 -50991 57167 -50957
rect 57251 -50978 57285 -50944
rect 53526 -51758 53614 -51724
rect 53858 -51934 53892 -51846
rect 54768 -51934 54802 -51846
rect 55046 -52016 55080 -51982
rect 55556 -52016 55590 -51982
rect 53526 -52668 53614 -52634
rect 53988 -52688 54022 -52650
rect 54916 -52688 54950 -52650
rect 55324 -52608 55358 -52574
rect 55882 -51804 55970 -51770
rect 55882 -52714 55970 -52680
rect 56492 -51240 56530 -51206
rect 56492 -52168 56530 -52134
rect 59103 -51112 59137 -51078
rect 59103 -51640 59137 -51606
rect 59874 -51062 59908 -51028
rect 60384 -51062 60418 -51028
rect 78579 -50943 78613 -50909
rect 77609 -51167 77643 -51133
rect 59546 -51332 59580 -51298
rect 59546 -51642 59580 -51608
rect 59862 -51332 59896 -51298
rect 59862 -51642 59896 -51608
rect 77755 -51167 77789 -51133
rect 77861 -51167 77895 -51133
rect 77957 -51167 77991 -51133
rect 78068 -51167 78102 -51133
rect 78357 -51167 78391 -51133
rect 78483 -51167 78517 -51133
rect 78659 -51167 78693 -51133
rect 78755 -51167 78789 -51133
rect 60359 -51599 60393 -51565
rect 61059 -51599 61093 -51565
rect 60359 -51691 60393 -51657
rect 61059 -51691 61093 -51657
rect 59103 -51842 59137 -51808
rect 57133 -52431 57167 -52397
rect 57251 -52444 57285 -52410
rect 59103 -52370 59137 -52336
rect 77609 -51703 77643 -51669
rect 77755 -51703 77789 -51669
rect 77861 -51703 77895 -51669
rect 77957 -51703 77991 -51669
rect 78068 -51703 78102 -51669
rect 59545 -51845 59579 -51811
rect 59545 -52155 59579 -52121
rect 59861 -51845 59895 -51811
rect 60359 -51775 60393 -51741
rect 61059 -51775 61093 -51741
rect 59861 -52155 59895 -52121
rect 60359 -51859 60393 -51825
rect 61059 -51859 61093 -51825
rect 82904 -51727 82938 -51693
rect 83040 -51727 83074 -51693
rect 83143 -51727 83177 -51693
rect 83378 -51727 83412 -51693
rect 83611 -51727 83645 -51693
rect 83703 -51727 83737 -51693
rect 83787 -51727 83821 -51693
rect 83871 -51727 83905 -51693
rect 84076 -51727 84110 -51693
rect 84250 -51727 84284 -51693
rect 84418 -51727 84452 -51693
rect 84587 -51727 84621 -51693
rect 84754 -51727 84788 -51693
rect 84922 -51727 84956 -51693
rect 85089 -51727 85123 -51693
rect 85548 -51727 85582 -51693
rect 85722 -51727 85756 -51693
rect 85890 -51727 85924 -51693
rect 86059 -51727 86093 -51693
rect 86226 -51727 86260 -51693
rect 86394 -51727 86428 -51693
rect 86561 -51727 86595 -51693
rect 87020 -51727 87054 -51693
rect 87194 -51727 87228 -51693
rect 87362 -51727 87396 -51693
rect 87531 -51727 87565 -51693
rect 87698 -51727 87732 -51693
rect 87866 -51727 87900 -51693
rect 88033 -51727 88067 -51693
rect 88492 -51727 88526 -51693
rect 88666 -51727 88700 -51693
rect 88834 -51727 88868 -51693
rect 89003 -51727 89037 -51693
rect 89170 -51727 89204 -51693
rect 89338 -51727 89372 -51693
rect 89505 -51727 89539 -51693
rect 89964 -51727 89998 -51693
rect 90138 -51727 90172 -51693
rect 90306 -51727 90340 -51693
rect 90475 -51727 90509 -51693
rect 90642 -51727 90676 -51693
rect 90810 -51727 90844 -51693
rect 90977 -51727 91011 -51693
rect 59560 -52642 59594 -52608
rect 59032 -52750 59066 -52716
rect 53988 -53044 54022 -53006
rect 54916 -53044 54950 -53006
rect 59874 -52428 59908 -52394
rect 60384 -52428 60418 -52394
rect 77609 -52399 77643 -52365
rect 77755 -52399 77789 -52365
rect 77861 -52399 77895 -52365
rect 77957 -52399 77991 -52365
rect 78068 -52399 78102 -52365
rect 77609 -52937 77643 -52903
rect 77755 -52937 77789 -52903
rect 77861 -52937 77895 -52903
rect 77957 -52937 77991 -52903
rect 78068 -52937 78102 -52903
rect 55526 -53236 55560 -53202
rect 77751 -53410 77785 -53376
rect 77613 -53683 77647 -53649
rect 77823 -53643 77857 -53609
rect 77919 -53637 77953 -53603
rect 78112 -53637 78146 -53603
rect 78755 -53413 78789 -53379
rect 78253 -53637 78287 -53603
rect 78361 -53637 78395 -53603
rect 78533 -53637 78567 -53603
rect 78659 -53637 78693 -53603
rect 78835 -53637 78869 -53603
rect 78931 -53637 78965 -53603
rect 53998 -55772 54032 -55734
rect 54926 -55772 54960 -55734
rect 53526 -56140 53614 -56106
rect 53998 -56128 54032 -56090
rect 54926 -56128 54960 -56090
rect 55334 -56202 55368 -56168
rect 53526 -57050 53614 -57016
rect 53858 -56928 53892 -56840
rect 54768 -56928 54802 -56840
rect 55046 -56794 55080 -56760
rect 55556 -56794 55590 -56760
rect 55882 -56090 55970 -56056
rect 55882 -57000 55970 -56966
rect 59560 -56135 59594 -56101
rect 59032 -56243 59066 -56209
rect 57133 -56391 57167 -56357
rect 57251 -56378 57285 -56344
rect 53526 -57158 53614 -57124
rect 53858 -57334 53892 -57246
rect 54768 -57334 54802 -57246
rect 55046 -57416 55080 -57382
rect 55556 -57416 55590 -57382
rect 53526 -58068 53614 -58034
rect 53988 -58088 54022 -58050
rect 54916 -58088 54950 -58050
rect 55324 -58008 55358 -57974
rect 55882 -57204 55970 -57170
rect 55882 -58114 55970 -58080
rect 56492 -56640 56530 -56606
rect 56492 -57568 56530 -57534
rect 59103 -56512 59137 -56478
rect 59103 -57040 59137 -57006
rect 59874 -56462 59908 -56428
rect 60384 -56462 60418 -56428
rect 59546 -56732 59580 -56698
rect 59546 -57042 59580 -57008
rect 59862 -56732 59896 -56698
rect 59862 -57042 59896 -57008
rect 60359 -56999 60393 -56965
rect 61059 -56999 61093 -56965
rect 60359 -57091 60393 -57057
rect 61059 -57091 61093 -57057
rect 59103 -57242 59137 -57208
rect 57133 -57831 57167 -57797
rect 57251 -57844 57285 -57810
rect 59103 -57770 59137 -57736
rect 59545 -57245 59579 -57211
rect 59545 -57555 59579 -57521
rect 59861 -57245 59895 -57211
rect 60359 -57175 60393 -57141
rect 61059 -57175 61093 -57141
rect 59861 -57555 59895 -57521
rect 60359 -57259 60393 -57225
rect 61059 -57259 61093 -57225
rect 59560 -58042 59594 -58008
rect 59032 -58150 59066 -58116
rect 53988 -58444 54022 -58406
rect 54916 -58444 54950 -58406
rect 59874 -57828 59908 -57794
rect 60384 -57828 60418 -57794
rect 55526 -58636 55560 -58602
rect 53998 -61172 54032 -61134
rect 54926 -61172 54960 -61134
rect 53526 -61540 53614 -61506
rect 53998 -61528 54032 -61490
rect 54926 -61528 54960 -61490
rect 55334 -61602 55368 -61568
rect 53526 -62450 53614 -62416
rect 53858 -62328 53892 -62240
rect 54768 -62328 54802 -62240
rect 55046 -62194 55080 -62160
rect 55556 -62194 55590 -62160
rect 55882 -61490 55970 -61456
rect 55882 -62400 55970 -62366
rect 59560 -61535 59594 -61501
rect 59032 -61643 59066 -61609
rect 57133 -61791 57167 -61757
rect 57251 -61778 57285 -61744
rect 53526 -62558 53614 -62524
rect 53858 -62734 53892 -62646
rect 54768 -62734 54802 -62646
rect 55046 -62816 55080 -62782
rect 55556 -62816 55590 -62782
rect 53526 -63468 53614 -63434
rect 53988 -63488 54022 -63450
rect 54916 -63488 54950 -63450
rect 55324 -63408 55358 -63374
rect 55882 -62604 55970 -62570
rect 55882 -63514 55970 -63480
rect 56492 -62040 56530 -62006
rect 56492 -62968 56530 -62934
rect 59103 -61912 59137 -61878
rect 59103 -62440 59137 -62406
rect 59874 -61862 59908 -61828
rect 60384 -61862 60418 -61828
rect 59546 -62132 59580 -62098
rect 59546 -62442 59580 -62408
rect 59862 -62132 59896 -62098
rect 59862 -62442 59896 -62408
rect 60359 -62399 60393 -62365
rect 61059 -62399 61093 -62365
rect 60359 -62491 60393 -62457
rect 61059 -62491 61093 -62457
rect 59103 -62642 59137 -62608
rect 57133 -63231 57167 -63197
rect 57251 -63244 57285 -63210
rect 59103 -63170 59137 -63136
rect 59545 -62645 59579 -62611
rect 59545 -62955 59579 -62921
rect 59861 -62645 59895 -62611
rect 60359 -62575 60393 -62541
rect 61059 -62575 61093 -62541
rect 59861 -62955 59895 -62921
rect 60359 -62659 60393 -62625
rect 61059 -62659 61093 -62625
rect 59560 -63442 59594 -63408
rect 59032 -63550 59066 -63516
rect 53988 -63844 54022 -63806
rect 54916 -63844 54950 -63806
rect 59874 -63228 59908 -63194
rect 60384 -63228 60418 -63194
rect 55526 -64036 55560 -64002
rect 53998 -66572 54032 -66534
rect 54926 -66572 54960 -66534
rect 53526 -66940 53614 -66906
rect 53998 -66928 54032 -66890
rect 54926 -66928 54960 -66890
rect 55334 -67002 55368 -66968
rect 53526 -67850 53614 -67816
rect 53858 -67728 53892 -67640
rect 54768 -67728 54802 -67640
rect 55046 -67594 55080 -67560
rect 55556 -67594 55590 -67560
rect 55882 -66890 55970 -66856
rect 55882 -67800 55970 -67766
rect 59560 -66935 59594 -66901
rect 59032 -67043 59066 -67009
rect 57133 -67191 57167 -67157
rect 57251 -67178 57285 -67144
rect 53526 -67958 53614 -67924
rect 53858 -68134 53892 -68046
rect 54768 -68134 54802 -68046
rect 55046 -68216 55080 -68182
rect 55556 -68216 55590 -68182
rect 53526 -68868 53614 -68834
rect 53988 -68888 54022 -68850
rect 54916 -68888 54950 -68850
rect 55324 -68808 55358 -68774
rect 55882 -68004 55970 -67970
rect 55882 -68914 55970 -68880
rect 56492 -67440 56530 -67406
rect 56492 -68368 56530 -68334
rect 59103 -67312 59137 -67278
rect 59103 -67840 59137 -67806
rect 59874 -67262 59908 -67228
rect 60384 -67262 60418 -67228
rect 59546 -67532 59580 -67498
rect 59546 -67842 59580 -67808
rect 59862 -67532 59896 -67498
rect 59862 -67842 59896 -67808
rect 60359 -67799 60393 -67765
rect 61059 -67799 61093 -67765
rect 60359 -67891 60393 -67857
rect 61059 -67891 61093 -67857
rect 59103 -68042 59137 -68008
rect 57133 -68631 57167 -68597
rect 57251 -68644 57285 -68610
rect 59103 -68570 59137 -68536
rect 59545 -68045 59579 -68011
rect 59545 -68355 59579 -68321
rect 59861 -68045 59895 -68011
rect 60359 -67975 60393 -67941
rect 61059 -67975 61093 -67941
rect 59861 -68355 59895 -68321
rect 60359 -68059 60393 -68025
rect 61059 -68059 61093 -68025
rect 59560 -68842 59594 -68808
rect 59032 -68950 59066 -68916
rect 53988 -69244 54022 -69206
rect 54916 -69244 54950 -69206
rect 59874 -68628 59908 -68594
rect 60384 -68628 60418 -68594
rect 55526 -69436 55560 -69402
rect 53998 -71972 54032 -71934
rect 54926 -71972 54960 -71934
rect 53526 -72340 53614 -72306
rect 53998 -72328 54032 -72290
rect 54926 -72328 54960 -72290
rect 55334 -72402 55368 -72368
rect 53526 -73250 53614 -73216
rect 53858 -73128 53892 -73040
rect 54768 -73128 54802 -73040
rect 55046 -72994 55080 -72960
rect 55556 -72994 55590 -72960
rect 55882 -72290 55970 -72256
rect 55882 -73200 55970 -73166
rect 59560 -72335 59594 -72301
rect 59032 -72443 59066 -72409
rect 57133 -72591 57167 -72557
rect 57251 -72578 57285 -72544
rect 53526 -73358 53614 -73324
rect 53858 -73534 53892 -73446
rect 54768 -73534 54802 -73446
rect 55046 -73616 55080 -73582
rect 55556 -73616 55590 -73582
rect 53526 -74268 53614 -74234
rect 53988 -74288 54022 -74250
rect 54916 -74288 54950 -74250
rect 55324 -74208 55358 -74174
rect 55882 -73404 55970 -73370
rect 55882 -74314 55970 -74280
rect 56492 -72840 56530 -72806
rect 56492 -73768 56530 -73734
rect 59103 -72712 59137 -72678
rect 59103 -73240 59137 -73206
rect 59874 -72662 59908 -72628
rect 60384 -72662 60418 -72628
rect 59546 -72932 59580 -72898
rect 59546 -73242 59580 -73208
rect 59862 -72932 59896 -72898
rect 59862 -73242 59896 -73208
rect 60359 -73199 60393 -73165
rect 61059 -73199 61093 -73165
rect 60359 -73291 60393 -73257
rect 61059 -73291 61093 -73257
rect 59103 -73442 59137 -73408
rect 57133 -74031 57167 -73997
rect 57251 -74044 57285 -74010
rect 59103 -73970 59137 -73936
rect 59545 -73445 59579 -73411
rect 59545 -73755 59579 -73721
rect 59861 -73445 59895 -73411
rect 60359 -73375 60393 -73341
rect 61059 -73375 61093 -73341
rect 59861 -73755 59895 -73721
rect 60359 -73459 60393 -73425
rect 61059 -73459 61093 -73425
rect 59560 -74242 59594 -74208
rect 59032 -74350 59066 -74316
rect 53988 -74644 54022 -74606
rect 54916 -74644 54950 -74606
rect 59874 -74028 59908 -73994
rect 60384 -74028 60418 -73994
rect 55526 -74836 55560 -74802
rect 53998 -77372 54032 -77334
rect 54926 -77372 54960 -77334
rect 53526 -77740 53614 -77706
rect 53998 -77728 54032 -77690
rect 54926 -77728 54960 -77690
rect 55334 -77802 55368 -77768
rect 53526 -78650 53614 -78616
rect 53858 -78528 53892 -78440
rect 54768 -78528 54802 -78440
rect 55046 -78394 55080 -78360
rect 55556 -78394 55590 -78360
rect 55882 -77690 55970 -77656
rect 55882 -78600 55970 -78566
rect 59560 -77735 59594 -77701
rect 59032 -77843 59066 -77809
rect 57133 -77991 57167 -77957
rect 57251 -77978 57285 -77944
rect 53526 -78758 53614 -78724
rect 53858 -78934 53892 -78846
rect 54768 -78934 54802 -78846
rect 55046 -79016 55080 -78982
rect 55556 -79016 55590 -78982
rect 53526 -79668 53614 -79634
rect 53988 -79688 54022 -79650
rect 54916 -79688 54950 -79650
rect 55324 -79608 55358 -79574
rect 55882 -78804 55970 -78770
rect 55882 -79714 55970 -79680
rect 56492 -78240 56530 -78206
rect 56492 -79168 56530 -79134
rect 59103 -78112 59137 -78078
rect 59103 -78640 59137 -78606
rect 59874 -78062 59908 -78028
rect 60384 -78062 60418 -78028
rect 59546 -78332 59580 -78298
rect 59546 -78642 59580 -78608
rect 59862 -78332 59896 -78298
rect 59862 -78642 59896 -78608
rect 60359 -78599 60393 -78565
rect 61059 -78599 61093 -78565
rect 60359 -78691 60393 -78657
rect 61059 -78691 61093 -78657
rect 59103 -78842 59137 -78808
rect 57133 -79431 57167 -79397
rect 57251 -79444 57285 -79410
rect 59103 -79370 59137 -79336
rect 59545 -78845 59579 -78811
rect 59545 -79155 59579 -79121
rect 59861 -78845 59895 -78811
rect 60359 -78775 60393 -78741
rect 61059 -78775 61093 -78741
rect 59861 -79155 59895 -79121
rect 60359 -78859 60393 -78825
rect 61059 -78859 61093 -78825
rect 59560 -79642 59594 -79608
rect 59032 -79750 59066 -79716
rect 53988 -80044 54022 -80006
rect 54916 -80044 54950 -80006
rect 59874 -79428 59908 -79394
rect 60384 -79428 60418 -79394
rect 55526 -80236 55560 -80202
rect 53998 -82772 54032 -82734
rect 54926 -82772 54960 -82734
rect 53526 -83140 53614 -83106
rect 53998 -83128 54032 -83090
rect 54926 -83128 54960 -83090
rect 55334 -83202 55368 -83168
rect 53526 -84050 53614 -84016
rect 53858 -83928 53892 -83840
rect 54768 -83928 54802 -83840
rect 55046 -83794 55080 -83760
rect 55556 -83794 55590 -83760
rect 55882 -83090 55970 -83056
rect 55882 -84000 55970 -83966
rect 59560 -83135 59594 -83101
rect 59032 -83243 59066 -83209
rect 57133 -83391 57167 -83357
rect 57251 -83378 57285 -83344
rect 53526 -84158 53614 -84124
rect 53858 -84334 53892 -84246
rect 54768 -84334 54802 -84246
rect 55046 -84416 55080 -84382
rect 55556 -84416 55590 -84382
rect 53526 -85068 53614 -85034
rect 53988 -85088 54022 -85050
rect 54916 -85088 54950 -85050
rect 55324 -85008 55358 -84974
rect 55882 -84204 55970 -84170
rect 55882 -85114 55970 -85080
rect 56492 -83640 56530 -83606
rect 56492 -84568 56530 -84534
rect 59103 -83512 59137 -83478
rect 59103 -84040 59137 -84006
rect 59874 -83462 59908 -83428
rect 60384 -83462 60418 -83428
rect 59546 -83732 59580 -83698
rect 59546 -84042 59580 -84008
rect 59862 -83732 59896 -83698
rect 59862 -84042 59896 -84008
rect 60359 -83999 60393 -83965
rect 61059 -83999 61093 -83965
rect 60359 -84091 60393 -84057
rect 61059 -84091 61093 -84057
rect 59103 -84242 59137 -84208
rect 57133 -84831 57167 -84797
rect 57251 -84844 57285 -84810
rect 59103 -84770 59137 -84736
rect 59545 -84245 59579 -84211
rect 59545 -84555 59579 -84521
rect 59861 -84245 59895 -84211
rect 60359 -84175 60393 -84141
rect 61059 -84175 61093 -84141
rect 59861 -84555 59895 -84521
rect 60359 -84259 60393 -84225
rect 61059 -84259 61093 -84225
rect 59560 -85042 59594 -85008
rect 59032 -85150 59066 -85116
rect 53988 -85444 54022 -85406
rect 54916 -85444 54950 -85406
rect 59874 -84828 59908 -84794
rect 60384 -84828 60418 -84794
rect 55526 -85636 55560 -85602
<< xpolycontact >>
rect 16566 -14662 16998 -13516
rect 34154 -14662 34586 -13516
rect 16566 -16034 16998 -14888
rect 34154 -16034 34586 -14888
rect 25868 -31560 27014 -31128
rect 25868 -32496 27014 -32064
rect 27110 -31560 28256 -31128
rect 27110 -32496 28256 -32064
rect 28352 -31560 29498 -31128
rect 28352 -32496 29498 -32064
rect 29594 -31560 30740 -31128
rect 29594 -32496 30740 -32064
rect 30836 -31560 31982 -31128
rect 30836 -32496 31982 -32064
rect 32078 -31560 33224 -31128
rect 32078 -32496 33224 -32064
rect 33320 -31560 34466 -31128
rect 33320 -32496 34466 -32064
rect 34562 -31560 35708 -31128
rect 34562 -32496 35708 -32064
rect 25866 -33158 27012 -32726
rect 25866 -34094 27012 -33662
rect 27108 -33158 28254 -32726
rect 27108 -34094 28254 -33662
rect 28350 -33158 29496 -32726
rect 28350 -34094 29496 -33662
rect 29592 -33158 30738 -32726
rect 29592 -34094 30738 -33662
rect 30834 -33158 31980 -32726
rect 30834 -34094 31980 -33662
rect 32076 -33158 33222 -32726
rect 32076 -34094 33222 -33662
rect 33318 -33158 34464 -32726
rect 33318 -34094 34464 -33662
rect 34560 -33158 35706 -32726
rect 34560 -34094 35706 -33662
rect 25866 -34756 27012 -34324
rect 25866 -35692 27012 -35260
rect 27108 -34756 28254 -34324
rect 27108 -35692 28254 -35260
rect 28350 -34756 29496 -34324
rect 28350 -35692 29496 -35260
rect 29592 -34756 30738 -34324
rect 29592 -35692 30738 -35260
rect 30834 -34756 31980 -34324
rect 30834 -35692 31980 -35260
rect 32076 -34756 33222 -34324
rect 32076 -35692 33222 -35260
rect 33318 -34756 34464 -34324
rect 33318 -35692 34464 -35260
rect 34560 -34756 35706 -34324
rect 34560 -35692 35706 -35260
rect 25866 -36358 27012 -35926
rect 25866 -37294 27012 -36862
rect 27108 -36358 28254 -35926
rect 27108 -37294 28254 -36862
rect 28350 -36358 29496 -35926
rect 28350 -37294 29496 -36862
rect 29592 -36358 30738 -35926
rect 29592 -37294 30738 -36862
rect 30834 -36358 31980 -35926
rect 30834 -37294 31980 -36862
rect 32076 -36358 33222 -35926
rect 32076 -37294 33222 -36862
rect 33318 -36358 34464 -35926
rect 33318 -37294 34464 -36862
rect 34560 -36358 35706 -35926
rect 34560 -37294 35706 -36862
rect 25866 -37958 27012 -37526
rect 25866 -38894 27012 -38462
rect 27108 -37958 28254 -37526
rect 27108 -38894 28254 -38462
rect 28350 -37958 29496 -37526
rect 28350 -38894 29496 -38462
rect 29592 -37958 30738 -37526
rect 29592 -38894 30738 -38462
rect 30834 -37958 31980 -37526
rect 30834 -38894 31980 -38462
rect 32076 -37958 33222 -37526
rect 32076 -38894 33222 -38462
rect 33318 -37958 34464 -37526
rect 33318 -38894 34464 -38462
rect 34560 -37958 35706 -37526
rect 34560 -38894 35706 -38462
rect 25868 -39560 27014 -39128
rect 25868 -40496 27014 -40064
rect 27110 -39560 28256 -39128
rect 27110 -40496 28256 -40064
rect 28352 -39560 29498 -39128
rect 28352 -40496 29498 -40064
rect 29594 -39560 30740 -39128
rect 29594 -40496 30740 -40064
rect 30836 -39560 31982 -39128
rect 30836 -40496 31982 -40064
rect 32078 -39560 33224 -39128
rect 32078 -40496 33224 -40064
rect 33320 -39560 34466 -39128
rect 33320 -40496 34466 -40064
rect 34562 -39560 35708 -39128
rect 34562 -40496 35708 -40064
rect 25866 -41158 27012 -40726
rect 25866 -42094 27012 -41662
rect 27108 -41158 28254 -40726
rect 27108 -42094 28254 -41662
rect 28350 -41158 29496 -40726
rect 28350 -42094 29496 -41662
rect 29592 -41158 30738 -40726
rect 29592 -42094 30738 -41662
rect 30834 -41158 31980 -40726
rect 30834 -42094 31980 -41662
rect 32076 -41158 33222 -40726
rect 32076 -42094 33222 -41662
rect 33318 -41158 34464 -40726
rect 33318 -42094 34464 -41662
rect 34560 -41158 35706 -40726
rect 34560 -42094 35706 -41662
rect 25866 -42756 27012 -42324
rect 25866 -43692 27012 -43260
rect 27108 -42756 28254 -42324
rect 27108 -43692 28254 -43260
rect 28350 -42756 29496 -42324
rect 28350 -43692 29496 -43260
rect 29592 -42756 30738 -42324
rect 29592 -43692 30738 -43260
rect 30834 -42756 31980 -42324
rect 30834 -43692 31980 -43260
rect 32076 -42756 33222 -42324
rect 32076 -43692 33222 -43260
rect 33318 -42756 34464 -42324
rect 33318 -43692 34464 -43260
rect 34560 -42756 35706 -42324
rect 34560 -43692 35706 -43260
rect 25866 -44358 27012 -43926
rect 25866 -45294 27012 -44862
rect 27108 -44358 28254 -43926
rect 27108 -45294 28254 -44862
rect 28350 -44358 29496 -43926
rect 28350 -45294 29496 -44862
rect 29592 -44358 30738 -43926
rect 29592 -45294 30738 -44862
rect 30834 -44358 31980 -43926
rect 30834 -45294 31980 -44862
rect 32076 -44358 33222 -43926
rect 32076 -45294 33222 -44862
rect 33318 -44358 34464 -43926
rect 33318 -45294 34464 -44862
rect 34560 -44358 35706 -43926
rect 34560 -45294 35706 -44862
rect 25866 -45956 27012 -45524
rect 25866 -46892 27012 -46460
rect 27108 -45956 28254 -45524
rect 27108 -46892 28254 -46460
rect 28350 -45956 29496 -45524
rect 28350 -46892 29496 -46460
rect 29592 -45956 30738 -45524
rect 29592 -46892 30738 -46460
rect 30834 -45956 31980 -45524
rect 30834 -46892 31980 -46460
rect 32076 -45956 33222 -45524
rect 32076 -46892 33222 -46460
rect 33318 -45956 34464 -45524
rect 33318 -46892 34464 -46460
rect 34560 -45956 35706 -45524
rect 34560 -46892 35706 -46460
rect 25866 -47550 27012 -47118
rect 25866 -48486 27012 -48054
rect 27108 -47550 28254 -47118
rect 27108 -48486 28254 -48054
rect 28350 -47550 29496 -47118
rect 28350 -48486 29496 -48054
rect 29592 -47550 30738 -47118
rect 29592 -48486 30738 -48054
rect 30834 -47550 31980 -47118
rect 30834 -48486 31980 -48054
rect 32076 -47550 33222 -47118
rect 32076 -48486 33222 -48054
rect 33318 -47550 34464 -47118
rect 33318 -48486 34464 -48054
rect 34560 -47550 35706 -47118
rect 34560 -48486 35706 -48054
rect 25866 -49148 27012 -48716
rect 25866 -50084 27012 -49652
rect 27108 -49148 28254 -48716
rect 27108 -50084 28254 -49652
rect 28350 -49148 29496 -48716
rect 28350 -50084 29496 -49652
rect 29592 -49148 30738 -48716
rect 29592 -50084 30738 -49652
rect 30834 -49148 31980 -48716
rect 30834 -50084 31980 -49652
rect 32076 -49148 33222 -48716
rect 32076 -50084 33222 -49652
rect 33318 -49148 34464 -48716
rect 33318 -50084 34464 -49652
rect 34560 -49148 35706 -48716
rect 34560 -50084 35706 -49652
rect 25866 -50750 27012 -50318
rect 25866 -51686 27012 -51254
rect 27108 -50750 28254 -50318
rect 27108 -51686 28254 -51254
rect 28350 -50750 29496 -50318
rect 28350 -51686 29496 -51254
rect 29592 -50750 30738 -50318
rect 29592 -51686 30738 -51254
rect 30834 -50750 31980 -50318
rect 30834 -51686 31980 -51254
rect 32076 -50750 33222 -50318
rect 32076 -51686 33222 -51254
rect 33318 -50750 34464 -50318
rect 33318 -51686 34464 -51254
rect 34560 -50750 35706 -50318
rect 34560 -51686 35706 -51254
rect 25866 -52348 27012 -51916
rect 25866 -53284 27012 -52852
rect 27108 -52348 28254 -51916
rect 27108 -53284 28254 -52852
rect 28350 -52348 29496 -51916
rect 28350 -53284 29496 -52852
rect 29592 -52348 30738 -51916
rect 29592 -53284 30738 -52852
rect 30834 -52348 31980 -51916
rect 30834 -53284 31980 -52852
rect 32076 -52348 33222 -51916
rect 32076 -53284 33222 -52852
rect 33318 -52348 34464 -51916
rect 33318 -53284 34464 -52852
rect 34560 -52348 35706 -51916
rect 34560 -53284 35706 -52852
rect 25868 -53950 27014 -53518
rect 25868 -54886 27014 -54454
rect 27110 -53950 28256 -53518
rect 27110 -54886 28256 -54454
rect 28352 -53950 29498 -53518
rect 28352 -54886 29498 -54454
rect 29594 -53950 30740 -53518
rect 29594 -54886 30740 -54454
rect 30836 -53950 31982 -53518
rect 30836 -54886 31982 -54454
rect 32078 -53950 33224 -53518
rect 32078 -54886 33224 -54454
rect 33320 -53950 34466 -53518
rect 33320 -54886 34466 -54454
rect 34562 -53950 35708 -53518
rect 34562 -54886 35708 -54454
rect 25866 -55548 27012 -55116
rect 25866 -56484 27012 -56052
rect 27108 -55548 28254 -55116
rect 27108 -56484 28254 -56052
rect 28350 -55548 29496 -55116
rect 28350 -56484 29496 -56052
rect 29592 -55548 30738 -55116
rect 29592 -56484 30738 -56052
rect 30834 -55548 31980 -55116
rect 30834 -56484 31980 -56052
rect 32076 -55548 33222 -55116
rect 32076 -56484 33222 -56052
rect 33318 -55548 34464 -55116
rect 33318 -56484 34464 -56052
rect 34560 -55548 35706 -55116
rect 34560 -56484 35706 -56052
rect 25866 -57148 27012 -56716
rect 25866 -58084 27012 -57652
rect 27108 -57148 28254 -56716
rect 27108 -58084 28254 -57652
rect 28350 -57148 29496 -56716
rect 28350 -58084 29496 -57652
rect 29592 -57148 30738 -56716
rect 29592 -58084 30738 -57652
rect 30834 -57148 31980 -56716
rect 30834 -58084 31980 -57652
rect 32076 -57148 33222 -56716
rect 32076 -58084 33222 -57652
rect 33318 -57148 34464 -56716
rect 33318 -58084 34464 -57652
rect 34560 -57148 35706 -56716
rect 34560 -58084 35706 -57652
<< xpolyres >>
rect 16998 -14662 34154 -13516
rect 16998 -16034 34154 -14888
rect 25868 -32064 27014 -31560
rect 27110 -32064 28256 -31560
rect 28352 -32064 29498 -31560
rect 29594 -32064 30740 -31560
rect 30836 -32064 31982 -31560
rect 32078 -32064 33224 -31560
rect 33320 -32064 34466 -31560
rect 34562 -32064 35708 -31560
rect 25866 -33662 27012 -33158
rect 27108 -33662 28254 -33158
rect 28350 -33662 29496 -33158
rect 29592 -33662 30738 -33158
rect 30834 -33662 31980 -33158
rect 32076 -33662 33222 -33158
rect 33318 -33662 34464 -33158
rect 34560 -33662 35706 -33158
rect 25866 -35260 27012 -34756
rect 27108 -35260 28254 -34756
rect 28350 -35260 29496 -34756
rect 29592 -35260 30738 -34756
rect 30834 -35260 31980 -34756
rect 32076 -35260 33222 -34756
rect 33318 -35260 34464 -34756
rect 34560 -35260 35706 -34756
rect 25866 -36862 27012 -36358
rect 27108 -36862 28254 -36358
rect 28350 -36862 29496 -36358
rect 29592 -36862 30738 -36358
rect 30834 -36862 31980 -36358
rect 32076 -36862 33222 -36358
rect 33318 -36862 34464 -36358
rect 34560 -36862 35706 -36358
rect 25866 -38462 27012 -37958
rect 27108 -38462 28254 -37958
rect 28350 -38462 29496 -37958
rect 29592 -38462 30738 -37958
rect 30834 -38462 31980 -37958
rect 32076 -38462 33222 -37958
rect 33318 -38462 34464 -37958
rect 34560 -38462 35706 -37958
rect 25868 -40064 27014 -39560
rect 27110 -40064 28256 -39560
rect 28352 -40064 29498 -39560
rect 29594 -40064 30740 -39560
rect 30836 -40064 31982 -39560
rect 32078 -40064 33224 -39560
rect 33320 -40064 34466 -39560
rect 34562 -40064 35708 -39560
rect 25866 -41662 27012 -41158
rect 27108 -41662 28254 -41158
rect 28350 -41662 29496 -41158
rect 29592 -41662 30738 -41158
rect 30834 -41662 31980 -41158
rect 32076 -41662 33222 -41158
rect 33318 -41662 34464 -41158
rect 34560 -41662 35706 -41158
rect 25866 -43260 27012 -42756
rect 27108 -43260 28254 -42756
rect 28350 -43260 29496 -42756
rect 29592 -43260 30738 -42756
rect 30834 -43260 31980 -42756
rect 32076 -43260 33222 -42756
rect 33318 -43260 34464 -42756
rect 34560 -43260 35706 -42756
rect 25866 -44862 27012 -44358
rect 27108 -44862 28254 -44358
rect 28350 -44862 29496 -44358
rect 29592 -44862 30738 -44358
rect 30834 -44862 31980 -44358
rect 32076 -44862 33222 -44358
rect 33318 -44862 34464 -44358
rect 34560 -44862 35706 -44358
rect 25866 -46460 27012 -45956
rect 27108 -46460 28254 -45956
rect 28350 -46460 29496 -45956
rect 29592 -46460 30738 -45956
rect 30834 -46460 31980 -45956
rect 32076 -46460 33222 -45956
rect 33318 -46460 34464 -45956
rect 34560 -46460 35706 -45956
rect 25866 -48054 27012 -47550
rect 27108 -48054 28254 -47550
rect 28350 -48054 29496 -47550
rect 29592 -48054 30738 -47550
rect 30834 -48054 31980 -47550
rect 32076 -48054 33222 -47550
rect 33318 -48054 34464 -47550
rect 34560 -48054 35706 -47550
rect 25866 -49652 27012 -49148
rect 27108 -49652 28254 -49148
rect 28350 -49652 29496 -49148
rect 29592 -49652 30738 -49148
rect 30834 -49652 31980 -49148
rect 32076 -49652 33222 -49148
rect 33318 -49652 34464 -49148
rect 34560 -49652 35706 -49148
rect 25866 -51254 27012 -50750
rect 27108 -51254 28254 -50750
rect 28350 -51254 29496 -50750
rect 29592 -51254 30738 -50750
rect 30834 -51254 31980 -50750
rect 32076 -51254 33222 -50750
rect 33318 -51254 34464 -50750
rect 34560 -51254 35706 -50750
rect 25866 -52852 27012 -52348
rect 27108 -52852 28254 -52348
rect 28350 -52852 29496 -52348
rect 29592 -52852 30738 -52348
rect 30834 -52852 31980 -52348
rect 32076 -52852 33222 -52348
rect 33318 -52852 34464 -52348
rect 34560 -52852 35706 -52348
rect 25868 -54454 27014 -53950
rect 27110 -54454 28256 -53950
rect 28352 -54454 29498 -53950
rect 29594 -54454 30740 -53950
rect 30836 -54454 31982 -53950
rect 32078 -54454 33224 -53950
rect 33320 -54454 34466 -53950
rect 34562 -54454 35708 -53950
rect 25866 -56052 27012 -55548
rect 27108 -56052 28254 -55548
rect 28350 -56052 29496 -55548
rect 29592 -56052 30738 -55548
rect 30834 -56052 31980 -55548
rect 32076 -56052 33222 -55548
rect 33318 -56052 34464 -55548
rect 34560 -56052 35706 -55548
rect 25866 -57652 27012 -57148
rect 27108 -57652 28254 -57148
rect 28350 -57652 29496 -57148
rect 29592 -57652 30738 -57148
rect 30834 -57652 31980 -57148
rect 32076 -57652 33222 -57148
rect 33318 -57652 34464 -57148
rect 34560 -57652 35706 -57148
<< locali >>
rect 53896 -1592 53992 -1558
rect 54966 -1592 55062 -1558
rect 53896 -1654 53930 -1592
rect 55028 -1654 55062 -1592
rect 54075 -1706 54091 -1672
rect 54867 -1706 54883 -1672
rect 53998 -1734 54032 -1718
rect 53998 -1788 54032 -1772
rect 54926 -1734 54960 -1718
rect 54926 -1788 54960 -1772
rect 54075 -1834 54091 -1800
rect 54867 -1834 54883 -1800
rect 53896 -1914 53930 -1852
rect 55028 -1914 55062 -1852
rect 55960 -1908 56040 -1898
rect 53896 -1948 53992 -1914
rect 54966 -1948 55062 -1914
rect 53350 -2038 53790 -2004
rect 53350 -2100 53384 -2038
rect 53510 -2140 53526 -2106
rect 53614 -2140 53630 -2106
rect 53464 -2190 53498 -2174
rect 53464 -2982 53498 -2966
rect 53642 -2190 53676 -2174
rect 53642 -2982 53676 -2966
rect 53756 -2664 53790 -2038
rect 53896 -2010 53930 -1948
rect 55028 -2010 55062 -1948
rect 55710 -1954 56040 -1908
rect 54075 -2062 54091 -2028
rect 54867 -2062 54883 -2028
rect 53998 -2090 54032 -2074
rect 53998 -2144 54032 -2128
rect 54926 -2090 54960 -2074
rect 54926 -2144 54960 -2128
rect 54075 -2190 54091 -2156
rect 54867 -2190 54883 -2156
rect 53896 -2270 53930 -2208
rect 55706 -1988 55802 -1954
rect 56050 -1988 56146 -1954
rect 55706 -2050 55740 -1988
rect 55028 -2270 55062 -2208
rect 53896 -2304 53992 -2270
rect 54966 -2304 55062 -2270
rect 55176 -2100 55272 -2066
rect 55430 -2100 55526 -2066
rect 55176 -2162 55210 -2100
rect 55492 -2162 55526 -2100
rect 55318 -2202 55334 -2168
rect 55368 -2202 55384 -2168
rect 55290 -2252 55324 -2236
rect 55290 -2444 55324 -2428
rect 55378 -2252 55412 -2236
rect 55378 -2444 55412 -2428
rect 55176 -2518 55210 -2456
rect 55492 -2518 55526 -2456
rect 54870 -2552 55272 -2518
rect 55430 -2552 55706 -2518
rect 54870 -2558 55706 -2552
rect 54870 -2664 54904 -2558
rect 53756 -2698 53852 -2664
rect 54808 -2698 54904 -2664
rect 53756 -2760 53790 -2698
rect 54870 -2760 54904 -2698
rect 55126 -2708 55142 -2674
rect 55494 -2708 55510 -2674
rect 53926 -2812 53942 -2778
rect 54718 -2812 54734 -2778
rect 53858 -2840 53892 -2824
rect 53858 -2944 53892 -2928
rect 54768 -2840 54802 -2824
rect 54768 -2944 54802 -2928
rect 53926 -2990 53942 -2956
rect 54718 -2990 54734 -2956
rect 53510 -3050 53526 -3016
rect 53614 -3050 53630 -3016
rect 53756 -3070 53790 -3008
rect 55046 -2760 55080 -2744
rect 55046 -2810 55080 -2794
rect 55556 -2760 55590 -2744
rect 55556 -2810 55590 -2794
rect 55126 -2880 55142 -2846
rect 55494 -2880 55510 -2846
rect 54870 -3038 54904 -3008
rect 55700 -3006 55706 -2558
rect 56112 -2050 56146 -1988
rect 58930 -1967 59026 -1933
rect 59600 -1967 59696 -1933
rect 58930 -2010 58964 -1967
rect 58926 -2020 58966 -2010
rect 55866 -2090 55882 -2056
rect 55970 -2090 55986 -2056
rect 55820 -2140 55854 -2124
rect 55820 -2932 55854 -2916
rect 55998 -2140 56032 -2124
rect 55998 -2932 56032 -2916
rect 55866 -3000 55882 -2966
rect 55970 -3000 55986 -2966
rect 55700 -3038 55740 -3006
rect 57096 -2079 57125 -2045
rect 57159 -2079 57217 -2045
rect 57251 -2079 57309 -2045
rect 57343 -2079 57372 -2045
rect 57129 -2129 57165 -2113
rect 57129 -2163 57131 -2129
rect 57129 -2197 57165 -2163
rect 57129 -2231 57131 -2197
rect 57201 -2129 57267 -2079
rect 57201 -2163 57217 -2129
rect 57251 -2163 57267 -2129
rect 57201 -2197 57267 -2163
rect 57201 -2231 57217 -2197
rect 57251 -2231 57267 -2197
rect 57301 -2129 57355 -2113
rect 57301 -2163 57303 -2129
rect 57337 -2163 57355 -2129
rect 57301 -2210 57355 -2163
rect 57129 -2265 57165 -2231
rect 57301 -2244 57303 -2210
rect 57337 -2244 57355 -2210
rect 57129 -2299 57264 -2265
rect 57301 -2294 57355 -2244
rect 57230 -2328 57264 -2299
rect 57117 -2344 57185 -2335
rect 57117 -2394 57118 -2344
rect 57178 -2394 57185 -2344
rect 57117 -2409 57185 -2394
rect 57230 -2344 57285 -2328
rect 57230 -2378 57251 -2344
rect 57230 -2394 57285 -2378
rect 57319 -2340 57355 -2294
rect 59662 -2029 59696 -1967
rect 59109 -2081 59125 -2047
rect 59501 -2081 59517 -2047
rect 59560 -2101 59594 -2085
rect 59560 -2151 59594 -2135
rect 59109 -2189 59125 -2155
rect 59501 -2189 59517 -2155
rect 59032 -2209 59066 -2193
rect 59032 -2259 59066 -2243
rect 59109 -2297 59125 -2263
rect 59501 -2297 59517 -2263
rect 58926 -2340 58966 -2320
rect 57319 -2380 57326 -2340
rect 58930 -2376 58964 -2340
rect 57230 -2445 57264 -2394
rect 57131 -2479 57264 -2445
rect 57319 -2454 57355 -2380
rect 57131 -2500 57165 -2479
rect 56316 -2518 56412 -2504
rect 54830 -3048 55830 -3038
rect 54830 -3070 55030 -3048
rect 53756 -3104 53852 -3070
rect 54808 -3104 55030 -3070
rect 53510 -3158 53526 -3124
rect 53614 -3158 53630 -3124
rect 53756 -3166 53790 -3104
rect 54830 -3128 55030 -3104
rect 55110 -3068 55740 -3048
rect 55810 -3068 55830 -3048
rect 56112 -3068 56146 -3006
rect 55110 -3108 55160 -3068
rect 55600 -3108 55740 -3068
rect 56050 -3102 56146 -3068
rect 55110 -3128 55740 -3108
rect 55810 -3128 55830 -3102
rect 54830 -3138 55830 -3128
rect 53464 -3208 53498 -3192
rect 53464 -4000 53498 -3984
rect 53642 -3208 53676 -3192
rect 53642 -4000 53676 -3984
rect 54870 -3166 54904 -3138
rect 53926 -3218 53942 -3184
rect 54718 -3218 54734 -3184
rect 53858 -3246 53892 -3230
rect 53858 -3350 53892 -3334
rect 54768 -3246 54802 -3230
rect 54768 -3350 54802 -3334
rect 53926 -3396 53942 -3362
rect 54718 -3396 54734 -3362
rect 53756 -3476 53790 -3414
rect 55700 -3164 55740 -3138
rect 55126 -3330 55142 -3296
rect 55494 -3330 55510 -3296
rect 54870 -3476 54904 -3414
rect 55046 -3382 55080 -3366
rect 55046 -3432 55080 -3416
rect 55556 -3382 55590 -3366
rect 55556 -3432 55590 -3416
rect 53756 -3510 53852 -3476
rect 54808 -3510 54904 -3476
rect 55126 -3502 55142 -3468
rect 55494 -3502 55510 -3468
rect 53510 -4068 53526 -4034
rect 53614 -4068 53630 -4034
rect 53350 -4136 53384 -4074
rect 53756 -4136 53790 -3510
rect 54870 -3618 54904 -3510
rect 55700 -3618 55706 -3164
rect 54870 -3624 55706 -3618
rect 54870 -3658 55262 -3624
rect 55420 -3658 55706 -3624
rect 55166 -3720 55200 -3658
rect 53350 -4170 53446 -4136
rect 53694 -4170 53790 -4136
rect 53886 -3908 53982 -3874
rect 54956 -3908 55052 -3874
rect 53886 -3970 53920 -3908
rect 55018 -3970 55052 -3908
rect 54065 -4022 54081 -3988
rect 54857 -4022 54873 -3988
rect 53988 -4050 54022 -4034
rect 53988 -4104 54022 -4088
rect 54916 -4050 54950 -4034
rect 54916 -4104 54950 -4088
rect 54065 -4150 54081 -4116
rect 54857 -4150 54873 -4116
rect 53886 -4230 53920 -4168
rect 55482 -3720 55516 -3658
rect 55280 -3748 55314 -3732
rect 55280 -3940 55314 -3924
rect 55368 -3748 55402 -3732
rect 55368 -3940 55402 -3924
rect 55308 -4008 55324 -3974
rect 55358 -4008 55374 -3974
rect 55166 -4076 55200 -4014
rect 55482 -4076 55516 -4014
rect 55166 -4110 55262 -4076
rect 55420 -4110 55516 -4076
rect 55018 -4230 55052 -4168
rect 56112 -3164 56146 -3102
rect 56350 -2538 56412 -2518
rect 56610 -2538 56706 -2504
rect 56672 -2600 56706 -2538
rect 57303 -2483 57355 -2454
rect 57131 -2555 57165 -2534
rect 57201 -2547 57217 -2513
rect 57251 -2547 57267 -2513
rect 57201 -2589 57267 -2547
rect 57337 -2517 57355 -2483
rect 57303 -2555 57355 -2517
rect 58930 -2410 59026 -2376
rect 59214 -2377 59310 -2376
rect 59662 -2377 59696 -2320
rect 59772 -2294 59866 -2260
rect 60426 -2294 60520 -2260
rect 59772 -2350 59806 -2294
rect 59214 -2410 59696 -2377
rect 58930 -2411 59696 -2410
rect 58930 -2472 58964 -2411
rect 59276 -2472 59310 -2411
rect 59087 -2512 59103 -2478
rect 59137 -2512 59153 -2478
rect 56476 -2640 56492 -2606
rect 56530 -2640 56546 -2606
rect 55866 -3204 55882 -3170
rect 55970 -3204 55986 -3170
rect 55820 -3254 55854 -3238
rect 55820 -4046 55854 -4030
rect 55998 -3254 56032 -3238
rect 55998 -4046 56032 -4030
rect 55866 -4114 55882 -4080
rect 55970 -4114 55986 -4080
rect 55706 -4182 55740 -4120
rect 56430 -2699 56464 -2683
rect 56430 -3491 56464 -3475
rect 56558 -2699 56592 -2683
rect 56558 -3491 56592 -3475
rect 56476 -3568 56492 -3534
rect 56530 -3568 56546 -3534
rect 56316 -3636 56350 -3574
rect 57096 -2623 57125 -2589
rect 57159 -2623 57217 -2589
rect 57251 -2623 57309 -2589
rect 57343 -2623 57372 -2589
rect 59044 -2571 59078 -2555
rect 59044 -2963 59078 -2947
rect 59162 -2571 59196 -2555
rect 59162 -2963 59196 -2947
rect 59087 -3040 59103 -3006
rect 59137 -3040 59153 -3006
rect 60486 -2356 60520 -2294
rect 59942 -2408 59958 -2374
rect 60334 -2408 60350 -2374
rect 59874 -2428 59908 -2412
rect 59874 -2478 59908 -2462
rect 60384 -2428 60418 -2412
rect 60384 -2478 60418 -2462
rect 59942 -2516 59958 -2482
rect 60334 -2516 60350 -2482
rect 59772 -2596 59806 -2540
rect 60486 -2596 60520 -2534
rect 59388 -2630 59476 -2596
rect 59656 -2630 59800 -2596
rect 59958 -2630 60520 -2596
rect 59388 -2690 59422 -2630
rect 59276 -3106 59310 -3046
rect 59530 -2732 59546 -2698
rect 59580 -2732 59596 -2698
rect 59502 -2782 59536 -2766
rect 59502 -2974 59536 -2958
rect 59590 -2782 59624 -2766
rect 59590 -2974 59624 -2958
rect 59530 -3042 59546 -3008
rect 59580 -3042 59596 -3008
rect 58966 -3142 59310 -3106
rect 59388 -3109 59422 -3050
rect 59704 -3109 59738 -2630
rect 60020 -2692 60054 -2630
rect 59846 -2732 59862 -2698
rect 59896 -2732 59912 -2698
rect 59818 -2782 59852 -2766
rect 59818 -2974 59852 -2958
rect 59906 -2782 59940 -2766
rect 59906 -2974 59940 -2958
rect 59846 -3042 59862 -3008
rect 59896 -3042 59912 -3008
rect 61186 -2800 61286 -2790
rect 61186 -2880 61196 -2800
rect 61186 -2890 61286 -2880
rect 60020 -3109 60054 -3048
rect 56672 -3636 56706 -3574
rect 57096 -3599 57125 -3565
rect 57159 -3599 57217 -3565
rect 57251 -3599 57309 -3565
rect 57343 -3599 57372 -3565
rect 56316 -3670 56412 -3636
rect 56610 -3670 56706 -3636
rect 57131 -3654 57165 -3633
rect 57201 -3641 57267 -3599
rect 57201 -3675 57217 -3641
rect 57251 -3675 57267 -3641
rect 57303 -3671 57355 -3633
rect 57131 -3709 57165 -3688
rect 57337 -3705 57355 -3671
rect 59276 -3202 59310 -3142
rect 59387 -3144 60054 -3109
rect 60127 -2954 60161 -2928
rect 60127 -2957 60253 -2954
rect 60161 -2973 60253 -2957
rect 60161 -2991 60203 -2973
rect 60127 -3007 60203 -2991
rect 60237 -3007 60253 -2973
rect 60359 -2960 60409 -2949
rect 60671 -2954 60705 -2928
rect 60359 -2965 60366 -2960
rect 60359 -3000 60366 -2999
rect 60406 -3000 60409 -2960
rect 60127 -3049 60161 -3007
rect 60127 -3141 60161 -3083
rect 60195 -3057 60325 -3041
rect 60195 -3091 60211 -3057
rect 60245 -3091 60325 -3057
rect 60195 -3107 60325 -3091
rect 59387 -3200 59421 -3144
rect 59087 -3242 59103 -3208
rect 59137 -3242 59153 -3208
rect 59044 -3301 59078 -3285
rect 57131 -3743 57264 -3709
rect 57303 -3734 57355 -3705
rect 57117 -3794 57185 -3779
rect 57117 -3844 57118 -3794
rect 57168 -3844 57185 -3794
rect 57117 -3853 57185 -3844
rect 57230 -3794 57264 -3743
rect 57319 -3770 57355 -3734
rect 57230 -3810 57285 -3794
rect 57230 -3844 57251 -3810
rect 57230 -3860 57285 -3844
rect 57319 -3810 57326 -3770
rect 59044 -3693 59078 -3677
rect 59162 -3301 59196 -3285
rect 59162 -3693 59196 -3677
rect 59087 -3770 59103 -3736
rect 59137 -3770 59153 -3736
rect 57230 -3889 57264 -3860
rect 57129 -3923 57264 -3889
rect 57319 -3894 57355 -3810
rect 57129 -3957 57165 -3923
rect 57301 -3944 57355 -3894
rect 58930 -3838 58964 -3776
rect 59529 -3245 59545 -3211
rect 59579 -3245 59595 -3211
rect 59501 -3295 59535 -3279
rect 59501 -3487 59535 -3471
rect 59589 -3295 59623 -3279
rect 59589 -3487 59623 -3471
rect 59529 -3555 59545 -3521
rect 59579 -3555 59595 -3521
rect 59387 -3623 59421 -3570
rect 59703 -3623 59737 -3144
rect 60019 -3205 60053 -3144
rect 59845 -3245 59861 -3211
rect 59895 -3245 59911 -3211
rect 59817 -3295 59851 -3279
rect 59817 -3487 59851 -3471
rect 59905 -3295 59939 -3279
rect 59905 -3487 59939 -3471
rect 59845 -3555 59861 -3521
rect 59895 -3555 59911 -3521
rect 60161 -3175 60203 -3141
rect 60237 -3175 60253 -3141
rect 60127 -3233 60161 -3175
rect 60289 -3209 60325 -3107
rect 60127 -3309 60161 -3267
rect 60195 -3225 60325 -3209
rect 60195 -3259 60211 -3225
rect 60245 -3259 60325 -3225
rect 60195 -3275 60325 -3259
rect 60359 -3050 60409 -3000
rect 60443 -2957 60705 -2954
rect 60443 -2973 60671 -2957
rect 60443 -3007 60459 -2973
rect 60493 -3007 60527 -2973
rect 60561 -3007 60595 -2973
rect 60629 -2991 60671 -2973
rect 60629 -3007 60705 -2991
rect 60359 -3057 60366 -3050
rect 60406 -3090 60409 -3050
rect 60393 -3091 60409 -3090
rect 60359 -3140 60409 -3091
rect 60359 -3141 60366 -3140
rect 60359 -3180 60366 -3175
rect 60406 -3180 60409 -3140
rect 60359 -3220 60409 -3180
rect 60359 -3225 60366 -3220
rect 60359 -3260 60366 -3259
rect 60406 -3260 60409 -3220
rect 60359 -3275 60409 -3260
rect 60443 -3057 60637 -3041
rect 60443 -3091 60459 -3057
rect 60493 -3091 60527 -3057
rect 60561 -3091 60595 -3057
rect 60629 -3091 60637 -3057
rect 60443 -3107 60637 -3091
rect 60671 -3049 60705 -3007
rect 60443 -3209 60477 -3107
rect 60671 -3141 60705 -3083
rect 60511 -3175 60527 -3141
rect 60561 -3175 60595 -3141
rect 60629 -3175 60671 -3141
rect 60443 -3225 60637 -3209
rect 60443 -3259 60459 -3225
rect 60493 -3259 60527 -3225
rect 60561 -3259 60595 -3225
rect 60629 -3259 60637 -3225
rect 60443 -3275 60637 -3259
rect 60671 -3233 60705 -3175
rect 60289 -3309 60325 -3275
rect 60443 -3309 60481 -3275
rect 60671 -3309 60705 -3267
rect 60127 -3325 60204 -3309
rect 60161 -3343 60204 -3325
rect 60238 -3343 60254 -3309
rect 60161 -3359 60254 -3343
rect 60289 -3325 60481 -3309
rect 60289 -3359 60297 -3325
rect 60331 -3359 60369 -3325
rect 60405 -3359 60449 -3325
rect 60579 -3343 60595 -3309
rect 60629 -3325 60705 -3309
rect 60629 -3343 60671 -3325
rect 60579 -3351 60671 -3343
rect 60127 -3388 60161 -3359
rect 60289 -3362 60481 -3359
rect 60671 -3388 60705 -3359
rect 60747 -2954 60781 -2928
rect 60747 -2957 61009 -2954
rect 60781 -2973 61009 -2957
rect 60781 -2991 60823 -2973
rect 60747 -3007 60823 -2991
rect 60857 -3007 60891 -2973
rect 60925 -3007 60959 -2973
rect 60993 -3007 61009 -2973
rect 61043 -2960 61093 -2949
rect 61291 -2954 61325 -2928
rect 61043 -3000 61046 -2960
rect 61086 -2965 61093 -2960
rect 61086 -3000 61093 -2999
rect 60747 -3049 60781 -3007
rect 60747 -3141 60781 -3083
rect 60815 -3057 61009 -3041
rect 60815 -3091 60823 -3057
rect 60857 -3091 60891 -3057
rect 60925 -3091 60959 -3057
rect 60993 -3091 61009 -3057
rect 60815 -3107 61009 -3091
rect 60781 -3175 60823 -3141
rect 60857 -3175 60891 -3141
rect 60925 -3175 60941 -3141
rect 60747 -3233 60781 -3175
rect 60975 -3209 61009 -3107
rect 60747 -3309 60781 -3267
rect 60815 -3225 61009 -3209
rect 60815 -3259 60823 -3225
rect 60857 -3259 60891 -3225
rect 60925 -3259 60959 -3225
rect 60993 -3259 61009 -3225
rect 60815 -3275 61009 -3259
rect 61043 -3050 61093 -3000
rect 61199 -2957 61325 -2954
rect 61199 -2973 61291 -2957
rect 61199 -3007 61215 -2973
rect 61249 -2991 61291 -2973
rect 61249 -3007 61325 -2991
rect 61043 -3090 61046 -3050
rect 61086 -3057 61093 -3050
rect 61043 -3091 61059 -3090
rect 61043 -3140 61093 -3091
rect 61043 -3180 61046 -3140
rect 61086 -3141 61093 -3140
rect 61086 -3180 61093 -3175
rect 61043 -3220 61093 -3180
rect 61043 -3260 61046 -3220
rect 61086 -3225 61093 -3220
rect 61086 -3260 61093 -3259
rect 61043 -3275 61093 -3260
rect 61127 -3057 61257 -3041
rect 61127 -3091 61207 -3057
rect 61241 -3091 61257 -3057
rect 61127 -3107 61257 -3091
rect 61291 -3049 61325 -3007
rect 61127 -3209 61163 -3107
rect 61291 -3141 61325 -3083
rect 61199 -3175 61215 -3141
rect 61249 -3175 61291 -3141
rect 61127 -3225 61257 -3209
rect 61127 -3259 61207 -3225
rect 61241 -3259 61257 -3225
rect 61127 -3275 61257 -3259
rect 61291 -3233 61325 -3175
rect 60971 -3309 61009 -3275
rect 61127 -3309 61163 -3275
rect 61291 -3309 61325 -3267
rect 60747 -3325 60823 -3309
rect 60781 -3343 60823 -3325
rect 60857 -3343 60873 -3309
rect 60781 -3351 60873 -3343
rect 60971 -3324 61163 -3309
rect 60971 -3325 61129 -3324
rect 60747 -3388 60781 -3359
rect 60971 -3359 60980 -3325
rect 61015 -3359 61053 -3325
rect 61088 -3358 61129 -3325
rect 61198 -3343 61214 -3309
rect 61248 -3325 61325 -3309
rect 61248 -3343 61291 -3325
rect 61088 -3359 61163 -3358
rect 61198 -3359 61291 -3343
rect 60971 -3362 61163 -3359
rect 61291 -3388 61325 -3359
rect 60466 -3460 60546 -3440
rect 60466 -3500 60486 -3460
rect 60526 -3500 60546 -3460
rect 60466 -3520 60546 -3500
rect 60606 -3460 60686 -3440
rect 60606 -3500 60626 -3460
rect 60666 -3500 60686 -3460
rect 60606 -3520 60686 -3500
rect 60746 -3460 60826 -3440
rect 60746 -3500 60766 -3460
rect 60806 -3500 60826 -3460
rect 60746 -3520 60826 -3500
rect 60886 -3460 60966 -3440
rect 60886 -3500 60906 -3460
rect 60946 -3500 60966 -3460
rect 60886 -3520 60966 -3500
rect 60019 -3623 60053 -3561
rect 59387 -3657 59476 -3623
rect 59646 -3657 59799 -3623
rect 59957 -3626 60053 -3623
rect 59957 -3657 60520 -3626
rect 59772 -3660 60520 -3657
rect 59772 -3720 59806 -3660
rect 59276 -3838 59310 -3776
rect 58930 -3872 59026 -3838
rect 59214 -3840 59310 -3838
rect 59214 -3872 59696 -3840
rect 58930 -3874 59696 -3872
rect 58930 -3910 58964 -3874
rect 57129 -3991 57131 -3957
rect 57129 -4025 57165 -3991
rect 57129 -4059 57131 -4025
rect 57129 -4075 57165 -4059
rect 57201 -3991 57217 -3957
rect 57251 -3991 57267 -3957
rect 57201 -4025 57267 -3991
rect 57201 -4059 57217 -4025
rect 57251 -4059 57267 -4025
rect 57201 -4109 57267 -4059
rect 57301 -3978 57303 -3944
rect 57337 -3978 57355 -3944
rect 57301 -4025 57355 -3978
rect 57301 -4059 57303 -4025
rect 57337 -4059 57355 -4025
rect 57301 -4075 57355 -4059
rect 59662 -3930 59696 -3874
rect 60486 -3722 60520 -3660
rect 59942 -3774 59958 -3740
rect 60334 -3774 60350 -3740
rect 59874 -3794 59908 -3778
rect 59874 -3844 59908 -3828
rect 60384 -3794 60418 -3778
rect 60384 -3844 60418 -3828
rect 59942 -3882 59958 -3848
rect 60334 -3882 60350 -3848
rect 56112 -4182 56146 -4120
rect 57096 -4143 57125 -4109
rect 57159 -4143 57217 -4109
rect 57251 -4143 57309 -4109
rect 57343 -4143 57372 -4109
rect 55706 -4216 55802 -4182
rect 56050 -4216 56146 -4182
rect 53886 -4264 53982 -4230
rect 54956 -4264 55052 -4230
rect 53886 -4326 53920 -4264
rect 55018 -4326 55052 -4264
rect 55720 -4258 56090 -4216
rect 55720 -4268 56020 -4258
rect 54065 -4378 54081 -4344
rect 54857 -4378 54873 -4344
rect 53988 -4406 54022 -4390
rect 53988 -4460 54022 -4444
rect 54916 -4406 54950 -4390
rect 54916 -4460 54950 -4444
rect 54065 -4506 54081 -4472
rect 54857 -4506 54873 -4472
rect 53886 -4586 53920 -4524
rect 56010 -4408 56020 -4268
rect 56080 -4408 56090 -4258
rect 59109 -3988 59125 -3954
rect 59501 -3988 59517 -3954
rect 59560 -4008 59594 -3992
rect 59560 -4058 59594 -4042
rect 59109 -4096 59125 -4062
rect 59501 -4096 59517 -4062
rect 59032 -4116 59066 -4100
rect 59032 -4166 59066 -4150
rect 59109 -4204 59125 -4170
rect 59501 -4204 59517 -4170
rect 56010 -4418 56090 -4408
rect 59772 -3962 59806 -3900
rect 60486 -3962 60520 -3900
rect 59772 -3996 59866 -3962
rect 60426 -3996 60520 -3962
rect 59662 -4284 59696 -4230
rect 58966 -4300 59026 -4284
rect 58930 -4318 59026 -4300
rect 59600 -4318 59696 -4284
rect 55018 -4586 55052 -4524
rect 53886 -4620 53982 -4586
rect 54956 -4620 55052 -4586
rect 55176 -4478 55272 -4444
rect 55566 -4478 55662 -4444
rect 55176 -4540 55210 -4478
rect 55628 -4540 55662 -4478
rect 55284 -4592 55300 -4558
rect 55476 -4592 55492 -4558
rect 55526 -4602 55560 -4586
rect 55284 -4680 55300 -4646
rect 55476 -4680 55492 -4646
rect 55526 -4652 55560 -4636
rect 55176 -4760 55210 -4698
rect 55628 -4760 55662 -4698
rect 55176 -4794 55272 -4760
rect 55566 -4794 55662 -4760
rect 53896 -6992 53992 -6958
rect 54966 -6992 55062 -6958
rect 53896 -7054 53930 -6992
rect 55028 -7054 55062 -6992
rect 54075 -7106 54091 -7072
rect 54867 -7106 54883 -7072
rect 53998 -7134 54032 -7118
rect 53998 -7188 54032 -7172
rect 54926 -7134 54960 -7118
rect 54926 -7188 54960 -7172
rect 54075 -7234 54091 -7200
rect 54867 -7234 54883 -7200
rect 53896 -7314 53930 -7252
rect 55028 -7314 55062 -7252
rect 55960 -7308 56040 -7298
rect 53896 -7348 53992 -7314
rect 54966 -7348 55062 -7314
rect 53350 -7438 53790 -7404
rect 53350 -7500 53384 -7438
rect 53510 -7540 53526 -7506
rect 53614 -7540 53630 -7506
rect 20732 -7707 20828 -7673
rect 21156 -7707 21314 -7673
rect 21642 -7707 21800 -7673
rect 22128 -7707 22224 -7673
rect 20732 -7769 20766 -7707
rect 21218 -7769 21252 -7707
rect 20892 -7809 20908 -7775
rect 21076 -7809 21092 -7775
rect 20846 -7868 20880 -7852
rect 20846 -11660 20880 -11644
rect 21104 -7868 21138 -7852
rect 21704 -7769 21738 -7707
rect 21378 -7809 21394 -7775
rect 21562 -7809 21578 -7775
rect 21332 -7868 21366 -7852
rect 21104 -11660 21138 -11644
rect 20892 -11737 20908 -11703
rect 21076 -11737 21092 -11703
rect 20732 -11805 20766 -11743
rect 21332 -11660 21366 -11644
rect 21590 -7868 21624 -7852
rect 21590 -11660 21624 -11644
rect 22190 -7769 22224 -7707
rect 21864 -7809 21880 -7775
rect 22048 -7809 22064 -7775
rect 21818 -7868 21852 -7852
rect 21378 -11737 21394 -11703
rect 21562 -11737 21578 -11703
rect 21218 -11805 21252 -11743
rect 21818 -11660 21852 -11644
rect 22076 -7868 22110 -7852
rect 22076 -11660 22110 -11644
rect 21864 -11737 21880 -11703
rect 22048 -11737 22064 -11703
rect 21704 -11805 21738 -11743
rect 53464 -7590 53498 -7574
rect 53464 -8382 53498 -8366
rect 53642 -7590 53676 -7574
rect 53642 -8382 53676 -8366
rect 53756 -8064 53790 -7438
rect 53896 -7410 53930 -7348
rect 55028 -7410 55062 -7348
rect 55710 -7354 56040 -7308
rect 54075 -7462 54091 -7428
rect 54867 -7462 54883 -7428
rect 53998 -7490 54032 -7474
rect 53998 -7544 54032 -7528
rect 54926 -7490 54960 -7474
rect 54926 -7544 54960 -7528
rect 54075 -7590 54091 -7556
rect 54867 -7590 54883 -7556
rect 53896 -7670 53930 -7608
rect 55706 -7388 55802 -7354
rect 56050 -7388 56146 -7354
rect 55706 -7450 55740 -7388
rect 55028 -7670 55062 -7608
rect 53896 -7704 53992 -7670
rect 54966 -7704 55062 -7670
rect 55176 -7500 55272 -7466
rect 55430 -7500 55526 -7466
rect 55176 -7562 55210 -7500
rect 55492 -7562 55526 -7500
rect 55318 -7602 55334 -7568
rect 55368 -7602 55384 -7568
rect 55290 -7652 55324 -7636
rect 55290 -7844 55324 -7828
rect 55378 -7652 55412 -7636
rect 55378 -7844 55412 -7828
rect 55176 -7918 55210 -7856
rect 55492 -7918 55526 -7856
rect 54870 -7952 55272 -7918
rect 55430 -7952 55706 -7918
rect 54870 -7958 55706 -7952
rect 54870 -8064 54904 -7958
rect 53756 -8098 53852 -8064
rect 54808 -8098 54904 -8064
rect 53756 -8160 53790 -8098
rect 54870 -8160 54904 -8098
rect 55126 -8108 55142 -8074
rect 55494 -8108 55510 -8074
rect 53926 -8212 53942 -8178
rect 54718 -8212 54734 -8178
rect 53858 -8240 53892 -8224
rect 53858 -8344 53892 -8328
rect 54768 -8240 54802 -8224
rect 54768 -8344 54802 -8328
rect 53926 -8390 53942 -8356
rect 54718 -8390 54734 -8356
rect 53510 -8450 53526 -8416
rect 53614 -8450 53630 -8416
rect 53756 -8470 53790 -8408
rect 55046 -8160 55080 -8144
rect 55046 -8210 55080 -8194
rect 55556 -8160 55590 -8144
rect 55556 -8210 55590 -8194
rect 55126 -8280 55142 -8246
rect 55494 -8280 55510 -8246
rect 54870 -8438 54904 -8408
rect 55700 -8406 55706 -7958
rect 56112 -7450 56146 -7388
rect 58930 -7367 59026 -7333
rect 59600 -7367 59696 -7333
rect 58930 -7410 58964 -7367
rect 58926 -7420 58966 -7410
rect 55866 -7490 55882 -7456
rect 55970 -7490 55986 -7456
rect 55820 -7540 55854 -7524
rect 55820 -8332 55854 -8316
rect 55998 -7540 56032 -7524
rect 55998 -8332 56032 -8316
rect 55866 -8400 55882 -8366
rect 55970 -8400 55986 -8366
rect 55700 -8438 55740 -8406
rect 57096 -7479 57125 -7445
rect 57159 -7479 57217 -7445
rect 57251 -7479 57309 -7445
rect 57343 -7479 57372 -7445
rect 57129 -7529 57165 -7513
rect 57129 -7563 57131 -7529
rect 57129 -7597 57165 -7563
rect 57129 -7631 57131 -7597
rect 57201 -7529 57267 -7479
rect 57201 -7563 57217 -7529
rect 57251 -7563 57267 -7529
rect 57201 -7597 57267 -7563
rect 57201 -7631 57217 -7597
rect 57251 -7631 57267 -7597
rect 57301 -7529 57355 -7513
rect 57301 -7563 57303 -7529
rect 57337 -7563 57355 -7529
rect 57301 -7610 57355 -7563
rect 57129 -7665 57165 -7631
rect 57301 -7644 57303 -7610
rect 57337 -7644 57355 -7610
rect 57129 -7699 57264 -7665
rect 57301 -7694 57355 -7644
rect 57230 -7728 57264 -7699
rect 57117 -7744 57185 -7735
rect 57117 -7794 57118 -7744
rect 57178 -7794 57185 -7744
rect 57117 -7809 57185 -7794
rect 57230 -7744 57285 -7728
rect 57230 -7778 57251 -7744
rect 57230 -7794 57285 -7778
rect 57319 -7740 57355 -7694
rect 59662 -7429 59696 -7367
rect 59109 -7481 59125 -7447
rect 59501 -7481 59517 -7447
rect 59560 -7501 59594 -7485
rect 59560 -7551 59594 -7535
rect 59109 -7589 59125 -7555
rect 59501 -7589 59517 -7555
rect 59032 -7609 59066 -7593
rect 59032 -7659 59066 -7643
rect 59109 -7697 59125 -7663
rect 59501 -7697 59517 -7663
rect 58926 -7740 58966 -7720
rect 57319 -7780 57326 -7740
rect 58930 -7776 58964 -7740
rect 57230 -7845 57264 -7794
rect 57131 -7879 57264 -7845
rect 57319 -7854 57355 -7780
rect 57131 -7900 57165 -7879
rect 56316 -7918 56412 -7904
rect 54830 -8448 55830 -8438
rect 54830 -8470 55030 -8448
rect 53756 -8504 53852 -8470
rect 54808 -8504 55030 -8470
rect 53510 -8558 53526 -8524
rect 53614 -8558 53630 -8524
rect 53756 -8566 53790 -8504
rect 54830 -8528 55030 -8504
rect 55110 -8468 55740 -8448
rect 55810 -8468 55830 -8448
rect 56112 -8468 56146 -8406
rect 55110 -8508 55160 -8468
rect 55600 -8508 55740 -8468
rect 56050 -8502 56146 -8468
rect 55110 -8528 55740 -8508
rect 55810 -8528 55830 -8502
rect 54830 -8538 55830 -8528
rect 53464 -8608 53498 -8592
rect 53464 -9400 53498 -9384
rect 53642 -8608 53676 -8592
rect 53642 -9400 53676 -9384
rect 54870 -8566 54904 -8538
rect 53926 -8618 53942 -8584
rect 54718 -8618 54734 -8584
rect 53858 -8646 53892 -8630
rect 53858 -8750 53892 -8734
rect 54768 -8646 54802 -8630
rect 54768 -8750 54802 -8734
rect 53926 -8796 53942 -8762
rect 54718 -8796 54734 -8762
rect 53756 -8876 53790 -8814
rect 55700 -8564 55740 -8538
rect 55126 -8730 55142 -8696
rect 55494 -8730 55510 -8696
rect 54870 -8876 54904 -8814
rect 55046 -8782 55080 -8766
rect 55046 -8832 55080 -8816
rect 55556 -8782 55590 -8766
rect 55556 -8832 55590 -8816
rect 53756 -8910 53852 -8876
rect 54808 -8910 54904 -8876
rect 55126 -8902 55142 -8868
rect 55494 -8902 55510 -8868
rect 53510 -9468 53526 -9434
rect 53614 -9468 53630 -9434
rect 53350 -9536 53384 -9474
rect 53756 -9536 53790 -8910
rect 54870 -9018 54904 -8910
rect 55700 -9018 55706 -8564
rect 54870 -9024 55706 -9018
rect 54870 -9058 55262 -9024
rect 55420 -9058 55706 -9024
rect 55166 -9120 55200 -9058
rect 53350 -9570 53446 -9536
rect 53694 -9570 53790 -9536
rect 53886 -9308 53982 -9274
rect 54956 -9308 55052 -9274
rect 53886 -9370 53920 -9308
rect 55018 -9370 55052 -9308
rect 54065 -9422 54081 -9388
rect 54857 -9422 54873 -9388
rect 53988 -9450 54022 -9434
rect 53988 -9504 54022 -9488
rect 54916 -9450 54950 -9434
rect 54916 -9504 54950 -9488
rect 54065 -9550 54081 -9516
rect 54857 -9550 54873 -9516
rect 53886 -9630 53920 -9568
rect 55482 -9120 55516 -9058
rect 55280 -9148 55314 -9132
rect 55280 -9340 55314 -9324
rect 55368 -9148 55402 -9132
rect 55368 -9340 55402 -9324
rect 55308 -9408 55324 -9374
rect 55358 -9408 55374 -9374
rect 55166 -9476 55200 -9414
rect 55482 -9476 55516 -9414
rect 55166 -9510 55262 -9476
rect 55420 -9510 55516 -9476
rect 55018 -9630 55052 -9568
rect 56112 -8564 56146 -8502
rect 56350 -7938 56412 -7918
rect 56610 -7938 56706 -7904
rect 56672 -8000 56706 -7938
rect 57303 -7883 57355 -7854
rect 57131 -7955 57165 -7934
rect 57201 -7947 57217 -7913
rect 57251 -7947 57267 -7913
rect 57201 -7989 57267 -7947
rect 57337 -7917 57355 -7883
rect 57303 -7955 57355 -7917
rect 58930 -7810 59026 -7776
rect 59214 -7777 59310 -7776
rect 59662 -7777 59696 -7720
rect 59772 -7694 59866 -7660
rect 60426 -7694 60520 -7660
rect 59772 -7750 59806 -7694
rect 59214 -7810 59696 -7777
rect 58930 -7811 59696 -7810
rect 58930 -7872 58964 -7811
rect 59276 -7872 59310 -7811
rect 59087 -7912 59103 -7878
rect 59137 -7912 59153 -7878
rect 56476 -8040 56492 -8006
rect 56530 -8040 56546 -8006
rect 55866 -8604 55882 -8570
rect 55970 -8604 55986 -8570
rect 55820 -8654 55854 -8638
rect 55820 -9446 55854 -9430
rect 55998 -8654 56032 -8638
rect 55998 -9446 56032 -9430
rect 55866 -9514 55882 -9480
rect 55970 -9514 55986 -9480
rect 55706 -9582 55740 -9520
rect 56430 -8099 56464 -8083
rect 56430 -8891 56464 -8875
rect 56558 -8099 56592 -8083
rect 56558 -8891 56592 -8875
rect 56476 -8968 56492 -8934
rect 56530 -8968 56546 -8934
rect 56316 -9036 56350 -8974
rect 57096 -8023 57125 -7989
rect 57159 -8023 57217 -7989
rect 57251 -8023 57309 -7989
rect 57343 -8023 57372 -7989
rect 59044 -7971 59078 -7955
rect 59044 -8363 59078 -8347
rect 59162 -7971 59196 -7955
rect 59162 -8363 59196 -8347
rect 59087 -8440 59103 -8406
rect 59137 -8440 59153 -8406
rect 60486 -7756 60520 -7694
rect 59942 -7808 59958 -7774
rect 60334 -7808 60350 -7774
rect 59874 -7828 59908 -7812
rect 59874 -7878 59908 -7862
rect 60384 -7828 60418 -7812
rect 60384 -7878 60418 -7862
rect 59942 -7916 59958 -7882
rect 60334 -7916 60350 -7882
rect 59772 -7996 59806 -7940
rect 60486 -7996 60520 -7934
rect 59388 -8030 59476 -7996
rect 59656 -8030 59800 -7996
rect 59958 -8030 60520 -7996
rect 59388 -8090 59422 -8030
rect 59276 -8506 59310 -8446
rect 59530 -8132 59546 -8098
rect 59580 -8132 59596 -8098
rect 59502 -8182 59536 -8166
rect 59502 -8374 59536 -8358
rect 59590 -8182 59624 -8166
rect 59590 -8374 59624 -8358
rect 59530 -8442 59546 -8408
rect 59580 -8442 59596 -8408
rect 58966 -8542 59310 -8506
rect 59388 -8509 59422 -8450
rect 59704 -8509 59738 -8030
rect 60020 -8092 60054 -8030
rect 59846 -8132 59862 -8098
rect 59896 -8132 59912 -8098
rect 59818 -8182 59852 -8166
rect 59818 -8374 59852 -8358
rect 59906 -8182 59940 -8166
rect 59906 -8374 59940 -8358
rect 59846 -8442 59862 -8408
rect 59896 -8442 59912 -8408
rect 61186 -8200 61286 -8190
rect 61186 -8280 61196 -8200
rect 61186 -8290 61286 -8280
rect 60020 -8509 60054 -8448
rect 56672 -9036 56706 -8974
rect 57096 -8999 57125 -8965
rect 57159 -8999 57217 -8965
rect 57251 -8999 57309 -8965
rect 57343 -8999 57372 -8965
rect 56316 -9070 56412 -9036
rect 56610 -9070 56706 -9036
rect 57131 -9054 57165 -9033
rect 57201 -9041 57267 -8999
rect 57201 -9075 57217 -9041
rect 57251 -9075 57267 -9041
rect 57303 -9071 57355 -9033
rect 57131 -9109 57165 -9088
rect 57337 -9105 57355 -9071
rect 59276 -8602 59310 -8542
rect 59387 -8544 60054 -8509
rect 60127 -8354 60161 -8328
rect 60127 -8357 60253 -8354
rect 60161 -8373 60253 -8357
rect 60161 -8391 60203 -8373
rect 60127 -8407 60203 -8391
rect 60237 -8407 60253 -8373
rect 60359 -8360 60409 -8349
rect 60671 -8354 60705 -8328
rect 60359 -8365 60366 -8360
rect 60359 -8400 60366 -8399
rect 60406 -8400 60409 -8360
rect 60127 -8449 60161 -8407
rect 60127 -8541 60161 -8483
rect 60195 -8457 60325 -8441
rect 60195 -8491 60211 -8457
rect 60245 -8491 60325 -8457
rect 60195 -8507 60325 -8491
rect 59387 -8600 59421 -8544
rect 59087 -8642 59103 -8608
rect 59137 -8642 59153 -8608
rect 59044 -8701 59078 -8685
rect 57131 -9143 57264 -9109
rect 57303 -9134 57355 -9105
rect 57117 -9194 57185 -9179
rect 57117 -9244 57118 -9194
rect 57168 -9244 57185 -9194
rect 57117 -9253 57185 -9244
rect 57230 -9194 57264 -9143
rect 57319 -9170 57355 -9134
rect 57230 -9210 57285 -9194
rect 57230 -9244 57251 -9210
rect 57230 -9260 57285 -9244
rect 57319 -9210 57326 -9170
rect 59044 -9093 59078 -9077
rect 59162 -8701 59196 -8685
rect 59162 -9093 59196 -9077
rect 59087 -9170 59103 -9136
rect 59137 -9170 59153 -9136
rect 57230 -9289 57264 -9260
rect 57129 -9323 57264 -9289
rect 57319 -9294 57355 -9210
rect 57129 -9357 57165 -9323
rect 57301 -9344 57355 -9294
rect 58930 -9238 58964 -9176
rect 59529 -8645 59545 -8611
rect 59579 -8645 59595 -8611
rect 59501 -8695 59535 -8679
rect 59501 -8887 59535 -8871
rect 59589 -8695 59623 -8679
rect 59589 -8887 59623 -8871
rect 59529 -8955 59545 -8921
rect 59579 -8955 59595 -8921
rect 59387 -9023 59421 -8970
rect 59703 -9023 59737 -8544
rect 60019 -8605 60053 -8544
rect 59845 -8645 59861 -8611
rect 59895 -8645 59911 -8611
rect 59817 -8695 59851 -8679
rect 59817 -8887 59851 -8871
rect 59905 -8695 59939 -8679
rect 59905 -8887 59939 -8871
rect 59845 -8955 59861 -8921
rect 59895 -8955 59911 -8921
rect 60161 -8575 60203 -8541
rect 60237 -8575 60253 -8541
rect 60127 -8633 60161 -8575
rect 60289 -8609 60325 -8507
rect 60127 -8709 60161 -8667
rect 60195 -8625 60325 -8609
rect 60195 -8659 60211 -8625
rect 60245 -8659 60325 -8625
rect 60195 -8675 60325 -8659
rect 60359 -8450 60409 -8400
rect 60443 -8357 60705 -8354
rect 60443 -8373 60671 -8357
rect 60443 -8407 60459 -8373
rect 60493 -8407 60527 -8373
rect 60561 -8407 60595 -8373
rect 60629 -8391 60671 -8373
rect 60629 -8407 60705 -8391
rect 60359 -8457 60366 -8450
rect 60406 -8490 60409 -8450
rect 60393 -8491 60409 -8490
rect 60359 -8540 60409 -8491
rect 60359 -8541 60366 -8540
rect 60359 -8580 60366 -8575
rect 60406 -8580 60409 -8540
rect 60359 -8620 60409 -8580
rect 60359 -8625 60366 -8620
rect 60359 -8660 60366 -8659
rect 60406 -8660 60409 -8620
rect 60359 -8675 60409 -8660
rect 60443 -8457 60637 -8441
rect 60443 -8491 60459 -8457
rect 60493 -8491 60527 -8457
rect 60561 -8491 60595 -8457
rect 60629 -8491 60637 -8457
rect 60443 -8507 60637 -8491
rect 60671 -8449 60705 -8407
rect 60443 -8609 60477 -8507
rect 60671 -8541 60705 -8483
rect 60511 -8575 60527 -8541
rect 60561 -8575 60595 -8541
rect 60629 -8575 60671 -8541
rect 60443 -8625 60637 -8609
rect 60443 -8659 60459 -8625
rect 60493 -8659 60527 -8625
rect 60561 -8659 60595 -8625
rect 60629 -8659 60637 -8625
rect 60443 -8675 60637 -8659
rect 60671 -8633 60705 -8575
rect 60289 -8709 60325 -8675
rect 60443 -8709 60481 -8675
rect 60671 -8709 60705 -8667
rect 60127 -8725 60204 -8709
rect 60161 -8743 60204 -8725
rect 60238 -8743 60254 -8709
rect 60161 -8759 60254 -8743
rect 60289 -8725 60481 -8709
rect 60289 -8759 60297 -8725
rect 60331 -8759 60369 -8725
rect 60405 -8759 60449 -8725
rect 60579 -8743 60595 -8709
rect 60629 -8725 60705 -8709
rect 60629 -8743 60671 -8725
rect 60579 -8751 60671 -8743
rect 60127 -8788 60161 -8759
rect 60289 -8762 60481 -8759
rect 60671 -8788 60705 -8759
rect 60747 -8354 60781 -8328
rect 60747 -8357 61009 -8354
rect 60781 -8373 61009 -8357
rect 60781 -8391 60823 -8373
rect 60747 -8407 60823 -8391
rect 60857 -8407 60891 -8373
rect 60925 -8407 60959 -8373
rect 60993 -8407 61009 -8373
rect 61043 -8360 61093 -8349
rect 61291 -8354 61325 -8328
rect 61043 -8400 61046 -8360
rect 61086 -8365 61093 -8360
rect 61086 -8400 61093 -8399
rect 60747 -8449 60781 -8407
rect 60747 -8541 60781 -8483
rect 60815 -8457 61009 -8441
rect 60815 -8491 60823 -8457
rect 60857 -8491 60891 -8457
rect 60925 -8491 60959 -8457
rect 60993 -8491 61009 -8457
rect 60815 -8507 61009 -8491
rect 60781 -8575 60823 -8541
rect 60857 -8575 60891 -8541
rect 60925 -8575 60941 -8541
rect 60747 -8633 60781 -8575
rect 60975 -8609 61009 -8507
rect 60747 -8709 60781 -8667
rect 60815 -8625 61009 -8609
rect 60815 -8659 60823 -8625
rect 60857 -8659 60891 -8625
rect 60925 -8659 60959 -8625
rect 60993 -8659 61009 -8625
rect 60815 -8675 61009 -8659
rect 61043 -8450 61093 -8400
rect 61199 -8357 61325 -8354
rect 61199 -8373 61291 -8357
rect 61199 -8407 61215 -8373
rect 61249 -8391 61291 -8373
rect 61249 -8407 61325 -8391
rect 61043 -8490 61046 -8450
rect 61086 -8457 61093 -8450
rect 61043 -8491 61059 -8490
rect 61043 -8540 61093 -8491
rect 61043 -8580 61046 -8540
rect 61086 -8541 61093 -8540
rect 61086 -8580 61093 -8575
rect 61043 -8620 61093 -8580
rect 61043 -8660 61046 -8620
rect 61086 -8625 61093 -8620
rect 61086 -8660 61093 -8659
rect 61043 -8675 61093 -8660
rect 61127 -8457 61257 -8441
rect 61127 -8491 61207 -8457
rect 61241 -8491 61257 -8457
rect 61127 -8507 61257 -8491
rect 61291 -8449 61325 -8407
rect 61127 -8609 61163 -8507
rect 61291 -8541 61325 -8483
rect 61199 -8575 61215 -8541
rect 61249 -8575 61291 -8541
rect 61127 -8625 61257 -8609
rect 61127 -8659 61207 -8625
rect 61241 -8659 61257 -8625
rect 61127 -8675 61257 -8659
rect 61291 -8633 61325 -8575
rect 60971 -8709 61009 -8675
rect 61127 -8709 61163 -8675
rect 61291 -8709 61325 -8667
rect 60747 -8725 60823 -8709
rect 60781 -8743 60823 -8725
rect 60857 -8743 60873 -8709
rect 60781 -8751 60873 -8743
rect 60971 -8724 61163 -8709
rect 60971 -8725 61129 -8724
rect 60747 -8788 60781 -8759
rect 60971 -8759 60980 -8725
rect 61015 -8759 61053 -8725
rect 61088 -8758 61129 -8725
rect 61198 -8743 61214 -8709
rect 61248 -8725 61325 -8709
rect 61248 -8743 61291 -8725
rect 61088 -8759 61163 -8758
rect 61198 -8759 61291 -8743
rect 60971 -8762 61163 -8759
rect 61291 -8788 61325 -8759
rect 60466 -8860 60546 -8840
rect 60466 -8900 60486 -8860
rect 60526 -8900 60546 -8860
rect 60466 -8920 60546 -8900
rect 60606 -8860 60686 -8840
rect 60606 -8900 60626 -8860
rect 60666 -8900 60686 -8860
rect 60606 -8920 60686 -8900
rect 60746 -8860 60826 -8840
rect 60746 -8900 60766 -8860
rect 60806 -8900 60826 -8860
rect 60746 -8920 60826 -8900
rect 60886 -8860 60966 -8840
rect 60886 -8900 60906 -8860
rect 60946 -8900 60966 -8860
rect 60886 -8920 60966 -8900
rect 60019 -9023 60053 -8961
rect 59387 -9057 59476 -9023
rect 59646 -9057 59799 -9023
rect 59957 -9026 60053 -9023
rect 59957 -9057 60520 -9026
rect 59772 -9060 60520 -9057
rect 59772 -9120 59806 -9060
rect 59276 -9238 59310 -9176
rect 58930 -9272 59026 -9238
rect 59214 -9240 59310 -9238
rect 59214 -9272 59696 -9240
rect 58930 -9274 59696 -9272
rect 58930 -9310 58964 -9274
rect 57129 -9391 57131 -9357
rect 57129 -9425 57165 -9391
rect 57129 -9459 57131 -9425
rect 57129 -9475 57165 -9459
rect 57201 -9391 57217 -9357
rect 57251 -9391 57267 -9357
rect 57201 -9425 57267 -9391
rect 57201 -9459 57217 -9425
rect 57251 -9459 57267 -9425
rect 57201 -9509 57267 -9459
rect 57301 -9378 57303 -9344
rect 57337 -9378 57355 -9344
rect 57301 -9425 57355 -9378
rect 57301 -9459 57303 -9425
rect 57337 -9459 57355 -9425
rect 57301 -9475 57355 -9459
rect 59662 -9330 59696 -9274
rect 60486 -9122 60520 -9060
rect 59942 -9174 59958 -9140
rect 60334 -9174 60350 -9140
rect 59874 -9194 59908 -9178
rect 59874 -9244 59908 -9228
rect 60384 -9194 60418 -9178
rect 60384 -9244 60418 -9228
rect 59942 -9282 59958 -9248
rect 60334 -9282 60350 -9248
rect 56112 -9582 56146 -9520
rect 57096 -9543 57125 -9509
rect 57159 -9543 57217 -9509
rect 57251 -9543 57309 -9509
rect 57343 -9543 57372 -9509
rect 55706 -9616 55802 -9582
rect 56050 -9616 56146 -9582
rect 53886 -9664 53982 -9630
rect 54956 -9664 55052 -9630
rect 53886 -9726 53920 -9664
rect 55018 -9726 55052 -9664
rect 55720 -9658 56090 -9616
rect 55720 -9668 56020 -9658
rect 54065 -9778 54081 -9744
rect 54857 -9778 54873 -9744
rect 53988 -9806 54022 -9790
rect 53988 -9860 54022 -9844
rect 54916 -9806 54950 -9790
rect 54916 -9860 54950 -9844
rect 54065 -9906 54081 -9872
rect 54857 -9906 54873 -9872
rect 53886 -9986 53920 -9924
rect 56010 -9808 56020 -9668
rect 56080 -9808 56090 -9658
rect 59109 -9388 59125 -9354
rect 59501 -9388 59517 -9354
rect 59560 -9408 59594 -9392
rect 59560 -9458 59594 -9442
rect 59109 -9496 59125 -9462
rect 59501 -9496 59517 -9462
rect 59032 -9516 59066 -9500
rect 59032 -9566 59066 -9550
rect 59109 -9604 59125 -9570
rect 59501 -9604 59517 -9570
rect 56010 -9818 56090 -9808
rect 59772 -9362 59806 -9300
rect 60486 -9362 60520 -9300
rect 59772 -9396 59866 -9362
rect 60426 -9396 60520 -9362
rect 59662 -9684 59696 -9630
rect 58966 -9700 59026 -9684
rect 58930 -9718 59026 -9700
rect 59600 -9718 59696 -9684
rect 55018 -9986 55052 -9924
rect 53886 -10020 53982 -9986
rect 54956 -10020 55052 -9986
rect 55176 -9878 55272 -9844
rect 55566 -9878 55662 -9844
rect 55176 -9940 55210 -9878
rect 55628 -9940 55662 -9878
rect 55284 -9992 55300 -9958
rect 55476 -9992 55492 -9958
rect 55526 -10002 55560 -9986
rect 55284 -10080 55300 -10046
rect 55476 -10080 55492 -10046
rect 55526 -10052 55560 -10036
rect 55176 -10160 55210 -10098
rect 55628 -10160 55662 -10098
rect 55176 -10194 55272 -10160
rect 55566 -10194 55662 -10160
rect 22190 -11805 22224 -11743
rect 20156 -11850 20252 -11816
rect 20430 -11850 20526 -11816
rect 20732 -11839 20828 -11805
rect 21156 -11839 21314 -11805
rect 21642 -11839 21800 -11805
rect 22128 -11839 22224 -11805
rect 20156 -11912 20190 -11850
rect 20492 -11912 20526 -11850
rect 20264 -11964 20280 -11930
rect 20340 -11964 20356 -11930
rect 20390 -11974 20424 -11958
rect 20264 -12052 20280 -12018
rect 20340 -12052 20356 -12018
rect 20390 -12024 20424 -12008
rect 20156 -12122 20190 -12070
rect 20492 -12122 20526 -12070
rect 16439 -12182 16440 -12143
rect 16439 -12239 16473 -12182
rect 16845 -12239 16879 -12182
rect 16599 -12279 16615 -12245
rect 16703 -12279 16719 -12245
rect 16553 -12329 16587 -12313
rect 16553 -13121 16587 -13105
rect 16731 -12329 16765 -12313
rect 16731 -13121 16765 -13105
rect 16599 -13189 16615 -13155
rect 16703 -13189 16719 -13155
rect 16439 -13254 16473 -13195
rect 17251 -12239 17285 -12182
rect 17005 -12279 17021 -12245
rect 17109 -12279 17125 -12245
rect 16959 -12329 16993 -12313
rect 16959 -13121 16993 -13105
rect 17137 -12329 17171 -12313
rect 17137 -13121 17171 -13105
rect 17005 -13189 17021 -13155
rect 17109 -13189 17125 -13155
rect 16845 -13254 16879 -13195
rect 17657 -12239 17691 -12182
rect 17411 -12279 17427 -12245
rect 17515 -12279 17531 -12245
rect 17365 -12329 17399 -12313
rect 17365 -13121 17399 -13105
rect 17543 -12329 17577 -12313
rect 17543 -13121 17577 -13105
rect 17411 -13189 17427 -13155
rect 17515 -13189 17531 -13155
rect 17251 -13254 17285 -13195
rect 18063 -12239 18097 -12182
rect 17817 -12279 17833 -12245
rect 17921 -12279 17937 -12245
rect 17771 -12329 17805 -12313
rect 17771 -13121 17805 -13105
rect 17949 -12329 17983 -12313
rect 17949 -13121 17983 -13105
rect 17817 -13189 17833 -13155
rect 17921 -13189 17937 -13155
rect 17657 -13254 17691 -13195
rect 18469 -12239 18503 -12182
rect 18223 -12279 18239 -12245
rect 18327 -12279 18343 -12245
rect 18177 -12329 18211 -12313
rect 18177 -13121 18211 -13105
rect 18355 -12329 18389 -12313
rect 18355 -13121 18389 -13105
rect 18223 -13189 18239 -13155
rect 18327 -13189 18343 -13155
rect 18063 -13254 18097 -13195
rect 18875 -12239 18909 -12182
rect 18629 -12279 18645 -12245
rect 18733 -12279 18749 -12245
rect 18583 -12329 18617 -12313
rect 18583 -13121 18617 -13105
rect 18761 -12329 18795 -12313
rect 18761 -13121 18795 -13105
rect 18629 -13189 18645 -13155
rect 18733 -13189 18749 -13155
rect 18469 -13254 18503 -13195
rect 19281 -12239 19315 -12182
rect 19035 -12279 19051 -12245
rect 19139 -12279 19155 -12245
rect 18989 -12329 19023 -12313
rect 18989 -13121 19023 -13105
rect 19167 -12329 19201 -12313
rect 19167 -13121 19201 -13105
rect 19035 -13189 19051 -13155
rect 19139 -13189 19155 -13155
rect 18875 -13254 18909 -13195
rect 19687 -12239 19721 -12182
rect 19441 -12279 19457 -12245
rect 19545 -12279 19561 -12245
rect 19395 -12329 19429 -12313
rect 19395 -13121 19429 -13105
rect 19573 -12329 19607 -12313
rect 19573 -13121 19607 -13105
rect 19441 -13189 19457 -13155
rect 19545 -13189 19561 -13155
rect 19281 -13254 19315 -13195
rect 20093 -12239 20127 -12182
rect 19847 -12279 19863 -12245
rect 19951 -12279 19967 -12245
rect 19801 -12329 19835 -12313
rect 19801 -13121 19835 -13105
rect 19979 -12329 20013 -12313
rect 19979 -13121 20013 -13105
rect 19847 -13189 19863 -13155
rect 19951 -13189 19967 -13155
rect 19687 -13254 19721 -13195
rect 20499 -12239 20533 -12182
rect 20253 -12279 20269 -12245
rect 20357 -12279 20373 -12245
rect 20207 -12329 20241 -12313
rect 20207 -13121 20241 -13105
rect 20385 -12329 20419 -12313
rect 20385 -13121 20419 -13105
rect 20253 -13189 20269 -13155
rect 20357 -13189 20373 -13155
rect 20093 -13254 20127 -13195
rect 20905 -12239 20939 -12182
rect 20659 -12279 20675 -12245
rect 20763 -12279 20779 -12245
rect 20613 -12329 20647 -12313
rect 20613 -13121 20647 -13105
rect 20791 -12329 20825 -12313
rect 20791 -13121 20825 -13105
rect 20659 -13189 20675 -13155
rect 20763 -13189 20779 -13155
rect 20499 -13254 20533 -13195
rect 21311 -12239 21345 -12182
rect 21065 -12279 21081 -12245
rect 21169 -12279 21185 -12245
rect 21019 -12329 21053 -12313
rect 21019 -13121 21053 -13105
rect 21197 -12329 21231 -12313
rect 21197 -13121 21231 -13105
rect 21065 -13189 21081 -13155
rect 21169 -13189 21185 -13155
rect 20905 -13254 20939 -13195
rect 21717 -12239 21751 -12182
rect 21471 -12279 21487 -12245
rect 21575 -12279 21591 -12245
rect 21425 -12329 21459 -12313
rect 21425 -13121 21459 -13105
rect 21603 -12329 21637 -12313
rect 21603 -13121 21637 -13105
rect 21471 -13189 21487 -13155
rect 21575 -13189 21591 -13155
rect 21311 -13254 21345 -13195
rect 22123 -12239 22157 -12182
rect 21877 -12279 21893 -12245
rect 21981 -12279 21997 -12245
rect 21831 -12329 21865 -12313
rect 21831 -13121 21865 -13105
rect 22009 -12329 22043 -12313
rect 22009 -13121 22043 -13105
rect 21877 -13189 21893 -13155
rect 21981 -13189 21997 -13155
rect 21717 -13254 21751 -13195
rect 22529 -12239 22563 -12182
rect 22283 -12279 22299 -12245
rect 22387 -12279 22403 -12245
rect 22237 -12329 22271 -12313
rect 22237 -13121 22271 -13105
rect 22415 -12329 22449 -12313
rect 22415 -13121 22449 -13105
rect 22283 -13189 22299 -13155
rect 22387 -13189 22403 -13155
rect 22123 -13254 22157 -13195
rect 22935 -12239 22969 -12182
rect 22689 -12279 22705 -12245
rect 22793 -12279 22809 -12245
rect 22643 -12329 22677 -12313
rect 22643 -13121 22677 -13105
rect 22821 -12329 22855 -12313
rect 22821 -13121 22855 -13105
rect 22689 -13189 22705 -13155
rect 22793 -13189 22809 -13155
rect 22529 -13254 22563 -13195
rect 23341 -12239 23375 -12182
rect 23095 -12279 23111 -12245
rect 23199 -12279 23215 -12245
rect 23049 -12329 23083 -12313
rect 23049 -13121 23083 -13105
rect 23227 -12329 23261 -12313
rect 23227 -13121 23261 -13105
rect 23095 -13189 23111 -13155
rect 23199 -13189 23215 -13155
rect 22935 -13254 22969 -13195
rect 23747 -12239 23781 -12182
rect 23501 -12279 23517 -12245
rect 23605 -12279 23621 -12245
rect 23455 -12329 23489 -12313
rect 23455 -13121 23489 -13105
rect 23633 -12329 23667 -12313
rect 23633 -13121 23667 -13105
rect 23501 -13189 23517 -13155
rect 23605 -13189 23621 -13155
rect 23341 -13254 23375 -13195
rect 24153 -12239 24187 -12182
rect 23907 -12279 23923 -12245
rect 24011 -12279 24027 -12245
rect 23861 -12329 23895 -12313
rect 23861 -13121 23895 -13105
rect 24039 -12329 24073 -12313
rect 24039 -13121 24073 -13105
rect 23907 -13189 23923 -13155
rect 24011 -13189 24027 -13155
rect 23747 -13254 23781 -13195
rect 24559 -12239 24593 -12182
rect 24313 -12279 24329 -12245
rect 24417 -12279 24433 -12245
rect 24267 -12329 24301 -12313
rect 24267 -13121 24301 -13105
rect 24445 -12329 24479 -12313
rect 24445 -13121 24479 -13105
rect 24313 -13189 24329 -13155
rect 24417 -13189 24433 -13155
rect 24153 -13254 24187 -13195
rect 24965 -12239 24999 -12182
rect 24719 -12279 24735 -12245
rect 24823 -12279 24839 -12245
rect 24673 -12329 24707 -12313
rect 24673 -13121 24707 -13105
rect 24851 -12329 24885 -12313
rect 24851 -13121 24885 -13105
rect 24719 -13189 24735 -13155
rect 24823 -13189 24839 -13155
rect 24559 -13254 24593 -13195
rect 25125 -12279 25141 -12245
rect 25229 -12279 25245 -12245
rect 25079 -12329 25113 -12313
rect 25079 -13121 25113 -13105
rect 25257 -12329 25291 -12313
rect 25257 -13121 25291 -13105
rect 25360 -13149 25362 -12276
rect 25125 -13189 25141 -13155
rect 25229 -13189 25245 -13155
rect 24965 -13254 24999 -13195
rect 25360 -13219 25361 -13149
rect 53896 -12392 53992 -12358
rect 54966 -12392 55062 -12358
rect 53896 -12454 53930 -12392
rect 55028 -12454 55062 -12392
rect 54075 -12506 54091 -12472
rect 54867 -12506 54883 -12472
rect 53998 -12534 54032 -12518
rect 53998 -12588 54032 -12572
rect 54926 -12534 54960 -12518
rect 54926 -12588 54960 -12572
rect 54075 -12634 54091 -12600
rect 54867 -12634 54883 -12600
rect 53896 -12714 53930 -12652
rect 55028 -12714 55062 -12652
rect 55960 -12708 56040 -12698
rect 53896 -12748 53992 -12714
rect 54966 -12748 55062 -12714
rect 53350 -12838 53790 -12804
rect 53350 -12900 53384 -12838
rect 53510 -12940 53526 -12906
rect 53614 -12940 53630 -12906
rect 16439 -13291 16448 -13254
rect 53464 -12990 53498 -12974
rect 53464 -13782 53498 -13766
rect 53642 -12990 53676 -12974
rect 53642 -13782 53676 -13766
rect 53756 -13464 53790 -12838
rect 53896 -12810 53930 -12748
rect 55028 -12810 55062 -12748
rect 55710 -12754 56040 -12708
rect 54075 -12862 54091 -12828
rect 54867 -12862 54883 -12828
rect 53998 -12890 54032 -12874
rect 53998 -12944 54032 -12928
rect 54926 -12890 54960 -12874
rect 54926 -12944 54960 -12928
rect 54075 -12990 54091 -12956
rect 54867 -12990 54883 -12956
rect 53896 -13070 53930 -13008
rect 55706 -12788 55802 -12754
rect 56050 -12788 56146 -12754
rect 55706 -12850 55740 -12788
rect 55028 -13070 55062 -13008
rect 53896 -13104 53992 -13070
rect 54966 -13104 55062 -13070
rect 55176 -12900 55272 -12866
rect 55430 -12900 55526 -12866
rect 55176 -12962 55210 -12900
rect 55492 -12962 55526 -12900
rect 55318 -13002 55334 -12968
rect 55368 -13002 55384 -12968
rect 55290 -13052 55324 -13036
rect 55290 -13244 55324 -13228
rect 55378 -13052 55412 -13036
rect 55378 -13244 55412 -13228
rect 55176 -13318 55210 -13256
rect 55492 -13318 55526 -13256
rect 54870 -13352 55272 -13318
rect 55430 -13352 55706 -13318
rect 54870 -13358 55706 -13352
rect 54870 -13464 54904 -13358
rect 53756 -13498 53852 -13464
rect 54808 -13498 54904 -13464
rect 53756 -13560 53790 -13498
rect 54870 -13560 54904 -13498
rect 55126 -13508 55142 -13474
rect 55494 -13508 55510 -13474
rect 53926 -13612 53942 -13578
rect 54718 -13612 54734 -13578
rect 53858 -13640 53892 -13624
rect 53858 -13744 53892 -13728
rect 54768 -13640 54802 -13624
rect 54768 -13744 54802 -13728
rect 53926 -13790 53942 -13756
rect 54718 -13790 54734 -13756
rect 53510 -13850 53526 -13816
rect 53614 -13850 53630 -13816
rect 53756 -13870 53790 -13808
rect 55046 -13560 55080 -13544
rect 55046 -13610 55080 -13594
rect 55556 -13560 55590 -13544
rect 55556 -13610 55590 -13594
rect 55126 -13680 55142 -13646
rect 55494 -13680 55510 -13646
rect 54870 -13838 54904 -13808
rect 55700 -13806 55706 -13358
rect 56112 -12850 56146 -12788
rect 58930 -12767 59026 -12733
rect 59600 -12767 59696 -12733
rect 58930 -12810 58964 -12767
rect 58926 -12820 58966 -12810
rect 55866 -12890 55882 -12856
rect 55970 -12890 55986 -12856
rect 55820 -12940 55854 -12924
rect 55820 -13732 55854 -13716
rect 55998 -12940 56032 -12924
rect 55998 -13732 56032 -13716
rect 55866 -13800 55882 -13766
rect 55970 -13800 55986 -13766
rect 55700 -13838 55740 -13806
rect 57096 -12879 57125 -12845
rect 57159 -12879 57217 -12845
rect 57251 -12879 57309 -12845
rect 57343 -12879 57372 -12845
rect 57129 -12929 57165 -12913
rect 57129 -12963 57131 -12929
rect 57129 -12997 57165 -12963
rect 57129 -13031 57131 -12997
rect 57201 -12929 57267 -12879
rect 57201 -12963 57217 -12929
rect 57251 -12963 57267 -12929
rect 57201 -12997 57267 -12963
rect 57201 -13031 57217 -12997
rect 57251 -13031 57267 -12997
rect 57301 -12929 57355 -12913
rect 57301 -12963 57303 -12929
rect 57337 -12963 57355 -12929
rect 57301 -13010 57355 -12963
rect 57129 -13065 57165 -13031
rect 57301 -13044 57303 -13010
rect 57337 -13044 57355 -13010
rect 57129 -13099 57264 -13065
rect 57301 -13094 57355 -13044
rect 57230 -13128 57264 -13099
rect 57117 -13144 57185 -13135
rect 57117 -13194 57118 -13144
rect 57178 -13194 57185 -13144
rect 57117 -13209 57185 -13194
rect 57230 -13144 57285 -13128
rect 57230 -13178 57251 -13144
rect 57230 -13194 57285 -13178
rect 57319 -13140 57355 -13094
rect 59662 -12829 59696 -12767
rect 59109 -12881 59125 -12847
rect 59501 -12881 59517 -12847
rect 59560 -12901 59594 -12885
rect 59560 -12951 59594 -12935
rect 59109 -12989 59125 -12955
rect 59501 -12989 59517 -12955
rect 59032 -13009 59066 -12993
rect 59032 -13059 59066 -13043
rect 59109 -13097 59125 -13063
rect 59501 -13097 59517 -13063
rect 58926 -13140 58966 -13120
rect 57319 -13180 57326 -13140
rect 58930 -13176 58964 -13140
rect 57230 -13245 57264 -13194
rect 57131 -13279 57264 -13245
rect 57319 -13254 57355 -13180
rect 57131 -13300 57165 -13279
rect 56316 -13318 56412 -13304
rect 54830 -13848 55830 -13838
rect 54830 -13870 55030 -13848
rect 53756 -13904 53852 -13870
rect 54808 -13904 55030 -13870
rect 53510 -13958 53526 -13924
rect 53614 -13958 53630 -13924
rect 53756 -13966 53790 -13904
rect 54830 -13928 55030 -13904
rect 55110 -13868 55740 -13848
rect 55810 -13868 55830 -13848
rect 56112 -13868 56146 -13806
rect 55110 -13908 55160 -13868
rect 55600 -13908 55740 -13868
rect 56050 -13902 56146 -13868
rect 55110 -13928 55740 -13908
rect 55810 -13928 55830 -13902
rect 54830 -13938 55830 -13928
rect 53464 -14008 53498 -13992
rect 53464 -14800 53498 -14784
rect 53642 -14008 53676 -13992
rect 53642 -14800 53676 -14784
rect 54870 -13966 54904 -13938
rect 53926 -14018 53942 -13984
rect 54718 -14018 54734 -13984
rect 53858 -14046 53892 -14030
rect 53858 -14150 53892 -14134
rect 54768 -14046 54802 -14030
rect 54768 -14150 54802 -14134
rect 53926 -14196 53942 -14162
rect 54718 -14196 54734 -14162
rect 53756 -14276 53790 -14214
rect 55700 -13964 55740 -13938
rect 55126 -14130 55142 -14096
rect 55494 -14130 55510 -14096
rect 54870 -14276 54904 -14214
rect 55046 -14182 55080 -14166
rect 55046 -14232 55080 -14216
rect 55556 -14182 55590 -14166
rect 55556 -14232 55590 -14216
rect 53756 -14310 53852 -14276
rect 54808 -14310 54904 -14276
rect 55126 -14302 55142 -14268
rect 55494 -14302 55510 -14268
rect 53510 -14868 53526 -14834
rect 53614 -14868 53630 -14834
rect 53350 -14936 53384 -14874
rect 53756 -14936 53790 -14310
rect 54870 -14418 54904 -14310
rect 55700 -14418 55706 -13964
rect 54870 -14424 55706 -14418
rect 54870 -14458 55262 -14424
rect 55420 -14458 55706 -14424
rect 55166 -14520 55200 -14458
rect 53350 -14970 53446 -14936
rect 53694 -14970 53790 -14936
rect 53886 -14708 53982 -14674
rect 54956 -14708 55052 -14674
rect 53886 -14770 53920 -14708
rect 55018 -14770 55052 -14708
rect 54065 -14822 54081 -14788
rect 54857 -14822 54873 -14788
rect 53988 -14850 54022 -14834
rect 53988 -14904 54022 -14888
rect 54916 -14850 54950 -14834
rect 54916 -14904 54950 -14888
rect 54065 -14950 54081 -14916
rect 54857 -14950 54873 -14916
rect 53886 -15030 53920 -14968
rect 55482 -14520 55516 -14458
rect 55280 -14548 55314 -14532
rect 55280 -14740 55314 -14724
rect 55368 -14548 55402 -14532
rect 55368 -14740 55402 -14724
rect 55308 -14808 55324 -14774
rect 55358 -14808 55374 -14774
rect 55166 -14876 55200 -14814
rect 55482 -14876 55516 -14814
rect 55166 -14910 55262 -14876
rect 55420 -14910 55516 -14876
rect 55018 -15030 55052 -14968
rect 56112 -13964 56146 -13902
rect 56350 -13338 56412 -13318
rect 56610 -13338 56706 -13304
rect 56672 -13400 56706 -13338
rect 57303 -13283 57355 -13254
rect 57131 -13355 57165 -13334
rect 57201 -13347 57217 -13313
rect 57251 -13347 57267 -13313
rect 57201 -13389 57267 -13347
rect 57337 -13317 57355 -13283
rect 57303 -13355 57355 -13317
rect 58930 -13210 59026 -13176
rect 59214 -13177 59310 -13176
rect 59662 -13177 59696 -13120
rect 59772 -13094 59866 -13060
rect 60426 -13094 60520 -13060
rect 59772 -13150 59806 -13094
rect 59214 -13210 59696 -13177
rect 58930 -13211 59696 -13210
rect 58930 -13272 58964 -13211
rect 59276 -13272 59310 -13211
rect 59087 -13312 59103 -13278
rect 59137 -13312 59153 -13278
rect 56476 -13440 56492 -13406
rect 56530 -13440 56546 -13406
rect 55866 -14004 55882 -13970
rect 55970 -14004 55986 -13970
rect 55820 -14054 55854 -14038
rect 55820 -14846 55854 -14830
rect 55998 -14054 56032 -14038
rect 55998 -14846 56032 -14830
rect 55866 -14914 55882 -14880
rect 55970 -14914 55986 -14880
rect 55706 -14982 55740 -14920
rect 56430 -13499 56464 -13483
rect 56430 -14291 56464 -14275
rect 56558 -13499 56592 -13483
rect 56558 -14291 56592 -14275
rect 56476 -14368 56492 -14334
rect 56530 -14368 56546 -14334
rect 56316 -14436 56350 -14374
rect 57096 -13423 57125 -13389
rect 57159 -13423 57217 -13389
rect 57251 -13423 57309 -13389
rect 57343 -13423 57372 -13389
rect 59044 -13371 59078 -13355
rect 59044 -13763 59078 -13747
rect 59162 -13371 59196 -13355
rect 59162 -13763 59196 -13747
rect 59087 -13840 59103 -13806
rect 59137 -13840 59153 -13806
rect 60486 -13156 60520 -13094
rect 59942 -13208 59958 -13174
rect 60334 -13208 60350 -13174
rect 59874 -13228 59908 -13212
rect 59874 -13278 59908 -13262
rect 60384 -13228 60418 -13212
rect 60384 -13278 60418 -13262
rect 59942 -13316 59958 -13282
rect 60334 -13316 60350 -13282
rect 59772 -13396 59806 -13340
rect 60486 -13396 60520 -13334
rect 59388 -13430 59476 -13396
rect 59656 -13430 59800 -13396
rect 59958 -13430 60520 -13396
rect 59388 -13490 59422 -13430
rect 59276 -13906 59310 -13846
rect 59530 -13532 59546 -13498
rect 59580 -13532 59596 -13498
rect 59502 -13582 59536 -13566
rect 59502 -13774 59536 -13758
rect 59590 -13582 59624 -13566
rect 59590 -13774 59624 -13758
rect 59530 -13842 59546 -13808
rect 59580 -13842 59596 -13808
rect 58966 -13942 59310 -13906
rect 59388 -13909 59422 -13850
rect 59704 -13909 59738 -13430
rect 60020 -13492 60054 -13430
rect 59846 -13532 59862 -13498
rect 59896 -13532 59912 -13498
rect 59818 -13582 59852 -13566
rect 59818 -13774 59852 -13758
rect 59906 -13582 59940 -13566
rect 59906 -13774 59940 -13758
rect 59846 -13842 59862 -13808
rect 59896 -13842 59912 -13808
rect 61186 -13600 61286 -13590
rect 61186 -13680 61196 -13600
rect 61186 -13690 61286 -13680
rect 60020 -13909 60054 -13848
rect 56672 -14436 56706 -14374
rect 57096 -14399 57125 -14365
rect 57159 -14399 57217 -14365
rect 57251 -14399 57309 -14365
rect 57343 -14399 57372 -14365
rect 56316 -14470 56412 -14436
rect 56610 -14470 56706 -14436
rect 57131 -14454 57165 -14433
rect 57201 -14441 57267 -14399
rect 57201 -14475 57217 -14441
rect 57251 -14475 57267 -14441
rect 57303 -14471 57355 -14433
rect 57131 -14509 57165 -14488
rect 57337 -14505 57355 -14471
rect 59276 -14002 59310 -13942
rect 59387 -13944 60054 -13909
rect 60127 -13754 60161 -13728
rect 60127 -13757 60253 -13754
rect 60161 -13773 60253 -13757
rect 60161 -13791 60203 -13773
rect 60127 -13807 60203 -13791
rect 60237 -13807 60253 -13773
rect 60359 -13760 60409 -13749
rect 60671 -13754 60705 -13728
rect 60359 -13765 60366 -13760
rect 60359 -13800 60366 -13799
rect 60406 -13800 60409 -13760
rect 60127 -13849 60161 -13807
rect 60127 -13941 60161 -13883
rect 60195 -13857 60325 -13841
rect 60195 -13891 60211 -13857
rect 60245 -13891 60325 -13857
rect 60195 -13907 60325 -13891
rect 59387 -14000 59421 -13944
rect 59087 -14042 59103 -14008
rect 59137 -14042 59153 -14008
rect 59044 -14101 59078 -14085
rect 57131 -14543 57264 -14509
rect 57303 -14534 57355 -14505
rect 57117 -14594 57185 -14579
rect 57117 -14644 57118 -14594
rect 57168 -14644 57185 -14594
rect 57117 -14653 57185 -14644
rect 57230 -14594 57264 -14543
rect 57319 -14570 57355 -14534
rect 57230 -14610 57285 -14594
rect 57230 -14644 57251 -14610
rect 57230 -14660 57285 -14644
rect 57319 -14610 57326 -14570
rect 59044 -14493 59078 -14477
rect 59162 -14101 59196 -14085
rect 59162 -14493 59196 -14477
rect 59087 -14570 59103 -14536
rect 59137 -14570 59153 -14536
rect 57230 -14689 57264 -14660
rect 57129 -14723 57264 -14689
rect 57319 -14694 57355 -14610
rect 57129 -14757 57165 -14723
rect 57301 -14744 57355 -14694
rect 58930 -14638 58964 -14576
rect 59529 -14045 59545 -14011
rect 59579 -14045 59595 -14011
rect 59501 -14095 59535 -14079
rect 59501 -14287 59535 -14271
rect 59589 -14095 59623 -14079
rect 59589 -14287 59623 -14271
rect 59529 -14355 59545 -14321
rect 59579 -14355 59595 -14321
rect 59387 -14423 59421 -14370
rect 59703 -14423 59737 -13944
rect 60019 -14005 60053 -13944
rect 59845 -14045 59861 -14011
rect 59895 -14045 59911 -14011
rect 59817 -14095 59851 -14079
rect 59817 -14287 59851 -14271
rect 59905 -14095 59939 -14079
rect 59905 -14287 59939 -14271
rect 59845 -14355 59861 -14321
rect 59895 -14355 59911 -14321
rect 60161 -13975 60203 -13941
rect 60237 -13975 60253 -13941
rect 60127 -14033 60161 -13975
rect 60289 -14009 60325 -13907
rect 60127 -14109 60161 -14067
rect 60195 -14025 60325 -14009
rect 60195 -14059 60211 -14025
rect 60245 -14059 60325 -14025
rect 60195 -14075 60325 -14059
rect 60359 -13850 60409 -13800
rect 60443 -13757 60705 -13754
rect 60443 -13773 60671 -13757
rect 60443 -13807 60459 -13773
rect 60493 -13807 60527 -13773
rect 60561 -13807 60595 -13773
rect 60629 -13791 60671 -13773
rect 60629 -13807 60705 -13791
rect 60359 -13857 60366 -13850
rect 60406 -13890 60409 -13850
rect 60393 -13891 60409 -13890
rect 60359 -13940 60409 -13891
rect 60359 -13941 60366 -13940
rect 60359 -13980 60366 -13975
rect 60406 -13980 60409 -13940
rect 60359 -14020 60409 -13980
rect 60359 -14025 60366 -14020
rect 60359 -14060 60366 -14059
rect 60406 -14060 60409 -14020
rect 60359 -14075 60409 -14060
rect 60443 -13857 60637 -13841
rect 60443 -13891 60459 -13857
rect 60493 -13891 60527 -13857
rect 60561 -13891 60595 -13857
rect 60629 -13891 60637 -13857
rect 60443 -13907 60637 -13891
rect 60671 -13849 60705 -13807
rect 60443 -14009 60477 -13907
rect 60671 -13941 60705 -13883
rect 60511 -13975 60527 -13941
rect 60561 -13975 60595 -13941
rect 60629 -13975 60671 -13941
rect 60443 -14025 60637 -14009
rect 60443 -14059 60459 -14025
rect 60493 -14059 60527 -14025
rect 60561 -14059 60595 -14025
rect 60629 -14059 60637 -14025
rect 60443 -14075 60637 -14059
rect 60671 -14033 60705 -13975
rect 60289 -14109 60325 -14075
rect 60443 -14109 60481 -14075
rect 60671 -14109 60705 -14067
rect 60127 -14125 60204 -14109
rect 60161 -14143 60204 -14125
rect 60238 -14143 60254 -14109
rect 60161 -14159 60254 -14143
rect 60289 -14125 60481 -14109
rect 60289 -14159 60297 -14125
rect 60331 -14159 60369 -14125
rect 60405 -14159 60449 -14125
rect 60579 -14143 60595 -14109
rect 60629 -14125 60705 -14109
rect 60629 -14143 60671 -14125
rect 60579 -14151 60671 -14143
rect 60127 -14188 60161 -14159
rect 60289 -14162 60481 -14159
rect 60671 -14188 60705 -14159
rect 60747 -13754 60781 -13728
rect 60747 -13757 61009 -13754
rect 60781 -13773 61009 -13757
rect 60781 -13791 60823 -13773
rect 60747 -13807 60823 -13791
rect 60857 -13807 60891 -13773
rect 60925 -13807 60959 -13773
rect 60993 -13807 61009 -13773
rect 61043 -13760 61093 -13749
rect 61291 -13754 61325 -13728
rect 61043 -13800 61046 -13760
rect 61086 -13765 61093 -13760
rect 61086 -13800 61093 -13799
rect 60747 -13849 60781 -13807
rect 60747 -13941 60781 -13883
rect 60815 -13857 61009 -13841
rect 60815 -13891 60823 -13857
rect 60857 -13891 60891 -13857
rect 60925 -13891 60959 -13857
rect 60993 -13891 61009 -13857
rect 60815 -13907 61009 -13891
rect 60781 -13975 60823 -13941
rect 60857 -13975 60891 -13941
rect 60925 -13975 60941 -13941
rect 60747 -14033 60781 -13975
rect 60975 -14009 61009 -13907
rect 60747 -14109 60781 -14067
rect 60815 -14025 61009 -14009
rect 60815 -14059 60823 -14025
rect 60857 -14059 60891 -14025
rect 60925 -14059 60959 -14025
rect 60993 -14059 61009 -14025
rect 60815 -14075 61009 -14059
rect 61043 -13850 61093 -13800
rect 61199 -13757 61325 -13754
rect 61199 -13773 61291 -13757
rect 61199 -13807 61215 -13773
rect 61249 -13791 61291 -13773
rect 61249 -13807 61325 -13791
rect 61043 -13890 61046 -13850
rect 61086 -13857 61093 -13850
rect 61043 -13891 61059 -13890
rect 61043 -13940 61093 -13891
rect 61043 -13980 61046 -13940
rect 61086 -13941 61093 -13940
rect 61086 -13980 61093 -13975
rect 61043 -14020 61093 -13980
rect 61043 -14060 61046 -14020
rect 61086 -14025 61093 -14020
rect 61086 -14060 61093 -14059
rect 61043 -14075 61093 -14060
rect 61127 -13857 61257 -13841
rect 61127 -13891 61207 -13857
rect 61241 -13891 61257 -13857
rect 61127 -13907 61257 -13891
rect 61291 -13849 61325 -13807
rect 61127 -14009 61163 -13907
rect 61291 -13941 61325 -13883
rect 61199 -13975 61215 -13941
rect 61249 -13975 61291 -13941
rect 61127 -14025 61257 -14009
rect 61127 -14059 61207 -14025
rect 61241 -14059 61257 -14025
rect 61127 -14075 61257 -14059
rect 61291 -14033 61325 -13975
rect 60971 -14109 61009 -14075
rect 61127 -14109 61163 -14075
rect 61291 -14109 61325 -14067
rect 60747 -14125 60823 -14109
rect 60781 -14143 60823 -14125
rect 60857 -14143 60873 -14109
rect 60781 -14151 60873 -14143
rect 60971 -14124 61163 -14109
rect 60971 -14125 61129 -14124
rect 60747 -14188 60781 -14159
rect 60971 -14159 60980 -14125
rect 61015 -14159 61053 -14125
rect 61088 -14158 61129 -14125
rect 61198 -14143 61214 -14109
rect 61248 -14125 61325 -14109
rect 61248 -14143 61291 -14125
rect 61088 -14159 61163 -14158
rect 61198 -14159 61291 -14143
rect 60971 -14162 61163 -14159
rect 61291 -14188 61325 -14159
rect 60466 -14260 60546 -14240
rect 60466 -14300 60486 -14260
rect 60526 -14300 60546 -14260
rect 60466 -14320 60546 -14300
rect 60606 -14260 60686 -14240
rect 60606 -14300 60626 -14260
rect 60666 -14300 60686 -14260
rect 60606 -14320 60686 -14300
rect 60746 -14260 60826 -14240
rect 60746 -14300 60766 -14260
rect 60806 -14300 60826 -14260
rect 60746 -14320 60826 -14300
rect 60886 -14260 60966 -14240
rect 60886 -14300 60906 -14260
rect 60946 -14300 60966 -14260
rect 60886 -14320 60966 -14300
rect 60019 -14423 60053 -14361
rect 59387 -14457 59476 -14423
rect 59646 -14457 59799 -14423
rect 59957 -14426 60053 -14423
rect 59957 -14457 60520 -14426
rect 59772 -14460 60520 -14457
rect 59772 -14520 59806 -14460
rect 59276 -14638 59310 -14576
rect 58930 -14672 59026 -14638
rect 59214 -14640 59310 -14638
rect 59214 -14672 59696 -14640
rect 58930 -14674 59696 -14672
rect 58930 -14710 58964 -14674
rect 57129 -14791 57131 -14757
rect 57129 -14825 57165 -14791
rect 57129 -14859 57131 -14825
rect 57129 -14875 57165 -14859
rect 57201 -14791 57217 -14757
rect 57251 -14791 57267 -14757
rect 57201 -14825 57267 -14791
rect 57201 -14859 57217 -14825
rect 57251 -14859 57267 -14825
rect 57201 -14909 57267 -14859
rect 57301 -14778 57303 -14744
rect 57337 -14778 57355 -14744
rect 57301 -14825 57355 -14778
rect 57301 -14859 57303 -14825
rect 57337 -14859 57355 -14825
rect 57301 -14875 57355 -14859
rect 59662 -14730 59696 -14674
rect 60486 -14522 60520 -14460
rect 59942 -14574 59958 -14540
rect 60334 -14574 60350 -14540
rect 59874 -14594 59908 -14578
rect 59874 -14644 59908 -14628
rect 60384 -14594 60418 -14578
rect 60384 -14644 60418 -14628
rect 59942 -14682 59958 -14648
rect 60334 -14682 60350 -14648
rect 56112 -14982 56146 -14920
rect 57096 -14943 57125 -14909
rect 57159 -14943 57217 -14909
rect 57251 -14943 57309 -14909
rect 57343 -14943 57372 -14909
rect 55706 -15016 55802 -14982
rect 56050 -15016 56146 -14982
rect 53886 -15064 53982 -15030
rect 54956 -15064 55052 -15030
rect 53886 -15126 53920 -15064
rect 55018 -15126 55052 -15064
rect 55720 -15058 56090 -15016
rect 55720 -15068 56020 -15058
rect 54065 -15178 54081 -15144
rect 54857 -15178 54873 -15144
rect 53988 -15206 54022 -15190
rect 53988 -15260 54022 -15244
rect 54916 -15206 54950 -15190
rect 54916 -15260 54950 -15244
rect 54065 -15306 54081 -15272
rect 54857 -15306 54873 -15272
rect 53886 -15386 53920 -15324
rect 56010 -15208 56020 -15068
rect 56080 -15208 56090 -15058
rect 59109 -14788 59125 -14754
rect 59501 -14788 59517 -14754
rect 59560 -14808 59594 -14792
rect 59560 -14858 59594 -14842
rect 59109 -14896 59125 -14862
rect 59501 -14896 59517 -14862
rect 59032 -14916 59066 -14900
rect 59032 -14966 59066 -14950
rect 59109 -15004 59125 -14970
rect 59501 -15004 59517 -14970
rect 56010 -15218 56090 -15208
rect 59772 -14762 59806 -14700
rect 60486 -14762 60520 -14700
rect 59772 -14796 59866 -14762
rect 60426 -14796 60520 -14762
rect 59662 -15084 59696 -15030
rect 58966 -15100 59026 -15084
rect 58930 -15118 59026 -15100
rect 59600 -15118 59696 -15084
rect 55018 -15386 55052 -15324
rect 53886 -15420 53982 -15386
rect 54956 -15420 55052 -15386
rect 55176 -15278 55272 -15244
rect 55566 -15278 55662 -15244
rect 55176 -15340 55210 -15278
rect 55628 -15340 55662 -15278
rect 55284 -15392 55300 -15358
rect 55476 -15392 55492 -15358
rect 55526 -15402 55560 -15386
rect 55284 -15480 55300 -15446
rect 55476 -15480 55492 -15446
rect 55526 -15452 55560 -15436
rect 55176 -15560 55210 -15498
rect 55628 -15560 55662 -15498
rect 55176 -15594 55272 -15560
rect 55566 -15594 55662 -15560
rect 53896 -17792 53992 -17758
rect 54966 -17792 55062 -17758
rect 53896 -17854 53930 -17792
rect 55028 -17854 55062 -17792
rect 54075 -17906 54091 -17872
rect 54867 -17906 54883 -17872
rect 53998 -17934 54032 -17918
rect 53998 -17988 54032 -17972
rect 54926 -17934 54960 -17918
rect 54926 -17988 54960 -17972
rect 54075 -18034 54091 -18000
rect 54867 -18034 54883 -18000
rect 53896 -18114 53930 -18052
rect 55028 -18114 55062 -18052
rect 55960 -18108 56040 -18098
rect 53896 -18148 53992 -18114
rect 54966 -18148 55062 -18114
rect 53350 -18238 53790 -18204
rect 53350 -18300 53384 -18238
rect 53510 -18340 53526 -18306
rect 53614 -18340 53630 -18306
rect 53464 -18390 53498 -18374
rect 53464 -19182 53498 -19166
rect 53642 -18390 53676 -18374
rect 53642 -19182 53676 -19166
rect 53756 -18864 53790 -18238
rect 53896 -18210 53930 -18148
rect 55028 -18210 55062 -18148
rect 55710 -18154 56040 -18108
rect 54075 -18262 54091 -18228
rect 54867 -18262 54883 -18228
rect 53998 -18290 54032 -18274
rect 53998 -18344 54032 -18328
rect 54926 -18290 54960 -18274
rect 54926 -18344 54960 -18328
rect 54075 -18390 54091 -18356
rect 54867 -18390 54883 -18356
rect 53896 -18470 53930 -18408
rect 55706 -18188 55802 -18154
rect 56050 -18188 56146 -18154
rect 55706 -18250 55740 -18188
rect 55028 -18470 55062 -18408
rect 53896 -18504 53992 -18470
rect 54966 -18504 55062 -18470
rect 55176 -18300 55272 -18266
rect 55430 -18300 55526 -18266
rect 55176 -18362 55210 -18300
rect 55492 -18362 55526 -18300
rect 55318 -18402 55334 -18368
rect 55368 -18402 55384 -18368
rect 55290 -18452 55324 -18436
rect 55290 -18644 55324 -18628
rect 55378 -18452 55412 -18436
rect 55378 -18644 55412 -18628
rect 55176 -18718 55210 -18656
rect 55492 -18718 55526 -18656
rect 54870 -18752 55272 -18718
rect 55430 -18752 55706 -18718
rect 54870 -18758 55706 -18752
rect 54870 -18864 54904 -18758
rect 53756 -18898 53852 -18864
rect 54808 -18898 54904 -18864
rect 53756 -18960 53790 -18898
rect 54870 -18960 54904 -18898
rect 55126 -18908 55142 -18874
rect 55494 -18908 55510 -18874
rect 53926 -19012 53942 -18978
rect 54718 -19012 54734 -18978
rect 53858 -19040 53892 -19024
rect 53858 -19144 53892 -19128
rect 54768 -19040 54802 -19024
rect 54768 -19144 54802 -19128
rect 53926 -19190 53942 -19156
rect 54718 -19190 54734 -19156
rect 53510 -19250 53526 -19216
rect 53614 -19250 53630 -19216
rect 53756 -19270 53790 -19208
rect 55046 -18960 55080 -18944
rect 55046 -19010 55080 -18994
rect 55556 -18960 55590 -18944
rect 55556 -19010 55590 -18994
rect 55126 -19080 55142 -19046
rect 55494 -19080 55510 -19046
rect 54870 -19238 54904 -19208
rect 55700 -19206 55706 -18758
rect 56112 -18250 56146 -18188
rect 58930 -18167 59026 -18133
rect 59600 -18167 59696 -18133
rect 58930 -18210 58964 -18167
rect 58926 -18220 58966 -18210
rect 55866 -18290 55882 -18256
rect 55970 -18290 55986 -18256
rect 55820 -18340 55854 -18324
rect 55820 -19132 55854 -19116
rect 55998 -18340 56032 -18324
rect 55998 -19132 56032 -19116
rect 55866 -19200 55882 -19166
rect 55970 -19200 55986 -19166
rect 55700 -19238 55740 -19206
rect 57096 -18279 57125 -18245
rect 57159 -18279 57217 -18245
rect 57251 -18279 57309 -18245
rect 57343 -18279 57372 -18245
rect 57129 -18329 57165 -18313
rect 57129 -18363 57131 -18329
rect 57129 -18397 57165 -18363
rect 57129 -18431 57131 -18397
rect 57201 -18329 57267 -18279
rect 57201 -18363 57217 -18329
rect 57251 -18363 57267 -18329
rect 57201 -18397 57267 -18363
rect 57201 -18431 57217 -18397
rect 57251 -18431 57267 -18397
rect 57301 -18329 57355 -18313
rect 57301 -18363 57303 -18329
rect 57337 -18363 57355 -18329
rect 57301 -18410 57355 -18363
rect 57129 -18465 57165 -18431
rect 57301 -18444 57303 -18410
rect 57337 -18444 57355 -18410
rect 57129 -18499 57264 -18465
rect 57301 -18494 57355 -18444
rect 57230 -18528 57264 -18499
rect 57117 -18544 57185 -18535
rect 57117 -18594 57118 -18544
rect 57178 -18594 57185 -18544
rect 57117 -18609 57185 -18594
rect 57230 -18544 57285 -18528
rect 57230 -18578 57251 -18544
rect 57230 -18594 57285 -18578
rect 57319 -18540 57355 -18494
rect 59662 -18229 59696 -18167
rect 59109 -18281 59125 -18247
rect 59501 -18281 59517 -18247
rect 59560 -18301 59594 -18285
rect 59560 -18351 59594 -18335
rect 59109 -18389 59125 -18355
rect 59501 -18389 59517 -18355
rect 59032 -18409 59066 -18393
rect 59032 -18459 59066 -18443
rect 59109 -18497 59125 -18463
rect 59501 -18497 59517 -18463
rect 58926 -18540 58966 -18520
rect 57319 -18580 57326 -18540
rect 58930 -18576 58964 -18540
rect 57230 -18645 57264 -18594
rect 57131 -18679 57264 -18645
rect 57319 -18654 57355 -18580
rect 57131 -18700 57165 -18679
rect 56316 -18718 56412 -18704
rect 54830 -19248 55830 -19238
rect 54830 -19270 55030 -19248
rect 53756 -19304 53852 -19270
rect 54808 -19304 55030 -19270
rect 53510 -19358 53526 -19324
rect 53614 -19358 53630 -19324
rect 53756 -19366 53790 -19304
rect 54830 -19328 55030 -19304
rect 55110 -19268 55740 -19248
rect 55810 -19268 55830 -19248
rect 56112 -19268 56146 -19206
rect 55110 -19308 55160 -19268
rect 55600 -19308 55740 -19268
rect 56050 -19302 56146 -19268
rect 55110 -19328 55740 -19308
rect 55810 -19328 55830 -19302
rect 54830 -19338 55830 -19328
rect 53464 -19408 53498 -19392
rect 53464 -20200 53498 -20184
rect 53642 -19408 53676 -19392
rect 53642 -20200 53676 -20184
rect 54870 -19366 54904 -19338
rect 53926 -19418 53942 -19384
rect 54718 -19418 54734 -19384
rect 53858 -19446 53892 -19430
rect 53858 -19550 53892 -19534
rect 54768 -19446 54802 -19430
rect 54768 -19550 54802 -19534
rect 53926 -19596 53942 -19562
rect 54718 -19596 54734 -19562
rect 53756 -19676 53790 -19614
rect 55700 -19364 55740 -19338
rect 55126 -19530 55142 -19496
rect 55494 -19530 55510 -19496
rect 54870 -19676 54904 -19614
rect 55046 -19582 55080 -19566
rect 55046 -19632 55080 -19616
rect 55556 -19582 55590 -19566
rect 55556 -19632 55590 -19616
rect 53756 -19710 53852 -19676
rect 54808 -19710 54904 -19676
rect 55126 -19702 55142 -19668
rect 55494 -19702 55510 -19668
rect 53510 -20268 53526 -20234
rect 53614 -20268 53630 -20234
rect 53350 -20336 53384 -20274
rect 53756 -20336 53790 -19710
rect 54870 -19818 54904 -19710
rect 55700 -19818 55706 -19364
rect 54870 -19824 55706 -19818
rect 54870 -19858 55262 -19824
rect 55420 -19858 55706 -19824
rect 55166 -19920 55200 -19858
rect 53350 -20370 53446 -20336
rect 53694 -20370 53790 -20336
rect 53886 -20108 53982 -20074
rect 54956 -20108 55052 -20074
rect 53886 -20170 53920 -20108
rect 55018 -20170 55052 -20108
rect 54065 -20222 54081 -20188
rect 54857 -20222 54873 -20188
rect 53988 -20250 54022 -20234
rect 53988 -20304 54022 -20288
rect 54916 -20250 54950 -20234
rect 54916 -20304 54950 -20288
rect 54065 -20350 54081 -20316
rect 54857 -20350 54873 -20316
rect 53886 -20430 53920 -20368
rect 55482 -19920 55516 -19858
rect 55280 -19948 55314 -19932
rect 55280 -20140 55314 -20124
rect 55368 -19948 55402 -19932
rect 55368 -20140 55402 -20124
rect 55308 -20208 55324 -20174
rect 55358 -20208 55374 -20174
rect 55166 -20276 55200 -20214
rect 55482 -20276 55516 -20214
rect 55166 -20310 55262 -20276
rect 55420 -20310 55516 -20276
rect 55018 -20430 55052 -20368
rect 56112 -19364 56146 -19302
rect 56350 -18738 56412 -18718
rect 56610 -18738 56706 -18704
rect 56672 -18800 56706 -18738
rect 57303 -18683 57355 -18654
rect 57131 -18755 57165 -18734
rect 57201 -18747 57217 -18713
rect 57251 -18747 57267 -18713
rect 57201 -18789 57267 -18747
rect 57337 -18717 57355 -18683
rect 57303 -18755 57355 -18717
rect 58930 -18610 59026 -18576
rect 59214 -18577 59310 -18576
rect 59662 -18577 59696 -18520
rect 59772 -18494 59866 -18460
rect 60426 -18494 60520 -18460
rect 59772 -18550 59806 -18494
rect 59214 -18610 59696 -18577
rect 58930 -18611 59696 -18610
rect 58930 -18672 58964 -18611
rect 59276 -18672 59310 -18611
rect 59087 -18712 59103 -18678
rect 59137 -18712 59153 -18678
rect 56476 -18840 56492 -18806
rect 56530 -18840 56546 -18806
rect 55866 -19404 55882 -19370
rect 55970 -19404 55986 -19370
rect 55820 -19454 55854 -19438
rect 55820 -20246 55854 -20230
rect 55998 -19454 56032 -19438
rect 55998 -20246 56032 -20230
rect 55866 -20314 55882 -20280
rect 55970 -20314 55986 -20280
rect 55706 -20382 55740 -20320
rect 56430 -18899 56464 -18883
rect 56430 -19691 56464 -19675
rect 56558 -18899 56592 -18883
rect 56558 -19691 56592 -19675
rect 56476 -19768 56492 -19734
rect 56530 -19768 56546 -19734
rect 56316 -19836 56350 -19774
rect 57096 -18823 57125 -18789
rect 57159 -18823 57217 -18789
rect 57251 -18823 57309 -18789
rect 57343 -18823 57372 -18789
rect 59044 -18771 59078 -18755
rect 59044 -19163 59078 -19147
rect 59162 -18771 59196 -18755
rect 59162 -19163 59196 -19147
rect 59087 -19240 59103 -19206
rect 59137 -19240 59153 -19206
rect 60486 -18556 60520 -18494
rect 59942 -18608 59958 -18574
rect 60334 -18608 60350 -18574
rect 59874 -18628 59908 -18612
rect 59874 -18678 59908 -18662
rect 60384 -18628 60418 -18612
rect 60384 -18678 60418 -18662
rect 59942 -18716 59958 -18682
rect 60334 -18716 60350 -18682
rect 59772 -18796 59806 -18740
rect 60486 -18796 60520 -18734
rect 59388 -18830 59476 -18796
rect 59656 -18830 59800 -18796
rect 59958 -18830 60520 -18796
rect 59388 -18890 59422 -18830
rect 59276 -19306 59310 -19246
rect 59530 -18932 59546 -18898
rect 59580 -18932 59596 -18898
rect 59502 -18982 59536 -18966
rect 59502 -19174 59536 -19158
rect 59590 -18982 59624 -18966
rect 59590 -19174 59624 -19158
rect 59530 -19242 59546 -19208
rect 59580 -19242 59596 -19208
rect 58966 -19342 59310 -19306
rect 59388 -19309 59422 -19250
rect 59704 -19309 59738 -18830
rect 60020 -18892 60054 -18830
rect 59846 -18932 59862 -18898
rect 59896 -18932 59912 -18898
rect 59818 -18982 59852 -18966
rect 59818 -19174 59852 -19158
rect 59906 -18982 59940 -18966
rect 59906 -19174 59940 -19158
rect 59846 -19242 59862 -19208
rect 59896 -19242 59912 -19208
rect 61186 -19000 61286 -18990
rect 61186 -19080 61196 -19000
rect 61186 -19090 61286 -19080
rect 60020 -19309 60054 -19248
rect 56672 -19836 56706 -19774
rect 57096 -19799 57125 -19765
rect 57159 -19799 57217 -19765
rect 57251 -19799 57309 -19765
rect 57343 -19799 57372 -19765
rect 56316 -19870 56412 -19836
rect 56610 -19870 56706 -19836
rect 57131 -19854 57165 -19833
rect 57201 -19841 57267 -19799
rect 57201 -19875 57217 -19841
rect 57251 -19875 57267 -19841
rect 57303 -19871 57355 -19833
rect 57131 -19909 57165 -19888
rect 57337 -19905 57355 -19871
rect 59276 -19402 59310 -19342
rect 59387 -19344 60054 -19309
rect 60127 -19154 60161 -19128
rect 60127 -19157 60253 -19154
rect 60161 -19173 60253 -19157
rect 60161 -19191 60203 -19173
rect 60127 -19207 60203 -19191
rect 60237 -19207 60253 -19173
rect 60359 -19160 60409 -19149
rect 60671 -19154 60705 -19128
rect 60359 -19165 60366 -19160
rect 60359 -19200 60366 -19199
rect 60406 -19200 60409 -19160
rect 60127 -19249 60161 -19207
rect 60127 -19341 60161 -19283
rect 60195 -19257 60325 -19241
rect 60195 -19291 60211 -19257
rect 60245 -19291 60325 -19257
rect 60195 -19307 60325 -19291
rect 59387 -19400 59421 -19344
rect 59087 -19442 59103 -19408
rect 59137 -19442 59153 -19408
rect 59044 -19501 59078 -19485
rect 57131 -19943 57264 -19909
rect 57303 -19934 57355 -19905
rect 57117 -19994 57185 -19979
rect 57117 -20044 57118 -19994
rect 57168 -20044 57185 -19994
rect 57117 -20053 57185 -20044
rect 57230 -19994 57264 -19943
rect 57319 -19970 57355 -19934
rect 57230 -20010 57285 -19994
rect 57230 -20044 57251 -20010
rect 57230 -20060 57285 -20044
rect 57319 -20010 57326 -19970
rect 59044 -19893 59078 -19877
rect 59162 -19501 59196 -19485
rect 59162 -19893 59196 -19877
rect 59087 -19970 59103 -19936
rect 59137 -19970 59153 -19936
rect 57230 -20089 57264 -20060
rect 57129 -20123 57264 -20089
rect 57319 -20094 57355 -20010
rect 57129 -20157 57165 -20123
rect 57301 -20144 57355 -20094
rect 58930 -20038 58964 -19976
rect 59529 -19445 59545 -19411
rect 59579 -19445 59595 -19411
rect 59501 -19495 59535 -19479
rect 59501 -19687 59535 -19671
rect 59589 -19495 59623 -19479
rect 59589 -19687 59623 -19671
rect 59529 -19755 59545 -19721
rect 59579 -19755 59595 -19721
rect 59387 -19823 59421 -19770
rect 59703 -19823 59737 -19344
rect 60019 -19405 60053 -19344
rect 59845 -19445 59861 -19411
rect 59895 -19445 59911 -19411
rect 59817 -19495 59851 -19479
rect 59817 -19687 59851 -19671
rect 59905 -19495 59939 -19479
rect 59905 -19687 59939 -19671
rect 59845 -19755 59861 -19721
rect 59895 -19755 59911 -19721
rect 60161 -19375 60203 -19341
rect 60237 -19375 60253 -19341
rect 60127 -19433 60161 -19375
rect 60289 -19409 60325 -19307
rect 60127 -19509 60161 -19467
rect 60195 -19425 60325 -19409
rect 60195 -19459 60211 -19425
rect 60245 -19459 60325 -19425
rect 60195 -19475 60325 -19459
rect 60359 -19250 60409 -19200
rect 60443 -19157 60705 -19154
rect 60443 -19173 60671 -19157
rect 60443 -19207 60459 -19173
rect 60493 -19207 60527 -19173
rect 60561 -19207 60595 -19173
rect 60629 -19191 60671 -19173
rect 60629 -19207 60705 -19191
rect 60359 -19257 60366 -19250
rect 60406 -19290 60409 -19250
rect 60393 -19291 60409 -19290
rect 60359 -19340 60409 -19291
rect 60359 -19341 60366 -19340
rect 60359 -19380 60366 -19375
rect 60406 -19380 60409 -19340
rect 60359 -19420 60409 -19380
rect 60359 -19425 60366 -19420
rect 60359 -19460 60366 -19459
rect 60406 -19460 60409 -19420
rect 60359 -19475 60409 -19460
rect 60443 -19257 60637 -19241
rect 60443 -19291 60459 -19257
rect 60493 -19291 60527 -19257
rect 60561 -19291 60595 -19257
rect 60629 -19291 60637 -19257
rect 60443 -19307 60637 -19291
rect 60671 -19249 60705 -19207
rect 60443 -19409 60477 -19307
rect 60671 -19341 60705 -19283
rect 60511 -19375 60527 -19341
rect 60561 -19375 60595 -19341
rect 60629 -19375 60671 -19341
rect 60443 -19425 60637 -19409
rect 60443 -19459 60459 -19425
rect 60493 -19459 60527 -19425
rect 60561 -19459 60595 -19425
rect 60629 -19459 60637 -19425
rect 60443 -19475 60637 -19459
rect 60671 -19433 60705 -19375
rect 60289 -19509 60325 -19475
rect 60443 -19509 60481 -19475
rect 60671 -19509 60705 -19467
rect 60127 -19525 60204 -19509
rect 60161 -19543 60204 -19525
rect 60238 -19543 60254 -19509
rect 60161 -19559 60254 -19543
rect 60289 -19525 60481 -19509
rect 60289 -19559 60297 -19525
rect 60331 -19559 60369 -19525
rect 60405 -19559 60449 -19525
rect 60579 -19543 60595 -19509
rect 60629 -19525 60705 -19509
rect 60629 -19543 60671 -19525
rect 60579 -19551 60671 -19543
rect 60127 -19588 60161 -19559
rect 60289 -19562 60481 -19559
rect 60671 -19588 60705 -19559
rect 60747 -19154 60781 -19128
rect 60747 -19157 61009 -19154
rect 60781 -19173 61009 -19157
rect 60781 -19191 60823 -19173
rect 60747 -19207 60823 -19191
rect 60857 -19207 60891 -19173
rect 60925 -19207 60959 -19173
rect 60993 -19207 61009 -19173
rect 61043 -19160 61093 -19149
rect 61291 -19154 61325 -19128
rect 61043 -19200 61046 -19160
rect 61086 -19165 61093 -19160
rect 61086 -19200 61093 -19199
rect 60747 -19249 60781 -19207
rect 60747 -19341 60781 -19283
rect 60815 -19257 61009 -19241
rect 60815 -19291 60823 -19257
rect 60857 -19291 60891 -19257
rect 60925 -19291 60959 -19257
rect 60993 -19291 61009 -19257
rect 60815 -19307 61009 -19291
rect 60781 -19375 60823 -19341
rect 60857 -19375 60891 -19341
rect 60925 -19375 60941 -19341
rect 60747 -19433 60781 -19375
rect 60975 -19409 61009 -19307
rect 60747 -19509 60781 -19467
rect 60815 -19425 61009 -19409
rect 60815 -19459 60823 -19425
rect 60857 -19459 60891 -19425
rect 60925 -19459 60959 -19425
rect 60993 -19459 61009 -19425
rect 60815 -19475 61009 -19459
rect 61043 -19250 61093 -19200
rect 61199 -19157 61325 -19154
rect 61199 -19173 61291 -19157
rect 61199 -19207 61215 -19173
rect 61249 -19191 61291 -19173
rect 61249 -19207 61325 -19191
rect 61043 -19290 61046 -19250
rect 61086 -19257 61093 -19250
rect 61043 -19291 61059 -19290
rect 61043 -19340 61093 -19291
rect 61043 -19380 61046 -19340
rect 61086 -19341 61093 -19340
rect 61086 -19380 61093 -19375
rect 61043 -19420 61093 -19380
rect 61043 -19460 61046 -19420
rect 61086 -19425 61093 -19420
rect 61086 -19460 61093 -19459
rect 61043 -19475 61093 -19460
rect 61127 -19257 61257 -19241
rect 61127 -19291 61207 -19257
rect 61241 -19291 61257 -19257
rect 61127 -19307 61257 -19291
rect 61291 -19249 61325 -19207
rect 61127 -19409 61163 -19307
rect 61291 -19341 61325 -19283
rect 61199 -19375 61215 -19341
rect 61249 -19375 61291 -19341
rect 61127 -19425 61257 -19409
rect 61127 -19459 61207 -19425
rect 61241 -19459 61257 -19425
rect 61127 -19475 61257 -19459
rect 61291 -19433 61325 -19375
rect 60971 -19509 61009 -19475
rect 61127 -19509 61163 -19475
rect 61291 -19509 61325 -19467
rect 60747 -19525 60823 -19509
rect 60781 -19543 60823 -19525
rect 60857 -19543 60873 -19509
rect 60781 -19551 60873 -19543
rect 60971 -19524 61163 -19509
rect 60971 -19525 61129 -19524
rect 60747 -19588 60781 -19559
rect 60971 -19559 60980 -19525
rect 61015 -19559 61053 -19525
rect 61088 -19558 61129 -19525
rect 61198 -19543 61214 -19509
rect 61248 -19525 61325 -19509
rect 61248 -19543 61291 -19525
rect 61088 -19559 61163 -19558
rect 61198 -19559 61291 -19543
rect 60971 -19562 61163 -19559
rect 61291 -19588 61325 -19559
rect 60466 -19660 60546 -19640
rect 60466 -19700 60486 -19660
rect 60526 -19700 60546 -19660
rect 60466 -19720 60546 -19700
rect 60606 -19660 60686 -19640
rect 60606 -19700 60626 -19660
rect 60666 -19700 60686 -19660
rect 60606 -19720 60686 -19700
rect 60746 -19660 60826 -19640
rect 60746 -19700 60766 -19660
rect 60806 -19700 60826 -19660
rect 60746 -19720 60826 -19700
rect 60886 -19660 60966 -19640
rect 60886 -19700 60906 -19660
rect 60946 -19700 60966 -19660
rect 60886 -19720 60966 -19700
rect 60019 -19823 60053 -19761
rect 59387 -19857 59476 -19823
rect 59646 -19857 59799 -19823
rect 59957 -19826 60053 -19823
rect 59957 -19857 60520 -19826
rect 59772 -19860 60520 -19857
rect 59772 -19920 59806 -19860
rect 59276 -20038 59310 -19976
rect 58930 -20072 59026 -20038
rect 59214 -20040 59310 -20038
rect 59214 -20072 59696 -20040
rect 58930 -20074 59696 -20072
rect 58930 -20110 58964 -20074
rect 57129 -20191 57131 -20157
rect 57129 -20225 57165 -20191
rect 57129 -20259 57131 -20225
rect 57129 -20275 57165 -20259
rect 57201 -20191 57217 -20157
rect 57251 -20191 57267 -20157
rect 57201 -20225 57267 -20191
rect 57201 -20259 57217 -20225
rect 57251 -20259 57267 -20225
rect 57201 -20309 57267 -20259
rect 57301 -20178 57303 -20144
rect 57337 -20178 57355 -20144
rect 57301 -20225 57355 -20178
rect 57301 -20259 57303 -20225
rect 57337 -20259 57355 -20225
rect 57301 -20275 57355 -20259
rect 59662 -20130 59696 -20074
rect 60486 -19922 60520 -19860
rect 59942 -19974 59958 -19940
rect 60334 -19974 60350 -19940
rect 59874 -19994 59908 -19978
rect 59874 -20044 59908 -20028
rect 60384 -19994 60418 -19978
rect 60384 -20044 60418 -20028
rect 59942 -20082 59958 -20048
rect 60334 -20082 60350 -20048
rect 56112 -20382 56146 -20320
rect 57096 -20343 57125 -20309
rect 57159 -20343 57217 -20309
rect 57251 -20343 57309 -20309
rect 57343 -20343 57372 -20309
rect 55706 -20416 55802 -20382
rect 56050 -20416 56146 -20382
rect 53886 -20464 53982 -20430
rect 54956 -20464 55052 -20430
rect 53886 -20526 53920 -20464
rect 55018 -20526 55052 -20464
rect 55720 -20458 56090 -20416
rect 55720 -20468 56020 -20458
rect 54065 -20578 54081 -20544
rect 54857 -20578 54873 -20544
rect 53988 -20606 54022 -20590
rect 53988 -20660 54022 -20644
rect 54916 -20606 54950 -20590
rect 54916 -20660 54950 -20644
rect 54065 -20706 54081 -20672
rect 54857 -20706 54873 -20672
rect 53886 -20786 53920 -20724
rect 56010 -20608 56020 -20468
rect 56080 -20608 56090 -20458
rect 59109 -20188 59125 -20154
rect 59501 -20188 59517 -20154
rect 59560 -20208 59594 -20192
rect 59560 -20258 59594 -20242
rect 59109 -20296 59125 -20262
rect 59501 -20296 59517 -20262
rect 59032 -20316 59066 -20300
rect 59032 -20366 59066 -20350
rect 59109 -20404 59125 -20370
rect 59501 -20404 59517 -20370
rect 56010 -20618 56090 -20608
rect 59772 -20162 59806 -20100
rect 60486 -20162 60520 -20100
rect 59772 -20196 59866 -20162
rect 60426 -20196 60520 -20162
rect 59662 -20484 59696 -20430
rect 58966 -20500 59026 -20484
rect 58930 -20518 59026 -20500
rect 59600 -20518 59696 -20484
rect 55018 -20786 55052 -20724
rect 53886 -20820 53982 -20786
rect 54956 -20820 55052 -20786
rect 55176 -20678 55272 -20644
rect 55566 -20678 55662 -20644
rect 55176 -20740 55210 -20678
rect 55628 -20740 55662 -20678
rect 55284 -20792 55300 -20758
rect 55476 -20792 55492 -20758
rect 55526 -20802 55560 -20786
rect 55284 -20880 55300 -20846
rect 55476 -20880 55492 -20846
rect 55526 -20852 55560 -20836
rect 55176 -20960 55210 -20898
rect 55628 -20960 55662 -20898
rect 55176 -20994 55272 -20960
rect 55566 -20994 55662 -20960
rect 53896 -23192 53992 -23158
rect 54966 -23192 55062 -23158
rect 53896 -23254 53930 -23192
rect 55028 -23254 55062 -23192
rect 54075 -23306 54091 -23272
rect 54867 -23306 54883 -23272
rect 53998 -23334 54032 -23318
rect 53998 -23388 54032 -23372
rect 54926 -23334 54960 -23318
rect 54926 -23388 54960 -23372
rect 54075 -23434 54091 -23400
rect 54867 -23434 54883 -23400
rect 53896 -23514 53930 -23452
rect 55028 -23514 55062 -23452
rect 55960 -23508 56040 -23498
rect 53896 -23548 53992 -23514
rect 54966 -23548 55062 -23514
rect 53350 -23638 53790 -23604
rect 53350 -23700 53384 -23638
rect 53510 -23740 53526 -23706
rect 53614 -23740 53630 -23706
rect 53464 -23790 53498 -23774
rect 53464 -24582 53498 -24566
rect 53642 -23790 53676 -23774
rect 53642 -24582 53676 -24566
rect 53756 -24264 53790 -23638
rect 53896 -23610 53930 -23548
rect 55028 -23610 55062 -23548
rect 55710 -23554 56040 -23508
rect 54075 -23662 54091 -23628
rect 54867 -23662 54883 -23628
rect 53998 -23690 54032 -23674
rect 53998 -23744 54032 -23728
rect 54926 -23690 54960 -23674
rect 54926 -23744 54960 -23728
rect 54075 -23790 54091 -23756
rect 54867 -23790 54883 -23756
rect 53896 -23870 53930 -23808
rect 55706 -23588 55802 -23554
rect 56050 -23588 56146 -23554
rect 55706 -23650 55740 -23588
rect 55028 -23870 55062 -23808
rect 53896 -23904 53992 -23870
rect 54966 -23904 55062 -23870
rect 55176 -23700 55272 -23666
rect 55430 -23700 55526 -23666
rect 55176 -23762 55210 -23700
rect 55492 -23762 55526 -23700
rect 55318 -23802 55334 -23768
rect 55368 -23802 55384 -23768
rect 55290 -23852 55324 -23836
rect 55290 -24044 55324 -24028
rect 55378 -23852 55412 -23836
rect 55378 -24044 55412 -24028
rect 55176 -24118 55210 -24056
rect 55492 -24118 55526 -24056
rect 54870 -24152 55272 -24118
rect 55430 -24152 55706 -24118
rect 54870 -24158 55706 -24152
rect 54870 -24264 54904 -24158
rect 53756 -24298 53852 -24264
rect 54808 -24298 54904 -24264
rect 53756 -24360 53790 -24298
rect 54870 -24360 54904 -24298
rect 55126 -24308 55142 -24274
rect 55494 -24308 55510 -24274
rect 53926 -24412 53942 -24378
rect 54718 -24412 54734 -24378
rect 53858 -24440 53892 -24424
rect 53858 -24544 53892 -24528
rect 54768 -24440 54802 -24424
rect 54768 -24544 54802 -24528
rect 53926 -24590 53942 -24556
rect 54718 -24590 54734 -24556
rect 53510 -24650 53526 -24616
rect 53614 -24650 53630 -24616
rect 53756 -24670 53790 -24608
rect 55046 -24360 55080 -24344
rect 55046 -24410 55080 -24394
rect 55556 -24360 55590 -24344
rect 55556 -24410 55590 -24394
rect 55126 -24480 55142 -24446
rect 55494 -24480 55510 -24446
rect 54870 -24638 54904 -24608
rect 55700 -24606 55706 -24158
rect 56112 -23650 56146 -23588
rect 58930 -23567 59026 -23533
rect 59600 -23567 59696 -23533
rect 58930 -23610 58964 -23567
rect 58926 -23620 58966 -23610
rect 55866 -23690 55882 -23656
rect 55970 -23690 55986 -23656
rect 55820 -23740 55854 -23724
rect 55820 -24532 55854 -24516
rect 55998 -23740 56032 -23724
rect 55998 -24532 56032 -24516
rect 55866 -24600 55882 -24566
rect 55970 -24600 55986 -24566
rect 55700 -24638 55740 -24606
rect 57096 -23679 57125 -23645
rect 57159 -23679 57217 -23645
rect 57251 -23679 57309 -23645
rect 57343 -23679 57372 -23645
rect 57129 -23729 57165 -23713
rect 57129 -23763 57131 -23729
rect 57129 -23797 57165 -23763
rect 57129 -23831 57131 -23797
rect 57201 -23729 57267 -23679
rect 57201 -23763 57217 -23729
rect 57251 -23763 57267 -23729
rect 57201 -23797 57267 -23763
rect 57201 -23831 57217 -23797
rect 57251 -23831 57267 -23797
rect 57301 -23729 57355 -23713
rect 57301 -23763 57303 -23729
rect 57337 -23763 57355 -23729
rect 57301 -23810 57355 -23763
rect 57129 -23865 57165 -23831
rect 57301 -23844 57303 -23810
rect 57337 -23844 57355 -23810
rect 57129 -23899 57264 -23865
rect 57301 -23894 57355 -23844
rect 57230 -23928 57264 -23899
rect 57117 -23944 57185 -23935
rect 57117 -23994 57118 -23944
rect 57178 -23994 57185 -23944
rect 57117 -24009 57185 -23994
rect 57230 -23944 57285 -23928
rect 57230 -23978 57251 -23944
rect 57230 -23994 57285 -23978
rect 57319 -23940 57355 -23894
rect 59662 -23629 59696 -23567
rect 59109 -23681 59125 -23647
rect 59501 -23681 59517 -23647
rect 59560 -23701 59594 -23685
rect 59560 -23751 59594 -23735
rect 59109 -23789 59125 -23755
rect 59501 -23789 59517 -23755
rect 59032 -23809 59066 -23793
rect 59032 -23859 59066 -23843
rect 59109 -23897 59125 -23863
rect 59501 -23897 59517 -23863
rect 58926 -23940 58966 -23920
rect 57319 -23980 57326 -23940
rect 58930 -23976 58964 -23940
rect 57230 -24045 57264 -23994
rect 57131 -24079 57264 -24045
rect 57319 -24054 57355 -23980
rect 57131 -24100 57165 -24079
rect 56316 -24118 56412 -24104
rect 54830 -24648 55830 -24638
rect 54830 -24670 55030 -24648
rect 53756 -24704 53852 -24670
rect 54808 -24704 55030 -24670
rect 53510 -24758 53526 -24724
rect 53614 -24758 53630 -24724
rect 53756 -24766 53790 -24704
rect 54830 -24728 55030 -24704
rect 55110 -24668 55740 -24648
rect 55810 -24668 55830 -24648
rect 56112 -24668 56146 -24606
rect 55110 -24708 55160 -24668
rect 55600 -24708 55740 -24668
rect 56050 -24702 56146 -24668
rect 55110 -24728 55740 -24708
rect 55810 -24728 55830 -24702
rect 54830 -24738 55830 -24728
rect 53464 -24808 53498 -24792
rect 53464 -25600 53498 -25584
rect 53642 -24808 53676 -24792
rect 53642 -25600 53676 -25584
rect 54870 -24766 54904 -24738
rect 53926 -24818 53942 -24784
rect 54718 -24818 54734 -24784
rect 53858 -24846 53892 -24830
rect 53858 -24950 53892 -24934
rect 54768 -24846 54802 -24830
rect 54768 -24950 54802 -24934
rect 53926 -24996 53942 -24962
rect 54718 -24996 54734 -24962
rect 53756 -25076 53790 -25014
rect 55700 -24764 55740 -24738
rect 55126 -24930 55142 -24896
rect 55494 -24930 55510 -24896
rect 54870 -25076 54904 -25014
rect 55046 -24982 55080 -24966
rect 55046 -25032 55080 -25016
rect 55556 -24982 55590 -24966
rect 55556 -25032 55590 -25016
rect 53756 -25110 53852 -25076
rect 54808 -25110 54904 -25076
rect 55126 -25102 55142 -25068
rect 55494 -25102 55510 -25068
rect 53510 -25668 53526 -25634
rect 53614 -25668 53630 -25634
rect 53350 -25736 53384 -25674
rect 53756 -25736 53790 -25110
rect 54870 -25218 54904 -25110
rect 55700 -25218 55706 -24764
rect 54870 -25224 55706 -25218
rect 54870 -25258 55262 -25224
rect 55420 -25258 55706 -25224
rect 55166 -25320 55200 -25258
rect 53350 -25770 53446 -25736
rect 53694 -25770 53790 -25736
rect 53886 -25508 53982 -25474
rect 54956 -25508 55052 -25474
rect 53886 -25570 53920 -25508
rect 55018 -25570 55052 -25508
rect 54065 -25622 54081 -25588
rect 54857 -25622 54873 -25588
rect 53988 -25650 54022 -25634
rect 53988 -25704 54022 -25688
rect 54916 -25650 54950 -25634
rect 54916 -25704 54950 -25688
rect 54065 -25750 54081 -25716
rect 54857 -25750 54873 -25716
rect 53886 -25830 53920 -25768
rect 55482 -25320 55516 -25258
rect 55280 -25348 55314 -25332
rect 55280 -25540 55314 -25524
rect 55368 -25348 55402 -25332
rect 55368 -25540 55402 -25524
rect 55308 -25608 55324 -25574
rect 55358 -25608 55374 -25574
rect 55166 -25676 55200 -25614
rect 55482 -25676 55516 -25614
rect 55166 -25710 55262 -25676
rect 55420 -25710 55516 -25676
rect 55018 -25830 55052 -25768
rect 56112 -24764 56146 -24702
rect 56350 -24138 56412 -24118
rect 56610 -24138 56706 -24104
rect 56672 -24200 56706 -24138
rect 57303 -24083 57355 -24054
rect 57131 -24155 57165 -24134
rect 57201 -24147 57217 -24113
rect 57251 -24147 57267 -24113
rect 57201 -24189 57267 -24147
rect 57337 -24117 57355 -24083
rect 57303 -24155 57355 -24117
rect 58930 -24010 59026 -23976
rect 59214 -23977 59310 -23976
rect 59662 -23977 59696 -23920
rect 59772 -23894 59866 -23860
rect 60426 -23894 60520 -23860
rect 59772 -23950 59806 -23894
rect 59214 -24010 59696 -23977
rect 58930 -24011 59696 -24010
rect 58930 -24072 58964 -24011
rect 59276 -24072 59310 -24011
rect 59087 -24112 59103 -24078
rect 59137 -24112 59153 -24078
rect 56476 -24240 56492 -24206
rect 56530 -24240 56546 -24206
rect 55866 -24804 55882 -24770
rect 55970 -24804 55986 -24770
rect 55820 -24854 55854 -24838
rect 55820 -25646 55854 -25630
rect 55998 -24854 56032 -24838
rect 55998 -25646 56032 -25630
rect 55866 -25714 55882 -25680
rect 55970 -25714 55986 -25680
rect 55706 -25782 55740 -25720
rect 56430 -24299 56464 -24283
rect 56430 -25091 56464 -25075
rect 56558 -24299 56592 -24283
rect 56558 -25091 56592 -25075
rect 56476 -25168 56492 -25134
rect 56530 -25168 56546 -25134
rect 56316 -25236 56350 -25174
rect 57096 -24223 57125 -24189
rect 57159 -24223 57217 -24189
rect 57251 -24223 57309 -24189
rect 57343 -24223 57372 -24189
rect 59044 -24171 59078 -24155
rect 59044 -24563 59078 -24547
rect 59162 -24171 59196 -24155
rect 59162 -24563 59196 -24547
rect 59087 -24640 59103 -24606
rect 59137 -24640 59153 -24606
rect 60486 -23956 60520 -23894
rect 59942 -24008 59958 -23974
rect 60334 -24008 60350 -23974
rect 59874 -24028 59908 -24012
rect 59874 -24078 59908 -24062
rect 60384 -24028 60418 -24012
rect 60384 -24078 60418 -24062
rect 59942 -24116 59958 -24082
rect 60334 -24116 60350 -24082
rect 59772 -24196 59806 -24140
rect 60486 -24196 60520 -24134
rect 59388 -24230 59476 -24196
rect 59656 -24230 59800 -24196
rect 59958 -24230 60520 -24196
rect 59388 -24290 59422 -24230
rect 59276 -24706 59310 -24646
rect 59530 -24332 59546 -24298
rect 59580 -24332 59596 -24298
rect 59502 -24382 59536 -24366
rect 59502 -24574 59536 -24558
rect 59590 -24382 59624 -24366
rect 59590 -24574 59624 -24558
rect 59530 -24642 59546 -24608
rect 59580 -24642 59596 -24608
rect 58966 -24742 59310 -24706
rect 59388 -24709 59422 -24650
rect 59704 -24709 59738 -24230
rect 60020 -24292 60054 -24230
rect 59846 -24332 59862 -24298
rect 59896 -24332 59912 -24298
rect 59818 -24382 59852 -24366
rect 59818 -24574 59852 -24558
rect 59906 -24382 59940 -24366
rect 59906 -24574 59940 -24558
rect 59846 -24642 59862 -24608
rect 59896 -24642 59912 -24608
rect 61186 -24400 61286 -24390
rect 61186 -24480 61196 -24400
rect 61186 -24490 61286 -24480
rect 60020 -24709 60054 -24648
rect 56672 -25236 56706 -25174
rect 57096 -25199 57125 -25165
rect 57159 -25199 57217 -25165
rect 57251 -25199 57309 -25165
rect 57343 -25199 57372 -25165
rect 56316 -25270 56412 -25236
rect 56610 -25270 56706 -25236
rect 57131 -25254 57165 -25233
rect 57201 -25241 57267 -25199
rect 57201 -25275 57217 -25241
rect 57251 -25275 57267 -25241
rect 57303 -25271 57355 -25233
rect 57131 -25309 57165 -25288
rect 57337 -25305 57355 -25271
rect 59276 -24802 59310 -24742
rect 59387 -24744 60054 -24709
rect 60127 -24554 60161 -24528
rect 60127 -24557 60253 -24554
rect 60161 -24573 60253 -24557
rect 60161 -24591 60203 -24573
rect 60127 -24607 60203 -24591
rect 60237 -24607 60253 -24573
rect 60359 -24560 60409 -24549
rect 60671 -24554 60705 -24528
rect 60359 -24565 60366 -24560
rect 60359 -24600 60366 -24599
rect 60406 -24600 60409 -24560
rect 60127 -24649 60161 -24607
rect 60127 -24741 60161 -24683
rect 60195 -24657 60325 -24641
rect 60195 -24691 60211 -24657
rect 60245 -24691 60325 -24657
rect 60195 -24707 60325 -24691
rect 59387 -24800 59421 -24744
rect 59087 -24842 59103 -24808
rect 59137 -24842 59153 -24808
rect 59044 -24901 59078 -24885
rect 57131 -25343 57264 -25309
rect 57303 -25334 57355 -25305
rect 57117 -25394 57185 -25379
rect 57117 -25444 57118 -25394
rect 57168 -25444 57185 -25394
rect 57117 -25453 57185 -25444
rect 57230 -25394 57264 -25343
rect 57319 -25370 57355 -25334
rect 57230 -25410 57285 -25394
rect 57230 -25444 57251 -25410
rect 57230 -25460 57285 -25444
rect 57319 -25410 57326 -25370
rect 59044 -25293 59078 -25277
rect 59162 -24901 59196 -24885
rect 59162 -25293 59196 -25277
rect 59087 -25370 59103 -25336
rect 59137 -25370 59153 -25336
rect 57230 -25489 57264 -25460
rect 57129 -25523 57264 -25489
rect 57319 -25494 57355 -25410
rect 57129 -25557 57165 -25523
rect 57301 -25544 57355 -25494
rect 58930 -25438 58964 -25376
rect 59529 -24845 59545 -24811
rect 59579 -24845 59595 -24811
rect 59501 -24895 59535 -24879
rect 59501 -25087 59535 -25071
rect 59589 -24895 59623 -24879
rect 59589 -25087 59623 -25071
rect 59529 -25155 59545 -25121
rect 59579 -25155 59595 -25121
rect 59387 -25223 59421 -25170
rect 59703 -25223 59737 -24744
rect 60019 -24805 60053 -24744
rect 59845 -24845 59861 -24811
rect 59895 -24845 59911 -24811
rect 59817 -24895 59851 -24879
rect 59817 -25087 59851 -25071
rect 59905 -24895 59939 -24879
rect 59905 -25087 59939 -25071
rect 59845 -25155 59861 -25121
rect 59895 -25155 59911 -25121
rect 60161 -24775 60203 -24741
rect 60237 -24775 60253 -24741
rect 60127 -24833 60161 -24775
rect 60289 -24809 60325 -24707
rect 60127 -24909 60161 -24867
rect 60195 -24825 60325 -24809
rect 60195 -24859 60211 -24825
rect 60245 -24859 60325 -24825
rect 60195 -24875 60325 -24859
rect 60359 -24650 60409 -24600
rect 60443 -24557 60705 -24554
rect 60443 -24573 60671 -24557
rect 60443 -24607 60459 -24573
rect 60493 -24607 60527 -24573
rect 60561 -24607 60595 -24573
rect 60629 -24591 60671 -24573
rect 60629 -24607 60705 -24591
rect 60359 -24657 60366 -24650
rect 60406 -24690 60409 -24650
rect 60393 -24691 60409 -24690
rect 60359 -24740 60409 -24691
rect 60359 -24741 60366 -24740
rect 60359 -24780 60366 -24775
rect 60406 -24780 60409 -24740
rect 60359 -24820 60409 -24780
rect 60359 -24825 60366 -24820
rect 60359 -24860 60366 -24859
rect 60406 -24860 60409 -24820
rect 60359 -24875 60409 -24860
rect 60443 -24657 60637 -24641
rect 60443 -24691 60459 -24657
rect 60493 -24691 60527 -24657
rect 60561 -24691 60595 -24657
rect 60629 -24691 60637 -24657
rect 60443 -24707 60637 -24691
rect 60671 -24649 60705 -24607
rect 60443 -24809 60477 -24707
rect 60671 -24741 60705 -24683
rect 60511 -24775 60527 -24741
rect 60561 -24775 60595 -24741
rect 60629 -24775 60671 -24741
rect 60443 -24825 60637 -24809
rect 60443 -24859 60459 -24825
rect 60493 -24859 60527 -24825
rect 60561 -24859 60595 -24825
rect 60629 -24859 60637 -24825
rect 60443 -24875 60637 -24859
rect 60671 -24833 60705 -24775
rect 60289 -24909 60325 -24875
rect 60443 -24909 60481 -24875
rect 60671 -24909 60705 -24867
rect 60127 -24925 60204 -24909
rect 60161 -24943 60204 -24925
rect 60238 -24943 60254 -24909
rect 60161 -24959 60254 -24943
rect 60289 -24925 60481 -24909
rect 60289 -24959 60297 -24925
rect 60331 -24959 60369 -24925
rect 60405 -24959 60449 -24925
rect 60579 -24943 60595 -24909
rect 60629 -24925 60705 -24909
rect 60629 -24943 60671 -24925
rect 60579 -24951 60671 -24943
rect 60127 -24988 60161 -24959
rect 60289 -24962 60481 -24959
rect 60671 -24988 60705 -24959
rect 60747 -24554 60781 -24528
rect 60747 -24557 61009 -24554
rect 60781 -24573 61009 -24557
rect 60781 -24591 60823 -24573
rect 60747 -24607 60823 -24591
rect 60857 -24607 60891 -24573
rect 60925 -24607 60959 -24573
rect 60993 -24607 61009 -24573
rect 61043 -24560 61093 -24549
rect 61291 -24554 61325 -24528
rect 61043 -24600 61046 -24560
rect 61086 -24565 61093 -24560
rect 61086 -24600 61093 -24599
rect 60747 -24649 60781 -24607
rect 60747 -24741 60781 -24683
rect 60815 -24657 61009 -24641
rect 60815 -24691 60823 -24657
rect 60857 -24691 60891 -24657
rect 60925 -24691 60959 -24657
rect 60993 -24691 61009 -24657
rect 60815 -24707 61009 -24691
rect 60781 -24775 60823 -24741
rect 60857 -24775 60891 -24741
rect 60925 -24775 60941 -24741
rect 60747 -24833 60781 -24775
rect 60975 -24809 61009 -24707
rect 60747 -24909 60781 -24867
rect 60815 -24825 61009 -24809
rect 60815 -24859 60823 -24825
rect 60857 -24859 60891 -24825
rect 60925 -24859 60959 -24825
rect 60993 -24859 61009 -24825
rect 60815 -24875 61009 -24859
rect 61043 -24650 61093 -24600
rect 61199 -24557 61325 -24554
rect 61199 -24573 61291 -24557
rect 61199 -24607 61215 -24573
rect 61249 -24591 61291 -24573
rect 61249 -24607 61325 -24591
rect 61043 -24690 61046 -24650
rect 61086 -24657 61093 -24650
rect 61043 -24691 61059 -24690
rect 61043 -24740 61093 -24691
rect 61043 -24780 61046 -24740
rect 61086 -24741 61093 -24740
rect 61086 -24780 61093 -24775
rect 61043 -24820 61093 -24780
rect 61043 -24860 61046 -24820
rect 61086 -24825 61093 -24820
rect 61086 -24860 61093 -24859
rect 61043 -24875 61093 -24860
rect 61127 -24657 61257 -24641
rect 61127 -24691 61207 -24657
rect 61241 -24691 61257 -24657
rect 61127 -24707 61257 -24691
rect 61291 -24649 61325 -24607
rect 61127 -24809 61163 -24707
rect 61291 -24741 61325 -24683
rect 61199 -24775 61215 -24741
rect 61249 -24775 61291 -24741
rect 61127 -24825 61257 -24809
rect 61127 -24859 61207 -24825
rect 61241 -24859 61257 -24825
rect 61127 -24875 61257 -24859
rect 61291 -24833 61325 -24775
rect 60971 -24909 61009 -24875
rect 61127 -24909 61163 -24875
rect 61291 -24909 61325 -24867
rect 60747 -24925 60823 -24909
rect 60781 -24943 60823 -24925
rect 60857 -24943 60873 -24909
rect 60781 -24951 60873 -24943
rect 60971 -24924 61163 -24909
rect 60971 -24925 61129 -24924
rect 60747 -24988 60781 -24959
rect 60971 -24959 60980 -24925
rect 61015 -24959 61053 -24925
rect 61088 -24958 61129 -24925
rect 61198 -24943 61214 -24909
rect 61248 -24925 61325 -24909
rect 61248 -24943 61291 -24925
rect 61088 -24959 61163 -24958
rect 61198 -24959 61291 -24943
rect 60971 -24962 61163 -24959
rect 61291 -24988 61325 -24959
rect 60466 -25060 60546 -25040
rect 60466 -25100 60486 -25060
rect 60526 -25100 60546 -25060
rect 60466 -25120 60546 -25100
rect 60606 -25060 60686 -25040
rect 60606 -25100 60626 -25060
rect 60666 -25100 60686 -25060
rect 60606 -25120 60686 -25100
rect 60746 -25060 60826 -25040
rect 60746 -25100 60766 -25060
rect 60806 -25100 60826 -25060
rect 60746 -25120 60826 -25100
rect 60886 -25060 60966 -25040
rect 60886 -25100 60906 -25060
rect 60946 -25100 60966 -25060
rect 60886 -25120 60966 -25100
rect 60019 -25223 60053 -25161
rect 59387 -25257 59476 -25223
rect 59646 -25257 59799 -25223
rect 59957 -25226 60053 -25223
rect 59957 -25257 60520 -25226
rect 59772 -25260 60520 -25257
rect 59772 -25320 59806 -25260
rect 59276 -25438 59310 -25376
rect 58930 -25472 59026 -25438
rect 59214 -25440 59310 -25438
rect 59214 -25472 59696 -25440
rect 58930 -25474 59696 -25472
rect 58930 -25510 58964 -25474
rect 57129 -25591 57131 -25557
rect 57129 -25625 57165 -25591
rect 57129 -25659 57131 -25625
rect 57129 -25675 57165 -25659
rect 57201 -25591 57217 -25557
rect 57251 -25591 57267 -25557
rect 57201 -25625 57267 -25591
rect 57201 -25659 57217 -25625
rect 57251 -25659 57267 -25625
rect 57201 -25709 57267 -25659
rect 57301 -25578 57303 -25544
rect 57337 -25578 57355 -25544
rect 57301 -25625 57355 -25578
rect 57301 -25659 57303 -25625
rect 57337 -25659 57355 -25625
rect 57301 -25675 57355 -25659
rect 59662 -25530 59696 -25474
rect 60486 -25322 60520 -25260
rect 59942 -25374 59958 -25340
rect 60334 -25374 60350 -25340
rect 59874 -25394 59908 -25378
rect 59874 -25444 59908 -25428
rect 60384 -25394 60418 -25378
rect 60384 -25444 60418 -25428
rect 59942 -25482 59958 -25448
rect 60334 -25482 60350 -25448
rect 56112 -25782 56146 -25720
rect 57096 -25743 57125 -25709
rect 57159 -25743 57217 -25709
rect 57251 -25743 57309 -25709
rect 57343 -25743 57372 -25709
rect 55706 -25816 55802 -25782
rect 56050 -25816 56146 -25782
rect 53886 -25864 53982 -25830
rect 54956 -25864 55052 -25830
rect 53886 -25926 53920 -25864
rect 55018 -25926 55052 -25864
rect 55720 -25858 56090 -25816
rect 55720 -25868 56020 -25858
rect 54065 -25978 54081 -25944
rect 54857 -25978 54873 -25944
rect 53988 -26006 54022 -25990
rect 53988 -26060 54022 -26044
rect 54916 -26006 54950 -25990
rect 54916 -26060 54950 -26044
rect 54065 -26106 54081 -26072
rect 54857 -26106 54873 -26072
rect 53886 -26186 53920 -26124
rect 56010 -26008 56020 -25868
rect 56080 -26008 56090 -25858
rect 59109 -25588 59125 -25554
rect 59501 -25588 59517 -25554
rect 59560 -25608 59594 -25592
rect 59560 -25658 59594 -25642
rect 59109 -25696 59125 -25662
rect 59501 -25696 59517 -25662
rect 59032 -25716 59066 -25700
rect 59032 -25766 59066 -25750
rect 59109 -25804 59125 -25770
rect 59501 -25804 59517 -25770
rect 56010 -26018 56090 -26008
rect 59772 -25562 59806 -25500
rect 60486 -25562 60520 -25500
rect 59772 -25596 59866 -25562
rect 60426 -25596 60520 -25562
rect 59662 -25884 59696 -25830
rect 58966 -25900 59026 -25884
rect 58930 -25918 59026 -25900
rect 59600 -25918 59696 -25884
rect 55018 -26186 55052 -26124
rect 53886 -26220 53982 -26186
rect 54956 -26220 55052 -26186
rect 55176 -26078 55272 -26044
rect 55566 -26078 55662 -26044
rect 55176 -26140 55210 -26078
rect 55628 -26140 55662 -26078
rect 55284 -26192 55300 -26158
rect 55476 -26192 55492 -26158
rect 55526 -26202 55560 -26186
rect 55284 -26280 55300 -26246
rect 55476 -26280 55492 -26246
rect 55526 -26252 55560 -26236
rect 55176 -26360 55210 -26298
rect 55628 -26360 55662 -26298
rect 55176 -26394 55272 -26360
rect 55566 -26394 55662 -26360
rect 53896 -28592 53992 -28558
rect 54966 -28592 55062 -28558
rect 53896 -28654 53930 -28592
rect 55028 -28654 55062 -28592
rect 54075 -28706 54091 -28672
rect 54867 -28706 54883 -28672
rect 53998 -28734 54032 -28718
rect 53998 -28788 54032 -28772
rect 54926 -28734 54960 -28718
rect 54926 -28788 54960 -28772
rect 54075 -28834 54091 -28800
rect 54867 -28834 54883 -28800
rect 53896 -28914 53930 -28852
rect 55028 -28914 55062 -28852
rect 55960 -28908 56040 -28898
rect 53896 -28948 53992 -28914
rect 54966 -28948 55062 -28914
rect 53350 -29038 53790 -29004
rect 53350 -29100 53384 -29038
rect 53510 -29140 53526 -29106
rect 53614 -29140 53630 -29106
rect 53464 -29190 53498 -29174
rect 53464 -29982 53498 -29966
rect 53642 -29190 53676 -29174
rect 53642 -29982 53676 -29966
rect 53756 -29664 53790 -29038
rect 53896 -29010 53930 -28948
rect 55028 -29010 55062 -28948
rect 55710 -28954 56040 -28908
rect 54075 -29062 54091 -29028
rect 54867 -29062 54883 -29028
rect 53998 -29090 54032 -29074
rect 53998 -29144 54032 -29128
rect 54926 -29090 54960 -29074
rect 54926 -29144 54960 -29128
rect 54075 -29190 54091 -29156
rect 54867 -29190 54883 -29156
rect 53896 -29270 53930 -29208
rect 55706 -28988 55802 -28954
rect 56050 -28988 56146 -28954
rect 55706 -29050 55740 -28988
rect 55028 -29270 55062 -29208
rect 53896 -29304 53992 -29270
rect 54966 -29304 55062 -29270
rect 55176 -29100 55272 -29066
rect 55430 -29100 55526 -29066
rect 55176 -29162 55210 -29100
rect 55492 -29162 55526 -29100
rect 55318 -29202 55334 -29168
rect 55368 -29202 55384 -29168
rect 55290 -29252 55324 -29236
rect 55290 -29444 55324 -29428
rect 55378 -29252 55412 -29236
rect 55378 -29444 55412 -29428
rect 55176 -29518 55210 -29456
rect 55492 -29518 55526 -29456
rect 54870 -29552 55272 -29518
rect 55430 -29552 55706 -29518
rect 54870 -29558 55706 -29552
rect 54870 -29664 54904 -29558
rect 53756 -29698 53852 -29664
rect 54808 -29698 54904 -29664
rect 53756 -29760 53790 -29698
rect 54870 -29760 54904 -29698
rect 55126 -29708 55142 -29674
rect 55494 -29708 55510 -29674
rect 53926 -29812 53942 -29778
rect 54718 -29812 54734 -29778
rect 53858 -29840 53892 -29824
rect 53858 -29944 53892 -29928
rect 54768 -29840 54802 -29824
rect 54768 -29944 54802 -29928
rect 53926 -29990 53942 -29956
rect 54718 -29990 54734 -29956
rect 53510 -30050 53526 -30016
rect 53614 -30050 53630 -30016
rect 53756 -30070 53790 -30008
rect 55046 -29760 55080 -29744
rect 55046 -29810 55080 -29794
rect 55556 -29760 55590 -29744
rect 55556 -29810 55590 -29794
rect 55126 -29880 55142 -29846
rect 55494 -29880 55510 -29846
rect 54870 -30038 54904 -30008
rect 55700 -30006 55706 -29558
rect 56112 -29050 56146 -28988
rect 58930 -28967 59026 -28933
rect 59600 -28967 59696 -28933
rect 58930 -29010 58964 -28967
rect 58926 -29020 58966 -29010
rect 55866 -29090 55882 -29056
rect 55970 -29090 55986 -29056
rect 55820 -29140 55854 -29124
rect 55820 -29932 55854 -29916
rect 55998 -29140 56032 -29124
rect 55998 -29932 56032 -29916
rect 55866 -30000 55882 -29966
rect 55970 -30000 55986 -29966
rect 55700 -30038 55740 -30006
rect 57096 -29079 57125 -29045
rect 57159 -29079 57217 -29045
rect 57251 -29079 57309 -29045
rect 57343 -29079 57372 -29045
rect 57129 -29129 57165 -29113
rect 57129 -29163 57131 -29129
rect 57129 -29197 57165 -29163
rect 57129 -29231 57131 -29197
rect 57201 -29129 57267 -29079
rect 57201 -29163 57217 -29129
rect 57251 -29163 57267 -29129
rect 57201 -29197 57267 -29163
rect 57201 -29231 57217 -29197
rect 57251 -29231 57267 -29197
rect 57301 -29129 57355 -29113
rect 57301 -29163 57303 -29129
rect 57337 -29163 57355 -29129
rect 57301 -29210 57355 -29163
rect 57129 -29265 57165 -29231
rect 57301 -29244 57303 -29210
rect 57337 -29244 57355 -29210
rect 57129 -29299 57264 -29265
rect 57301 -29294 57355 -29244
rect 57230 -29328 57264 -29299
rect 57117 -29344 57185 -29335
rect 57117 -29394 57118 -29344
rect 57178 -29394 57185 -29344
rect 57117 -29409 57185 -29394
rect 57230 -29344 57285 -29328
rect 57230 -29378 57251 -29344
rect 57230 -29394 57285 -29378
rect 57319 -29340 57355 -29294
rect 59662 -29029 59696 -28967
rect 59109 -29081 59125 -29047
rect 59501 -29081 59517 -29047
rect 59560 -29101 59594 -29085
rect 59560 -29151 59594 -29135
rect 59109 -29189 59125 -29155
rect 59501 -29189 59517 -29155
rect 59032 -29209 59066 -29193
rect 59032 -29259 59066 -29243
rect 59109 -29297 59125 -29263
rect 59501 -29297 59517 -29263
rect 58926 -29340 58966 -29320
rect 57319 -29380 57326 -29340
rect 58930 -29376 58964 -29340
rect 57230 -29445 57264 -29394
rect 57131 -29479 57264 -29445
rect 57319 -29454 57355 -29380
rect 57131 -29500 57165 -29479
rect 56316 -29518 56412 -29504
rect 54830 -30048 55830 -30038
rect 54830 -30070 55030 -30048
rect 53756 -30104 53852 -30070
rect 54808 -30104 55030 -30070
rect 53510 -30158 53526 -30124
rect 53614 -30158 53630 -30124
rect 53756 -30166 53790 -30104
rect 54830 -30128 55030 -30104
rect 55110 -30068 55740 -30048
rect 55810 -30068 55830 -30048
rect 56112 -30068 56146 -30006
rect 55110 -30108 55160 -30068
rect 55600 -30108 55740 -30068
rect 56050 -30102 56146 -30068
rect 55110 -30128 55740 -30108
rect 55810 -30128 55830 -30102
rect 54830 -30138 55830 -30128
rect 53464 -30208 53498 -30192
rect 25738 -31020 35838 -30998
rect 25780 -31032 35838 -31020
rect 35804 -31094 35838 -31032
rect 53464 -31000 53498 -30984
rect 53642 -30208 53676 -30192
rect 53642 -31000 53676 -30984
rect 54870 -30166 54904 -30138
rect 53926 -30218 53942 -30184
rect 54718 -30218 54734 -30184
rect 53858 -30246 53892 -30230
rect 53858 -30350 53892 -30334
rect 54768 -30246 54802 -30230
rect 54768 -30350 54802 -30334
rect 53926 -30396 53942 -30362
rect 54718 -30396 54734 -30362
rect 53756 -30476 53790 -30414
rect 55700 -30164 55740 -30138
rect 55126 -30330 55142 -30296
rect 55494 -30330 55510 -30296
rect 54870 -30476 54904 -30414
rect 55046 -30382 55080 -30366
rect 55046 -30432 55080 -30416
rect 55556 -30382 55590 -30366
rect 55556 -30432 55590 -30416
rect 53756 -30510 53852 -30476
rect 54808 -30510 54904 -30476
rect 55126 -30502 55142 -30468
rect 55494 -30502 55510 -30468
rect 53510 -31068 53526 -31034
rect 53614 -31068 53630 -31034
rect 53350 -31136 53384 -31074
rect 53756 -31136 53790 -30510
rect 54870 -30618 54904 -30510
rect 55700 -30618 55706 -30164
rect 54870 -30624 55706 -30618
rect 54870 -30658 55262 -30624
rect 55420 -30658 55706 -30624
rect 55166 -30720 55200 -30658
rect 53350 -31170 53446 -31136
rect 53694 -31170 53790 -31136
rect 53886 -30908 53982 -30874
rect 54956 -30908 55052 -30874
rect 53886 -30970 53920 -30908
rect 55018 -30970 55052 -30908
rect 54065 -31022 54081 -30988
rect 54857 -31022 54873 -30988
rect 53988 -31050 54022 -31034
rect 53988 -31104 54022 -31088
rect 54916 -31050 54950 -31034
rect 54916 -31104 54950 -31088
rect 54065 -31150 54081 -31116
rect 54857 -31150 54873 -31116
rect 53886 -31230 53920 -31168
rect 55482 -30720 55516 -30658
rect 55280 -30748 55314 -30732
rect 55280 -30940 55314 -30924
rect 55368 -30748 55402 -30732
rect 55368 -30940 55402 -30924
rect 55308 -31008 55324 -30974
rect 55358 -31008 55374 -30974
rect 55166 -31076 55200 -31014
rect 55482 -31076 55516 -31014
rect 55166 -31110 55262 -31076
rect 55420 -31110 55516 -31076
rect 55018 -31230 55052 -31168
rect 56112 -30164 56146 -30102
rect 56350 -29538 56412 -29518
rect 56610 -29538 56706 -29504
rect 56672 -29600 56706 -29538
rect 57303 -29483 57355 -29454
rect 57131 -29555 57165 -29534
rect 57201 -29547 57217 -29513
rect 57251 -29547 57267 -29513
rect 57201 -29589 57267 -29547
rect 57337 -29517 57355 -29483
rect 57303 -29555 57355 -29517
rect 58930 -29410 59026 -29376
rect 59214 -29377 59310 -29376
rect 59662 -29377 59696 -29320
rect 59772 -29294 59866 -29260
rect 60426 -29294 60520 -29260
rect 59772 -29350 59806 -29294
rect 59214 -29410 59696 -29377
rect 58930 -29411 59696 -29410
rect 58930 -29472 58964 -29411
rect 59276 -29472 59310 -29411
rect 59087 -29512 59103 -29478
rect 59137 -29512 59153 -29478
rect 56476 -29640 56492 -29606
rect 56530 -29640 56546 -29606
rect 55866 -30204 55882 -30170
rect 55970 -30204 55986 -30170
rect 55820 -30254 55854 -30238
rect 55820 -31046 55854 -31030
rect 55998 -30254 56032 -30238
rect 55998 -31046 56032 -31030
rect 55866 -31114 55882 -31080
rect 55970 -31114 55986 -31080
rect 55706 -31182 55740 -31120
rect 56430 -29699 56464 -29683
rect 56430 -30491 56464 -30475
rect 56558 -29699 56592 -29683
rect 56558 -30491 56592 -30475
rect 56476 -30568 56492 -30534
rect 56530 -30568 56546 -30534
rect 56316 -30636 56350 -30574
rect 57096 -29623 57125 -29589
rect 57159 -29623 57217 -29589
rect 57251 -29623 57309 -29589
rect 57343 -29623 57372 -29589
rect 59044 -29571 59078 -29555
rect 59044 -29963 59078 -29947
rect 59162 -29571 59196 -29555
rect 59162 -29963 59196 -29947
rect 59087 -30040 59103 -30006
rect 59137 -30040 59153 -30006
rect 60486 -29356 60520 -29294
rect 59942 -29408 59958 -29374
rect 60334 -29408 60350 -29374
rect 59874 -29428 59908 -29412
rect 59874 -29478 59908 -29462
rect 60384 -29428 60418 -29412
rect 60384 -29478 60418 -29462
rect 59942 -29516 59958 -29482
rect 60334 -29516 60350 -29482
rect 59772 -29596 59806 -29540
rect 60486 -29596 60520 -29534
rect 59388 -29630 59476 -29596
rect 59656 -29630 59800 -29596
rect 59958 -29630 60520 -29596
rect 59388 -29690 59422 -29630
rect 59276 -30106 59310 -30046
rect 59530 -29732 59546 -29698
rect 59580 -29732 59596 -29698
rect 59502 -29782 59536 -29766
rect 59502 -29974 59536 -29958
rect 59590 -29782 59624 -29766
rect 59590 -29974 59624 -29958
rect 59530 -30042 59546 -30008
rect 59580 -30042 59596 -30008
rect 58966 -30142 59310 -30106
rect 59388 -30109 59422 -30050
rect 59704 -30109 59738 -29630
rect 60020 -29692 60054 -29630
rect 59846 -29732 59862 -29698
rect 59896 -29732 59912 -29698
rect 59818 -29782 59852 -29766
rect 59818 -29974 59852 -29958
rect 59906 -29782 59940 -29766
rect 59906 -29974 59940 -29958
rect 59846 -30042 59862 -30008
rect 59896 -30042 59912 -30008
rect 61186 -29800 61286 -29790
rect 61186 -29880 61196 -29800
rect 61186 -29890 61286 -29880
rect 60020 -30109 60054 -30048
rect 56672 -30636 56706 -30574
rect 57096 -30599 57125 -30565
rect 57159 -30599 57217 -30565
rect 57251 -30599 57309 -30565
rect 57343 -30599 57372 -30565
rect 56316 -30670 56412 -30636
rect 56610 -30670 56706 -30636
rect 57131 -30654 57165 -30633
rect 57201 -30641 57267 -30599
rect 57201 -30675 57217 -30641
rect 57251 -30675 57267 -30641
rect 57303 -30671 57355 -30633
rect 57131 -30709 57165 -30688
rect 57337 -30705 57355 -30671
rect 59276 -30202 59310 -30142
rect 59387 -30144 60054 -30109
rect 60127 -29954 60161 -29928
rect 60127 -29957 60253 -29954
rect 60161 -29973 60253 -29957
rect 60161 -29991 60203 -29973
rect 60127 -30007 60203 -29991
rect 60237 -30007 60253 -29973
rect 60359 -29960 60409 -29949
rect 60671 -29954 60705 -29928
rect 60359 -29965 60366 -29960
rect 60359 -30000 60366 -29999
rect 60406 -30000 60409 -29960
rect 60127 -30049 60161 -30007
rect 60127 -30141 60161 -30083
rect 60195 -30057 60325 -30041
rect 60195 -30091 60211 -30057
rect 60245 -30091 60325 -30057
rect 60195 -30107 60325 -30091
rect 59387 -30200 59421 -30144
rect 59087 -30242 59103 -30208
rect 59137 -30242 59153 -30208
rect 59044 -30301 59078 -30285
rect 57131 -30743 57264 -30709
rect 57303 -30734 57355 -30705
rect 57117 -30794 57185 -30779
rect 57117 -30844 57118 -30794
rect 57168 -30844 57185 -30794
rect 57117 -30853 57185 -30844
rect 57230 -30794 57264 -30743
rect 57319 -30770 57355 -30734
rect 57230 -30810 57285 -30794
rect 57230 -30844 57251 -30810
rect 57230 -30860 57285 -30844
rect 57319 -30810 57326 -30770
rect 59044 -30693 59078 -30677
rect 59162 -30301 59196 -30285
rect 59162 -30693 59196 -30677
rect 59087 -30770 59103 -30736
rect 59137 -30770 59153 -30736
rect 57230 -30889 57264 -30860
rect 57129 -30923 57264 -30889
rect 57319 -30894 57355 -30810
rect 57129 -30957 57165 -30923
rect 57301 -30944 57355 -30894
rect 58930 -30838 58964 -30776
rect 59529 -30245 59545 -30211
rect 59579 -30245 59595 -30211
rect 59501 -30295 59535 -30279
rect 59501 -30487 59535 -30471
rect 59589 -30295 59623 -30279
rect 59589 -30487 59623 -30471
rect 59529 -30555 59545 -30521
rect 59579 -30555 59595 -30521
rect 59387 -30623 59421 -30570
rect 59703 -30623 59737 -30144
rect 60019 -30205 60053 -30144
rect 59845 -30245 59861 -30211
rect 59895 -30245 59911 -30211
rect 59817 -30295 59851 -30279
rect 59817 -30487 59851 -30471
rect 59905 -30295 59939 -30279
rect 59905 -30487 59939 -30471
rect 59845 -30555 59861 -30521
rect 59895 -30555 59911 -30521
rect 60161 -30175 60203 -30141
rect 60237 -30175 60253 -30141
rect 60127 -30233 60161 -30175
rect 60289 -30209 60325 -30107
rect 60127 -30309 60161 -30267
rect 60195 -30225 60325 -30209
rect 60195 -30259 60211 -30225
rect 60245 -30259 60325 -30225
rect 60195 -30275 60325 -30259
rect 60359 -30050 60409 -30000
rect 60443 -29957 60705 -29954
rect 60443 -29973 60671 -29957
rect 60443 -30007 60459 -29973
rect 60493 -30007 60527 -29973
rect 60561 -30007 60595 -29973
rect 60629 -29991 60671 -29973
rect 60629 -30007 60705 -29991
rect 60359 -30057 60366 -30050
rect 60406 -30090 60409 -30050
rect 60393 -30091 60409 -30090
rect 60359 -30140 60409 -30091
rect 60359 -30141 60366 -30140
rect 60359 -30180 60366 -30175
rect 60406 -30180 60409 -30140
rect 60359 -30220 60409 -30180
rect 60359 -30225 60366 -30220
rect 60359 -30260 60366 -30259
rect 60406 -30260 60409 -30220
rect 60359 -30275 60409 -30260
rect 60443 -30057 60637 -30041
rect 60443 -30091 60459 -30057
rect 60493 -30091 60527 -30057
rect 60561 -30091 60595 -30057
rect 60629 -30091 60637 -30057
rect 60443 -30107 60637 -30091
rect 60671 -30049 60705 -30007
rect 60443 -30209 60477 -30107
rect 60671 -30141 60705 -30083
rect 60511 -30175 60527 -30141
rect 60561 -30175 60595 -30141
rect 60629 -30175 60671 -30141
rect 60443 -30225 60637 -30209
rect 60443 -30259 60459 -30225
rect 60493 -30259 60527 -30225
rect 60561 -30259 60595 -30225
rect 60629 -30259 60637 -30225
rect 60443 -30275 60637 -30259
rect 60671 -30233 60705 -30175
rect 60289 -30309 60325 -30275
rect 60443 -30309 60481 -30275
rect 60671 -30309 60705 -30267
rect 60127 -30325 60204 -30309
rect 60161 -30343 60204 -30325
rect 60238 -30343 60254 -30309
rect 60161 -30359 60254 -30343
rect 60289 -30325 60481 -30309
rect 60289 -30359 60297 -30325
rect 60331 -30359 60369 -30325
rect 60405 -30359 60449 -30325
rect 60579 -30343 60595 -30309
rect 60629 -30325 60705 -30309
rect 60629 -30343 60671 -30325
rect 60579 -30351 60671 -30343
rect 60127 -30388 60161 -30359
rect 60289 -30362 60481 -30359
rect 60671 -30388 60705 -30359
rect 60747 -29954 60781 -29928
rect 60747 -29957 61009 -29954
rect 60781 -29973 61009 -29957
rect 60781 -29991 60823 -29973
rect 60747 -30007 60823 -29991
rect 60857 -30007 60891 -29973
rect 60925 -30007 60959 -29973
rect 60993 -30007 61009 -29973
rect 61043 -29960 61093 -29949
rect 61291 -29954 61325 -29928
rect 61043 -30000 61046 -29960
rect 61086 -29965 61093 -29960
rect 61086 -30000 61093 -29999
rect 60747 -30049 60781 -30007
rect 60747 -30141 60781 -30083
rect 60815 -30057 61009 -30041
rect 60815 -30091 60823 -30057
rect 60857 -30091 60891 -30057
rect 60925 -30091 60959 -30057
rect 60993 -30091 61009 -30057
rect 60815 -30107 61009 -30091
rect 60781 -30175 60823 -30141
rect 60857 -30175 60891 -30141
rect 60925 -30175 60941 -30141
rect 60747 -30233 60781 -30175
rect 60975 -30209 61009 -30107
rect 60747 -30309 60781 -30267
rect 60815 -30225 61009 -30209
rect 60815 -30259 60823 -30225
rect 60857 -30259 60891 -30225
rect 60925 -30259 60959 -30225
rect 60993 -30259 61009 -30225
rect 60815 -30275 61009 -30259
rect 61043 -30050 61093 -30000
rect 61199 -29957 61325 -29954
rect 61199 -29973 61291 -29957
rect 61199 -30007 61215 -29973
rect 61249 -29991 61291 -29973
rect 61249 -30007 61325 -29991
rect 61043 -30090 61046 -30050
rect 61086 -30057 61093 -30050
rect 61043 -30091 61059 -30090
rect 61043 -30140 61093 -30091
rect 61043 -30180 61046 -30140
rect 61086 -30141 61093 -30140
rect 61086 -30180 61093 -30175
rect 61043 -30220 61093 -30180
rect 61043 -30260 61046 -30220
rect 61086 -30225 61093 -30220
rect 61086 -30260 61093 -30259
rect 61043 -30275 61093 -30260
rect 61127 -30057 61257 -30041
rect 61127 -30091 61207 -30057
rect 61241 -30091 61257 -30057
rect 61127 -30107 61257 -30091
rect 61291 -30049 61325 -30007
rect 61127 -30209 61163 -30107
rect 61291 -30141 61325 -30083
rect 61199 -30175 61215 -30141
rect 61249 -30175 61291 -30141
rect 61127 -30225 61257 -30209
rect 61127 -30259 61207 -30225
rect 61241 -30259 61257 -30225
rect 61127 -30275 61257 -30259
rect 61291 -30233 61325 -30175
rect 60971 -30309 61009 -30275
rect 61127 -30309 61163 -30275
rect 61291 -30309 61325 -30267
rect 60747 -30325 60823 -30309
rect 60781 -30343 60823 -30325
rect 60857 -30343 60873 -30309
rect 60781 -30351 60873 -30343
rect 60971 -30324 61163 -30309
rect 60971 -30325 61129 -30324
rect 60747 -30388 60781 -30359
rect 60971 -30359 60980 -30325
rect 61015 -30359 61053 -30325
rect 61088 -30358 61129 -30325
rect 61198 -30343 61214 -30309
rect 61248 -30325 61325 -30309
rect 61248 -30343 61291 -30325
rect 61088 -30359 61163 -30358
rect 61198 -30359 61291 -30343
rect 60971 -30362 61163 -30359
rect 61291 -30388 61325 -30359
rect 60466 -30460 60546 -30440
rect 60466 -30500 60486 -30460
rect 60526 -30500 60546 -30460
rect 60466 -30520 60546 -30500
rect 60606 -30460 60686 -30440
rect 60606 -30500 60626 -30460
rect 60666 -30500 60686 -30460
rect 60606 -30520 60686 -30500
rect 60746 -30460 60826 -30440
rect 60746 -30500 60766 -30460
rect 60806 -30500 60826 -30460
rect 60746 -30520 60826 -30500
rect 60886 -30460 60966 -30440
rect 60886 -30500 60906 -30460
rect 60946 -30500 60966 -30460
rect 60886 -30520 60966 -30500
rect 60019 -30623 60053 -30561
rect 59387 -30657 59476 -30623
rect 59646 -30657 59799 -30623
rect 59957 -30626 60053 -30623
rect 59957 -30657 60520 -30626
rect 59772 -30660 60520 -30657
rect 59772 -30720 59806 -30660
rect 59276 -30838 59310 -30776
rect 58930 -30872 59026 -30838
rect 59214 -30840 59310 -30838
rect 59214 -30872 59696 -30840
rect 58930 -30874 59696 -30872
rect 58930 -30910 58964 -30874
rect 57129 -30991 57131 -30957
rect 57129 -31025 57165 -30991
rect 57129 -31059 57131 -31025
rect 57129 -31075 57165 -31059
rect 57201 -30991 57217 -30957
rect 57251 -30991 57267 -30957
rect 57201 -31025 57267 -30991
rect 57201 -31059 57217 -31025
rect 57251 -31059 57267 -31025
rect 57201 -31109 57267 -31059
rect 57301 -30978 57303 -30944
rect 57337 -30978 57355 -30944
rect 57301 -31025 57355 -30978
rect 57301 -31059 57303 -31025
rect 57337 -31059 57355 -31025
rect 57301 -31075 57355 -31059
rect 59662 -30930 59696 -30874
rect 60486 -30722 60520 -30660
rect 59942 -30774 59958 -30740
rect 60334 -30774 60350 -30740
rect 59874 -30794 59908 -30778
rect 59874 -30844 59908 -30828
rect 60384 -30794 60418 -30778
rect 60384 -30844 60418 -30828
rect 59942 -30882 59958 -30848
rect 60334 -30882 60350 -30848
rect 56112 -31182 56146 -31120
rect 57096 -31143 57125 -31109
rect 57159 -31143 57217 -31109
rect 57251 -31143 57309 -31109
rect 57343 -31143 57372 -31109
rect 55706 -31216 55802 -31182
rect 56050 -31216 56146 -31182
rect 53886 -31264 53982 -31230
rect 54956 -31264 55052 -31230
rect 53886 -31326 53920 -31264
rect 55018 -31326 55052 -31264
rect 55720 -31258 56090 -31216
rect 55720 -31268 56020 -31258
rect 54065 -31378 54081 -31344
rect 54857 -31378 54873 -31344
rect 53988 -31406 54022 -31390
rect 53988 -31460 54022 -31444
rect 54916 -31406 54950 -31390
rect 54916 -31460 54950 -31444
rect 54065 -31506 54081 -31472
rect 54857 -31506 54873 -31472
rect 53886 -31586 53920 -31524
rect 56010 -31408 56020 -31268
rect 56080 -31408 56090 -31258
rect 59109 -30988 59125 -30954
rect 59501 -30988 59517 -30954
rect 59560 -31008 59594 -30992
rect 59560 -31058 59594 -31042
rect 59109 -31096 59125 -31062
rect 59501 -31096 59517 -31062
rect 59032 -31116 59066 -31100
rect 59032 -31166 59066 -31150
rect 59109 -31204 59125 -31170
rect 59501 -31204 59517 -31170
rect 56010 -31418 56090 -31408
rect 59772 -30962 59806 -30900
rect 60486 -30962 60520 -30900
rect 59772 -30996 59866 -30962
rect 60426 -30996 60520 -30962
rect 59662 -31284 59696 -31230
rect 58966 -31300 59026 -31284
rect 58930 -31318 59026 -31300
rect 59600 -31318 59696 -31284
rect 55018 -31586 55052 -31524
rect 53886 -31620 53982 -31586
rect 54956 -31620 55052 -31586
rect 55176 -31478 55272 -31444
rect 55566 -31478 55662 -31444
rect 55176 -31540 55210 -31478
rect 55628 -31540 55662 -31478
rect 55284 -31592 55300 -31558
rect 55476 -31592 55492 -31558
rect 55526 -31602 55560 -31586
rect 55284 -31680 55300 -31646
rect 55476 -31680 55492 -31646
rect 55526 -31652 55560 -31636
rect 55176 -31760 55210 -31698
rect 55628 -31760 55662 -31698
rect 55176 -31794 55272 -31760
rect 55566 -31794 55662 -31760
rect 35804 -32592 35838 -32530
rect 25780 -32626 35838 -32592
rect 25780 -32630 35836 -32626
rect 35802 -32692 35836 -32630
rect 35802 -34190 35836 -34128
rect 25780 -34228 35836 -34190
rect 35802 -34290 35836 -34228
rect 53896 -33992 53992 -33958
rect 54966 -33992 55062 -33958
rect 53896 -34054 53930 -33992
rect 55028 -34054 55062 -33992
rect 54075 -34106 54091 -34072
rect 54867 -34106 54883 -34072
rect 53998 -34134 54032 -34118
rect 53998 -34188 54032 -34172
rect 54926 -34134 54960 -34118
rect 54926 -34188 54960 -34172
rect 54075 -34234 54091 -34200
rect 54867 -34234 54883 -34200
rect 53896 -34314 53930 -34252
rect 55028 -34314 55062 -34252
rect 55960 -34308 56040 -34298
rect 53896 -34348 53992 -34314
rect 54966 -34348 55062 -34314
rect 53350 -34438 53790 -34404
rect 53350 -34500 53384 -34438
rect 53510 -34540 53526 -34506
rect 53614 -34540 53630 -34506
rect 35802 -35788 35836 -35726
rect 25780 -35830 35836 -35788
rect 35802 -35892 35836 -35830
rect 53464 -34590 53498 -34574
rect 53464 -35382 53498 -35366
rect 53642 -34590 53676 -34574
rect 53642 -35382 53676 -35366
rect 53756 -35064 53790 -34438
rect 53896 -34410 53930 -34348
rect 55028 -34410 55062 -34348
rect 55710 -34354 56040 -34308
rect 54075 -34462 54091 -34428
rect 54867 -34462 54883 -34428
rect 53998 -34490 54032 -34474
rect 53998 -34544 54032 -34528
rect 54926 -34490 54960 -34474
rect 54926 -34544 54960 -34528
rect 54075 -34590 54091 -34556
rect 54867 -34590 54883 -34556
rect 53896 -34670 53930 -34608
rect 55706 -34388 55802 -34354
rect 56050 -34388 56146 -34354
rect 55706 -34450 55740 -34388
rect 55028 -34670 55062 -34608
rect 53896 -34704 53992 -34670
rect 54966 -34704 55062 -34670
rect 55176 -34500 55272 -34466
rect 55430 -34500 55526 -34466
rect 55176 -34562 55210 -34500
rect 55492 -34562 55526 -34500
rect 55318 -34602 55334 -34568
rect 55368 -34602 55384 -34568
rect 55290 -34652 55324 -34636
rect 55290 -34844 55324 -34828
rect 55378 -34652 55412 -34636
rect 55378 -34844 55412 -34828
rect 55176 -34918 55210 -34856
rect 55492 -34918 55526 -34856
rect 54870 -34952 55272 -34918
rect 55430 -34952 55706 -34918
rect 54870 -34958 55706 -34952
rect 54870 -35064 54904 -34958
rect 53756 -35098 53852 -35064
rect 54808 -35098 54904 -35064
rect 53756 -35160 53790 -35098
rect 54870 -35160 54904 -35098
rect 55126 -35108 55142 -35074
rect 55494 -35108 55510 -35074
rect 53926 -35212 53942 -35178
rect 54718 -35212 54734 -35178
rect 53858 -35240 53892 -35224
rect 53858 -35344 53892 -35328
rect 54768 -35240 54802 -35224
rect 54768 -35344 54802 -35328
rect 53926 -35390 53942 -35356
rect 54718 -35390 54734 -35356
rect 53510 -35450 53526 -35416
rect 53614 -35450 53630 -35416
rect 53756 -35470 53790 -35408
rect 55046 -35160 55080 -35144
rect 55046 -35210 55080 -35194
rect 55556 -35160 55590 -35144
rect 55556 -35210 55590 -35194
rect 55126 -35280 55142 -35246
rect 55494 -35280 55510 -35246
rect 54870 -35438 54904 -35408
rect 55700 -35406 55706 -34958
rect 56112 -34450 56146 -34388
rect 58930 -34367 59026 -34333
rect 59600 -34367 59696 -34333
rect 58930 -34410 58964 -34367
rect 58926 -34420 58966 -34410
rect 55866 -34490 55882 -34456
rect 55970 -34490 55986 -34456
rect 55820 -34540 55854 -34524
rect 55820 -35332 55854 -35316
rect 55998 -34540 56032 -34524
rect 55998 -35332 56032 -35316
rect 55866 -35400 55882 -35366
rect 55970 -35400 55986 -35366
rect 55700 -35438 55740 -35406
rect 57096 -34479 57125 -34445
rect 57159 -34479 57217 -34445
rect 57251 -34479 57309 -34445
rect 57343 -34479 57372 -34445
rect 57129 -34529 57165 -34513
rect 57129 -34563 57131 -34529
rect 57129 -34597 57165 -34563
rect 57129 -34631 57131 -34597
rect 57201 -34529 57267 -34479
rect 57201 -34563 57217 -34529
rect 57251 -34563 57267 -34529
rect 57201 -34597 57267 -34563
rect 57201 -34631 57217 -34597
rect 57251 -34631 57267 -34597
rect 57301 -34529 57355 -34513
rect 57301 -34563 57303 -34529
rect 57337 -34563 57355 -34529
rect 57301 -34610 57355 -34563
rect 57129 -34665 57165 -34631
rect 57301 -34644 57303 -34610
rect 57337 -34644 57355 -34610
rect 57129 -34699 57264 -34665
rect 57301 -34694 57355 -34644
rect 57230 -34728 57264 -34699
rect 57117 -34744 57185 -34735
rect 57117 -34794 57118 -34744
rect 57178 -34794 57185 -34744
rect 57117 -34809 57185 -34794
rect 57230 -34744 57285 -34728
rect 57230 -34778 57251 -34744
rect 57230 -34794 57285 -34778
rect 57319 -34740 57355 -34694
rect 59662 -34429 59696 -34367
rect 59109 -34481 59125 -34447
rect 59501 -34481 59517 -34447
rect 59560 -34501 59594 -34485
rect 59560 -34551 59594 -34535
rect 59109 -34589 59125 -34555
rect 59501 -34589 59517 -34555
rect 59032 -34609 59066 -34593
rect 59032 -34659 59066 -34643
rect 59109 -34697 59125 -34663
rect 59501 -34697 59517 -34663
rect 58926 -34740 58966 -34720
rect 57319 -34780 57326 -34740
rect 58930 -34776 58964 -34740
rect 57230 -34845 57264 -34794
rect 57131 -34879 57264 -34845
rect 57319 -34854 57355 -34780
rect 57131 -34900 57165 -34879
rect 56316 -34918 56412 -34904
rect 54830 -35448 55830 -35438
rect 54830 -35470 55030 -35448
rect 53756 -35504 53852 -35470
rect 54808 -35504 55030 -35470
rect 53510 -35558 53526 -35524
rect 53614 -35558 53630 -35524
rect 53756 -35566 53790 -35504
rect 54830 -35528 55030 -35504
rect 55110 -35468 55740 -35448
rect 55810 -35468 55830 -35448
rect 56112 -35468 56146 -35406
rect 55110 -35508 55160 -35468
rect 55600 -35508 55740 -35468
rect 56050 -35502 56146 -35468
rect 55110 -35528 55740 -35508
rect 55810 -35528 55830 -35502
rect 54830 -35538 55830 -35528
rect 53464 -35608 53498 -35592
rect 53464 -36400 53498 -36384
rect 53642 -35608 53676 -35592
rect 53642 -36400 53676 -36384
rect 54870 -35566 54904 -35538
rect 53926 -35618 53942 -35584
rect 54718 -35618 54734 -35584
rect 53858 -35646 53892 -35630
rect 53858 -35750 53892 -35734
rect 54768 -35646 54802 -35630
rect 54768 -35750 54802 -35734
rect 53926 -35796 53942 -35762
rect 54718 -35796 54734 -35762
rect 53756 -35876 53790 -35814
rect 55700 -35564 55740 -35538
rect 55126 -35730 55142 -35696
rect 55494 -35730 55510 -35696
rect 54870 -35876 54904 -35814
rect 55046 -35782 55080 -35766
rect 55046 -35832 55080 -35816
rect 55556 -35782 55590 -35766
rect 55556 -35832 55590 -35816
rect 53756 -35910 53852 -35876
rect 54808 -35910 54904 -35876
rect 55126 -35902 55142 -35868
rect 55494 -35902 55510 -35868
rect 53510 -36468 53526 -36434
rect 53614 -36468 53630 -36434
rect 53350 -36536 53384 -36474
rect 53756 -36536 53790 -35910
rect 54870 -36018 54904 -35910
rect 55700 -36018 55706 -35564
rect 54870 -36024 55706 -36018
rect 54870 -36058 55262 -36024
rect 55420 -36058 55706 -36024
rect 55166 -36120 55200 -36058
rect 53350 -36570 53446 -36536
rect 53694 -36570 53790 -36536
rect 53886 -36308 53982 -36274
rect 54956 -36308 55052 -36274
rect 53886 -36370 53920 -36308
rect 55018 -36370 55052 -36308
rect 54065 -36422 54081 -36388
rect 54857 -36422 54873 -36388
rect 53988 -36450 54022 -36434
rect 53988 -36504 54022 -36488
rect 54916 -36450 54950 -36434
rect 54916 -36504 54950 -36488
rect 54065 -36550 54081 -36516
rect 54857 -36550 54873 -36516
rect 53886 -36630 53920 -36568
rect 55482 -36120 55516 -36058
rect 55280 -36148 55314 -36132
rect 55280 -36340 55314 -36324
rect 55368 -36148 55402 -36132
rect 55368 -36340 55402 -36324
rect 55308 -36408 55324 -36374
rect 55358 -36408 55374 -36374
rect 55166 -36476 55200 -36414
rect 55482 -36476 55516 -36414
rect 55166 -36510 55262 -36476
rect 55420 -36510 55516 -36476
rect 55018 -36630 55052 -36568
rect 56112 -35564 56146 -35502
rect 56350 -34938 56412 -34918
rect 56610 -34938 56706 -34904
rect 56672 -35000 56706 -34938
rect 57303 -34883 57355 -34854
rect 57131 -34955 57165 -34934
rect 57201 -34947 57217 -34913
rect 57251 -34947 57267 -34913
rect 57201 -34989 57267 -34947
rect 57337 -34917 57355 -34883
rect 57303 -34955 57355 -34917
rect 58930 -34810 59026 -34776
rect 59214 -34777 59310 -34776
rect 59662 -34777 59696 -34720
rect 59772 -34694 59866 -34660
rect 60426 -34694 60520 -34660
rect 59772 -34750 59806 -34694
rect 59214 -34810 59696 -34777
rect 58930 -34811 59696 -34810
rect 58930 -34872 58964 -34811
rect 59276 -34872 59310 -34811
rect 59087 -34912 59103 -34878
rect 59137 -34912 59153 -34878
rect 56476 -35040 56492 -35006
rect 56530 -35040 56546 -35006
rect 55866 -35604 55882 -35570
rect 55970 -35604 55986 -35570
rect 55820 -35654 55854 -35638
rect 55820 -36446 55854 -36430
rect 55998 -35654 56032 -35638
rect 55998 -36446 56032 -36430
rect 55866 -36514 55882 -36480
rect 55970 -36514 55986 -36480
rect 55706 -36582 55740 -36520
rect 56430 -35099 56464 -35083
rect 56430 -35891 56464 -35875
rect 56558 -35099 56592 -35083
rect 56558 -35891 56592 -35875
rect 56476 -35968 56492 -35934
rect 56530 -35968 56546 -35934
rect 56316 -36036 56350 -35974
rect 57096 -35023 57125 -34989
rect 57159 -35023 57217 -34989
rect 57251 -35023 57309 -34989
rect 57343 -35023 57372 -34989
rect 59044 -34971 59078 -34955
rect 59044 -35363 59078 -35347
rect 59162 -34971 59196 -34955
rect 59162 -35363 59196 -35347
rect 59087 -35440 59103 -35406
rect 59137 -35440 59153 -35406
rect 60486 -34756 60520 -34694
rect 59942 -34808 59958 -34774
rect 60334 -34808 60350 -34774
rect 59874 -34828 59908 -34812
rect 59874 -34878 59908 -34862
rect 60384 -34828 60418 -34812
rect 60384 -34878 60418 -34862
rect 59942 -34916 59958 -34882
rect 60334 -34916 60350 -34882
rect 59772 -34996 59806 -34940
rect 60486 -34996 60520 -34934
rect 59388 -35030 59476 -34996
rect 59656 -35030 59800 -34996
rect 59958 -35030 60520 -34996
rect 59388 -35090 59422 -35030
rect 59276 -35506 59310 -35446
rect 59530 -35132 59546 -35098
rect 59580 -35132 59596 -35098
rect 59502 -35182 59536 -35166
rect 59502 -35374 59536 -35358
rect 59590 -35182 59624 -35166
rect 59590 -35374 59624 -35358
rect 59530 -35442 59546 -35408
rect 59580 -35442 59596 -35408
rect 58966 -35542 59310 -35506
rect 59388 -35509 59422 -35450
rect 59704 -35509 59738 -35030
rect 60020 -35092 60054 -35030
rect 59846 -35132 59862 -35098
rect 59896 -35132 59912 -35098
rect 59818 -35182 59852 -35166
rect 59818 -35374 59852 -35358
rect 59906 -35182 59940 -35166
rect 59906 -35374 59940 -35358
rect 59846 -35442 59862 -35408
rect 59896 -35442 59912 -35408
rect 61186 -35200 61286 -35190
rect 61186 -35280 61196 -35200
rect 61186 -35290 61286 -35280
rect 60020 -35509 60054 -35448
rect 56672 -36036 56706 -35974
rect 57096 -35999 57125 -35965
rect 57159 -35999 57217 -35965
rect 57251 -35999 57309 -35965
rect 57343 -35999 57372 -35965
rect 56316 -36070 56412 -36036
rect 56610 -36070 56706 -36036
rect 57131 -36054 57165 -36033
rect 57201 -36041 57267 -35999
rect 57201 -36075 57217 -36041
rect 57251 -36075 57267 -36041
rect 57303 -36071 57355 -36033
rect 57131 -36109 57165 -36088
rect 57337 -36105 57355 -36071
rect 59276 -35602 59310 -35542
rect 59387 -35544 60054 -35509
rect 60127 -35354 60161 -35328
rect 60127 -35357 60253 -35354
rect 60161 -35373 60253 -35357
rect 60161 -35391 60203 -35373
rect 60127 -35407 60203 -35391
rect 60237 -35407 60253 -35373
rect 60359 -35360 60409 -35349
rect 60671 -35354 60705 -35328
rect 60359 -35365 60366 -35360
rect 60359 -35400 60366 -35399
rect 60406 -35400 60409 -35360
rect 60127 -35449 60161 -35407
rect 60127 -35541 60161 -35483
rect 60195 -35457 60325 -35441
rect 60195 -35491 60211 -35457
rect 60245 -35491 60325 -35457
rect 60195 -35507 60325 -35491
rect 59387 -35600 59421 -35544
rect 59087 -35642 59103 -35608
rect 59137 -35642 59153 -35608
rect 59044 -35701 59078 -35685
rect 57131 -36143 57264 -36109
rect 57303 -36134 57355 -36105
rect 57117 -36194 57185 -36179
rect 57117 -36244 57118 -36194
rect 57168 -36244 57185 -36194
rect 57117 -36253 57185 -36244
rect 57230 -36194 57264 -36143
rect 57319 -36170 57355 -36134
rect 57230 -36210 57285 -36194
rect 57230 -36244 57251 -36210
rect 57230 -36260 57285 -36244
rect 57319 -36210 57326 -36170
rect 59044 -36093 59078 -36077
rect 59162 -35701 59196 -35685
rect 59162 -36093 59196 -36077
rect 59087 -36170 59103 -36136
rect 59137 -36170 59153 -36136
rect 57230 -36289 57264 -36260
rect 57129 -36323 57264 -36289
rect 57319 -36294 57355 -36210
rect 57129 -36357 57165 -36323
rect 57301 -36344 57355 -36294
rect 58930 -36238 58964 -36176
rect 59529 -35645 59545 -35611
rect 59579 -35645 59595 -35611
rect 59501 -35695 59535 -35679
rect 59501 -35887 59535 -35871
rect 59589 -35695 59623 -35679
rect 59589 -35887 59623 -35871
rect 59529 -35955 59545 -35921
rect 59579 -35955 59595 -35921
rect 59387 -36023 59421 -35970
rect 59703 -36023 59737 -35544
rect 60019 -35605 60053 -35544
rect 59845 -35645 59861 -35611
rect 59895 -35645 59911 -35611
rect 59817 -35695 59851 -35679
rect 59817 -35887 59851 -35871
rect 59905 -35695 59939 -35679
rect 59905 -35887 59939 -35871
rect 59845 -35955 59861 -35921
rect 59895 -35955 59911 -35921
rect 60161 -35575 60203 -35541
rect 60237 -35575 60253 -35541
rect 60127 -35633 60161 -35575
rect 60289 -35609 60325 -35507
rect 60127 -35709 60161 -35667
rect 60195 -35625 60325 -35609
rect 60195 -35659 60211 -35625
rect 60245 -35659 60325 -35625
rect 60195 -35675 60325 -35659
rect 60359 -35450 60409 -35400
rect 60443 -35357 60705 -35354
rect 60443 -35373 60671 -35357
rect 60443 -35407 60459 -35373
rect 60493 -35407 60527 -35373
rect 60561 -35407 60595 -35373
rect 60629 -35391 60671 -35373
rect 60629 -35407 60705 -35391
rect 60359 -35457 60366 -35450
rect 60406 -35490 60409 -35450
rect 60393 -35491 60409 -35490
rect 60359 -35540 60409 -35491
rect 60359 -35541 60366 -35540
rect 60359 -35580 60366 -35575
rect 60406 -35580 60409 -35540
rect 60359 -35620 60409 -35580
rect 60359 -35625 60366 -35620
rect 60359 -35660 60366 -35659
rect 60406 -35660 60409 -35620
rect 60359 -35675 60409 -35660
rect 60443 -35457 60637 -35441
rect 60443 -35491 60459 -35457
rect 60493 -35491 60527 -35457
rect 60561 -35491 60595 -35457
rect 60629 -35491 60637 -35457
rect 60443 -35507 60637 -35491
rect 60671 -35449 60705 -35407
rect 60443 -35609 60477 -35507
rect 60671 -35541 60705 -35483
rect 60511 -35575 60527 -35541
rect 60561 -35575 60595 -35541
rect 60629 -35575 60671 -35541
rect 60443 -35625 60637 -35609
rect 60443 -35659 60459 -35625
rect 60493 -35659 60527 -35625
rect 60561 -35659 60595 -35625
rect 60629 -35659 60637 -35625
rect 60443 -35675 60637 -35659
rect 60671 -35633 60705 -35575
rect 60289 -35709 60325 -35675
rect 60443 -35709 60481 -35675
rect 60671 -35709 60705 -35667
rect 60127 -35725 60204 -35709
rect 60161 -35743 60204 -35725
rect 60238 -35743 60254 -35709
rect 60161 -35759 60254 -35743
rect 60289 -35725 60481 -35709
rect 60289 -35759 60297 -35725
rect 60331 -35759 60369 -35725
rect 60405 -35759 60449 -35725
rect 60579 -35743 60595 -35709
rect 60629 -35725 60705 -35709
rect 60629 -35743 60671 -35725
rect 60579 -35751 60671 -35743
rect 60127 -35788 60161 -35759
rect 60289 -35762 60481 -35759
rect 60671 -35788 60705 -35759
rect 60747 -35354 60781 -35328
rect 60747 -35357 61009 -35354
rect 60781 -35373 61009 -35357
rect 60781 -35391 60823 -35373
rect 60747 -35407 60823 -35391
rect 60857 -35407 60891 -35373
rect 60925 -35407 60959 -35373
rect 60993 -35407 61009 -35373
rect 61043 -35360 61093 -35349
rect 61291 -35354 61325 -35328
rect 61043 -35400 61046 -35360
rect 61086 -35365 61093 -35360
rect 61086 -35400 61093 -35399
rect 60747 -35449 60781 -35407
rect 60747 -35541 60781 -35483
rect 60815 -35457 61009 -35441
rect 60815 -35491 60823 -35457
rect 60857 -35491 60891 -35457
rect 60925 -35491 60959 -35457
rect 60993 -35491 61009 -35457
rect 60815 -35507 61009 -35491
rect 60781 -35575 60823 -35541
rect 60857 -35575 60891 -35541
rect 60925 -35575 60941 -35541
rect 60747 -35633 60781 -35575
rect 60975 -35609 61009 -35507
rect 60747 -35709 60781 -35667
rect 60815 -35625 61009 -35609
rect 60815 -35659 60823 -35625
rect 60857 -35659 60891 -35625
rect 60925 -35659 60959 -35625
rect 60993 -35659 61009 -35625
rect 60815 -35675 61009 -35659
rect 61043 -35450 61093 -35400
rect 61199 -35357 61325 -35354
rect 61199 -35373 61291 -35357
rect 61199 -35407 61215 -35373
rect 61249 -35391 61291 -35373
rect 61249 -35407 61325 -35391
rect 61043 -35490 61046 -35450
rect 61086 -35457 61093 -35450
rect 61043 -35491 61059 -35490
rect 61043 -35540 61093 -35491
rect 61043 -35580 61046 -35540
rect 61086 -35541 61093 -35540
rect 61086 -35580 61093 -35575
rect 61043 -35620 61093 -35580
rect 61043 -35660 61046 -35620
rect 61086 -35625 61093 -35620
rect 61086 -35660 61093 -35659
rect 61043 -35675 61093 -35660
rect 61127 -35457 61257 -35441
rect 61127 -35491 61207 -35457
rect 61241 -35491 61257 -35457
rect 61127 -35507 61257 -35491
rect 61291 -35449 61325 -35407
rect 61127 -35609 61163 -35507
rect 61291 -35541 61325 -35483
rect 61199 -35575 61215 -35541
rect 61249 -35575 61291 -35541
rect 61127 -35625 61257 -35609
rect 61127 -35659 61207 -35625
rect 61241 -35659 61257 -35625
rect 61127 -35675 61257 -35659
rect 61291 -35633 61325 -35575
rect 60971 -35709 61009 -35675
rect 61127 -35709 61163 -35675
rect 61291 -35709 61325 -35667
rect 60747 -35725 60823 -35709
rect 60781 -35743 60823 -35725
rect 60857 -35743 60873 -35709
rect 60781 -35751 60873 -35743
rect 60971 -35724 61163 -35709
rect 60971 -35725 61129 -35724
rect 60747 -35788 60781 -35759
rect 60971 -35759 60980 -35725
rect 61015 -35759 61053 -35725
rect 61088 -35758 61129 -35725
rect 61198 -35743 61214 -35709
rect 61248 -35725 61325 -35709
rect 61248 -35743 61291 -35725
rect 61088 -35759 61163 -35758
rect 61198 -35759 61291 -35743
rect 60971 -35762 61163 -35759
rect 61291 -35788 61325 -35759
rect 60466 -35860 60546 -35840
rect 60466 -35900 60486 -35860
rect 60526 -35900 60546 -35860
rect 60466 -35920 60546 -35900
rect 60606 -35860 60686 -35840
rect 60606 -35900 60626 -35860
rect 60666 -35900 60686 -35860
rect 60606 -35920 60686 -35900
rect 60746 -35860 60826 -35840
rect 60746 -35900 60766 -35860
rect 60806 -35900 60826 -35860
rect 60746 -35920 60826 -35900
rect 60886 -35860 60966 -35840
rect 60886 -35900 60906 -35860
rect 60946 -35900 60966 -35860
rect 60886 -35920 60966 -35900
rect 60019 -36023 60053 -35961
rect 59387 -36057 59476 -36023
rect 59646 -36057 59799 -36023
rect 59957 -36026 60053 -36023
rect 59957 -36057 60520 -36026
rect 59772 -36060 60520 -36057
rect 59772 -36120 59806 -36060
rect 59276 -36238 59310 -36176
rect 58930 -36272 59026 -36238
rect 59214 -36240 59310 -36238
rect 59214 -36272 59696 -36240
rect 58930 -36274 59696 -36272
rect 58930 -36310 58964 -36274
rect 57129 -36391 57131 -36357
rect 57129 -36425 57165 -36391
rect 57129 -36459 57131 -36425
rect 57129 -36475 57165 -36459
rect 57201 -36391 57217 -36357
rect 57251 -36391 57267 -36357
rect 57201 -36425 57267 -36391
rect 57201 -36459 57217 -36425
rect 57251 -36459 57267 -36425
rect 57201 -36509 57267 -36459
rect 57301 -36378 57303 -36344
rect 57337 -36378 57355 -36344
rect 57301 -36425 57355 -36378
rect 57301 -36459 57303 -36425
rect 57337 -36459 57355 -36425
rect 57301 -36475 57355 -36459
rect 59662 -36330 59696 -36274
rect 60486 -36122 60520 -36060
rect 59942 -36174 59958 -36140
rect 60334 -36174 60350 -36140
rect 59874 -36194 59908 -36178
rect 59874 -36244 59908 -36228
rect 60384 -36194 60418 -36178
rect 60384 -36244 60418 -36228
rect 59942 -36282 59958 -36248
rect 60334 -36282 60350 -36248
rect 56112 -36582 56146 -36520
rect 57096 -36543 57125 -36509
rect 57159 -36543 57217 -36509
rect 57251 -36543 57309 -36509
rect 57343 -36543 57372 -36509
rect 55706 -36616 55802 -36582
rect 56050 -36616 56146 -36582
rect 53886 -36664 53982 -36630
rect 54956 -36664 55052 -36630
rect 53886 -36726 53920 -36664
rect 55018 -36726 55052 -36664
rect 55720 -36658 56090 -36616
rect 55720 -36668 56020 -36658
rect 54065 -36778 54081 -36744
rect 54857 -36778 54873 -36744
rect 53988 -36806 54022 -36790
rect 53988 -36860 54022 -36844
rect 54916 -36806 54950 -36790
rect 54916 -36860 54950 -36844
rect 54065 -36906 54081 -36872
rect 54857 -36906 54873 -36872
rect 53886 -36986 53920 -36924
rect 56010 -36808 56020 -36668
rect 56080 -36808 56090 -36658
rect 59109 -36388 59125 -36354
rect 59501 -36388 59517 -36354
rect 59560 -36408 59594 -36392
rect 59560 -36458 59594 -36442
rect 59109 -36496 59125 -36462
rect 59501 -36496 59517 -36462
rect 59032 -36516 59066 -36500
rect 59032 -36566 59066 -36550
rect 59109 -36604 59125 -36570
rect 59501 -36604 59517 -36570
rect 56010 -36818 56090 -36808
rect 59772 -36362 59806 -36300
rect 60486 -36362 60520 -36300
rect 59772 -36396 59866 -36362
rect 60426 -36396 60520 -36362
rect 59662 -36684 59696 -36630
rect 58966 -36700 59026 -36684
rect 58930 -36718 59026 -36700
rect 59600 -36718 59696 -36684
rect 55018 -36986 55052 -36924
rect 53886 -37020 53982 -36986
rect 54956 -37020 55052 -36986
rect 55176 -36878 55272 -36844
rect 55566 -36878 55662 -36844
rect 55176 -36940 55210 -36878
rect 55628 -36940 55662 -36878
rect 55284 -36992 55300 -36958
rect 55476 -36992 55492 -36958
rect 55526 -37002 55560 -36986
rect 55284 -37080 55300 -37046
rect 55476 -37080 55492 -37046
rect 55526 -37052 55560 -37036
rect 55176 -37160 55210 -37098
rect 55628 -37160 55662 -37098
rect 55176 -37194 55272 -37160
rect 55566 -37194 55662 -37160
rect 35802 -37390 35836 -37328
rect 25780 -37430 35836 -37390
rect 35802 -37492 35836 -37430
rect 75506 -38405 75535 -38371
rect 75569 -38405 75627 -38371
rect 75661 -38405 75719 -38371
rect 75753 -38405 75811 -38371
rect 75845 -38405 75903 -38371
rect 75937 -38405 75995 -38371
rect 76029 -38405 76085 -38371
rect 76119 -38405 76177 -38371
rect 76211 -38405 76269 -38371
rect 76303 -38405 76361 -38371
rect 76395 -38405 76453 -38371
rect 76487 -38405 76545 -38371
rect 76579 -38405 76637 -38371
rect 76671 -38405 76729 -38371
rect 76763 -38405 76821 -38371
rect 76855 -38405 76884 -38371
rect 75570 -38451 75616 -38405
rect 75570 -38485 75582 -38451
rect 75570 -38519 75616 -38485
rect 75570 -38553 75582 -38519
rect 75570 -38569 75616 -38553
rect 75650 -38451 75716 -38439
rect 75650 -38485 75666 -38451
rect 75700 -38485 75716 -38451
rect 75650 -38517 75716 -38485
rect 75650 -38519 75670 -38517
rect 75650 -38553 75666 -38519
rect 75704 -38551 75716 -38517
rect 75700 -38553 75716 -38551
rect 75650 -38565 75716 -38553
rect 75570 -38610 75586 -38603
rect 75570 -38650 75580 -38610
rect 75620 -38650 75636 -38603
rect 75570 -38651 75636 -38650
rect 75670 -38609 75716 -38565
rect 75846 -38451 75892 -38405
rect 75846 -38485 75858 -38451
rect 75846 -38519 75892 -38485
rect 75846 -38553 75858 -38519
rect 75846 -38569 75892 -38553
rect 75926 -38451 75992 -38439
rect 75926 -38485 75942 -38451
rect 75976 -38485 75992 -38451
rect 75926 -38519 75992 -38485
rect 75926 -38554 75942 -38519
rect 75976 -38554 75992 -38519
rect 75926 -38565 75992 -38554
rect 75704 -38643 75716 -38609
rect 75670 -38685 75716 -38643
rect 75846 -38637 75862 -38603
rect 75896 -38637 75912 -38603
rect 75846 -38651 75912 -38637
rect 75946 -38609 75992 -38565
rect 76120 -38451 76166 -38405
rect 76120 -38485 76132 -38451
rect 76120 -38519 76166 -38485
rect 76120 -38553 76132 -38519
rect 76120 -38569 76166 -38553
rect 76200 -38451 76266 -38439
rect 76200 -38485 76216 -38451
rect 76250 -38485 76266 -38451
rect 76200 -38519 76266 -38485
rect 76200 -38553 76216 -38519
rect 76251 -38553 76266 -38519
rect 76200 -38565 76266 -38553
rect 75946 -38643 75947 -38609
rect 75981 -38643 75992 -38609
rect 75946 -38685 75992 -38643
rect 76120 -38610 76136 -38603
rect 76120 -38644 76128 -38610
rect 76170 -38637 76186 -38603
rect 76162 -38644 76186 -38637
rect 76120 -38651 76186 -38644
rect 76220 -38610 76266 -38565
rect 76396 -38451 76442 -38405
rect 76396 -38485 76408 -38451
rect 76396 -38519 76442 -38485
rect 76396 -38553 76408 -38519
rect 76396 -38569 76442 -38553
rect 76476 -38451 76542 -38439
rect 76476 -38485 76492 -38451
rect 76526 -38485 76542 -38451
rect 76476 -38519 76542 -38485
rect 76476 -38553 76492 -38519
rect 76526 -38553 76542 -38519
rect 76476 -38565 76542 -38553
rect 76220 -38644 76224 -38610
rect 76258 -38644 76266 -38610
rect 76220 -38685 76266 -38644
rect 76396 -38609 76412 -38603
rect 76396 -38643 76404 -38609
rect 76446 -38637 76462 -38603
rect 76438 -38643 76462 -38637
rect 76396 -38651 76462 -38643
rect 76496 -38609 76542 -38565
rect 76672 -38451 76718 -38405
rect 76672 -38485 76684 -38451
rect 76672 -38519 76718 -38485
rect 76672 -38553 76684 -38519
rect 76672 -38569 76718 -38553
rect 76752 -38451 76818 -38439
rect 76752 -38485 76768 -38451
rect 76802 -38485 76818 -38451
rect 76752 -38519 76818 -38485
rect 76752 -38555 76768 -38519
rect 76802 -38555 76818 -38519
rect 76752 -38565 76818 -38555
rect 76496 -38643 76497 -38609
rect 76531 -38643 76542 -38609
rect 76496 -38685 76542 -38643
rect 76672 -38609 76688 -38603
rect 76672 -38643 76680 -38609
rect 76722 -38637 76738 -38603
rect 76714 -38643 76738 -38637
rect 76672 -38651 76738 -38643
rect 76772 -38610 76818 -38565
rect 76806 -38644 76818 -38610
rect 76772 -38685 76818 -38644
rect 75574 -38703 75616 -38687
rect 75574 -38737 75582 -38703
rect 75574 -38771 75616 -38737
rect 75574 -38805 75582 -38771
rect 75574 -38839 75616 -38805
rect 75574 -38873 75582 -38839
rect 75574 -38915 75616 -38873
rect 75650 -38698 75716 -38685
rect 75650 -38703 75670 -38698
rect 75650 -38737 75666 -38703
rect 75704 -38732 75716 -38698
rect 75700 -38737 75716 -38732
rect 75650 -38771 75716 -38737
rect 75650 -38805 75666 -38771
rect 75700 -38805 75716 -38771
rect 75650 -38839 75716 -38805
rect 75650 -38873 75666 -38839
rect 75700 -38873 75716 -38839
rect 75650 -38881 75716 -38873
rect 75850 -38703 75892 -38687
rect 75850 -38737 75858 -38703
rect 75850 -38771 75892 -38737
rect 75850 -38805 75858 -38771
rect 75850 -38839 75892 -38805
rect 75850 -38873 75858 -38839
rect 75850 -38915 75892 -38873
rect 75926 -38703 75992 -38685
rect 75926 -38737 75942 -38703
rect 75977 -38737 75992 -38703
rect 75926 -38771 75992 -38737
rect 75926 -38805 75942 -38771
rect 75976 -38805 75992 -38771
rect 75926 -38839 75992 -38805
rect 75926 -38873 75942 -38839
rect 75976 -38873 75992 -38839
rect 75926 -38881 75992 -38873
rect 76124 -38703 76166 -38687
rect 76124 -38737 76132 -38703
rect 76124 -38771 76166 -38737
rect 76124 -38805 76132 -38771
rect 76124 -38839 76166 -38805
rect 76124 -38873 76132 -38839
rect 76124 -38915 76166 -38873
rect 76200 -38703 76266 -38685
rect 76200 -38704 76216 -38703
rect 76200 -38738 76215 -38704
rect 76250 -38737 76266 -38703
rect 76249 -38738 76266 -38737
rect 76200 -38771 76266 -38738
rect 76200 -38805 76216 -38771
rect 76250 -38776 76266 -38771
rect 76200 -38810 76218 -38805
rect 76252 -38810 76266 -38776
rect 76200 -38839 76266 -38810
rect 76200 -38873 76216 -38839
rect 76250 -38873 76266 -38839
rect 76200 -38881 76266 -38873
rect 76400 -38703 76442 -38687
rect 76400 -38737 76408 -38703
rect 76400 -38771 76442 -38737
rect 76400 -38805 76408 -38771
rect 76400 -38839 76442 -38805
rect 76400 -38873 76408 -38839
rect 76400 -38915 76442 -38873
rect 76476 -38703 76542 -38685
rect 76476 -38737 76492 -38703
rect 76526 -38737 76542 -38703
rect 76476 -38771 76542 -38737
rect 76476 -38805 76492 -38771
rect 76526 -38805 76542 -38771
rect 76476 -38839 76542 -38805
rect 76476 -38873 76492 -38839
rect 76526 -38873 76542 -38839
rect 76476 -38881 76542 -38873
rect 76676 -38703 76718 -38687
rect 76676 -38737 76684 -38703
rect 76676 -38771 76718 -38737
rect 76676 -38805 76684 -38771
rect 76676 -38839 76718 -38805
rect 76676 -38873 76684 -38839
rect 76676 -38915 76718 -38873
rect 76752 -38703 76818 -38685
rect 76752 -38737 76768 -38703
rect 76802 -38737 76818 -38703
rect 76752 -38771 76818 -38737
rect 76752 -38805 76768 -38771
rect 76802 -38805 76818 -38771
rect 76752 -38839 76818 -38805
rect 76752 -38873 76768 -38839
rect 76802 -38873 76818 -38839
rect 76752 -38881 76818 -38873
rect 35802 -38990 35836 -38928
rect 75506 -38949 75535 -38915
rect 75569 -38949 75627 -38915
rect 75661 -38949 75719 -38915
rect 75753 -38949 75811 -38915
rect 75845 -38949 75903 -38915
rect 75937 -38949 75995 -38915
rect 76029 -38949 76085 -38915
rect 76119 -38949 76177 -38915
rect 76211 -38949 76269 -38915
rect 76303 -38949 76361 -38915
rect 76395 -38949 76453 -38915
rect 76487 -38949 76545 -38915
rect 76579 -38949 76637 -38915
rect 76671 -38949 76729 -38915
rect 76763 -38949 76821 -38915
rect 76855 -38949 76884 -38915
rect 25780 -38998 35836 -38990
rect 25780 -39032 35838 -38998
rect 35804 -39094 35838 -39032
rect 77578 -39075 77607 -39041
rect 77641 -39075 77699 -39041
rect 77733 -39075 77791 -39041
rect 77825 -39075 77883 -39041
rect 77917 -39075 77975 -39041
rect 78009 -39075 78067 -39041
rect 78101 -39075 78159 -39041
rect 78193 -39075 78251 -39041
rect 78285 -39075 78343 -39041
rect 78377 -39075 78435 -39041
rect 78469 -39075 78527 -39041
rect 78561 -39075 78619 -39041
rect 78653 -39075 78711 -39041
rect 78745 -39075 78803 -39041
rect 78837 -39075 78895 -39041
rect 78929 -39075 78987 -39041
rect 79021 -39075 79050 -39041
rect 77961 -39117 78017 -39075
rect 77596 -39120 77927 -39119
rect 77410 -39129 77927 -39120
rect 77410 -39130 77835 -39129
rect 77410 -39170 77430 -39130
rect 77520 -39163 77835 -39130
rect 77869 -39163 77927 -39129
rect 77520 -39170 77927 -39163
rect 77410 -39180 77540 -39170
rect 77596 -39177 77927 -39170
rect 77961 -39151 77974 -39117
rect 78008 -39151 78017 -39117
rect 77961 -39185 78017 -39151
rect 77596 -39245 77914 -39211
rect 77961 -39219 77974 -39185
rect 78008 -39219 78017 -39185
rect 77961 -39235 78017 -39219
rect 78059 -39120 78113 -39109
rect 78419 -39117 78475 -39075
rect 78147 -39120 78385 -39119
rect 78059 -39129 78385 -39120
rect 78059 -39148 78293 -39129
rect 78093 -39163 78293 -39148
rect 78327 -39163 78385 -39129
rect 78093 -39170 78385 -39163
rect 78093 -39182 78113 -39170
rect 78147 -39177 78385 -39170
rect 78419 -39151 78432 -39117
rect 78466 -39151 78475 -39117
rect 78059 -39216 78113 -39182
rect 78419 -39185 78475 -39151
rect 77596 -39248 77660 -39245
rect 77596 -39282 77613 -39248
rect 77647 -39282 77660 -39248
rect 77880 -39269 77914 -39245
rect 78093 -39250 78113 -39216
rect 77596 -39303 77660 -39282
rect 77700 -39280 77842 -39279
rect 77700 -39320 77780 -39280
rect 77820 -39320 77842 -39280
rect 77880 -39303 78025 -39269
rect 78059 -39303 78113 -39250
rect 78151 -39245 78385 -39211
rect 78419 -39219 78432 -39185
rect 78466 -39219 78475 -39185
rect 78419 -39235 78475 -39219
rect 78517 -39148 78572 -39109
rect 78551 -39182 78572 -39148
rect 78517 -39216 78572 -39182
rect 78647 -39159 78703 -39075
rect 78837 -39117 78903 -39075
rect 78647 -39193 78661 -39159
rect 78695 -39193 78703 -39159
rect 78647 -39209 78703 -39193
rect 78737 -39159 78797 -39143
rect 78737 -39193 78745 -39159
rect 78779 -39193 78797 -39159
rect 78151 -39248 78216 -39245
rect 78151 -39282 78167 -39248
rect 78201 -39282 78216 -39248
rect 78351 -39269 78385 -39245
rect 78551 -39250 78572 -39216
rect 78517 -39260 78572 -39250
rect 78737 -39253 78797 -39193
rect 78837 -39151 78853 -39117
rect 78887 -39151 78903 -39117
rect 78837 -39185 78903 -39151
rect 78837 -39219 78853 -39185
rect 78887 -39219 78903 -39185
rect 78941 -39110 79033 -39109
rect 78941 -39117 79170 -39110
rect 78941 -39151 78957 -39117
rect 78991 -39151 79170 -39117
rect 80738 -39125 80767 -39091
rect 80801 -39125 80859 -39091
rect 80893 -39125 80951 -39091
rect 80985 -39125 81043 -39091
rect 81077 -39125 81135 -39091
rect 81169 -39125 81227 -39091
rect 81261 -39125 81319 -39091
rect 81353 -39125 81411 -39091
rect 81445 -39125 81503 -39091
rect 81537 -39125 81595 -39091
rect 81629 -39125 81687 -39091
rect 81721 -39125 81779 -39091
rect 81813 -39125 81871 -39091
rect 81905 -39125 81963 -39091
rect 81997 -39125 82055 -39091
rect 82089 -39125 82147 -39091
rect 82181 -39125 82239 -39091
rect 82273 -39125 82331 -39091
rect 82365 -39125 82423 -39091
rect 82457 -39125 82515 -39091
rect 82549 -39125 82607 -39091
rect 82641 -39125 82699 -39091
rect 82733 -39125 82791 -39091
rect 82825 -39125 82883 -39091
rect 82917 -39125 82975 -39091
rect 83009 -39125 83067 -39091
rect 83101 -39125 83159 -39091
rect 83193 -39125 83251 -39091
rect 83285 -39125 83343 -39091
rect 83377 -39125 83435 -39091
rect 83469 -39125 83527 -39091
rect 83561 -39125 83619 -39091
rect 83653 -39125 83711 -39091
rect 83745 -39125 83803 -39091
rect 83837 -39125 83895 -39091
rect 83929 -39125 83987 -39091
rect 84021 -39125 84079 -39091
rect 84113 -39125 84171 -39091
rect 84205 -39125 84263 -39091
rect 84297 -39125 84355 -39091
rect 84389 -39125 84447 -39091
rect 84481 -39125 84539 -39091
rect 84573 -39125 84631 -39091
rect 84665 -39125 84723 -39091
rect 84757 -39125 84815 -39091
rect 84849 -39125 84907 -39091
rect 84941 -39125 84999 -39091
rect 85033 -39125 85091 -39091
rect 85125 -39125 85183 -39091
rect 85217 -39125 85275 -39091
rect 85309 -39125 85367 -39091
rect 85401 -39125 85459 -39091
rect 85493 -39125 85551 -39091
rect 85585 -39125 85643 -39091
rect 85677 -39125 85735 -39091
rect 85769 -39125 85827 -39091
rect 85861 -39125 85919 -39091
rect 85953 -39125 86011 -39091
rect 86045 -39125 86103 -39091
rect 86137 -39125 86195 -39091
rect 86229 -39125 86287 -39091
rect 86321 -39125 86379 -39091
rect 86413 -39125 86471 -39091
rect 86505 -39125 86563 -39091
rect 86597 -39125 86655 -39091
rect 86689 -39125 86747 -39091
rect 86781 -39125 86839 -39091
rect 86873 -39125 86931 -39091
rect 86965 -39125 87023 -39091
rect 87057 -39125 87115 -39091
rect 87149 -39125 87207 -39091
rect 87241 -39125 87299 -39091
rect 87333 -39125 87391 -39091
rect 87425 -39125 87483 -39091
rect 87517 -39125 87575 -39091
rect 87609 -39125 87667 -39091
rect 87701 -39125 87759 -39091
rect 87793 -39125 87851 -39091
rect 87885 -39125 87943 -39091
rect 87977 -39125 88035 -39091
rect 88069 -39125 88127 -39091
rect 88161 -39125 88219 -39091
rect 88253 -39125 88311 -39091
rect 88345 -39125 88403 -39091
rect 88437 -39125 88495 -39091
rect 88529 -39125 88587 -39091
rect 88621 -39125 88679 -39091
rect 88713 -39125 88771 -39091
rect 88805 -39125 88834 -39091
rect 78941 -39185 79170 -39151
rect 78941 -39219 78957 -39185
rect 78991 -39219 79170 -39185
rect 78151 -39303 78216 -39282
rect 77596 -39340 77666 -39337
rect 77220 -39353 77666 -39340
rect 53896 -39392 53992 -39358
rect 54966 -39392 55062 -39358
rect 53896 -39454 53930 -39392
rect 55028 -39454 55062 -39392
rect 54075 -39506 54091 -39472
rect 54867 -39506 54883 -39472
rect 53998 -39534 54032 -39518
rect 53998 -39588 54032 -39572
rect 54926 -39534 54960 -39518
rect 54926 -39588 54960 -39572
rect 54075 -39634 54091 -39600
rect 54867 -39634 54883 -39600
rect 53896 -39714 53930 -39652
rect 77220 -39387 77613 -39353
rect 77647 -39387 77666 -39353
rect 77220 -39410 77666 -39387
rect 77700 -39353 77842 -39320
rect 77991 -39337 78025 -39303
rect 77700 -39387 77739 -39353
rect 77773 -39387 77842 -39353
rect 77700 -39403 77842 -39387
rect 77876 -39350 77957 -39337
rect 77876 -39390 77900 -39350
rect 77940 -39353 77957 -39350
rect 77949 -39387 77957 -39353
rect 77940 -39390 77957 -39387
rect 77876 -39403 77957 -39390
rect 77991 -39353 78045 -39337
rect 77991 -39387 78011 -39353
rect 77991 -39403 78045 -39387
rect 77220 -39450 77320 -39410
rect 77220 -39490 77240 -39450
rect 77300 -39490 77320 -39450
rect 77596 -39451 77666 -39410
rect 77991 -39437 78025 -39403
rect 77220 -39520 77320 -39490
rect 77703 -39471 78025 -39437
rect 78079 -39450 78113 -39303
rect 78250 -39337 78289 -39279
rect 78351 -39303 78483 -39269
rect 78517 -39303 78670 -39260
rect 78737 -39287 78925 -39253
rect 78449 -39337 78483 -39303
rect 78538 -39330 78670 -39303
rect 78147 -39350 78216 -39337
rect 78147 -39390 78160 -39350
rect 78200 -39390 78216 -39350
rect 78147 -39403 78216 -39390
rect 78250 -39350 78415 -39337
rect 78250 -39390 78290 -39350
rect 78330 -39390 78370 -39350
rect 78410 -39390 78415 -39350
rect 78250 -39403 78415 -39390
rect 78449 -39353 78504 -39337
rect 78449 -39387 78470 -39353
rect 78449 -39403 78504 -39387
rect 78538 -39370 78590 -39330
rect 78630 -39337 78670 -39330
rect 78891 -39337 78925 -39287
rect 78630 -39353 78745 -39337
rect 78630 -39370 78664 -39353
rect 78538 -39387 78664 -39370
rect 78698 -39387 78745 -39353
rect 78789 -39340 78857 -39337
rect 78789 -39380 78800 -39340
rect 78850 -39380 78857 -39340
rect 78789 -39387 78805 -39380
rect 78839 -39387 78857 -39380
rect 78891 -39353 78949 -39337
rect 78891 -39387 78913 -39353
rect 78947 -39387 78949 -39353
rect 78538 -39390 78610 -39387
rect 78449 -39437 78483 -39403
rect 78059 -39467 78113 -39450
rect 55028 -39714 55062 -39652
rect 77597 -39519 77613 -39485
rect 77647 -39519 77663 -39485
rect 77597 -39585 77663 -39519
rect 77703 -39491 77737 -39471
rect 77877 -39491 77911 -39471
rect 77703 -39541 77737 -39525
rect 77777 -39539 77793 -39505
rect 77827 -39539 77843 -39505
rect 77777 -39585 77843 -39539
rect 78093 -39501 78113 -39467
rect 77877 -39541 77911 -39525
rect 77945 -39539 77971 -39505
rect 78005 -39539 78021 -39505
rect 78059 -39519 78113 -39501
rect 78150 -39471 78483 -39437
rect 78538 -39450 78572 -39390
rect 78891 -39403 78949 -39387
rect 78983 -39340 79170 -39219
rect 80806 -39167 80848 -39125
rect 80806 -39201 80814 -39167
rect 80806 -39235 80848 -39201
rect 80806 -39269 80814 -39235
rect 80806 -39303 80848 -39269
rect 78983 -39400 79080 -39340
rect 79140 -39400 79170 -39340
rect 78891 -39421 78925 -39403
rect 78517 -39467 78572 -39450
rect 78150 -39491 78201 -39471
rect 77945 -39585 78021 -39539
rect 78150 -39525 78167 -39491
rect 78335 -39491 78369 -39471
rect 78150 -39541 78201 -39525
rect 78235 -39539 78251 -39505
rect 78285 -39539 78301 -39505
rect 78235 -39585 78301 -39539
rect 78551 -39501 78572 -39467
rect 78335 -39541 78369 -39525
rect 78403 -39539 78429 -39505
rect 78463 -39539 78479 -39505
rect 78517 -39519 78572 -39501
rect 78647 -39459 78925 -39421
rect 78983 -39450 79170 -39400
rect 78647 -39481 78713 -39459
rect 78647 -39515 78661 -39481
rect 78695 -39515 78713 -39481
rect 78983 -39493 79080 -39450
rect 78647 -39531 78713 -39515
rect 78837 -39509 78887 -39493
rect 78403 -39585 78479 -39539
rect 78837 -39543 78853 -39509
rect 78837 -39585 78887 -39543
rect 78921 -39509 79080 -39493
rect 78921 -39543 78937 -39509
rect 78971 -39510 79080 -39509
rect 79140 -39510 79170 -39450
rect 78971 -39543 79170 -39510
rect 80460 -39350 80750 -39330
rect 80460 -39510 80480 -39350
rect 80640 -39390 80750 -39350
rect 80806 -39337 80814 -39303
rect 80806 -39353 80848 -39337
rect 80882 -39167 80948 -39159
rect 80882 -39201 80898 -39167
rect 80932 -39201 80948 -39167
rect 80882 -39235 80948 -39201
rect 80882 -39269 80898 -39235
rect 80932 -39269 80948 -39235
rect 80882 -39303 80948 -39269
rect 80882 -39337 80898 -39303
rect 80932 -39337 80948 -39303
rect 80882 -39355 80948 -39337
rect 81040 -39167 81093 -39125
rect 81040 -39201 81059 -39167
rect 81040 -39235 81093 -39201
rect 81040 -39269 81059 -39235
rect 81040 -39303 81093 -39269
rect 81040 -39337 81059 -39303
rect 81040 -39353 81093 -39337
rect 81127 -39167 81193 -39159
rect 81127 -39201 81143 -39167
rect 81177 -39201 81193 -39167
rect 81127 -39235 81193 -39201
rect 81127 -39269 81143 -39235
rect 81177 -39269 81193 -39235
rect 81127 -39303 81193 -39269
rect 81227 -39167 81261 -39125
rect 81227 -39235 81261 -39201
rect 81227 -39285 81261 -39269
rect 81295 -39167 81361 -39159
rect 81295 -39201 81311 -39167
rect 81345 -39201 81361 -39167
rect 81295 -39235 81361 -39201
rect 81395 -39167 81437 -39125
rect 81429 -39201 81437 -39167
rect 81395 -39217 81437 -39201
rect 81514 -39167 81556 -39125
rect 81514 -39201 81522 -39167
rect 81295 -39269 81311 -39235
rect 81345 -39269 81361 -39235
rect 81127 -39337 81143 -39303
rect 81177 -39319 81193 -39303
rect 81295 -39303 81361 -39269
rect 81295 -39319 81311 -39303
rect 81177 -39337 81311 -39319
rect 81345 -39315 81361 -39303
rect 81514 -39235 81556 -39201
rect 81514 -39269 81522 -39235
rect 81514 -39305 81556 -39269
rect 81345 -39337 81448 -39315
rect 81127 -39353 81448 -39337
rect 80902 -39380 80948 -39355
rect 81395 -39380 81448 -39353
rect 81514 -39339 81522 -39305
rect 81514 -39355 81556 -39339
rect 81590 -39167 81656 -39159
rect 81590 -39201 81606 -39167
rect 81640 -39201 81656 -39167
rect 81590 -39235 81656 -39201
rect 81590 -39269 81606 -39235
rect 81640 -39269 81656 -39235
rect 81590 -39305 81656 -39269
rect 81690 -39167 81724 -39125
rect 81690 -39235 81724 -39201
rect 81690 -39285 81724 -39269
rect 81758 -39167 81824 -39159
rect 81758 -39201 81774 -39167
rect 81808 -39201 81824 -39167
rect 81758 -39235 81824 -39201
rect 81758 -39269 81774 -39235
rect 81808 -39269 81824 -39235
rect 81590 -39339 81606 -39305
rect 81640 -39319 81656 -39305
rect 81758 -39305 81824 -39269
rect 81858 -39167 81892 -39125
rect 81858 -39235 81892 -39201
rect 81858 -39285 81892 -39269
rect 81926 -39167 81992 -39159
rect 81926 -39201 81942 -39167
rect 81976 -39201 81992 -39167
rect 81926 -39235 81992 -39201
rect 81926 -39269 81942 -39235
rect 81976 -39269 81992 -39235
rect 81758 -39319 81774 -39305
rect 81640 -39339 81774 -39319
rect 81808 -39319 81824 -39305
rect 81926 -39305 81992 -39269
rect 82026 -39167 82060 -39125
rect 82026 -39235 82060 -39201
rect 82026 -39285 82060 -39269
rect 82094 -39167 82160 -39159
rect 82094 -39201 82110 -39167
rect 82144 -39201 82160 -39167
rect 82094 -39235 82160 -39201
rect 82094 -39269 82110 -39235
rect 82144 -39269 82160 -39235
rect 81926 -39319 81942 -39305
rect 81808 -39339 81942 -39319
rect 81976 -39319 81992 -39305
rect 82094 -39305 82160 -39269
rect 82194 -39167 82228 -39125
rect 82194 -39235 82228 -39201
rect 82194 -39285 82228 -39269
rect 82262 -39167 82328 -39159
rect 82262 -39201 82278 -39167
rect 82312 -39201 82328 -39167
rect 82262 -39235 82328 -39201
rect 82262 -39269 82278 -39235
rect 82312 -39269 82328 -39235
rect 82094 -39319 82110 -39305
rect 81976 -39339 82110 -39319
rect 82144 -39319 82160 -39305
rect 82262 -39305 82328 -39269
rect 82362 -39167 82396 -39125
rect 82362 -39235 82396 -39201
rect 82362 -39285 82396 -39269
rect 82430 -39167 82496 -39159
rect 82430 -39201 82446 -39167
rect 82480 -39201 82496 -39167
rect 82430 -39235 82496 -39201
rect 82430 -39269 82446 -39235
rect 82480 -39269 82496 -39235
rect 82262 -39319 82278 -39305
rect 82144 -39339 82278 -39319
rect 82312 -39319 82328 -39305
rect 82430 -39305 82496 -39269
rect 82530 -39167 82564 -39125
rect 82530 -39235 82564 -39201
rect 82530 -39285 82564 -39269
rect 82598 -39167 82664 -39159
rect 82598 -39201 82614 -39167
rect 82648 -39201 82664 -39167
rect 82598 -39235 82664 -39201
rect 82598 -39269 82614 -39235
rect 82648 -39269 82664 -39235
rect 82430 -39319 82446 -39305
rect 82312 -39339 82446 -39319
rect 82480 -39319 82496 -39305
rect 82598 -39305 82664 -39269
rect 82698 -39167 82732 -39125
rect 82698 -39235 82732 -39201
rect 82698 -39285 82732 -39269
rect 82766 -39167 82832 -39159
rect 82766 -39201 82782 -39167
rect 82816 -39201 82832 -39167
rect 82766 -39235 82832 -39201
rect 82766 -39240 82782 -39235
rect 82816 -39240 82832 -39235
rect 82766 -39280 82780 -39240
rect 82820 -39280 82832 -39240
rect 82598 -39319 82614 -39305
rect 82480 -39339 82614 -39319
rect 82648 -39319 82664 -39305
rect 82766 -39305 82832 -39280
rect 82866 -39167 82908 -39125
rect 82900 -39201 82908 -39167
rect 82866 -39235 82908 -39201
rect 82900 -39269 82908 -39235
rect 82866 -39285 82908 -39269
rect 82986 -39167 83028 -39125
rect 82986 -39201 82994 -39167
rect 82986 -39235 83028 -39201
rect 82986 -39269 82994 -39235
rect 82766 -39319 82782 -39305
rect 82648 -39320 82782 -39319
rect 82816 -39320 82832 -39305
rect 82648 -39339 82780 -39320
rect 81590 -39353 82780 -39339
rect 82766 -39360 82780 -39353
rect 82820 -39360 82832 -39320
rect 82986 -39305 83028 -39269
rect 82986 -39339 82994 -39305
rect 82986 -39355 83028 -39339
rect 83062 -39167 83128 -39159
rect 83062 -39201 83078 -39167
rect 83112 -39201 83128 -39167
rect 83062 -39235 83128 -39201
rect 83062 -39269 83078 -39235
rect 83112 -39269 83128 -39235
rect 83062 -39305 83128 -39269
rect 83162 -39167 83196 -39125
rect 83162 -39235 83196 -39201
rect 83162 -39285 83196 -39269
rect 83230 -39167 83296 -39159
rect 83230 -39201 83246 -39167
rect 83280 -39201 83296 -39167
rect 83230 -39235 83296 -39201
rect 83230 -39269 83246 -39235
rect 83280 -39269 83296 -39235
rect 83062 -39339 83078 -39305
rect 83112 -39319 83128 -39305
rect 83230 -39305 83296 -39269
rect 83330 -39167 83364 -39125
rect 83330 -39235 83364 -39201
rect 83330 -39285 83364 -39269
rect 83398 -39167 83464 -39159
rect 83398 -39201 83414 -39167
rect 83448 -39201 83464 -39167
rect 83398 -39235 83464 -39201
rect 83398 -39269 83414 -39235
rect 83448 -39269 83464 -39235
rect 83230 -39319 83246 -39305
rect 83112 -39339 83246 -39319
rect 83280 -39319 83296 -39305
rect 83398 -39305 83464 -39269
rect 83498 -39167 83532 -39125
rect 83498 -39235 83532 -39201
rect 83498 -39285 83532 -39269
rect 83566 -39167 83632 -39159
rect 83566 -39201 83582 -39167
rect 83616 -39201 83632 -39167
rect 83566 -39235 83632 -39201
rect 83566 -39269 83582 -39235
rect 83616 -39269 83632 -39235
rect 83398 -39319 83414 -39305
rect 83280 -39339 83414 -39319
rect 83448 -39319 83464 -39305
rect 83566 -39305 83632 -39269
rect 83666 -39167 83700 -39125
rect 83666 -39235 83700 -39201
rect 83666 -39285 83700 -39269
rect 83734 -39167 83800 -39159
rect 83734 -39201 83750 -39167
rect 83784 -39201 83800 -39167
rect 83734 -39235 83800 -39201
rect 83734 -39269 83750 -39235
rect 83784 -39269 83800 -39235
rect 83566 -39319 83582 -39305
rect 83448 -39339 83582 -39319
rect 83616 -39319 83632 -39305
rect 83734 -39305 83800 -39269
rect 83834 -39167 83868 -39125
rect 83834 -39235 83868 -39201
rect 83834 -39285 83868 -39269
rect 83902 -39167 83968 -39159
rect 83902 -39201 83918 -39167
rect 83952 -39201 83968 -39167
rect 83902 -39235 83968 -39201
rect 83902 -39269 83918 -39235
rect 83952 -39269 83968 -39235
rect 83734 -39319 83750 -39305
rect 83616 -39339 83750 -39319
rect 83784 -39319 83800 -39305
rect 83902 -39305 83968 -39269
rect 84002 -39167 84036 -39125
rect 84002 -39235 84036 -39201
rect 84002 -39285 84036 -39269
rect 84070 -39167 84136 -39159
rect 84070 -39201 84086 -39167
rect 84120 -39201 84136 -39167
rect 84070 -39235 84136 -39201
rect 84070 -39269 84086 -39235
rect 84120 -39269 84136 -39235
rect 83902 -39319 83918 -39305
rect 83784 -39339 83918 -39319
rect 83952 -39319 83968 -39305
rect 84070 -39305 84136 -39269
rect 84170 -39167 84204 -39125
rect 84170 -39235 84204 -39201
rect 84170 -39285 84204 -39269
rect 84238 -39167 84304 -39159
rect 84238 -39201 84254 -39167
rect 84288 -39201 84304 -39167
rect 84238 -39235 84304 -39201
rect 84238 -39260 84254 -39235
rect 84288 -39260 84304 -39235
rect 84070 -39319 84086 -39305
rect 83952 -39339 84086 -39319
rect 84120 -39319 84136 -39305
rect 84238 -39319 84250 -39260
rect 84120 -39339 84250 -39319
rect 83062 -39353 84250 -39339
rect 80802 -39390 80868 -39389
rect 80640 -39403 80868 -39390
rect 80640 -39430 80818 -39403
rect 80640 -39510 80750 -39430
rect 80802 -39437 80818 -39430
rect 80852 -39437 80868 -39403
rect 80902 -39390 80950 -39380
rect 81035 -39390 81361 -39387
rect 80902 -39403 81361 -39390
rect 80902 -39437 81051 -39403
rect 81085 -39437 81143 -39403
rect 81177 -39437 81227 -39403
rect 81261 -39437 81311 -39403
rect 81345 -39437 81361 -39403
rect 81395 -39390 81450 -39380
rect 81491 -39390 82579 -39389
rect 81395 -39403 82579 -39390
rect 81395 -39437 81516 -39403
rect 81550 -39437 81690 -39403
rect 81724 -39437 81858 -39403
rect 81892 -39437 82027 -39403
rect 82061 -39437 82194 -39403
rect 82228 -39437 82362 -39403
rect 82396 -39437 82529 -39403
rect 82563 -39437 82579 -39403
rect 82766 -39400 82832 -39360
rect 80902 -39440 81110 -39437
rect 81395 -39440 81560 -39437
rect 82766 -39440 82780 -39400
rect 82820 -39440 82832 -39400
rect 82963 -39394 84051 -39389
rect 82963 -39403 83368 -39394
rect 83773 -39403 84051 -39394
rect 82963 -39437 82988 -39403
rect 83022 -39437 83162 -39403
rect 83196 -39437 83330 -39403
rect 83364 -39434 83368 -39403
rect 83773 -39434 83834 -39403
rect 83364 -39437 83499 -39434
rect 83533 -39437 83666 -39434
rect 83700 -39437 83834 -39434
rect 83868 -39437 84001 -39403
rect 84035 -39437 84051 -39403
rect 80460 -39530 80750 -39510
rect 80802 -39487 80848 -39471
rect 80902 -39475 80948 -39440
rect 81395 -39471 81448 -39440
rect 82766 -39471 82832 -39440
rect 84238 -39471 84250 -39353
rect 80802 -39521 80814 -39487
rect 78921 -39550 79170 -39543
rect 78921 -39551 79033 -39550
rect 80802 -39555 80848 -39521
rect 77578 -39619 77607 -39585
rect 77641 -39619 77699 -39585
rect 77733 -39619 77791 -39585
rect 77825 -39619 77883 -39585
rect 77917 -39619 77975 -39585
rect 78009 -39619 78067 -39585
rect 78101 -39619 78159 -39585
rect 78193 -39619 78251 -39585
rect 78285 -39619 78343 -39585
rect 78377 -39619 78435 -39585
rect 78469 -39619 78527 -39585
rect 78561 -39619 78619 -39585
rect 78653 -39619 78711 -39585
rect 78745 -39619 78803 -39585
rect 78837 -39619 78895 -39585
rect 78929 -39619 78987 -39585
rect 79021 -39619 79050 -39585
rect 80802 -39589 80814 -39555
rect 80802 -39635 80848 -39589
rect 80882 -39487 80948 -39475
rect 80882 -39521 80898 -39487
rect 80932 -39521 80948 -39487
rect 80882 -39555 80948 -39521
rect 81127 -39507 81448 -39471
rect 81510 -39491 81556 -39475
rect 80882 -39589 80898 -39555
rect 80932 -39589 80948 -39555
rect 80882 -39601 80948 -39589
rect 81040 -39559 81093 -39543
rect 81040 -39593 81059 -39559
rect 81040 -39635 81093 -39593
rect 81127 -39551 81193 -39507
rect 81127 -39585 81143 -39551
rect 81177 -39585 81193 -39551
rect 81127 -39601 81193 -39585
rect 81227 -39559 81261 -39543
rect 81227 -39635 81261 -39593
rect 81295 -39551 81361 -39507
rect 81510 -39525 81522 -39491
rect 81295 -39585 81311 -39551
rect 81345 -39585 81361 -39551
rect 81295 -39601 81361 -39585
rect 81395 -39558 81445 -39542
rect 81429 -39592 81445 -39558
rect 81395 -39635 81445 -39592
rect 81510 -39559 81556 -39525
rect 81510 -39593 81522 -39559
rect 81510 -39635 81556 -39593
rect 81590 -39490 82832 -39471
rect 81590 -39491 82780 -39490
rect 81590 -39525 81606 -39491
rect 81640 -39509 81774 -39491
rect 81640 -39525 81656 -39509
rect 81590 -39559 81656 -39525
rect 81758 -39525 81774 -39509
rect 81808 -39509 81942 -39491
rect 81808 -39525 81824 -39509
rect 81590 -39593 81606 -39559
rect 81640 -39593 81656 -39559
rect 81590 -39601 81656 -39593
rect 81690 -39559 81724 -39543
rect 81690 -39635 81724 -39593
rect 81758 -39559 81824 -39525
rect 81926 -39525 81942 -39509
rect 81976 -39509 82110 -39491
rect 81976 -39525 81992 -39509
rect 81758 -39593 81774 -39559
rect 81808 -39593 81824 -39559
rect 81758 -39601 81824 -39593
rect 81858 -39559 81892 -39543
rect 81858 -39635 81892 -39593
rect 81926 -39559 81992 -39525
rect 82094 -39525 82110 -39509
rect 82144 -39509 82278 -39491
rect 82144 -39525 82160 -39509
rect 81926 -39593 81942 -39559
rect 81976 -39593 81992 -39559
rect 81926 -39601 81992 -39593
rect 82026 -39559 82060 -39543
rect 82026 -39635 82060 -39593
rect 82094 -39559 82160 -39525
rect 82262 -39525 82278 -39509
rect 82312 -39509 82446 -39491
rect 82312 -39525 82328 -39509
rect 82094 -39593 82110 -39559
rect 82144 -39593 82160 -39559
rect 82094 -39601 82160 -39593
rect 82194 -39559 82228 -39543
rect 82194 -39635 82228 -39593
rect 82262 -39559 82328 -39525
rect 82430 -39525 82446 -39509
rect 82480 -39509 82614 -39491
rect 82480 -39525 82496 -39509
rect 82262 -39593 82278 -39559
rect 82312 -39593 82328 -39559
rect 82262 -39601 82328 -39593
rect 82362 -39559 82396 -39543
rect 82362 -39635 82396 -39593
rect 82430 -39559 82496 -39525
rect 82598 -39525 82614 -39509
rect 82648 -39509 82780 -39491
rect 82648 -39525 82664 -39509
rect 82430 -39593 82446 -39559
rect 82480 -39593 82496 -39559
rect 82430 -39601 82496 -39593
rect 82530 -39559 82564 -39543
rect 82530 -39635 82564 -39593
rect 82598 -39559 82664 -39525
rect 82766 -39530 82780 -39509
rect 82820 -39530 82832 -39490
rect 82598 -39593 82614 -39559
rect 82648 -39593 82664 -39559
rect 82598 -39601 82664 -39593
rect 82698 -39559 82732 -39543
rect 82698 -39635 82732 -39593
rect 82766 -39559 82832 -39530
rect 82766 -39593 82782 -39559
rect 82816 -39593 82832 -39559
rect 82766 -39601 82832 -39593
rect 82866 -39491 82908 -39475
rect 82900 -39525 82908 -39491
rect 82866 -39559 82908 -39525
rect 82900 -39593 82908 -39559
rect 82866 -39635 82908 -39593
rect 82982 -39491 83028 -39475
rect 82982 -39525 82994 -39491
rect 82982 -39559 83028 -39525
rect 82982 -39593 82994 -39559
rect 82982 -39635 83028 -39593
rect 83062 -39491 84250 -39471
rect 83062 -39525 83078 -39491
rect 83112 -39509 83246 -39491
rect 83112 -39525 83128 -39509
rect 83062 -39559 83128 -39525
rect 83230 -39525 83246 -39509
rect 83280 -39509 83414 -39491
rect 83280 -39525 83296 -39509
rect 83062 -39593 83078 -39559
rect 83112 -39593 83128 -39559
rect 83062 -39601 83128 -39593
rect 83162 -39559 83196 -39543
rect 83162 -39635 83196 -39593
rect 83230 -39559 83296 -39525
rect 83398 -39525 83414 -39509
rect 83448 -39509 83582 -39491
rect 83448 -39525 83464 -39509
rect 83230 -39593 83246 -39559
rect 83280 -39593 83296 -39559
rect 83230 -39601 83296 -39593
rect 83330 -39559 83364 -39543
rect 83330 -39635 83364 -39593
rect 83398 -39559 83464 -39525
rect 83566 -39525 83582 -39509
rect 83616 -39509 83750 -39491
rect 83616 -39525 83632 -39509
rect 83398 -39593 83414 -39559
rect 83448 -39593 83464 -39559
rect 83398 -39601 83464 -39593
rect 83498 -39559 83532 -39543
rect 83498 -39635 83532 -39593
rect 83566 -39559 83632 -39525
rect 83734 -39525 83750 -39509
rect 83784 -39509 83918 -39491
rect 83784 -39525 83800 -39509
rect 83566 -39593 83582 -39559
rect 83616 -39593 83632 -39559
rect 83566 -39601 83632 -39593
rect 83666 -39559 83700 -39543
rect 83666 -39635 83700 -39593
rect 83734 -39559 83800 -39525
rect 83902 -39525 83918 -39509
rect 83952 -39509 84086 -39491
rect 83952 -39525 83968 -39509
rect 83734 -39593 83750 -39559
rect 83784 -39593 83800 -39559
rect 83734 -39601 83800 -39593
rect 83834 -39559 83868 -39543
rect 83834 -39635 83868 -39593
rect 83902 -39559 83968 -39525
rect 84070 -39525 84086 -39509
rect 84120 -39509 84250 -39491
rect 84120 -39525 84136 -39509
rect 83902 -39593 83918 -39559
rect 83952 -39593 83968 -39559
rect 83902 -39601 83968 -39593
rect 84002 -39559 84036 -39543
rect 84002 -39635 84036 -39593
rect 84070 -39559 84136 -39525
rect 84238 -39530 84250 -39509
rect 84290 -39530 84304 -39260
rect 84338 -39167 84380 -39125
rect 84372 -39201 84380 -39167
rect 84338 -39235 84380 -39201
rect 84372 -39269 84380 -39235
rect 84338 -39285 84380 -39269
rect 84458 -39167 84500 -39125
rect 84458 -39201 84466 -39167
rect 84458 -39235 84500 -39201
rect 84458 -39269 84466 -39235
rect 84458 -39305 84500 -39269
rect 84458 -39339 84466 -39305
rect 84458 -39355 84500 -39339
rect 84534 -39167 84600 -39159
rect 84534 -39201 84550 -39167
rect 84584 -39201 84600 -39167
rect 84534 -39235 84600 -39201
rect 84534 -39269 84550 -39235
rect 84584 -39269 84600 -39235
rect 84534 -39305 84600 -39269
rect 84634 -39167 84668 -39125
rect 84634 -39235 84668 -39201
rect 84634 -39285 84668 -39269
rect 84702 -39167 84768 -39159
rect 84702 -39201 84718 -39167
rect 84752 -39201 84768 -39167
rect 84702 -39235 84768 -39201
rect 84702 -39269 84718 -39235
rect 84752 -39269 84768 -39235
rect 84534 -39339 84550 -39305
rect 84584 -39319 84600 -39305
rect 84702 -39305 84768 -39269
rect 84802 -39167 84836 -39125
rect 84802 -39235 84836 -39201
rect 84802 -39285 84836 -39269
rect 84870 -39167 84936 -39159
rect 84870 -39201 84886 -39167
rect 84920 -39201 84936 -39167
rect 84870 -39235 84936 -39201
rect 84870 -39269 84886 -39235
rect 84920 -39269 84936 -39235
rect 84702 -39319 84718 -39305
rect 84584 -39339 84718 -39319
rect 84752 -39319 84768 -39305
rect 84870 -39305 84936 -39269
rect 84970 -39167 85004 -39125
rect 84970 -39235 85004 -39201
rect 84970 -39285 85004 -39269
rect 85038 -39167 85104 -39159
rect 85038 -39201 85054 -39167
rect 85088 -39201 85104 -39167
rect 85038 -39235 85104 -39201
rect 85038 -39269 85054 -39235
rect 85088 -39269 85104 -39235
rect 84870 -39319 84886 -39305
rect 84752 -39339 84886 -39319
rect 84920 -39319 84936 -39305
rect 85038 -39305 85104 -39269
rect 85138 -39167 85172 -39125
rect 85138 -39235 85172 -39201
rect 85138 -39285 85172 -39269
rect 85206 -39167 85272 -39159
rect 85206 -39201 85222 -39167
rect 85256 -39201 85272 -39167
rect 85206 -39235 85272 -39201
rect 85206 -39269 85222 -39235
rect 85256 -39269 85272 -39235
rect 85038 -39319 85054 -39305
rect 84920 -39339 85054 -39319
rect 85088 -39319 85104 -39305
rect 85206 -39305 85272 -39269
rect 85306 -39167 85340 -39125
rect 85306 -39235 85340 -39201
rect 85306 -39285 85340 -39269
rect 85374 -39167 85440 -39159
rect 85374 -39201 85390 -39167
rect 85424 -39201 85440 -39167
rect 85374 -39235 85440 -39201
rect 85374 -39269 85390 -39235
rect 85424 -39269 85440 -39235
rect 85206 -39319 85222 -39305
rect 85088 -39339 85222 -39319
rect 85256 -39319 85272 -39305
rect 85374 -39305 85440 -39269
rect 85474 -39167 85508 -39125
rect 85474 -39235 85508 -39201
rect 85474 -39285 85508 -39269
rect 85542 -39167 85608 -39159
rect 85542 -39201 85558 -39167
rect 85592 -39201 85608 -39167
rect 85542 -39235 85608 -39201
rect 85542 -39269 85558 -39235
rect 85592 -39269 85608 -39235
rect 85374 -39319 85390 -39305
rect 85256 -39339 85390 -39319
rect 85424 -39319 85440 -39305
rect 85542 -39305 85608 -39269
rect 85642 -39167 85676 -39125
rect 85642 -39235 85676 -39201
rect 85642 -39285 85676 -39269
rect 85710 -39167 85776 -39159
rect 85710 -39201 85726 -39167
rect 85760 -39201 85776 -39167
rect 85710 -39235 85776 -39201
rect 85710 -39269 85726 -39235
rect 85760 -39269 85776 -39235
rect 85710 -39270 85776 -39269
rect 85542 -39319 85558 -39305
rect 85424 -39339 85558 -39319
rect 85592 -39319 85608 -39305
rect 85710 -39305 85730 -39270
rect 85710 -39319 85726 -39305
rect 85592 -39339 85726 -39319
rect 84534 -39353 85730 -39339
rect 84435 -39397 85523 -39389
rect 84435 -39403 84870 -39397
rect 85240 -39403 85523 -39397
rect 84435 -39437 84460 -39403
rect 84494 -39437 84634 -39403
rect 84668 -39437 84802 -39403
rect 84836 -39437 84870 -39403
rect 85240 -39437 85306 -39403
rect 85340 -39437 85473 -39403
rect 85507 -39437 85523 -39403
rect 85710 -39471 85730 -39353
rect 84070 -39593 84086 -39559
rect 84120 -39593 84136 -39559
rect 84070 -39601 84136 -39593
rect 84170 -39559 84204 -39543
rect 84170 -39635 84204 -39593
rect 84238 -39559 84304 -39530
rect 84238 -39593 84254 -39559
rect 84288 -39593 84304 -39559
rect 84238 -39601 84304 -39593
rect 84338 -39491 84380 -39475
rect 84372 -39525 84380 -39491
rect 84338 -39559 84380 -39525
rect 84372 -39593 84380 -39559
rect 84338 -39635 84380 -39593
rect 84454 -39491 84500 -39475
rect 84454 -39525 84466 -39491
rect 84454 -39559 84500 -39525
rect 84454 -39593 84466 -39559
rect 84454 -39635 84500 -39593
rect 84534 -39491 85730 -39471
rect 84534 -39525 84550 -39491
rect 84584 -39509 84718 -39491
rect 84584 -39525 84600 -39509
rect 84534 -39559 84600 -39525
rect 84702 -39525 84718 -39509
rect 84752 -39509 84886 -39491
rect 84752 -39525 84768 -39509
rect 84534 -39593 84550 -39559
rect 84584 -39593 84600 -39559
rect 84534 -39601 84600 -39593
rect 84634 -39559 84668 -39543
rect 84634 -39635 84668 -39593
rect 84702 -39559 84768 -39525
rect 84870 -39525 84886 -39509
rect 84920 -39509 85054 -39491
rect 84920 -39525 84936 -39509
rect 84702 -39593 84718 -39559
rect 84752 -39593 84768 -39559
rect 84702 -39601 84768 -39593
rect 84802 -39559 84836 -39543
rect 84802 -39635 84836 -39593
rect 84870 -39559 84936 -39525
rect 85038 -39525 85054 -39509
rect 85088 -39509 85222 -39491
rect 85088 -39525 85104 -39509
rect 84870 -39593 84886 -39559
rect 84920 -39593 84936 -39559
rect 84870 -39601 84936 -39593
rect 84970 -39559 85004 -39543
rect 84970 -39635 85004 -39593
rect 85038 -39559 85104 -39525
rect 85206 -39525 85222 -39509
rect 85256 -39509 85390 -39491
rect 85256 -39525 85272 -39509
rect 85038 -39593 85054 -39559
rect 85088 -39593 85104 -39559
rect 85038 -39601 85104 -39593
rect 85138 -39559 85172 -39543
rect 85138 -39635 85172 -39593
rect 85206 -39559 85272 -39525
rect 85374 -39525 85390 -39509
rect 85424 -39509 85558 -39491
rect 85424 -39525 85440 -39509
rect 85206 -39593 85222 -39559
rect 85256 -39593 85272 -39559
rect 85206 -39601 85272 -39593
rect 85306 -39559 85340 -39543
rect 85306 -39635 85340 -39593
rect 85374 -39559 85440 -39525
rect 85542 -39525 85558 -39509
rect 85592 -39509 85726 -39491
rect 85592 -39525 85608 -39509
rect 85374 -39593 85390 -39559
rect 85424 -39593 85440 -39559
rect 85374 -39601 85440 -39593
rect 85474 -39559 85508 -39543
rect 85474 -39635 85508 -39593
rect 85542 -39559 85608 -39525
rect 85710 -39525 85726 -39509
rect 85710 -39540 85730 -39525
rect 85770 -39540 85776 -39270
rect 85810 -39167 85852 -39125
rect 85844 -39201 85852 -39167
rect 85810 -39235 85852 -39201
rect 85844 -39269 85852 -39235
rect 85810 -39285 85852 -39269
rect 85930 -39167 85972 -39125
rect 85930 -39201 85938 -39167
rect 85930 -39235 85972 -39201
rect 85930 -39269 85938 -39235
rect 85930 -39305 85972 -39269
rect 85930 -39339 85938 -39305
rect 85930 -39355 85972 -39339
rect 86006 -39167 86072 -39159
rect 86006 -39201 86022 -39167
rect 86056 -39201 86072 -39167
rect 86006 -39235 86072 -39201
rect 86006 -39269 86022 -39235
rect 86056 -39269 86072 -39235
rect 86006 -39305 86072 -39269
rect 86106 -39167 86140 -39125
rect 86106 -39235 86140 -39201
rect 86106 -39285 86140 -39269
rect 86174 -39167 86240 -39159
rect 86174 -39201 86190 -39167
rect 86224 -39201 86240 -39167
rect 86174 -39235 86240 -39201
rect 86174 -39269 86190 -39235
rect 86224 -39269 86240 -39235
rect 86006 -39339 86022 -39305
rect 86056 -39319 86072 -39305
rect 86174 -39305 86240 -39269
rect 86274 -39167 86308 -39125
rect 86274 -39235 86308 -39201
rect 86274 -39285 86308 -39269
rect 86342 -39167 86408 -39159
rect 86342 -39201 86358 -39167
rect 86392 -39201 86408 -39167
rect 86342 -39235 86408 -39201
rect 86342 -39269 86358 -39235
rect 86392 -39269 86408 -39235
rect 86174 -39319 86190 -39305
rect 86056 -39339 86190 -39319
rect 86224 -39319 86240 -39305
rect 86342 -39305 86408 -39269
rect 86442 -39167 86476 -39125
rect 86442 -39235 86476 -39201
rect 86442 -39285 86476 -39269
rect 86510 -39167 86576 -39159
rect 86510 -39201 86526 -39167
rect 86560 -39201 86576 -39167
rect 86510 -39235 86576 -39201
rect 86510 -39269 86526 -39235
rect 86560 -39269 86576 -39235
rect 86342 -39319 86358 -39305
rect 86224 -39339 86358 -39319
rect 86392 -39319 86408 -39305
rect 86510 -39305 86576 -39269
rect 86610 -39167 86644 -39125
rect 86610 -39235 86644 -39201
rect 86610 -39285 86644 -39269
rect 86678 -39167 86744 -39159
rect 86678 -39201 86694 -39167
rect 86728 -39201 86744 -39167
rect 86678 -39235 86744 -39201
rect 86678 -39269 86694 -39235
rect 86728 -39269 86744 -39235
rect 86510 -39319 86526 -39305
rect 86392 -39339 86526 -39319
rect 86560 -39319 86576 -39305
rect 86678 -39305 86744 -39269
rect 86778 -39167 86812 -39125
rect 86778 -39235 86812 -39201
rect 86778 -39285 86812 -39269
rect 86846 -39167 86912 -39159
rect 86846 -39201 86862 -39167
rect 86896 -39201 86912 -39167
rect 86846 -39235 86912 -39201
rect 86846 -39269 86862 -39235
rect 86896 -39269 86912 -39235
rect 86678 -39319 86694 -39305
rect 86560 -39339 86694 -39319
rect 86728 -39319 86744 -39305
rect 86846 -39305 86912 -39269
rect 86946 -39167 86980 -39125
rect 86946 -39235 86980 -39201
rect 86946 -39285 86980 -39269
rect 87014 -39167 87080 -39159
rect 87014 -39201 87030 -39167
rect 87064 -39201 87080 -39167
rect 87014 -39235 87080 -39201
rect 87014 -39269 87030 -39235
rect 87064 -39269 87080 -39235
rect 86846 -39319 86862 -39305
rect 86728 -39339 86862 -39319
rect 86896 -39319 86912 -39305
rect 87014 -39305 87080 -39269
rect 87114 -39167 87148 -39125
rect 87114 -39235 87148 -39201
rect 87114 -39285 87148 -39269
rect 87182 -39167 87248 -39159
rect 87182 -39201 87198 -39167
rect 87232 -39201 87248 -39167
rect 87182 -39235 87248 -39201
rect 87182 -39269 87198 -39235
rect 87232 -39240 87248 -39235
rect 87014 -39319 87030 -39305
rect 86896 -39339 87030 -39319
rect 87064 -39319 87080 -39305
rect 87182 -39305 87200 -39269
rect 87182 -39319 87198 -39305
rect 87064 -39339 87198 -39319
rect 86006 -39353 87200 -39339
rect 85907 -39394 86995 -39389
rect 85907 -39403 86329 -39394
rect 86699 -39403 86995 -39394
rect 85907 -39437 85932 -39403
rect 85966 -39437 86106 -39403
rect 86140 -39437 86274 -39403
rect 86308 -39434 86329 -39403
rect 86699 -39434 86778 -39403
rect 86308 -39437 86443 -39434
rect 86477 -39437 86610 -39434
rect 86644 -39437 86778 -39434
rect 86812 -39437 86945 -39403
rect 86979 -39437 86995 -39403
rect 87182 -39471 87200 -39353
rect 85542 -39593 85558 -39559
rect 85592 -39593 85608 -39559
rect 85542 -39601 85608 -39593
rect 85642 -39559 85676 -39543
rect 85642 -39635 85676 -39593
rect 85710 -39559 85776 -39540
rect 85710 -39593 85726 -39559
rect 85760 -39593 85776 -39559
rect 85710 -39601 85776 -39593
rect 85810 -39491 85852 -39475
rect 85844 -39525 85852 -39491
rect 85810 -39559 85852 -39525
rect 85844 -39593 85852 -39559
rect 85810 -39635 85852 -39593
rect 85926 -39491 85972 -39475
rect 85926 -39525 85938 -39491
rect 85926 -39559 85972 -39525
rect 85926 -39593 85938 -39559
rect 85926 -39635 85972 -39593
rect 86006 -39491 87200 -39471
rect 86006 -39525 86022 -39491
rect 86056 -39509 86190 -39491
rect 86056 -39525 86072 -39509
rect 86006 -39559 86072 -39525
rect 86174 -39525 86190 -39509
rect 86224 -39509 86358 -39491
rect 86224 -39525 86240 -39509
rect 86006 -39593 86022 -39559
rect 86056 -39593 86072 -39559
rect 86006 -39601 86072 -39593
rect 86106 -39559 86140 -39543
rect 86106 -39635 86140 -39593
rect 86174 -39559 86240 -39525
rect 86342 -39525 86358 -39509
rect 86392 -39509 86526 -39491
rect 86392 -39525 86408 -39509
rect 86174 -39593 86190 -39559
rect 86224 -39593 86240 -39559
rect 86174 -39601 86240 -39593
rect 86274 -39559 86308 -39543
rect 86274 -39635 86308 -39593
rect 86342 -39559 86408 -39525
rect 86510 -39525 86526 -39509
rect 86560 -39509 86694 -39491
rect 86560 -39525 86576 -39509
rect 86342 -39593 86358 -39559
rect 86392 -39593 86408 -39559
rect 86342 -39601 86408 -39593
rect 86442 -39559 86476 -39543
rect 86442 -39635 86476 -39593
rect 86510 -39559 86576 -39525
rect 86678 -39525 86694 -39509
rect 86728 -39509 86862 -39491
rect 86728 -39525 86744 -39509
rect 86510 -39593 86526 -39559
rect 86560 -39593 86576 -39559
rect 86510 -39601 86576 -39593
rect 86610 -39559 86644 -39543
rect 86610 -39635 86644 -39593
rect 86678 -39559 86744 -39525
rect 86846 -39525 86862 -39509
rect 86896 -39509 87030 -39491
rect 86896 -39525 86912 -39509
rect 86678 -39593 86694 -39559
rect 86728 -39593 86744 -39559
rect 86678 -39601 86744 -39593
rect 86778 -39559 86812 -39543
rect 86778 -39635 86812 -39593
rect 86846 -39559 86912 -39525
rect 87014 -39525 87030 -39509
rect 87064 -39509 87198 -39491
rect 87064 -39525 87080 -39509
rect 86846 -39593 86862 -39559
rect 86896 -39593 86912 -39559
rect 86846 -39601 86912 -39593
rect 86946 -39559 86980 -39543
rect 86946 -39635 86980 -39593
rect 87014 -39559 87080 -39525
rect 87182 -39525 87198 -39509
rect 87240 -39510 87248 -39240
rect 87282 -39167 87324 -39125
rect 87316 -39201 87324 -39167
rect 87282 -39235 87324 -39201
rect 87316 -39269 87324 -39235
rect 87282 -39285 87324 -39269
rect 87402 -39167 87444 -39125
rect 87402 -39201 87410 -39167
rect 87402 -39235 87444 -39201
rect 87402 -39269 87410 -39235
rect 87402 -39305 87444 -39269
rect 87402 -39339 87410 -39305
rect 87402 -39355 87444 -39339
rect 87478 -39167 87544 -39159
rect 87478 -39201 87494 -39167
rect 87528 -39201 87544 -39167
rect 87478 -39235 87544 -39201
rect 87478 -39269 87494 -39235
rect 87528 -39269 87544 -39235
rect 87478 -39305 87544 -39269
rect 87578 -39167 87612 -39125
rect 87578 -39235 87612 -39201
rect 87578 -39285 87612 -39269
rect 87646 -39167 87712 -39159
rect 87646 -39201 87662 -39167
rect 87696 -39201 87712 -39167
rect 87646 -39235 87712 -39201
rect 87646 -39269 87662 -39235
rect 87696 -39269 87712 -39235
rect 87478 -39339 87494 -39305
rect 87528 -39319 87544 -39305
rect 87646 -39305 87712 -39269
rect 87746 -39167 87780 -39125
rect 87746 -39235 87780 -39201
rect 87746 -39285 87780 -39269
rect 87814 -39167 87880 -39159
rect 87814 -39201 87830 -39167
rect 87864 -39201 87880 -39167
rect 87814 -39235 87880 -39201
rect 87814 -39269 87830 -39235
rect 87864 -39269 87880 -39235
rect 87646 -39319 87662 -39305
rect 87528 -39339 87662 -39319
rect 87696 -39319 87712 -39305
rect 87814 -39305 87880 -39269
rect 87914 -39167 87948 -39125
rect 87914 -39235 87948 -39201
rect 87914 -39285 87948 -39269
rect 87982 -39167 88048 -39159
rect 87982 -39201 87998 -39167
rect 88032 -39201 88048 -39167
rect 87982 -39235 88048 -39201
rect 87982 -39269 87998 -39235
rect 88032 -39269 88048 -39235
rect 87814 -39319 87830 -39305
rect 87696 -39339 87830 -39319
rect 87864 -39319 87880 -39305
rect 87982 -39305 88048 -39269
rect 88082 -39167 88116 -39125
rect 88082 -39235 88116 -39201
rect 88082 -39285 88116 -39269
rect 88150 -39167 88216 -39159
rect 88150 -39201 88166 -39167
rect 88200 -39201 88216 -39167
rect 88150 -39235 88216 -39201
rect 88150 -39269 88166 -39235
rect 88200 -39269 88216 -39235
rect 87982 -39319 87998 -39305
rect 87864 -39339 87998 -39319
rect 88032 -39319 88048 -39305
rect 88150 -39305 88216 -39269
rect 88250 -39167 88284 -39125
rect 88250 -39235 88284 -39201
rect 88250 -39285 88284 -39269
rect 88318 -39167 88384 -39159
rect 88318 -39201 88334 -39167
rect 88368 -39201 88384 -39167
rect 88318 -39235 88384 -39201
rect 88318 -39269 88334 -39235
rect 88368 -39269 88384 -39235
rect 88150 -39319 88166 -39305
rect 88032 -39339 88166 -39319
rect 88200 -39319 88216 -39305
rect 88318 -39305 88384 -39269
rect 88418 -39167 88452 -39125
rect 88418 -39235 88452 -39201
rect 88418 -39285 88452 -39269
rect 88486 -39167 88552 -39159
rect 88486 -39201 88502 -39167
rect 88536 -39201 88552 -39167
rect 88486 -39235 88552 -39201
rect 88486 -39269 88502 -39235
rect 88536 -39269 88552 -39235
rect 88318 -39319 88334 -39305
rect 88200 -39339 88334 -39319
rect 88368 -39319 88384 -39305
rect 88486 -39305 88552 -39269
rect 88586 -39167 88620 -39125
rect 88586 -39235 88620 -39201
rect 88586 -39285 88620 -39269
rect 88654 -39167 88720 -39159
rect 88654 -39201 88670 -39167
rect 88704 -39201 88720 -39167
rect 88654 -39235 88720 -39201
rect 88486 -39319 88502 -39305
rect 88368 -39339 88502 -39319
rect 88536 -39319 88552 -39305
rect 88654 -39319 88670 -39235
rect 88704 -39260 88720 -39235
rect 88536 -39339 88670 -39319
rect 87478 -39353 88670 -39339
rect 87379 -39395 88467 -39389
rect 87379 -39403 87469 -39395
rect 87749 -39403 88467 -39395
rect 87379 -39437 87404 -39403
rect 87438 -39435 87469 -39403
rect 87438 -39437 87578 -39435
rect 87612 -39437 87746 -39435
rect 87780 -39437 87915 -39403
rect 87949 -39437 88082 -39403
rect 88116 -39437 88250 -39403
rect 88284 -39437 88417 -39403
rect 88451 -39437 88467 -39403
rect 88654 -39471 88670 -39353
rect 87232 -39525 87248 -39510
rect 87014 -39593 87030 -39559
rect 87064 -39593 87080 -39559
rect 87014 -39601 87080 -39593
rect 87114 -39559 87148 -39543
rect 87114 -39635 87148 -39593
rect 87182 -39559 87248 -39525
rect 87182 -39593 87198 -39559
rect 87232 -39593 87248 -39559
rect 87182 -39601 87248 -39593
rect 87282 -39491 87324 -39475
rect 87316 -39525 87324 -39491
rect 87282 -39559 87324 -39525
rect 87316 -39593 87324 -39559
rect 87282 -39635 87324 -39593
rect 87398 -39491 87444 -39475
rect 87398 -39525 87410 -39491
rect 87398 -39559 87444 -39525
rect 87398 -39593 87410 -39559
rect 87398 -39635 87444 -39593
rect 87478 -39491 88670 -39471
rect 87478 -39525 87494 -39491
rect 87528 -39509 87662 -39491
rect 87528 -39525 87544 -39509
rect 87478 -39559 87544 -39525
rect 87646 -39525 87662 -39509
rect 87696 -39509 87830 -39491
rect 87696 -39525 87712 -39509
rect 87478 -39593 87494 -39559
rect 87528 -39593 87544 -39559
rect 87478 -39601 87544 -39593
rect 87578 -39559 87612 -39543
rect 87578 -39635 87612 -39593
rect 87646 -39559 87712 -39525
rect 87814 -39525 87830 -39509
rect 87864 -39509 87998 -39491
rect 87864 -39525 87880 -39509
rect 87646 -39593 87662 -39559
rect 87696 -39593 87712 -39559
rect 87646 -39601 87712 -39593
rect 87746 -39559 87780 -39543
rect 87746 -39635 87780 -39593
rect 87814 -39559 87880 -39525
rect 87982 -39525 87998 -39509
rect 88032 -39509 88166 -39491
rect 88032 -39525 88048 -39509
rect 87814 -39593 87830 -39559
rect 87864 -39593 87880 -39559
rect 87814 -39601 87880 -39593
rect 87914 -39559 87948 -39543
rect 87914 -39635 87948 -39593
rect 87982 -39559 88048 -39525
rect 88150 -39525 88166 -39509
rect 88200 -39509 88334 -39491
rect 88200 -39525 88216 -39509
rect 87982 -39593 87998 -39559
rect 88032 -39593 88048 -39559
rect 87982 -39601 88048 -39593
rect 88082 -39559 88116 -39543
rect 88082 -39635 88116 -39593
rect 88150 -39559 88216 -39525
rect 88318 -39525 88334 -39509
rect 88368 -39509 88502 -39491
rect 88368 -39525 88384 -39509
rect 88150 -39593 88166 -39559
rect 88200 -39593 88216 -39559
rect 88150 -39601 88216 -39593
rect 88250 -39559 88284 -39543
rect 88250 -39635 88284 -39593
rect 88318 -39559 88384 -39525
rect 88486 -39525 88502 -39509
rect 88536 -39509 88670 -39491
rect 88536 -39525 88552 -39509
rect 88318 -39593 88334 -39559
rect 88368 -39593 88384 -39559
rect 88318 -39601 88384 -39593
rect 88418 -39559 88452 -39543
rect 88418 -39635 88452 -39593
rect 88486 -39559 88552 -39525
rect 88654 -39530 88670 -39509
rect 88710 -39530 88720 -39260
rect 88754 -39167 88796 -39125
rect 88788 -39201 88796 -39167
rect 88754 -39235 88796 -39201
rect 88788 -39269 88796 -39235
rect 88754 -39285 88796 -39269
rect 88486 -39593 88502 -39559
rect 88536 -39593 88552 -39559
rect 88486 -39601 88552 -39593
rect 88586 -39559 88620 -39543
rect 88586 -39635 88620 -39593
rect 88654 -39559 88720 -39530
rect 88654 -39593 88670 -39559
rect 88704 -39593 88720 -39559
rect 88654 -39601 88720 -39593
rect 88754 -39491 88796 -39475
rect 88788 -39525 88796 -39491
rect 88754 -39559 88796 -39525
rect 88788 -39593 88796 -39559
rect 88754 -39635 88796 -39593
rect 55960 -39708 56040 -39698
rect 53896 -39748 53992 -39714
rect 54966 -39748 55062 -39714
rect 53350 -39838 53790 -39804
rect 53350 -39900 53384 -39838
rect 53510 -39940 53526 -39906
rect 53614 -39940 53630 -39906
rect 35804 -40592 35838 -40530
rect 25780 -40626 35838 -40592
rect 25780 -40630 35836 -40626
rect 35802 -40692 35836 -40630
rect 53464 -39990 53498 -39974
rect 53464 -40782 53498 -40766
rect 53642 -39990 53676 -39974
rect 53642 -40782 53676 -40766
rect 53756 -40464 53790 -39838
rect 53896 -39810 53930 -39748
rect 55028 -39810 55062 -39748
rect 55710 -39754 56040 -39708
rect 54075 -39862 54091 -39828
rect 54867 -39862 54883 -39828
rect 53998 -39890 54032 -39874
rect 53998 -39944 54032 -39928
rect 54926 -39890 54960 -39874
rect 54926 -39944 54960 -39928
rect 54075 -39990 54091 -39956
rect 54867 -39990 54883 -39956
rect 53896 -40070 53930 -40008
rect 55706 -39788 55802 -39754
rect 56050 -39788 56146 -39754
rect 55706 -39850 55740 -39788
rect 55028 -40070 55062 -40008
rect 53896 -40104 53992 -40070
rect 54966 -40104 55062 -40070
rect 55176 -39900 55272 -39866
rect 55430 -39900 55526 -39866
rect 55176 -39962 55210 -39900
rect 55492 -39962 55526 -39900
rect 55318 -40002 55334 -39968
rect 55368 -40002 55384 -39968
rect 55290 -40052 55324 -40036
rect 55290 -40244 55324 -40228
rect 55378 -40052 55412 -40036
rect 55378 -40244 55412 -40228
rect 55176 -40318 55210 -40256
rect 55492 -40318 55526 -40256
rect 54870 -40352 55272 -40318
rect 55430 -40352 55706 -40318
rect 54870 -40358 55706 -40352
rect 54870 -40464 54904 -40358
rect 53756 -40498 53852 -40464
rect 54808 -40498 54904 -40464
rect 53756 -40560 53790 -40498
rect 54870 -40560 54904 -40498
rect 55126 -40508 55142 -40474
rect 55494 -40508 55510 -40474
rect 53926 -40612 53942 -40578
rect 54718 -40612 54734 -40578
rect 53858 -40640 53892 -40624
rect 53858 -40744 53892 -40728
rect 54768 -40640 54802 -40624
rect 54768 -40744 54802 -40728
rect 53926 -40790 53942 -40756
rect 54718 -40790 54734 -40756
rect 53510 -40850 53526 -40816
rect 53614 -40850 53630 -40816
rect 53756 -40870 53790 -40808
rect 55046 -40560 55080 -40544
rect 55046 -40610 55080 -40594
rect 55556 -40560 55590 -40544
rect 55556 -40610 55590 -40594
rect 55126 -40680 55142 -40646
rect 55494 -40680 55510 -40646
rect 54870 -40838 54904 -40808
rect 55700 -40806 55706 -40358
rect 56112 -39850 56146 -39788
rect 80738 -39669 80767 -39635
rect 80801 -39669 80859 -39635
rect 80893 -39669 80951 -39635
rect 80985 -39669 81043 -39635
rect 81077 -39669 81135 -39635
rect 81169 -39669 81227 -39635
rect 81261 -39669 81319 -39635
rect 81353 -39669 81411 -39635
rect 81445 -39669 81503 -39635
rect 81537 -39669 81595 -39635
rect 81629 -39669 81687 -39635
rect 81721 -39669 81779 -39635
rect 81813 -39669 81871 -39635
rect 81905 -39669 81963 -39635
rect 81997 -39669 82055 -39635
rect 82089 -39669 82147 -39635
rect 82181 -39669 82239 -39635
rect 82273 -39669 82331 -39635
rect 82365 -39669 82423 -39635
rect 82457 -39669 82515 -39635
rect 82549 -39669 82607 -39635
rect 82641 -39669 82699 -39635
rect 82733 -39669 82791 -39635
rect 82825 -39669 82883 -39635
rect 82917 -39669 82975 -39635
rect 83009 -39669 83067 -39635
rect 83101 -39669 83159 -39635
rect 83193 -39669 83251 -39635
rect 83285 -39669 83343 -39635
rect 83377 -39669 83435 -39635
rect 83469 -39669 83527 -39635
rect 83561 -39669 83619 -39635
rect 83653 -39669 83711 -39635
rect 83745 -39669 83803 -39635
rect 83837 -39669 83895 -39635
rect 83929 -39669 83987 -39635
rect 84021 -39669 84079 -39635
rect 84113 -39669 84171 -39635
rect 84205 -39669 84263 -39635
rect 84297 -39669 84355 -39635
rect 84389 -39669 84447 -39635
rect 84481 -39669 84539 -39635
rect 84573 -39669 84631 -39635
rect 84665 -39669 84723 -39635
rect 84757 -39669 84815 -39635
rect 84849 -39669 84907 -39635
rect 84941 -39669 84999 -39635
rect 85033 -39669 85091 -39635
rect 85125 -39669 85183 -39635
rect 85217 -39669 85275 -39635
rect 85309 -39669 85367 -39635
rect 85401 -39669 85459 -39635
rect 85493 -39669 85551 -39635
rect 85585 -39669 85643 -39635
rect 85677 -39669 85735 -39635
rect 85769 -39669 85827 -39635
rect 85861 -39669 85919 -39635
rect 85953 -39669 86011 -39635
rect 86045 -39669 86103 -39635
rect 86137 -39669 86195 -39635
rect 86229 -39669 86287 -39635
rect 86321 -39669 86379 -39635
rect 86413 -39669 86471 -39635
rect 86505 -39669 86563 -39635
rect 86597 -39669 86655 -39635
rect 86689 -39669 86747 -39635
rect 86781 -39669 86839 -39635
rect 86873 -39669 86931 -39635
rect 86965 -39669 87023 -39635
rect 87057 -39669 87115 -39635
rect 87149 -39669 87207 -39635
rect 87241 -39669 87299 -39635
rect 87333 -39669 87391 -39635
rect 87425 -39669 87483 -39635
rect 87517 -39669 87575 -39635
rect 87609 -39669 87667 -39635
rect 87701 -39669 87759 -39635
rect 87793 -39669 87851 -39635
rect 87885 -39669 87943 -39635
rect 87977 -39669 88035 -39635
rect 88069 -39669 88127 -39635
rect 88161 -39669 88219 -39635
rect 88253 -39669 88311 -39635
rect 88345 -39669 88403 -39635
rect 88437 -39669 88495 -39635
rect 88529 -39669 88587 -39635
rect 88621 -39669 88679 -39635
rect 88713 -39669 88771 -39635
rect 88805 -39669 88834 -39635
rect 58930 -39767 59026 -39733
rect 59600 -39767 59696 -39733
rect 77578 -39705 77607 -39671
rect 77641 -39705 77699 -39671
rect 77733 -39705 77791 -39671
rect 77825 -39705 77883 -39671
rect 77917 -39705 77975 -39671
rect 78009 -39705 78067 -39671
rect 78101 -39705 78130 -39671
rect 58930 -39810 58964 -39767
rect 58926 -39820 58966 -39810
rect 55866 -39890 55882 -39856
rect 55970 -39890 55986 -39856
rect 55820 -39940 55854 -39924
rect 55820 -40732 55854 -40716
rect 55998 -39940 56032 -39924
rect 55998 -40732 56032 -40716
rect 55866 -40800 55882 -40766
rect 55970 -40800 55986 -40766
rect 55700 -40838 55740 -40806
rect 57096 -39879 57125 -39845
rect 57159 -39879 57217 -39845
rect 57251 -39879 57309 -39845
rect 57343 -39879 57372 -39845
rect 57129 -39929 57165 -39913
rect 57129 -39963 57131 -39929
rect 57129 -39997 57165 -39963
rect 57129 -40031 57131 -39997
rect 57201 -39929 57267 -39879
rect 57201 -39963 57217 -39929
rect 57251 -39963 57267 -39929
rect 57201 -39997 57267 -39963
rect 57201 -40031 57217 -39997
rect 57251 -40031 57267 -39997
rect 57301 -39929 57355 -39913
rect 57301 -39963 57303 -39929
rect 57337 -39963 57355 -39929
rect 57301 -40010 57355 -39963
rect 57129 -40065 57165 -40031
rect 57301 -40044 57303 -40010
rect 57337 -40044 57355 -40010
rect 57129 -40099 57264 -40065
rect 57301 -40094 57355 -40044
rect 57230 -40128 57264 -40099
rect 57117 -40144 57185 -40135
rect 57117 -40194 57118 -40144
rect 57178 -40194 57185 -40144
rect 57117 -40209 57185 -40194
rect 57230 -40144 57285 -40128
rect 57230 -40178 57251 -40144
rect 57230 -40194 57285 -40178
rect 57319 -40140 57355 -40094
rect 59662 -39829 59696 -39767
rect 59109 -39881 59125 -39847
rect 59501 -39881 59517 -39847
rect 59560 -39901 59594 -39885
rect 59560 -39951 59594 -39935
rect 59109 -39989 59125 -39955
rect 59501 -39989 59517 -39955
rect 59032 -40009 59066 -39993
rect 59032 -40059 59066 -40043
rect 59109 -40097 59125 -40063
rect 59501 -40097 59517 -40063
rect 77150 -39790 77280 -39760
rect 77597 -39771 77663 -39705
rect 77150 -39840 77170 -39790
rect 77260 -39840 77280 -39790
rect 77597 -39805 77613 -39771
rect 77647 -39805 77663 -39771
rect 77703 -39765 77737 -39749
rect 77777 -39751 77843 -39705
rect 77777 -39785 77793 -39751
rect 77827 -39785 77843 -39751
rect 77877 -39765 77911 -39749
rect 77703 -39819 77737 -39799
rect 77945 -39751 78021 -39705
rect 80788 -39745 80817 -39711
rect 80851 -39745 80909 -39711
rect 80943 -39745 81001 -39711
rect 81035 -39745 81064 -39711
rect 77945 -39785 77971 -39751
rect 78005 -39785 78021 -39751
rect 78080 -39771 78220 -39770
rect 77877 -39819 77911 -39799
rect 78059 -39789 78220 -39771
rect 77596 -39840 77666 -39839
rect 77150 -39903 77666 -39840
rect 77703 -39853 78025 -39819
rect 78093 -39790 78220 -39789
rect 78093 -39823 78160 -39790
rect 78059 -39830 78160 -39823
rect 78200 -39830 78220 -39790
rect 78059 -39840 78220 -39830
rect 77991 -39887 78025 -39853
rect 77150 -39937 77613 -39903
rect 77647 -39937 77666 -39903
rect 77150 -39950 77666 -39937
rect 77596 -39953 77666 -39950
rect 77700 -39903 77842 -39887
rect 77700 -39937 77739 -39903
rect 77773 -39937 77842 -39903
rect 77700 -39960 77842 -39937
rect 77876 -39900 77957 -39887
rect 77876 -39940 77900 -39900
rect 77940 -39903 77957 -39900
rect 77949 -39937 77957 -39903
rect 77940 -39940 77957 -39937
rect 77876 -39953 77957 -39940
rect 77991 -39903 78045 -39887
rect 77991 -39937 78011 -39903
rect 77991 -39953 78045 -39937
rect 78079 -39900 78220 -39840
rect 78079 -39940 78160 -39900
rect 78200 -39940 78220 -39900
rect 77596 -40008 77660 -39987
rect 77596 -40042 77613 -40008
rect 77647 -40042 77660 -40008
rect 77700 -40000 77770 -39960
rect 77810 -40000 77842 -39960
rect 77991 -39987 78025 -39953
rect 78079 -39987 78220 -39940
rect 77700 -40011 77842 -40000
rect 77596 -40045 77660 -40042
rect 77880 -40021 78025 -39987
rect 78059 -40020 78220 -39987
rect 80460 -39800 80730 -39780
rect 80460 -39960 80480 -39800
rect 80640 -39950 80730 -39800
rect 80852 -39791 80898 -39745
rect 80852 -39825 80864 -39791
rect 80852 -39859 80898 -39825
rect 80852 -39893 80864 -39859
rect 80852 -39909 80898 -39893
rect 80932 -39791 80998 -39779
rect 80932 -39825 80948 -39791
rect 80982 -39825 80998 -39791
rect 80932 -39859 80998 -39825
rect 80932 -39893 80948 -39859
rect 80982 -39893 80998 -39859
rect 80932 -39905 80998 -39893
rect 80852 -39950 80868 -39943
rect 80640 -39960 80868 -39950
rect 80460 -39977 80868 -39960
rect 80902 -39977 80918 -39943
rect 80460 -39990 80918 -39977
rect 80852 -39991 80918 -39990
rect 77880 -40045 77914 -40021
rect 58926 -40140 58966 -40120
rect 57319 -40180 57326 -40140
rect 58930 -40176 58964 -40140
rect 57230 -40245 57264 -40194
rect 57131 -40279 57264 -40245
rect 57319 -40254 57355 -40180
rect 57131 -40300 57165 -40279
rect 56316 -40318 56412 -40304
rect 54830 -40848 55830 -40838
rect 54830 -40870 55030 -40848
rect 53756 -40904 53852 -40870
rect 54808 -40904 55030 -40870
rect 53510 -40958 53526 -40924
rect 53614 -40958 53630 -40924
rect 53756 -40966 53790 -40904
rect 54830 -40928 55030 -40904
rect 55110 -40868 55740 -40848
rect 55810 -40868 55830 -40848
rect 56112 -40868 56146 -40806
rect 55110 -40908 55160 -40868
rect 55600 -40908 55740 -40868
rect 56050 -40902 56146 -40868
rect 55110 -40928 55740 -40908
rect 55810 -40928 55830 -40902
rect 54830 -40938 55830 -40928
rect 53464 -41008 53498 -40992
rect 53464 -41800 53498 -41784
rect 53642 -41008 53676 -40992
rect 53642 -41800 53676 -41784
rect 54870 -40966 54904 -40938
rect 53926 -41018 53942 -40984
rect 54718 -41018 54734 -40984
rect 53858 -41046 53892 -41030
rect 53858 -41150 53892 -41134
rect 54768 -41046 54802 -41030
rect 54768 -41150 54802 -41134
rect 53926 -41196 53942 -41162
rect 54718 -41196 54734 -41162
rect 53756 -41276 53790 -41214
rect 55700 -40964 55740 -40938
rect 55126 -41130 55142 -41096
rect 55494 -41130 55510 -41096
rect 54870 -41276 54904 -41214
rect 55046 -41182 55080 -41166
rect 55046 -41232 55080 -41216
rect 55556 -41182 55590 -41166
rect 55556 -41232 55590 -41216
rect 53756 -41310 53852 -41276
rect 54808 -41310 54904 -41276
rect 55126 -41302 55142 -41268
rect 55494 -41302 55510 -41268
rect 53510 -41868 53526 -41834
rect 53614 -41868 53630 -41834
rect 53350 -41936 53384 -41874
rect 53756 -41936 53790 -41310
rect 54870 -41418 54904 -41310
rect 55700 -41418 55706 -40964
rect 54870 -41424 55706 -41418
rect 54870 -41458 55262 -41424
rect 55420 -41458 55706 -41424
rect 55166 -41520 55200 -41458
rect 53350 -41970 53446 -41936
rect 53694 -41970 53790 -41936
rect 53886 -41708 53982 -41674
rect 54956 -41708 55052 -41674
rect 53886 -41770 53920 -41708
rect 55018 -41770 55052 -41708
rect 54065 -41822 54081 -41788
rect 54857 -41822 54873 -41788
rect 53988 -41850 54022 -41834
rect 53988 -41904 54022 -41888
rect 54916 -41850 54950 -41834
rect 54916 -41904 54950 -41888
rect 54065 -41950 54081 -41916
rect 54857 -41950 54873 -41916
rect 35802 -42190 35836 -42128
rect 25780 -42228 35836 -42190
rect 35802 -42290 35836 -42228
rect 53886 -42030 53920 -41968
rect 55482 -41520 55516 -41458
rect 55280 -41548 55314 -41532
rect 55280 -41740 55314 -41724
rect 55368 -41548 55402 -41532
rect 55368 -41740 55402 -41724
rect 55308 -41808 55324 -41774
rect 55358 -41808 55374 -41774
rect 55166 -41876 55200 -41814
rect 55482 -41876 55516 -41814
rect 55166 -41910 55262 -41876
rect 55420 -41910 55516 -41876
rect 55018 -42030 55052 -41968
rect 56112 -40964 56146 -40902
rect 56350 -40338 56412 -40318
rect 56610 -40338 56706 -40304
rect 56672 -40400 56706 -40338
rect 57303 -40283 57355 -40254
rect 57131 -40355 57165 -40334
rect 57201 -40347 57217 -40313
rect 57251 -40347 57267 -40313
rect 57201 -40389 57267 -40347
rect 57337 -40317 57355 -40283
rect 57303 -40355 57355 -40317
rect 58930 -40210 59026 -40176
rect 59214 -40177 59310 -40176
rect 59662 -40177 59696 -40120
rect 59772 -40094 59866 -40060
rect 60426 -40094 60520 -40060
rect 77596 -40079 77914 -40045
rect 78059 -40040 78160 -40020
rect 77961 -40071 78017 -40055
rect 59772 -40150 59806 -40094
rect 59214 -40210 59696 -40177
rect 58930 -40211 59696 -40210
rect 58930 -40272 58964 -40211
rect 59276 -40272 59310 -40211
rect 59087 -40312 59103 -40278
rect 59137 -40312 59153 -40278
rect 56476 -40440 56492 -40406
rect 56530 -40440 56546 -40406
rect 55866 -41004 55882 -40970
rect 55970 -41004 55986 -40970
rect 55820 -41054 55854 -41038
rect 55820 -41846 55854 -41830
rect 55998 -41054 56032 -41038
rect 55998 -41846 56032 -41830
rect 55866 -41914 55882 -41880
rect 55970 -41914 55986 -41880
rect 55706 -41982 55740 -41920
rect 56430 -40499 56464 -40483
rect 56430 -41291 56464 -41275
rect 56558 -40499 56592 -40483
rect 56558 -41291 56592 -41275
rect 56476 -41368 56492 -41334
rect 56530 -41368 56546 -41334
rect 56316 -41436 56350 -41374
rect 57096 -40423 57125 -40389
rect 57159 -40423 57217 -40389
rect 57251 -40423 57309 -40389
rect 57343 -40423 57372 -40389
rect 59044 -40371 59078 -40355
rect 59044 -40763 59078 -40747
rect 59162 -40371 59196 -40355
rect 59162 -40763 59196 -40747
rect 59087 -40840 59103 -40806
rect 59137 -40840 59153 -40806
rect 60486 -40156 60520 -40094
rect 59942 -40208 59958 -40174
rect 60334 -40208 60350 -40174
rect 59874 -40228 59908 -40212
rect 59874 -40278 59908 -40262
rect 60384 -40228 60418 -40212
rect 60384 -40278 60418 -40262
rect 59942 -40316 59958 -40282
rect 60334 -40316 60350 -40282
rect 59772 -40396 59806 -40340
rect 77400 -40120 77490 -40100
rect 77961 -40105 77974 -40071
rect 78008 -40105 78017 -40071
rect 77596 -40120 77927 -40113
rect 77400 -40170 77420 -40120
rect 77470 -40127 77927 -40120
rect 77470 -40161 77835 -40127
rect 77869 -40161 77927 -40127
rect 77470 -40170 77927 -40161
rect 77400 -40190 77490 -40170
rect 77596 -40171 77927 -40170
rect 77961 -40139 78017 -40105
rect 77961 -40173 77974 -40139
rect 78008 -40173 78017 -40139
rect 77961 -40215 78017 -40173
rect 78093 -40060 78160 -40040
rect 78200 -40060 78220 -40020
rect 80952 -40025 80998 -39905
rect 78093 -40074 78220 -40060
rect 78059 -40100 78220 -40074
rect 80856 -40043 80898 -40027
rect 80856 -40077 80864 -40043
rect 78059 -40108 78113 -40100
rect 78093 -40142 78113 -40108
rect 78059 -40181 78113 -40142
rect 80856 -40111 80898 -40077
rect 80856 -40145 80864 -40111
rect 80856 -40179 80898 -40145
rect 80856 -40213 80864 -40179
rect 77578 -40249 77607 -40215
rect 77641 -40249 77699 -40215
rect 77733 -40249 77791 -40215
rect 77825 -40249 77883 -40215
rect 77917 -40249 77975 -40215
rect 78009 -40249 78067 -40215
rect 78101 -40249 78130 -40215
rect 77578 -40325 77607 -40291
rect 77641 -40325 77699 -40291
rect 77733 -40325 77791 -40291
rect 77825 -40325 77883 -40291
rect 77917 -40325 77975 -40291
rect 78009 -40325 78038 -40291
rect 60486 -40396 60520 -40334
rect 59388 -40430 59476 -40396
rect 59656 -40430 59800 -40396
rect 59958 -40430 60520 -40396
rect 77635 -40409 77691 -40325
rect 77825 -40367 77891 -40325
rect 80856 -40255 80898 -40213
rect 80932 -40043 80998 -40025
rect 80932 -40050 80948 -40043
rect 80982 -40050 80998 -40043
rect 80932 -40160 80940 -40050
rect 80990 -40160 80998 -40050
rect 80932 -40179 80998 -40160
rect 80932 -40213 80948 -40179
rect 80982 -40213 80998 -40179
rect 80932 -40221 80998 -40213
rect 80788 -40289 80817 -40255
rect 80851 -40289 80909 -40255
rect 80943 -40289 81001 -40255
rect 81035 -40289 81064 -40255
rect 59388 -40490 59422 -40430
rect 59276 -40906 59310 -40846
rect 59530 -40532 59546 -40498
rect 59580 -40532 59596 -40498
rect 59502 -40582 59536 -40566
rect 59502 -40774 59536 -40758
rect 59590 -40582 59624 -40566
rect 59590 -40774 59624 -40758
rect 59530 -40842 59546 -40808
rect 59580 -40842 59596 -40808
rect 58966 -40942 59310 -40906
rect 59388 -40909 59422 -40850
rect 59704 -40909 59738 -40430
rect 60020 -40492 60054 -40430
rect 77635 -40443 77649 -40409
rect 77683 -40443 77691 -40409
rect 77635 -40459 77691 -40443
rect 77725 -40409 77785 -40393
rect 77725 -40443 77733 -40409
rect 77767 -40443 77785 -40409
rect 59846 -40532 59862 -40498
rect 59896 -40532 59912 -40498
rect 59818 -40582 59852 -40566
rect 59818 -40774 59852 -40758
rect 59906 -40582 59940 -40566
rect 59906 -40774 59940 -40758
rect 59846 -40842 59862 -40808
rect 59896 -40842 59912 -40808
rect 77725 -40503 77785 -40443
rect 77825 -40401 77841 -40367
rect 77875 -40401 77891 -40367
rect 77825 -40435 77891 -40401
rect 77825 -40469 77841 -40435
rect 77875 -40469 77891 -40435
rect 77929 -40367 78021 -40359
rect 77929 -40401 77945 -40367
rect 77979 -40370 78021 -40367
rect 77979 -40401 78060 -40370
rect 77929 -40435 78060 -40401
rect 77929 -40469 77945 -40435
rect 77979 -40469 78060 -40435
rect 77598 -40520 77651 -40515
rect 77410 -40550 77651 -40520
rect 77725 -40537 77913 -40503
rect 61186 -40600 61286 -40590
rect 77410 -40600 77460 -40550
rect 77510 -40580 77651 -40550
rect 77510 -40600 77740 -40580
rect 77879 -40587 77913 -40537
rect 77971 -40530 78060 -40469
rect 77971 -40570 78000 -40530
rect 78040 -40570 78060 -40530
rect 61186 -40680 61196 -40600
rect 77410 -40603 77740 -40600
rect 77410 -40630 77652 -40603
rect 77598 -40637 77652 -40630
rect 77686 -40630 77740 -40603
rect 77777 -40590 77845 -40587
rect 77777 -40630 77790 -40590
rect 77830 -40630 77845 -40590
rect 77686 -40637 77733 -40630
rect 77777 -40637 77793 -40630
rect 77827 -40637 77845 -40630
rect 77879 -40603 77937 -40587
rect 77879 -40637 77901 -40603
rect 77935 -40637 77937 -40603
rect 77879 -40653 77937 -40637
rect 77971 -40620 78060 -40570
rect 77879 -40671 77913 -40653
rect 61186 -40690 61286 -40680
rect 60020 -40909 60054 -40848
rect 56672 -41436 56706 -41374
rect 57096 -41399 57125 -41365
rect 57159 -41399 57217 -41365
rect 57251 -41399 57309 -41365
rect 57343 -41399 57372 -41365
rect 56316 -41470 56412 -41436
rect 56610 -41470 56706 -41436
rect 57131 -41454 57165 -41433
rect 57201 -41441 57267 -41399
rect 57201 -41475 57217 -41441
rect 57251 -41475 57267 -41441
rect 57303 -41471 57355 -41433
rect 57131 -41509 57165 -41488
rect 57337 -41505 57355 -41471
rect 59276 -41002 59310 -40942
rect 59387 -40944 60054 -40909
rect 60127 -40754 60161 -40728
rect 60127 -40757 60253 -40754
rect 60161 -40773 60253 -40757
rect 60161 -40791 60203 -40773
rect 60127 -40807 60203 -40791
rect 60237 -40807 60253 -40773
rect 60359 -40760 60409 -40749
rect 60671 -40754 60705 -40728
rect 60359 -40765 60366 -40760
rect 60359 -40800 60366 -40799
rect 60406 -40800 60409 -40760
rect 60127 -40849 60161 -40807
rect 60127 -40941 60161 -40883
rect 60195 -40857 60325 -40841
rect 60195 -40891 60211 -40857
rect 60245 -40891 60325 -40857
rect 60195 -40907 60325 -40891
rect 59387 -41000 59421 -40944
rect 59087 -41042 59103 -41008
rect 59137 -41042 59153 -41008
rect 59044 -41101 59078 -41085
rect 57131 -41543 57264 -41509
rect 57303 -41534 57355 -41505
rect 57117 -41594 57185 -41579
rect 57117 -41644 57118 -41594
rect 57168 -41644 57185 -41594
rect 57117 -41653 57185 -41644
rect 57230 -41594 57264 -41543
rect 57319 -41570 57355 -41534
rect 57230 -41610 57285 -41594
rect 57230 -41644 57251 -41610
rect 57230 -41660 57285 -41644
rect 57319 -41610 57326 -41570
rect 59044 -41493 59078 -41477
rect 59162 -41101 59196 -41085
rect 59162 -41493 59196 -41477
rect 59087 -41570 59103 -41536
rect 59137 -41570 59153 -41536
rect 57230 -41689 57264 -41660
rect 57129 -41723 57264 -41689
rect 57319 -41694 57355 -41610
rect 57129 -41757 57165 -41723
rect 57301 -41744 57355 -41694
rect 58930 -41638 58964 -41576
rect 59529 -41045 59545 -41011
rect 59579 -41045 59595 -41011
rect 59501 -41095 59535 -41079
rect 59501 -41287 59535 -41271
rect 59589 -41095 59623 -41079
rect 59589 -41287 59623 -41271
rect 59529 -41355 59545 -41321
rect 59579 -41355 59595 -41321
rect 59387 -41423 59421 -41370
rect 59703 -41423 59737 -40944
rect 60019 -41005 60053 -40944
rect 59845 -41045 59861 -41011
rect 59895 -41045 59911 -41011
rect 59817 -41095 59851 -41079
rect 59817 -41287 59851 -41271
rect 59905 -41095 59939 -41079
rect 59905 -41287 59939 -41271
rect 59845 -41355 59861 -41321
rect 59895 -41355 59911 -41321
rect 60161 -40975 60203 -40941
rect 60237 -40975 60253 -40941
rect 60127 -41033 60161 -40975
rect 60289 -41009 60325 -40907
rect 60127 -41109 60161 -41067
rect 60195 -41025 60325 -41009
rect 60195 -41059 60211 -41025
rect 60245 -41059 60325 -41025
rect 60195 -41075 60325 -41059
rect 60359 -40850 60409 -40800
rect 60443 -40757 60705 -40754
rect 60443 -40773 60671 -40757
rect 60443 -40807 60459 -40773
rect 60493 -40807 60527 -40773
rect 60561 -40807 60595 -40773
rect 60629 -40791 60671 -40773
rect 60629 -40807 60705 -40791
rect 60359 -40857 60366 -40850
rect 60406 -40890 60409 -40850
rect 60393 -40891 60409 -40890
rect 60359 -40940 60409 -40891
rect 60359 -40941 60366 -40940
rect 60359 -40980 60366 -40975
rect 60406 -40980 60409 -40940
rect 60359 -41020 60409 -40980
rect 60359 -41025 60366 -41020
rect 60359 -41060 60366 -41059
rect 60406 -41060 60409 -41020
rect 60359 -41075 60409 -41060
rect 60443 -40857 60637 -40841
rect 60443 -40891 60459 -40857
rect 60493 -40891 60527 -40857
rect 60561 -40891 60595 -40857
rect 60629 -40891 60637 -40857
rect 60443 -40907 60637 -40891
rect 60671 -40849 60705 -40807
rect 60443 -41009 60477 -40907
rect 60671 -40941 60705 -40883
rect 60511 -40975 60527 -40941
rect 60561 -40975 60595 -40941
rect 60629 -40975 60671 -40941
rect 60443 -41025 60637 -41009
rect 60443 -41059 60459 -41025
rect 60493 -41059 60527 -41025
rect 60561 -41059 60595 -41025
rect 60629 -41059 60637 -41025
rect 60443 -41075 60637 -41059
rect 60671 -41033 60705 -40975
rect 60289 -41109 60325 -41075
rect 60443 -41109 60481 -41075
rect 60671 -41109 60705 -41067
rect 60127 -41125 60204 -41109
rect 60161 -41143 60204 -41125
rect 60238 -41143 60254 -41109
rect 60161 -41159 60254 -41143
rect 60289 -41125 60481 -41109
rect 60289 -41159 60297 -41125
rect 60331 -41159 60369 -41125
rect 60405 -41159 60449 -41125
rect 60579 -41143 60595 -41109
rect 60629 -41125 60705 -41109
rect 60629 -41143 60671 -41125
rect 60579 -41151 60671 -41143
rect 60127 -41188 60161 -41159
rect 60289 -41162 60481 -41159
rect 60671 -41188 60705 -41159
rect 60747 -40754 60781 -40728
rect 60747 -40757 61009 -40754
rect 60781 -40773 61009 -40757
rect 60781 -40791 60823 -40773
rect 60747 -40807 60823 -40791
rect 60857 -40807 60891 -40773
rect 60925 -40807 60959 -40773
rect 60993 -40807 61009 -40773
rect 61043 -40760 61093 -40749
rect 61291 -40754 61325 -40728
rect 61043 -40800 61046 -40760
rect 61086 -40765 61093 -40760
rect 61086 -40800 61093 -40799
rect 60747 -40849 60781 -40807
rect 60747 -40941 60781 -40883
rect 60815 -40857 61009 -40841
rect 60815 -40891 60823 -40857
rect 60857 -40891 60891 -40857
rect 60925 -40891 60959 -40857
rect 60993 -40891 61009 -40857
rect 60815 -40907 61009 -40891
rect 60781 -40975 60823 -40941
rect 60857 -40975 60891 -40941
rect 60925 -40975 60941 -40941
rect 60747 -41033 60781 -40975
rect 60975 -41009 61009 -40907
rect 60747 -41109 60781 -41067
rect 60815 -41025 61009 -41009
rect 60815 -41059 60823 -41025
rect 60857 -41059 60891 -41025
rect 60925 -41059 60959 -41025
rect 60993 -41059 61009 -41025
rect 60815 -41075 61009 -41059
rect 61043 -40850 61093 -40800
rect 61199 -40757 61325 -40754
rect 61199 -40773 61291 -40757
rect 61199 -40807 61215 -40773
rect 61249 -40791 61291 -40773
rect 61249 -40807 61325 -40791
rect 61043 -40890 61046 -40850
rect 61086 -40857 61093 -40850
rect 61043 -40891 61059 -40890
rect 61043 -40940 61093 -40891
rect 61043 -40980 61046 -40940
rect 61086 -40941 61093 -40940
rect 61086 -40980 61093 -40975
rect 61043 -41020 61093 -40980
rect 61043 -41060 61046 -41020
rect 61086 -41025 61093 -41020
rect 61086 -41060 61093 -41059
rect 61043 -41075 61093 -41060
rect 61127 -40857 61257 -40841
rect 61127 -40891 61207 -40857
rect 61241 -40891 61257 -40857
rect 61127 -40907 61257 -40891
rect 61291 -40849 61325 -40807
rect 77635 -40709 77913 -40671
rect 77971 -40660 78000 -40620
rect 78040 -40660 78060 -40620
rect 77971 -40700 78060 -40660
rect 77635 -40731 77701 -40709
rect 77635 -40765 77649 -40731
rect 77683 -40765 77701 -40731
rect 77971 -40740 78000 -40700
rect 78040 -40740 78060 -40700
rect 77971 -40743 78060 -40740
rect 77635 -40781 77701 -40765
rect 77825 -40759 77875 -40743
rect 77825 -40793 77841 -40759
rect 77825 -40835 77875 -40793
rect 77909 -40759 78060 -40743
rect 77909 -40793 77925 -40759
rect 77959 -40790 78060 -40759
rect 77959 -40793 78021 -40790
rect 77909 -40801 78021 -40793
rect 77578 -40869 77607 -40835
rect 77641 -40869 77699 -40835
rect 77733 -40869 77791 -40835
rect 77825 -40869 77883 -40835
rect 77917 -40869 77975 -40835
rect 78009 -40869 78038 -40835
rect 61127 -41009 61163 -40907
rect 61291 -40941 61325 -40883
rect 61199 -40975 61215 -40941
rect 61249 -40975 61291 -40941
rect 77578 -40945 77607 -40911
rect 77641 -40945 77699 -40911
rect 77733 -40945 77791 -40911
rect 77825 -40945 77883 -40911
rect 77917 -40945 77975 -40911
rect 78009 -40945 78067 -40911
rect 78101 -40945 78159 -40911
rect 78193 -40945 78251 -40911
rect 78285 -40945 78343 -40911
rect 78377 -40945 78435 -40911
rect 78469 -40945 78527 -40911
rect 78561 -40945 78590 -40911
rect 61127 -41025 61257 -41009
rect 61127 -41059 61207 -41025
rect 61241 -41059 61257 -41025
rect 61127 -41075 61257 -41059
rect 61291 -41033 61325 -40975
rect 60971 -41109 61009 -41075
rect 61127 -41109 61163 -41075
rect 61291 -41109 61325 -41067
rect 77825 -40987 77875 -40945
rect 77635 -41015 77701 -40999
rect 77635 -41049 77649 -41015
rect 77683 -41049 77701 -41015
rect 77825 -41021 77841 -40987
rect 77825 -41037 77875 -41021
rect 77909 -40987 78021 -40979
rect 77909 -41021 77925 -40987
rect 77959 -41021 78021 -40987
rect 77909 -41037 78021 -41021
rect 77635 -41071 77701 -41049
rect 77635 -41109 77913 -41071
rect 60747 -41125 60823 -41109
rect 60781 -41143 60823 -41125
rect 60857 -41143 60873 -41109
rect 60781 -41151 60873 -41143
rect 60971 -41124 61163 -41109
rect 60971 -41125 61129 -41124
rect 60747 -41188 60781 -41159
rect 60971 -41159 60980 -41125
rect 61015 -41159 61053 -41125
rect 61088 -41158 61129 -41125
rect 61198 -41143 61214 -41109
rect 61248 -41125 61325 -41109
rect 61248 -41143 61291 -41125
rect 61088 -41159 61163 -41158
rect 61198 -41159 61291 -41143
rect 77879 -41127 77913 -41109
rect 77879 -41143 77937 -41127
rect 77598 -41150 77652 -41143
rect 60971 -41162 61163 -41159
rect 61291 -41188 61325 -41159
rect 77430 -41177 77652 -41150
rect 77686 -41177 77733 -41143
rect 77430 -41180 77733 -41177
rect 77430 -41220 77470 -41180
rect 77510 -41193 77733 -41180
rect 77777 -41150 77793 -41143
rect 77827 -41150 77845 -41143
rect 77777 -41190 77790 -41150
rect 77830 -41190 77845 -41150
rect 77777 -41193 77845 -41190
rect 77879 -41177 77901 -41143
rect 77935 -41177 77937 -41143
rect 77879 -41193 77937 -41177
rect 77510 -41220 77651 -41193
rect 60466 -41260 60546 -41240
rect 60466 -41300 60486 -41260
rect 60526 -41300 60546 -41260
rect 60466 -41320 60546 -41300
rect 60606 -41260 60686 -41240
rect 60606 -41300 60626 -41260
rect 60666 -41300 60686 -41260
rect 60606 -41320 60686 -41300
rect 60746 -41260 60826 -41240
rect 60746 -41300 60766 -41260
rect 60806 -41300 60826 -41260
rect 60746 -41320 60826 -41300
rect 60886 -41260 60966 -41240
rect 77430 -41260 77651 -41220
rect 77879 -41243 77913 -41193
rect 60886 -41300 60906 -41260
rect 60946 -41300 60966 -41260
rect 77598 -41265 77651 -41260
rect 60886 -41320 60966 -41300
rect 77725 -41277 77913 -41243
rect 60019 -41423 60053 -41361
rect 59387 -41457 59476 -41423
rect 59646 -41457 59799 -41423
rect 59957 -41426 60053 -41423
rect 77635 -41337 77691 -41321
rect 77635 -41371 77649 -41337
rect 77683 -41371 77691 -41337
rect 59957 -41457 60520 -41426
rect 77635 -41455 77691 -41371
rect 77725 -41337 77785 -41277
rect 77971 -41311 78021 -41037
rect 78057 -41011 78123 -40945
rect 78057 -41045 78073 -41011
rect 78107 -41045 78123 -41011
rect 78163 -41005 78197 -40989
rect 78237 -40991 78303 -40945
rect 78237 -41025 78253 -40991
rect 78287 -41025 78303 -40991
rect 78337 -41005 78371 -40989
rect 78163 -41059 78197 -41039
rect 78405 -40991 78481 -40945
rect 78405 -41025 78431 -40991
rect 78465 -41025 78481 -40991
rect 78540 -41011 78660 -41010
rect 78337 -41059 78371 -41039
rect 78519 -41029 78660 -41011
rect 78056 -41090 78126 -41079
rect 78056 -41180 78070 -41090
rect 78110 -41180 78126 -41090
rect 78163 -41093 78485 -41059
rect 78553 -41030 78660 -41029
rect 78553 -41063 78570 -41030
rect 78519 -41080 78570 -41063
rect 78451 -41127 78485 -41093
rect 78539 -41100 78570 -41080
rect 78640 -41100 78660 -41030
rect 78056 -41193 78126 -41180
rect 78160 -41140 78302 -41127
rect 77725 -41371 77733 -41337
rect 77767 -41371 77785 -41337
rect 77725 -41387 77785 -41371
rect 77825 -41345 77841 -41311
rect 77875 -41345 77891 -41311
rect 77825 -41379 77891 -41345
rect 77825 -41413 77841 -41379
rect 77875 -41413 77891 -41379
rect 77825 -41455 77891 -41413
rect 77929 -41345 77945 -41311
rect 77979 -41345 78021 -41311
rect 78056 -41248 78120 -41227
rect 78056 -41282 78073 -41248
rect 78107 -41282 78120 -41248
rect 78160 -41230 78190 -41140
rect 78280 -41230 78302 -41140
rect 78336 -41140 78417 -41127
rect 78336 -41180 78360 -41140
rect 78400 -41143 78417 -41140
rect 78409 -41177 78417 -41143
rect 78400 -41180 78417 -41177
rect 78336 -41193 78417 -41180
rect 78451 -41143 78505 -41127
rect 78451 -41177 78471 -41143
rect 78451 -41193 78505 -41177
rect 78539 -41170 78660 -41100
rect 78451 -41227 78485 -41193
rect 78539 -41227 78570 -41170
rect 78160 -41251 78302 -41230
rect 78056 -41285 78120 -41282
rect 78340 -41261 78485 -41227
rect 78519 -41240 78570 -41227
rect 78640 -41240 78660 -41170
rect 78340 -41285 78374 -41261
rect 78056 -41319 78374 -41285
rect 78519 -41280 78660 -41240
rect 78421 -41311 78477 -41295
rect 77929 -41360 78021 -41345
rect 78421 -41345 78434 -41311
rect 78468 -41345 78477 -41311
rect 78056 -41360 78387 -41353
rect 77929 -41367 78387 -41360
rect 77929 -41379 78295 -41367
rect 77929 -41413 77945 -41379
rect 77979 -41401 78295 -41379
rect 78329 -41401 78387 -41367
rect 77979 -41411 78387 -41401
rect 78421 -41379 78477 -41345
rect 77979 -41413 78380 -41411
rect 77929 -41420 78380 -41413
rect 78421 -41413 78434 -41379
rect 78468 -41413 78477 -41379
rect 77929 -41421 78021 -41420
rect 78421 -41455 78477 -41413
rect 78553 -41310 78660 -41280
rect 78553 -41314 78570 -41310
rect 78519 -41348 78570 -41314
rect 78553 -41380 78570 -41348
rect 78640 -41380 78660 -41310
rect 78553 -41382 78660 -41380
rect 78519 -41420 78660 -41382
rect 78519 -41421 78573 -41420
rect 59772 -41460 60520 -41457
rect 59772 -41520 59806 -41460
rect 59276 -41638 59310 -41576
rect 58930 -41672 59026 -41638
rect 59214 -41640 59310 -41638
rect 59214 -41672 59696 -41640
rect 58930 -41674 59696 -41672
rect 58930 -41710 58964 -41674
rect 57129 -41791 57131 -41757
rect 57129 -41825 57165 -41791
rect 57129 -41859 57131 -41825
rect 57129 -41875 57165 -41859
rect 57201 -41791 57217 -41757
rect 57251 -41791 57267 -41757
rect 57201 -41825 57267 -41791
rect 57201 -41859 57217 -41825
rect 57251 -41859 57267 -41825
rect 57201 -41909 57267 -41859
rect 57301 -41778 57303 -41744
rect 57337 -41778 57355 -41744
rect 57301 -41825 57355 -41778
rect 57301 -41859 57303 -41825
rect 57337 -41859 57355 -41825
rect 57301 -41875 57355 -41859
rect 59662 -41730 59696 -41674
rect 60486 -41522 60520 -41460
rect 77578 -41489 77607 -41455
rect 77641 -41489 77699 -41455
rect 77733 -41489 77791 -41455
rect 77825 -41489 77883 -41455
rect 77917 -41489 77975 -41455
rect 78009 -41489 78067 -41455
rect 78101 -41489 78159 -41455
rect 78193 -41489 78251 -41455
rect 78285 -41489 78343 -41455
rect 78377 -41489 78435 -41455
rect 78469 -41489 78527 -41455
rect 78561 -41489 78590 -41455
rect 59942 -41574 59958 -41540
rect 60334 -41574 60350 -41540
rect 59874 -41594 59908 -41578
rect 59874 -41644 59908 -41628
rect 60384 -41594 60418 -41578
rect 60384 -41644 60418 -41628
rect 59942 -41682 59958 -41648
rect 60334 -41682 60350 -41648
rect 56112 -41982 56146 -41920
rect 57096 -41943 57125 -41909
rect 57159 -41943 57217 -41909
rect 57251 -41943 57309 -41909
rect 57343 -41943 57372 -41909
rect 55706 -42016 55802 -41982
rect 56050 -42016 56146 -41982
rect 53886 -42064 53982 -42030
rect 54956 -42064 55052 -42030
rect 53886 -42126 53920 -42064
rect 55018 -42126 55052 -42064
rect 55720 -42058 56090 -42016
rect 55720 -42068 56020 -42058
rect 54065 -42178 54081 -42144
rect 54857 -42178 54873 -42144
rect 53988 -42206 54022 -42190
rect 53988 -42260 54022 -42244
rect 54916 -42206 54950 -42190
rect 54916 -42260 54950 -42244
rect 54065 -42306 54081 -42272
rect 54857 -42306 54873 -42272
rect 53886 -42386 53920 -42324
rect 56010 -42208 56020 -42068
rect 56080 -42208 56090 -42058
rect 59109 -41788 59125 -41754
rect 59501 -41788 59517 -41754
rect 59560 -41808 59594 -41792
rect 59560 -41858 59594 -41842
rect 59109 -41896 59125 -41862
rect 59501 -41896 59517 -41862
rect 59032 -41916 59066 -41900
rect 59032 -41966 59066 -41950
rect 59109 -42004 59125 -41970
rect 59501 -42004 59517 -41970
rect 56010 -42218 56090 -42208
rect 59772 -41762 59806 -41700
rect 77578 -41565 77607 -41531
rect 77641 -41565 77699 -41531
rect 77733 -41565 77791 -41531
rect 77825 -41565 77883 -41531
rect 77917 -41565 77975 -41531
rect 78009 -41565 78038 -41531
rect 77635 -41649 77691 -41565
rect 77825 -41607 77891 -41565
rect 77635 -41683 77649 -41649
rect 77683 -41683 77691 -41649
rect 77635 -41699 77691 -41683
rect 77725 -41649 77785 -41633
rect 77725 -41683 77733 -41649
rect 77767 -41683 77785 -41649
rect 60486 -41762 60520 -41700
rect 77725 -41743 77785 -41683
rect 77825 -41641 77841 -41607
rect 77875 -41641 77891 -41607
rect 77825 -41675 77891 -41641
rect 77825 -41709 77841 -41675
rect 77875 -41709 77891 -41675
rect 77929 -41607 78021 -41599
rect 77929 -41641 77945 -41607
rect 77979 -41641 78021 -41607
rect 77929 -41675 78021 -41641
rect 77929 -41709 77945 -41675
rect 77979 -41709 78021 -41675
rect 77971 -41740 78021 -41709
rect 77598 -41760 77651 -41755
rect 59772 -41796 59866 -41762
rect 60426 -41796 60520 -41762
rect 77470 -41790 77690 -41760
rect 77725 -41777 77913 -41743
rect 77470 -41840 77510 -41790
rect 77560 -41827 77690 -41790
rect 77879 -41827 77913 -41777
rect 77971 -41780 77980 -41740
rect 78020 -41780 78021 -41740
rect 77560 -41840 77733 -41827
rect 77470 -41843 77733 -41840
rect 77470 -41870 77652 -41843
rect 77598 -41877 77652 -41870
rect 77686 -41877 77733 -41843
rect 77777 -41830 77845 -41827
rect 77777 -41870 77790 -41830
rect 77830 -41870 77845 -41830
rect 77777 -41877 77793 -41870
rect 77827 -41877 77845 -41870
rect 77879 -41843 77937 -41827
rect 77879 -41877 77901 -41843
rect 77935 -41877 77937 -41843
rect 77879 -41893 77937 -41877
rect 77971 -41860 78021 -41780
rect 77879 -41911 77913 -41893
rect 77635 -41949 77913 -41911
rect 77971 -41900 77980 -41860
rect 78020 -41900 78021 -41860
rect 59662 -42084 59696 -42030
rect 58966 -42100 59026 -42084
rect 58930 -42118 59026 -42100
rect 59600 -42118 59696 -42084
rect 77635 -41971 77701 -41949
rect 77635 -42005 77649 -41971
rect 77683 -42005 77701 -41971
rect 77971 -41960 78021 -41900
rect 77971 -41983 77980 -41960
rect 77635 -42021 77701 -42005
rect 77825 -41999 77875 -41983
rect 77825 -42033 77841 -41999
rect 77825 -42075 77875 -42033
rect 77909 -41999 77980 -41983
rect 77909 -42033 77925 -41999
rect 77959 -42000 77980 -41999
rect 78020 -42000 78021 -41960
rect 77959 -42033 78021 -42000
rect 77909 -42041 78021 -42033
rect 77578 -42109 77607 -42075
rect 77641 -42109 77699 -42075
rect 77733 -42109 77791 -42075
rect 77825 -42109 77883 -42075
rect 77917 -42109 77975 -42075
rect 78009 -42109 78038 -42075
rect 77580 -42199 77609 -42165
rect 77643 -42199 77701 -42165
rect 77735 -42199 77793 -42165
rect 77827 -42199 77885 -42165
rect 77919 -42199 77977 -42165
rect 78011 -42199 78040 -42165
rect 55018 -42386 55052 -42324
rect 53886 -42420 53982 -42386
rect 54956 -42420 55052 -42386
rect 55176 -42278 55272 -42244
rect 55566 -42278 55662 -42244
rect 77827 -42241 77877 -42199
rect 55176 -42340 55210 -42278
rect 55628 -42340 55662 -42278
rect 55284 -42392 55300 -42358
rect 55476 -42392 55492 -42358
rect 55526 -42402 55560 -42386
rect 55284 -42480 55300 -42446
rect 55476 -42480 55492 -42446
rect 55526 -42452 55560 -42436
rect 55176 -42560 55210 -42498
rect 77637 -42269 77703 -42253
rect 77637 -42303 77651 -42269
rect 77685 -42303 77703 -42269
rect 77827 -42275 77843 -42241
rect 77827 -42291 77877 -42275
rect 77911 -42241 78023 -42233
rect 77911 -42275 77927 -42241
rect 77961 -42275 78023 -42241
rect 77911 -42291 78023 -42275
rect 77637 -42325 77703 -42303
rect 77637 -42363 77915 -42325
rect 77881 -42381 77915 -42363
rect 77973 -42340 78023 -42291
rect 77973 -42380 77980 -42340
rect 78020 -42380 78023 -42340
rect 77881 -42397 77939 -42381
rect 77600 -42400 77654 -42397
rect 55628 -42560 55662 -42498
rect 77440 -42430 77654 -42400
rect 77440 -42480 77490 -42430
rect 77540 -42431 77654 -42430
rect 77688 -42431 77735 -42397
rect 77540 -42447 77735 -42431
rect 77779 -42400 77795 -42397
rect 77829 -42400 77847 -42397
rect 77779 -42440 77790 -42400
rect 77830 -42440 77847 -42400
rect 77779 -42447 77847 -42440
rect 77881 -42431 77903 -42397
rect 77937 -42431 77939 -42397
rect 77881 -42447 77939 -42431
rect 77973 -42420 78023 -42380
rect 77540 -42480 77690 -42447
rect 77440 -42510 77690 -42480
rect 77881 -42497 77915 -42447
rect 77600 -42519 77653 -42510
rect 55176 -42594 55272 -42560
rect 55566 -42594 55662 -42560
rect 77727 -42531 77915 -42497
rect 77973 -42460 77980 -42420
rect 78020 -42460 78023 -42420
rect 77973 -42520 78023 -42460
rect 77637 -42591 77693 -42575
rect 77637 -42625 77651 -42591
rect 77685 -42625 77693 -42591
rect 77637 -42709 77693 -42625
rect 77727 -42591 77787 -42531
rect 77973 -42560 77980 -42520
rect 78020 -42560 78023 -42520
rect 77973 -42565 78023 -42560
rect 77727 -42625 77735 -42591
rect 77769 -42625 77787 -42591
rect 77727 -42641 77787 -42625
rect 77827 -42599 77843 -42565
rect 77877 -42599 77893 -42565
rect 77827 -42633 77893 -42599
rect 77827 -42667 77843 -42633
rect 77877 -42667 77893 -42633
rect 77827 -42709 77893 -42667
rect 77931 -42599 77947 -42565
rect 77981 -42599 78023 -42565
rect 77931 -42600 78023 -42599
rect 77931 -42633 77980 -42600
rect 77931 -42667 77947 -42633
rect 78020 -42640 78023 -42600
rect 77981 -42667 78023 -42640
rect 77931 -42675 78023 -42667
rect 77580 -42743 77609 -42709
rect 77643 -42743 77701 -42709
rect 77735 -42743 77793 -42709
rect 77827 -42743 77885 -42709
rect 77919 -42743 77977 -42709
rect 78011 -42743 78040 -42709
rect 77578 -42815 77607 -42781
rect 77641 -42815 77699 -42781
rect 77733 -42815 77791 -42781
rect 77825 -42815 77883 -42781
rect 77917 -42815 77975 -42781
rect 78009 -42815 78067 -42781
rect 78101 -42815 78159 -42781
rect 78193 -42815 78222 -42781
rect 78322 -42815 78351 -42781
rect 78385 -42815 78443 -42781
rect 78477 -42815 78535 -42781
rect 78569 -42815 78627 -42781
rect 78661 -42815 78719 -42781
rect 78753 -42815 78811 -42781
rect 78845 -42815 78874 -42781
rect 77596 -42857 77663 -42815
rect 77596 -42891 77613 -42857
rect 77647 -42891 77663 -42857
rect 77697 -42865 77747 -42849
rect 77697 -42899 77705 -42865
rect 77739 -42899 77747 -42865
rect 77595 -42930 77643 -42927
rect 77570 -42940 77643 -42930
rect 77570 -42990 77580 -42940
rect 77630 -42990 77643 -42940
rect 77570 -43093 77643 -42990
rect 77697 -43009 77747 -42899
rect 77791 -42857 77857 -42815
rect 77791 -42891 77807 -42857
rect 77841 -42891 77857 -42857
rect 77791 -42959 77857 -42891
rect 77894 -42865 77944 -42849
rect 77894 -42899 77902 -42865
rect 77936 -42899 77944 -42865
rect 77894 -43009 77944 -42899
rect 78037 -42857 78103 -42815
rect 78037 -42891 78053 -42857
rect 78087 -42891 78103 -42857
rect 78037 -42925 78103 -42891
rect 78137 -42857 78205 -42849
rect 78137 -42891 78153 -42857
rect 78187 -42891 78205 -42857
rect 78137 -42901 78205 -42891
rect 78037 -42959 78053 -42925
rect 78087 -42959 78103 -42925
rect 78037 -42975 78103 -42959
rect 78153 -42925 78205 -42901
rect 78187 -42959 78205 -42925
rect 78240 -42859 78340 -42850
rect 78705 -42857 78761 -42815
rect 78240 -42869 78671 -42859
rect 78240 -42889 78579 -42869
rect 78240 -42923 78250 -42889
rect 78290 -42903 78579 -42889
rect 78613 -42903 78671 -42869
rect 78290 -42917 78671 -42903
rect 78705 -42891 78718 -42857
rect 78752 -42891 78761 -42857
rect 78290 -42920 78310 -42917
rect 78290 -42923 78300 -42920
rect 78240 -42950 78300 -42923
rect 78705 -42925 78761 -42891
rect 78153 -42993 78205 -42959
rect 77570 -43127 77609 -43093
rect 77570 -43189 77643 -43127
rect 77677 -43043 78115 -43009
rect 77570 -43190 77640 -43189
rect 77677 -43225 77711 -43043
rect 78052 -43077 78115 -43043
rect 78187 -43010 78205 -42993
rect 78340 -42985 78658 -42951
rect 78705 -42959 78718 -42925
rect 78752 -42959 78761 -42925
rect 78705 -42975 78761 -42959
rect 78803 -42850 78857 -42849
rect 78803 -42888 78920 -42850
rect 78837 -42920 78920 -42888
rect 78837 -42922 78850 -42920
rect 78803 -42956 78850 -42922
rect 78340 -42988 78404 -42985
rect 77612 -43241 77711 -43225
rect 77612 -43275 77613 -43241
rect 77647 -43275 77711 -43241
rect 77755 -43090 77825 -43077
rect 77755 -43093 77770 -43090
rect 77755 -43130 77770 -43127
rect 77810 -43130 77825 -43090
rect 77755 -43270 77825 -43130
rect 77861 -43093 77921 -43077
rect 77895 -43120 77921 -43093
rect 77861 -43160 77870 -43127
rect 77910 -43160 77921 -43120
rect 77861 -43200 77921 -43160
rect 77861 -43240 77870 -43200
rect 77910 -43240 77921 -43200
rect 77861 -43271 77921 -43240
rect 77957 -43093 78013 -43077
rect 77991 -43127 78013 -43093
rect 78052 -43093 78118 -43077
rect 78052 -43127 78068 -43093
rect 78102 -43127 78118 -43093
rect 77957 -43210 78013 -43127
rect 77957 -43250 77970 -43210
rect 78010 -43250 78013 -43210
rect 77957 -43271 78013 -43250
rect 78049 -43181 78103 -43165
rect 78153 -43180 78170 -43027
rect 78340 -43022 78357 -42988
rect 78391 -43022 78404 -42988
rect 78624 -43009 78658 -42985
rect 78837 -42970 78850 -42956
rect 78900 -42970 78920 -42920
rect 78837 -42990 78920 -42970
rect 78340 -43043 78404 -43022
rect 78444 -43040 78586 -43019
rect 78153 -43181 78220 -43180
rect 78049 -43215 78054 -43181
rect 78088 -43215 78103 -43181
rect 78049 -43249 78103 -43215
rect 77612 -43291 77711 -43275
rect 78049 -43283 78054 -43249
rect 78088 -43283 78103 -43249
rect 78137 -43215 78153 -43181
rect 78187 -43200 78220 -43181
rect 78340 -43093 78410 -43077
rect 78340 -43127 78357 -43093
rect 78391 -43127 78410 -43093
rect 78340 -43140 78410 -43127
rect 78340 -43180 78350 -43140
rect 78400 -43180 78410 -43140
rect 78444 -43090 78470 -43040
rect 78560 -43090 78586 -43040
rect 78624 -43043 78769 -43009
rect 78803 -43040 78920 -42990
rect 78803 -43043 78850 -43040
rect 78735 -43077 78769 -43043
rect 78444 -43093 78586 -43090
rect 78444 -43127 78483 -43093
rect 78517 -43127 78586 -43093
rect 78444 -43143 78586 -43127
rect 78620 -43090 78701 -43077
rect 78620 -43130 78640 -43090
rect 78690 -43093 78701 -43090
rect 78693 -43127 78701 -43093
rect 78690 -43130 78701 -43127
rect 78620 -43143 78701 -43130
rect 78735 -43093 78789 -43077
rect 78735 -43127 78755 -43093
rect 78735 -43143 78789 -43127
rect 78823 -43090 78850 -43043
rect 78900 -43090 78920 -43040
rect 78735 -43177 78769 -43143
rect 78340 -43191 78410 -43180
rect 78187 -43215 78205 -43200
rect 78137 -43249 78205 -43215
rect 78447 -43211 78769 -43177
rect 78823 -43160 78920 -43090
rect 78823 -43190 78850 -43160
rect 78803 -43207 78850 -43190
rect 78137 -43283 78153 -43249
rect 78187 -43283 78205 -43249
rect 78341 -43259 78357 -43225
rect 78391 -43259 78407 -43225
rect 78049 -43325 78103 -43283
rect 78341 -43325 78407 -43259
rect 78447 -43231 78481 -43211
rect 78621 -43231 78655 -43211
rect 78447 -43281 78481 -43265
rect 78521 -43279 78537 -43245
rect 78571 -43279 78587 -43245
rect 78521 -43325 78587 -43279
rect 78837 -43210 78850 -43207
rect 78900 -43210 78920 -43160
rect 78837 -43241 78920 -43210
rect 78621 -43281 78655 -43265
rect 78689 -43279 78715 -43245
rect 78749 -43279 78765 -43245
rect 78803 -43259 78920 -43241
rect 78830 -43260 78920 -43259
rect 78689 -43325 78765 -43279
rect 77578 -43359 77607 -43325
rect 77641 -43359 77699 -43325
rect 77733 -43359 77791 -43325
rect 77825 -43359 77883 -43325
rect 77917 -43359 77975 -43325
rect 78009 -43359 78067 -43325
rect 78101 -43359 78159 -43325
rect 78193 -43359 78222 -43325
rect 78322 -43359 78351 -43325
rect 78385 -43359 78443 -43325
rect 78477 -43359 78535 -43325
rect 78569 -43359 78627 -43325
rect 78661 -43359 78719 -43325
rect 78753 -43359 78811 -43325
rect 78845 -43359 78874 -43325
rect 77578 -43431 77607 -43397
rect 77641 -43431 77699 -43397
rect 77733 -43431 77791 -43397
rect 77825 -43431 77883 -43397
rect 77917 -43431 77975 -43397
rect 78009 -43431 78067 -43397
rect 78101 -43431 78159 -43397
rect 78193 -43431 78222 -43397
rect 77612 -43481 77711 -43465
rect 77612 -43515 77613 -43481
rect 77647 -43515 77711 -43481
rect 78049 -43473 78103 -43431
rect 77612 -43531 77711 -43515
rect 77595 -43629 77643 -43567
rect 77595 -43663 77609 -43629
rect 77595 -43700 77643 -43663
rect 35802 -43788 35836 -43726
rect 25780 -43830 35836 -43788
rect 35802 -43892 35836 -43830
rect 77420 -43770 77643 -43700
rect 77677 -43713 77711 -43531
rect 77755 -43520 77825 -43486
rect 77755 -43560 77770 -43520
rect 77810 -43560 77825 -43520
rect 77755 -43610 77825 -43560
rect 77755 -43629 77770 -43610
rect 77810 -43650 77825 -43610
rect 77789 -43663 77825 -43650
rect 77755 -43679 77825 -43663
rect 77861 -43540 77921 -43485
rect 77861 -43580 77870 -43540
rect 77910 -43580 77921 -43540
rect 77861 -43620 77921 -43580
rect 77861 -43629 77870 -43620
rect 77910 -43660 77921 -43620
rect 77895 -43663 77921 -43660
rect 77861 -43679 77921 -43663
rect 77957 -43629 78013 -43485
rect 78049 -43507 78054 -43473
rect 78088 -43507 78103 -43473
rect 78049 -43541 78103 -43507
rect 78049 -43575 78054 -43541
rect 78088 -43575 78103 -43541
rect 78137 -43507 78153 -43473
rect 78187 -43490 78205 -43473
rect 78187 -43507 78300 -43490
rect 78137 -43510 78300 -43507
rect 78137 -43541 78200 -43510
rect 78137 -43575 78153 -43541
rect 78187 -43560 78200 -43541
rect 78280 -43560 78300 -43510
rect 78187 -43575 78300 -43560
rect 78049 -43591 78103 -43575
rect 77991 -43630 78013 -43629
rect 77957 -43670 77970 -43663
rect 78010 -43670 78013 -43630
rect 77957 -43679 78013 -43670
rect 78052 -43663 78068 -43629
rect 78102 -43663 78118 -43629
rect 78052 -43679 78118 -43663
rect 78153 -43650 78300 -43575
rect 82838 -43625 82867 -43591
rect 82901 -43625 82959 -43591
rect 82993 -43625 83051 -43591
rect 83085 -43625 83143 -43591
rect 83177 -43625 83235 -43591
rect 83269 -43625 83327 -43591
rect 83361 -43625 83419 -43591
rect 83453 -43625 83511 -43591
rect 83545 -43625 83603 -43591
rect 83637 -43625 83695 -43591
rect 83729 -43625 83787 -43591
rect 83821 -43625 83879 -43591
rect 83913 -43625 83971 -43591
rect 84005 -43625 84063 -43591
rect 84097 -43625 84155 -43591
rect 84189 -43625 84247 -43591
rect 84281 -43625 84339 -43591
rect 84373 -43625 84431 -43591
rect 84465 -43625 84523 -43591
rect 84557 -43625 84615 -43591
rect 84649 -43625 84707 -43591
rect 84741 -43625 84799 -43591
rect 84833 -43625 84891 -43591
rect 84925 -43625 84983 -43591
rect 85017 -43625 85075 -43591
rect 85109 -43625 85167 -43591
rect 85201 -43625 85259 -43591
rect 85293 -43625 85351 -43591
rect 85385 -43625 85443 -43591
rect 85477 -43625 85535 -43591
rect 85569 -43625 85627 -43591
rect 85661 -43625 85719 -43591
rect 85753 -43625 85811 -43591
rect 85845 -43625 85903 -43591
rect 85937 -43625 85995 -43591
rect 86029 -43625 86087 -43591
rect 86121 -43625 86179 -43591
rect 86213 -43625 86271 -43591
rect 86305 -43625 86363 -43591
rect 86397 -43625 86455 -43591
rect 86489 -43625 86547 -43591
rect 86581 -43625 86639 -43591
rect 86673 -43625 86731 -43591
rect 86765 -43625 86823 -43591
rect 86857 -43625 86915 -43591
rect 86949 -43625 87007 -43591
rect 87041 -43625 87099 -43591
rect 87133 -43625 87191 -43591
rect 87225 -43625 87283 -43591
rect 87317 -43625 87375 -43591
rect 87409 -43625 87467 -43591
rect 87501 -43625 87559 -43591
rect 87593 -43625 87651 -43591
rect 87685 -43625 87743 -43591
rect 87777 -43625 87835 -43591
rect 87869 -43625 87927 -43591
rect 87961 -43625 88019 -43591
rect 88053 -43625 88111 -43591
rect 88145 -43625 88203 -43591
rect 88237 -43625 88295 -43591
rect 88329 -43625 88387 -43591
rect 88421 -43625 88479 -43591
rect 88513 -43625 88571 -43591
rect 88605 -43625 88663 -43591
rect 88697 -43625 88755 -43591
rect 88789 -43625 88847 -43591
rect 88881 -43625 88939 -43591
rect 88973 -43625 89031 -43591
rect 89065 -43625 89123 -43591
rect 89157 -43625 89215 -43591
rect 89249 -43625 89307 -43591
rect 89341 -43625 89399 -43591
rect 89433 -43625 89491 -43591
rect 89525 -43625 89583 -43591
rect 89617 -43625 89675 -43591
rect 89709 -43625 89767 -43591
rect 89801 -43625 89859 -43591
rect 89893 -43625 89951 -43591
rect 89985 -43625 90043 -43591
rect 90077 -43625 90135 -43591
rect 90169 -43625 90227 -43591
rect 90261 -43625 90319 -43591
rect 90353 -43625 90411 -43591
rect 90445 -43625 90503 -43591
rect 90537 -43625 90595 -43591
rect 90629 -43625 90687 -43591
rect 90721 -43625 90779 -43591
rect 90813 -43625 90871 -43591
rect 90905 -43625 90963 -43591
rect 90997 -43625 91055 -43591
rect 91089 -43625 91147 -43591
rect 91181 -43625 91239 -43591
rect 91273 -43625 91331 -43591
rect 91365 -43625 91394 -43591
rect 78052 -43713 78115 -43679
rect 77677 -43747 78115 -43713
rect 78153 -43700 78200 -43650
rect 78280 -43700 78300 -43650
rect 78153 -43729 78300 -43700
rect 77420 -43820 77440 -43770
rect 77490 -43820 77643 -43770
rect 77420 -43840 77530 -43820
rect 77595 -43829 77643 -43820
rect 77697 -43857 77747 -43747
rect 77596 -43899 77613 -43865
rect 77647 -43899 77663 -43865
rect 77596 -43941 77663 -43899
rect 77697 -43891 77705 -43857
rect 77739 -43891 77747 -43857
rect 77697 -43907 77747 -43891
rect 77791 -43865 77857 -43797
rect 77791 -43899 77807 -43865
rect 77841 -43899 77857 -43865
rect 77791 -43941 77857 -43899
rect 77894 -43857 77944 -43747
rect 78187 -43763 78300 -43729
rect 77894 -43891 77902 -43857
rect 77936 -43891 77944 -43857
rect 77894 -43907 77944 -43891
rect 78037 -43797 78103 -43781
rect 78037 -43831 78053 -43797
rect 78087 -43831 78103 -43797
rect 78037 -43865 78103 -43831
rect 78153 -43790 78300 -43763
rect 83067 -43683 83133 -43625
rect 83067 -43717 83083 -43683
rect 83117 -43717 83133 -43683
rect 83067 -43751 83133 -43717
rect 78153 -43797 78200 -43790
rect 78187 -43831 78200 -43797
rect 78153 -43840 78200 -43831
rect 78280 -43840 78300 -43790
rect 78153 -43855 78300 -43840
rect 82892 -43803 82970 -43784
rect 83067 -43785 83083 -43751
rect 83117 -43785 83133 -43751
rect 83167 -43667 83274 -43659
rect 83167 -43701 83183 -43667
rect 83217 -43701 83274 -43667
rect 83167 -43735 83274 -43701
rect 83167 -43769 83183 -43735
rect 83217 -43769 83274 -43735
rect 83167 -43783 83274 -43769
rect 82892 -43837 82914 -43803
rect 82948 -43819 82970 -43803
rect 82948 -43837 83177 -43819
rect 82892 -43853 83177 -43837
rect 78037 -43899 78053 -43865
rect 78087 -43899 78103 -43865
rect 78037 -43941 78103 -43899
rect 78137 -43865 78300 -43855
rect 78137 -43899 78153 -43865
rect 78187 -43880 78300 -43865
rect 78187 -43899 78205 -43880
rect 78137 -43907 78205 -43899
rect 82867 -43900 82938 -43887
rect 77578 -43975 77607 -43941
rect 77641 -43975 77699 -43941
rect 77733 -43975 77791 -43941
rect 77825 -43975 77883 -43941
rect 77917 -43975 77975 -43941
rect 78009 -43975 78067 -43941
rect 78101 -43975 78159 -43941
rect 78193 -43975 78222 -43941
rect 77578 -44047 77607 -44013
rect 77641 -44047 77699 -44013
rect 77733 -44047 77791 -44013
rect 77825 -44047 77883 -44013
rect 77917 -44047 77975 -44013
rect 78009 -44047 78067 -44013
rect 78101 -44047 78159 -44013
rect 78193 -44047 78222 -44013
rect 77596 -44089 77663 -44047
rect 77596 -44123 77613 -44089
rect 77647 -44123 77663 -44089
rect 77697 -44097 77747 -44081
rect 77697 -44131 77705 -44097
rect 77739 -44131 77747 -44097
rect 77450 -44160 77530 -44150
rect 77595 -44160 77643 -44159
rect 77450 -44170 77643 -44160
rect 77450 -44220 77470 -44170
rect 77510 -44220 77643 -44170
rect 77450 -44230 77643 -44220
rect 77450 -44240 77530 -44230
rect 77595 -44325 77643 -44230
rect 77697 -44241 77747 -44131
rect 77791 -44089 77857 -44047
rect 77791 -44123 77807 -44089
rect 77841 -44123 77857 -44089
rect 77791 -44191 77857 -44123
rect 77894 -44097 77944 -44081
rect 77894 -44131 77902 -44097
rect 77936 -44131 77944 -44097
rect 77894 -44241 77944 -44131
rect 78037 -44089 78103 -44047
rect 82867 -43990 82880 -43900
rect 82930 -43903 82938 -43900
rect 82930 -43990 82938 -43937
rect 82867 -43999 82938 -43990
rect 82972 -44033 83006 -43853
rect 83040 -43903 83093 -43887
rect 83074 -43910 83093 -43903
rect 83040 -43990 83050 -43937
rect 83090 -43990 83093 -43910
rect 83143 -43903 83177 -43853
rect 83143 -43953 83177 -43937
rect 83211 -43870 83274 -43783
rect 83366 -43667 83408 -43625
rect 83366 -43701 83374 -43667
rect 83366 -43735 83408 -43701
rect 83366 -43769 83374 -43735
rect 83366 -43803 83408 -43769
rect 83366 -43837 83374 -43803
rect 83366 -43853 83408 -43837
rect 83442 -43667 83508 -43659
rect 83442 -43701 83458 -43667
rect 83492 -43701 83508 -43667
rect 83442 -43735 83508 -43701
rect 83442 -43769 83458 -43735
rect 83492 -43769 83508 -43735
rect 83442 -43803 83508 -43769
rect 83442 -43837 83458 -43803
rect 83492 -43837 83508 -43803
rect 83442 -43855 83508 -43837
rect 83600 -43667 83653 -43625
rect 83600 -43701 83619 -43667
rect 83600 -43735 83653 -43701
rect 83600 -43769 83619 -43735
rect 83600 -43803 83653 -43769
rect 83600 -43837 83619 -43803
rect 83600 -43853 83653 -43837
rect 83687 -43667 83753 -43659
rect 83687 -43701 83703 -43667
rect 83737 -43701 83753 -43667
rect 83687 -43735 83753 -43701
rect 83687 -43769 83703 -43735
rect 83737 -43769 83753 -43735
rect 83687 -43803 83753 -43769
rect 83787 -43667 83821 -43625
rect 83787 -43735 83821 -43701
rect 83787 -43785 83821 -43769
rect 83855 -43667 83921 -43659
rect 83855 -43701 83871 -43667
rect 83905 -43701 83921 -43667
rect 83855 -43735 83921 -43701
rect 83955 -43667 83997 -43625
rect 83989 -43701 83997 -43667
rect 83955 -43717 83997 -43701
rect 84074 -43667 84116 -43625
rect 84074 -43701 84082 -43667
rect 83855 -43769 83871 -43735
rect 83905 -43769 83921 -43735
rect 83687 -43837 83703 -43803
rect 83737 -43819 83753 -43803
rect 83855 -43803 83921 -43769
rect 83855 -43819 83871 -43803
rect 83737 -43837 83871 -43819
rect 83905 -43815 83921 -43803
rect 84074 -43735 84116 -43701
rect 84074 -43769 84082 -43735
rect 84074 -43805 84116 -43769
rect 83905 -43837 84008 -43815
rect 83687 -43853 84008 -43837
rect 83211 -43890 83320 -43870
rect 83362 -43890 83428 -43889
rect 83211 -43903 83428 -43890
rect 83211 -43930 83378 -43903
rect 83211 -43950 83320 -43930
rect 83362 -43937 83378 -43930
rect 83412 -43937 83428 -43903
rect 83462 -43890 83508 -43855
rect 83595 -43890 83921 -43887
rect 83462 -43903 83921 -43890
rect 83462 -43937 83611 -43903
rect 83645 -43937 83703 -43903
rect 83737 -43937 83787 -43903
rect 83821 -43937 83871 -43903
rect 83905 -43937 83921 -43903
rect 83955 -43890 84008 -43853
rect 84074 -43839 84082 -43805
rect 84074 -43855 84116 -43839
rect 84150 -43667 84216 -43659
rect 84150 -43701 84166 -43667
rect 84200 -43701 84216 -43667
rect 84150 -43735 84216 -43701
rect 84150 -43769 84166 -43735
rect 84200 -43769 84216 -43735
rect 84150 -43805 84216 -43769
rect 84250 -43667 84284 -43625
rect 84250 -43735 84284 -43701
rect 84250 -43785 84284 -43769
rect 84318 -43667 84384 -43659
rect 84318 -43701 84334 -43667
rect 84368 -43701 84384 -43667
rect 84318 -43735 84384 -43701
rect 84318 -43769 84334 -43735
rect 84368 -43769 84384 -43735
rect 84150 -43839 84166 -43805
rect 84200 -43819 84216 -43805
rect 84318 -43805 84384 -43769
rect 84418 -43667 84452 -43625
rect 84418 -43735 84452 -43701
rect 84418 -43785 84452 -43769
rect 84486 -43667 84552 -43659
rect 84486 -43701 84502 -43667
rect 84536 -43701 84552 -43667
rect 84486 -43735 84552 -43701
rect 84486 -43769 84502 -43735
rect 84536 -43769 84552 -43735
rect 84318 -43819 84334 -43805
rect 84200 -43839 84334 -43819
rect 84368 -43819 84384 -43805
rect 84486 -43805 84552 -43769
rect 84586 -43667 84620 -43625
rect 84586 -43735 84620 -43701
rect 84586 -43785 84620 -43769
rect 84654 -43667 84720 -43659
rect 84654 -43701 84670 -43667
rect 84704 -43701 84720 -43667
rect 84654 -43735 84720 -43701
rect 84654 -43769 84670 -43735
rect 84704 -43769 84720 -43735
rect 84486 -43819 84502 -43805
rect 84368 -43839 84502 -43819
rect 84536 -43819 84552 -43805
rect 84654 -43805 84720 -43769
rect 84754 -43667 84788 -43625
rect 84754 -43735 84788 -43701
rect 84754 -43785 84788 -43769
rect 84822 -43667 84888 -43659
rect 84822 -43701 84838 -43667
rect 84872 -43701 84888 -43667
rect 84822 -43735 84888 -43701
rect 84822 -43769 84838 -43735
rect 84872 -43769 84888 -43735
rect 84654 -43819 84670 -43805
rect 84536 -43839 84670 -43819
rect 84704 -43819 84720 -43805
rect 84822 -43805 84888 -43769
rect 84922 -43667 84956 -43625
rect 84922 -43735 84956 -43701
rect 84922 -43785 84956 -43769
rect 84990 -43667 85056 -43659
rect 84990 -43701 85006 -43667
rect 85040 -43701 85056 -43667
rect 84990 -43735 85056 -43701
rect 84990 -43769 85006 -43735
rect 85040 -43769 85056 -43735
rect 84822 -43819 84838 -43805
rect 84704 -43839 84838 -43819
rect 84872 -43819 84888 -43805
rect 84990 -43805 85056 -43769
rect 85090 -43667 85124 -43625
rect 85090 -43735 85124 -43701
rect 85090 -43785 85124 -43769
rect 85158 -43667 85224 -43659
rect 85158 -43701 85174 -43667
rect 85208 -43701 85224 -43667
rect 85158 -43735 85224 -43701
rect 85158 -43769 85174 -43735
rect 85208 -43769 85224 -43735
rect 84990 -43819 85006 -43805
rect 84872 -43839 85006 -43819
rect 85040 -43819 85056 -43805
rect 85158 -43805 85224 -43769
rect 85258 -43667 85292 -43625
rect 85258 -43735 85292 -43701
rect 85258 -43785 85292 -43769
rect 85326 -43667 85392 -43659
rect 85326 -43701 85342 -43667
rect 85376 -43701 85392 -43667
rect 85326 -43735 85392 -43701
rect 85326 -43769 85342 -43735
rect 85376 -43769 85392 -43735
rect 85158 -43819 85174 -43805
rect 85040 -43839 85174 -43819
rect 85208 -43819 85224 -43805
rect 85326 -43805 85392 -43769
rect 85426 -43667 85468 -43625
rect 85460 -43701 85468 -43667
rect 85426 -43735 85468 -43701
rect 85460 -43769 85468 -43735
rect 85426 -43785 85468 -43769
rect 85546 -43667 85588 -43625
rect 85546 -43701 85554 -43667
rect 85546 -43735 85588 -43701
rect 85546 -43769 85554 -43735
rect 85326 -43819 85342 -43805
rect 85208 -43820 85342 -43819
rect 85376 -43820 85392 -43805
rect 85208 -43839 85330 -43820
rect 84150 -43853 85330 -43839
rect 84051 -43890 85139 -43889
rect 83955 -43903 85139 -43890
rect 83955 -43937 84076 -43903
rect 84110 -43937 84250 -43903
rect 84284 -43937 84418 -43903
rect 84452 -43937 84587 -43903
rect 84621 -43937 84754 -43903
rect 84788 -43937 84922 -43903
rect 84956 -43937 85089 -43903
rect 85123 -43937 85139 -43903
rect 83462 -43940 83640 -43937
rect 83955 -43940 84100 -43937
rect 83211 -43987 83274 -43950
rect 83040 -43999 83093 -43990
rect 83151 -43989 83274 -43987
rect 83151 -44023 83167 -43989
rect 83201 -44023 83274 -43989
rect 82888 -44049 82936 -44033
rect 78037 -44123 78053 -44089
rect 78087 -44123 78103 -44089
rect 78037 -44157 78103 -44123
rect 78137 -44089 78205 -44081
rect 78137 -44123 78153 -44089
rect 78187 -44090 78205 -44089
rect 82888 -44083 82902 -44049
rect 78187 -44123 78310 -44090
rect 78137 -44133 78310 -44123
rect 78037 -44191 78053 -44157
rect 78087 -44191 78103 -44157
rect 78037 -44207 78103 -44191
rect 78153 -44140 78310 -44133
rect 82888 -44135 82936 -44083
rect 82972 -44049 83028 -44033
rect 82972 -44083 82986 -44049
rect 83020 -44083 83028 -44049
rect 82972 -44099 83028 -44083
rect 83074 -44049 83117 -44033
rect 83074 -44083 83082 -44049
rect 83116 -44083 83117 -44049
rect 83074 -44135 83117 -44083
rect 83151 -44057 83274 -44023
rect 83151 -44091 83167 -44057
rect 83201 -44091 83274 -44057
rect 83151 -44101 83274 -44091
rect 83362 -43987 83408 -43971
rect 83462 -43975 83508 -43940
rect 83955 -43971 84008 -43940
rect 85326 -43971 85330 -43853
rect 83362 -44021 83374 -43987
rect 83362 -44055 83408 -44021
rect 83362 -44089 83374 -44055
rect 83362 -44135 83408 -44089
rect 83442 -43987 83508 -43975
rect 83442 -44021 83458 -43987
rect 83492 -44021 83508 -43987
rect 83442 -44055 83508 -44021
rect 83687 -44007 84008 -43971
rect 84070 -43991 84116 -43975
rect 83442 -44089 83458 -44055
rect 83492 -44089 83508 -44055
rect 83442 -44101 83508 -44089
rect 83600 -44059 83653 -44043
rect 83600 -44093 83619 -44059
rect 83600 -44135 83653 -44093
rect 83687 -44051 83753 -44007
rect 83687 -44085 83703 -44051
rect 83737 -44085 83753 -44051
rect 83687 -44101 83753 -44085
rect 83787 -44059 83821 -44043
rect 83787 -44135 83821 -44093
rect 83855 -44051 83921 -44007
rect 84070 -44025 84082 -43991
rect 83855 -44085 83871 -44051
rect 83905 -44085 83921 -44051
rect 83855 -44101 83921 -44085
rect 83955 -44058 84005 -44042
rect 83989 -44092 84005 -44058
rect 83955 -44135 84005 -44092
rect 84070 -44059 84116 -44025
rect 84070 -44093 84082 -44059
rect 84070 -44135 84116 -44093
rect 84150 -43990 85330 -43971
rect 85380 -43990 85392 -43820
rect 85546 -43805 85588 -43769
rect 85546 -43839 85554 -43805
rect 85546 -43855 85588 -43839
rect 85622 -43667 85688 -43659
rect 85622 -43701 85638 -43667
rect 85672 -43701 85688 -43667
rect 85622 -43735 85688 -43701
rect 85622 -43769 85638 -43735
rect 85672 -43769 85688 -43735
rect 85622 -43805 85688 -43769
rect 85722 -43667 85756 -43625
rect 85722 -43735 85756 -43701
rect 85722 -43785 85756 -43769
rect 85790 -43667 85856 -43659
rect 85790 -43701 85806 -43667
rect 85840 -43701 85856 -43667
rect 85790 -43735 85856 -43701
rect 85790 -43769 85806 -43735
rect 85840 -43769 85856 -43735
rect 85622 -43839 85638 -43805
rect 85672 -43819 85688 -43805
rect 85790 -43805 85856 -43769
rect 85890 -43667 85924 -43625
rect 85890 -43735 85924 -43701
rect 85890 -43785 85924 -43769
rect 85958 -43667 86024 -43659
rect 85958 -43701 85974 -43667
rect 86008 -43701 86024 -43667
rect 85958 -43735 86024 -43701
rect 85958 -43769 85974 -43735
rect 86008 -43769 86024 -43735
rect 85790 -43819 85806 -43805
rect 85672 -43839 85806 -43819
rect 85840 -43819 85856 -43805
rect 85958 -43805 86024 -43769
rect 86058 -43667 86092 -43625
rect 86058 -43735 86092 -43701
rect 86058 -43785 86092 -43769
rect 86126 -43667 86192 -43659
rect 86126 -43701 86142 -43667
rect 86176 -43701 86192 -43667
rect 86126 -43735 86192 -43701
rect 86126 -43769 86142 -43735
rect 86176 -43769 86192 -43735
rect 85958 -43819 85974 -43805
rect 85840 -43839 85974 -43819
rect 86008 -43819 86024 -43805
rect 86126 -43805 86192 -43769
rect 86226 -43667 86260 -43625
rect 86226 -43735 86260 -43701
rect 86226 -43785 86260 -43769
rect 86294 -43667 86360 -43659
rect 86294 -43701 86310 -43667
rect 86344 -43701 86360 -43667
rect 86294 -43735 86360 -43701
rect 86294 -43769 86310 -43735
rect 86344 -43769 86360 -43735
rect 86126 -43819 86142 -43805
rect 86008 -43839 86142 -43819
rect 86176 -43819 86192 -43805
rect 86294 -43805 86360 -43769
rect 86394 -43667 86428 -43625
rect 86394 -43735 86428 -43701
rect 86394 -43785 86428 -43769
rect 86462 -43667 86528 -43659
rect 86462 -43701 86478 -43667
rect 86512 -43701 86528 -43667
rect 86462 -43735 86528 -43701
rect 86462 -43769 86478 -43735
rect 86512 -43769 86528 -43735
rect 86294 -43819 86310 -43805
rect 86176 -43839 86310 -43819
rect 86344 -43819 86360 -43805
rect 86462 -43805 86528 -43769
rect 86562 -43667 86596 -43625
rect 86562 -43735 86596 -43701
rect 86562 -43785 86596 -43769
rect 86630 -43667 86696 -43659
rect 86630 -43701 86646 -43667
rect 86680 -43701 86696 -43667
rect 86630 -43735 86696 -43701
rect 86630 -43769 86646 -43735
rect 86680 -43769 86696 -43735
rect 86462 -43819 86478 -43805
rect 86344 -43839 86478 -43819
rect 86512 -43819 86528 -43805
rect 86630 -43805 86696 -43769
rect 86730 -43667 86764 -43625
rect 86730 -43735 86764 -43701
rect 86730 -43785 86764 -43769
rect 86798 -43667 86864 -43659
rect 86798 -43701 86814 -43667
rect 86848 -43701 86864 -43667
rect 86798 -43735 86864 -43701
rect 86798 -43769 86814 -43735
rect 86848 -43769 86864 -43735
rect 86630 -43819 86646 -43805
rect 86512 -43839 86646 -43819
rect 86680 -43819 86696 -43805
rect 86798 -43800 86864 -43769
rect 86898 -43667 86940 -43625
rect 86932 -43701 86940 -43667
rect 86898 -43735 86940 -43701
rect 86932 -43769 86940 -43735
rect 86898 -43785 86940 -43769
rect 87018 -43667 87060 -43625
rect 87018 -43701 87026 -43667
rect 87018 -43735 87060 -43701
rect 87018 -43769 87026 -43735
rect 86798 -43819 86810 -43800
rect 86680 -43839 86810 -43819
rect 85622 -43853 86810 -43839
rect 85523 -43897 86611 -43889
rect 85523 -43903 85610 -43897
rect 86471 -43903 86611 -43897
rect 85523 -43937 85548 -43903
rect 85582 -43931 85610 -43903
rect 86471 -43931 86561 -43903
rect 85582 -43937 85722 -43931
rect 85756 -43937 85890 -43931
rect 85924 -43937 86059 -43931
rect 86093 -43937 86226 -43931
rect 86260 -43937 86394 -43931
rect 86428 -43937 86561 -43931
rect 86595 -43937 86611 -43903
rect 86798 -43971 86810 -43853
rect 84150 -43991 85392 -43990
rect 84150 -44025 84166 -43991
rect 84200 -44009 84334 -43991
rect 84200 -44025 84216 -44009
rect 84150 -44059 84216 -44025
rect 84318 -44025 84334 -44009
rect 84368 -44009 84502 -43991
rect 84368 -44025 84384 -44009
rect 84150 -44093 84166 -44059
rect 84200 -44093 84216 -44059
rect 84150 -44101 84216 -44093
rect 84250 -44059 84284 -44043
rect 84250 -44135 84284 -44093
rect 84318 -44059 84384 -44025
rect 84486 -44025 84502 -44009
rect 84536 -44009 84670 -43991
rect 84536 -44025 84552 -44009
rect 84318 -44093 84334 -44059
rect 84368 -44093 84384 -44059
rect 84318 -44101 84384 -44093
rect 84418 -44059 84452 -44043
rect 84418 -44135 84452 -44093
rect 84486 -44059 84552 -44025
rect 84654 -44025 84670 -44009
rect 84704 -44009 84838 -43991
rect 84704 -44025 84720 -44009
rect 84486 -44093 84502 -44059
rect 84536 -44093 84552 -44059
rect 84486 -44101 84552 -44093
rect 84586 -44059 84620 -44043
rect 84586 -44135 84620 -44093
rect 84654 -44059 84720 -44025
rect 84822 -44025 84838 -44009
rect 84872 -44009 85006 -43991
rect 84872 -44025 84888 -44009
rect 84654 -44093 84670 -44059
rect 84704 -44093 84720 -44059
rect 84654 -44101 84720 -44093
rect 84754 -44059 84788 -44043
rect 84754 -44135 84788 -44093
rect 84822 -44059 84888 -44025
rect 84990 -44025 85006 -44009
rect 85040 -44009 85174 -43991
rect 85040 -44025 85056 -44009
rect 84822 -44093 84838 -44059
rect 84872 -44093 84888 -44059
rect 84822 -44101 84888 -44093
rect 84922 -44059 84956 -44043
rect 84922 -44135 84956 -44093
rect 84990 -44059 85056 -44025
rect 85158 -44025 85174 -44009
rect 85208 -44009 85342 -43991
rect 85208 -44025 85224 -44009
rect 84990 -44093 85006 -44059
rect 85040 -44093 85056 -44059
rect 84990 -44101 85056 -44093
rect 85090 -44059 85124 -44043
rect 85090 -44135 85124 -44093
rect 85158 -44059 85224 -44025
rect 85326 -44025 85342 -44009
rect 85376 -44025 85392 -43991
rect 85158 -44093 85174 -44059
rect 85208 -44093 85224 -44059
rect 85158 -44101 85224 -44093
rect 85258 -44059 85292 -44043
rect 85258 -44135 85292 -44093
rect 85326 -44059 85392 -44025
rect 85326 -44093 85342 -44059
rect 85376 -44093 85392 -44059
rect 85326 -44101 85392 -44093
rect 85426 -43991 85468 -43975
rect 85460 -44025 85468 -43991
rect 85426 -44059 85468 -44025
rect 85460 -44093 85468 -44059
rect 85426 -44135 85468 -44093
rect 85542 -43991 85588 -43975
rect 85542 -44025 85554 -43991
rect 85542 -44059 85588 -44025
rect 85542 -44093 85554 -44059
rect 85542 -44135 85588 -44093
rect 85622 -43990 86810 -43971
rect 86860 -43990 86864 -43800
rect 87018 -43805 87060 -43769
rect 87018 -43839 87026 -43805
rect 87018 -43855 87060 -43839
rect 87094 -43667 87160 -43659
rect 87094 -43701 87110 -43667
rect 87144 -43701 87160 -43667
rect 87094 -43735 87160 -43701
rect 87094 -43769 87110 -43735
rect 87144 -43769 87160 -43735
rect 87094 -43805 87160 -43769
rect 87194 -43667 87228 -43625
rect 87194 -43735 87228 -43701
rect 87194 -43785 87228 -43769
rect 87262 -43667 87328 -43659
rect 87262 -43701 87278 -43667
rect 87312 -43701 87328 -43667
rect 87262 -43735 87328 -43701
rect 87262 -43769 87278 -43735
rect 87312 -43769 87328 -43735
rect 87094 -43839 87110 -43805
rect 87144 -43819 87160 -43805
rect 87262 -43805 87328 -43769
rect 87362 -43667 87396 -43625
rect 87362 -43735 87396 -43701
rect 87362 -43785 87396 -43769
rect 87430 -43667 87496 -43659
rect 87430 -43701 87446 -43667
rect 87480 -43701 87496 -43667
rect 87430 -43735 87496 -43701
rect 87430 -43769 87446 -43735
rect 87480 -43769 87496 -43735
rect 87262 -43819 87278 -43805
rect 87144 -43839 87278 -43819
rect 87312 -43819 87328 -43805
rect 87430 -43805 87496 -43769
rect 87530 -43667 87564 -43625
rect 87530 -43735 87564 -43701
rect 87530 -43785 87564 -43769
rect 87598 -43667 87664 -43659
rect 87598 -43701 87614 -43667
rect 87648 -43701 87664 -43667
rect 87598 -43735 87664 -43701
rect 87598 -43769 87614 -43735
rect 87648 -43769 87664 -43735
rect 87430 -43819 87446 -43805
rect 87312 -43839 87446 -43819
rect 87480 -43819 87496 -43805
rect 87598 -43805 87664 -43769
rect 87698 -43667 87732 -43625
rect 87698 -43735 87732 -43701
rect 87698 -43785 87732 -43769
rect 87766 -43667 87832 -43659
rect 87766 -43701 87782 -43667
rect 87816 -43701 87832 -43667
rect 87766 -43735 87832 -43701
rect 87766 -43769 87782 -43735
rect 87816 -43769 87832 -43735
rect 87598 -43819 87614 -43805
rect 87480 -43839 87614 -43819
rect 87648 -43819 87664 -43805
rect 87766 -43805 87832 -43769
rect 87866 -43667 87900 -43625
rect 87866 -43735 87900 -43701
rect 87866 -43785 87900 -43769
rect 87934 -43667 88000 -43659
rect 87934 -43701 87950 -43667
rect 87984 -43701 88000 -43667
rect 87934 -43735 88000 -43701
rect 87934 -43769 87950 -43735
rect 87984 -43769 88000 -43735
rect 87766 -43819 87782 -43805
rect 87648 -43839 87782 -43819
rect 87816 -43819 87832 -43805
rect 87934 -43805 88000 -43769
rect 88034 -43667 88068 -43625
rect 88034 -43735 88068 -43701
rect 88034 -43785 88068 -43769
rect 88102 -43667 88168 -43659
rect 88102 -43701 88118 -43667
rect 88152 -43701 88168 -43667
rect 88102 -43735 88168 -43701
rect 88102 -43769 88118 -43735
rect 88152 -43769 88168 -43735
rect 87934 -43819 87950 -43805
rect 87816 -43839 87950 -43819
rect 87984 -43819 88000 -43805
rect 88102 -43805 88168 -43769
rect 88202 -43667 88236 -43625
rect 88202 -43735 88236 -43701
rect 88202 -43785 88236 -43769
rect 88270 -43667 88336 -43659
rect 88270 -43701 88286 -43667
rect 88320 -43701 88336 -43667
rect 88270 -43735 88336 -43701
rect 88270 -43769 88286 -43735
rect 88320 -43769 88336 -43735
rect 88102 -43819 88118 -43805
rect 87984 -43839 88118 -43819
rect 88152 -43819 88168 -43805
rect 88270 -43805 88336 -43769
rect 88370 -43667 88412 -43625
rect 88404 -43701 88412 -43667
rect 88370 -43735 88412 -43701
rect 88404 -43769 88412 -43735
rect 88370 -43785 88412 -43769
rect 88490 -43667 88532 -43625
rect 88490 -43701 88498 -43667
rect 88490 -43735 88532 -43701
rect 88490 -43769 88498 -43735
rect 88270 -43810 88286 -43805
rect 88320 -43810 88336 -43805
rect 88270 -43819 88280 -43810
rect 88152 -43839 88280 -43819
rect 87094 -43853 88280 -43839
rect 86995 -43896 88083 -43889
rect 86995 -43903 87044 -43896
rect 87905 -43903 88083 -43896
rect 86995 -43937 87020 -43903
rect 87905 -43930 88033 -43903
rect 87054 -43937 87194 -43930
rect 87228 -43937 87362 -43930
rect 87396 -43937 87531 -43930
rect 87565 -43937 87698 -43930
rect 87732 -43937 87866 -43930
rect 87900 -43937 88033 -43930
rect 88067 -43937 88083 -43903
rect 88270 -43971 88280 -43853
rect 85622 -43991 86864 -43990
rect 85622 -44025 85638 -43991
rect 85672 -44009 85806 -43991
rect 85672 -44025 85688 -44009
rect 85622 -44059 85688 -44025
rect 85790 -44025 85806 -44009
rect 85840 -44009 85974 -43991
rect 85840 -44025 85856 -44009
rect 85622 -44093 85638 -44059
rect 85672 -44093 85688 -44059
rect 85622 -44101 85688 -44093
rect 85722 -44059 85756 -44043
rect 85722 -44135 85756 -44093
rect 85790 -44059 85856 -44025
rect 85958 -44025 85974 -44009
rect 86008 -44009 86142 -43991
rect 86008 -44025 86024 -44009
rect 85790 -44093 85806 -44059
rect 85840 -44093 85856 -44059
rect 85790 -44101 85856 -44093
rect 85890 -44059 85924 -44043
rect 85890 -44135 85924 -44093
rect 85958 -44059 86024 -44025
rect 86126 -44025 86142 -44009
rect 86176 -44009 86310 -43991
rect 86176 -44025 86192 -44009
rect 85958 -44093 85974 -44059
rect 86008 -44093 86024 -44059
rect 85958 -44101 86024 -44093
rect 86058 -44059 86092 -44043
rect 86058 -44135 86092 -44093
rect 86126 -44059 86192 -44025
rect 86294 -44025 86310 -44009
rect 86344 -44009 86478 -43991
rect 86344 -44025 86360 -44009
rect 86126 -44093 86142 -44059
rect 86176 -44093 86192 -44059
rect 86126 -44101 86192 -44093
rect 86226 -44059 86260 -44043
rect 86226 -44135 86260 -44093
rect 86294 -44059 86360 -44025
rect 86462 -44025 86478 -44009
rect 86512 -44009 86646 -43991
rect 86512 -44025 86528 -44009
rect 86294 -44093 86310 -44059
rect 86344 -44093 86360 -44059
rect 86294 -44101 86360 -44093
rect 86394 -44059 86428 -44043
rect 86394 -44135 86428 -44093
rect 86462 -44059 86528 -44025
rect 86630 -44025 86646 -44009
rect 86680 -44009 86814 -43991
rect 86680 -44025 86696 -44009
rect 86462 -44093 86478 -44059
rect 86512 -44093 86528 -44059
rect 86462 -44101 86528 -44093
rect 86562 -44059 86596 -44043
rect 86562 -44135 86596 -44093
rect 86630 -44059 86696 -44025
rect 86798 -44025 86814 -44009
rect 86848 -44025 86864 -43991
rect 86630 -44093 86646 -44059
rect 86680 -44093 86696 -44059
rect 86630 -44101 86696 -44093
rect 86730 -44059 86764 -44043
rect 86730 -44135 86764 -44093
rect 86798 -44059 86864 -44025
rect 86798 -44093 86814 -44059
rect 86848 -44093 86864 -44059
rect 86798 -44101 86864 -44093
rect 86898 -43991 86940 -43975
rect 86932 -44025 86940 -43991
rect 86898 -44059 86940 -44025
rect 86932 -44093 86940 -44059
rect 86898 -44135 86940 -44093
rect 87014 -43991 87060 -43975
rect 87014 -44025 87026 -43991
rect 87014 -44059 87060 -44025
rect 87014 -44093 87026 -44059
rect 87014 -44135 87060 -44093
rect 87094 -43990 88280 -43971
rect 88330 -43990 88336 -43810
rect 88490 -43805 88532 -43769
rect 88490 -43839 88498 -43805
rect 88490 -43855 88532 -43839
rect 88566 -43667 88632 -43659
rect 88566 -43701 88582 -43667
rect 88616 -43701 88632 -43667
rect 88566 -43735 88632 -43701
rect 88566 -43769 88582 -43735
rect 88616 -43769 88632 -43735
rect 88566 -43805 88632 -43769
rect 88666 -43667 88700 -43625
rect 88666 -43735 88700 -43701
rect 88666 -43785 88700 -43769
rect 88734 -43667 88800 -43659
rect 88734 -43701 88750 -43667
rect 88784 -43701 88800 -43667
rect 88734 -43735 88800 -43701
rect 88734 -43769 88750 -43735
rect 88784 -43769 88800 -43735
rect 88566 -43839 88582 -43805
rect 88616 -43819 88632 -43805
rect 88734 -43805 88800 -43769
rect 88834 -43667 88868 -43625
rect 88834 -43735 88868 -43701
rect 88834 -43785 88868 -43769
rect 88902 -43667 88968 -43659
rect 88902 -43701 88918 -43667
rect 88952 -43701 88968 -43667
rect 88902 -43735 88968 -43701
rect 88902 -43769 88918 -43735
rect 88952 -43769 88968 -43735
rect 88734 -43819 88750 -43805
rect 88616 -43839 88750 -43819
rect 88784 -43819 88800 -43805
rect 88902 -43805 88968 -43769
rect 89002 -43667 89036 -43625
rect 89002 -43735 89036 -43701
rect 89002 -43785 89036 -43769
rect 89070 -43667 89136 -43659
rect 89070 -43701 89086 -43667
rect 89120 -43701 89136 -43667
rect 89070 -43735 89136 -43701
rect 89070 -43769 89086 -43735
rect 89120 -43769 89136 -43735
rect 88902 -43819 88918 -43805
rect 88784 -43839 88918 -43819
rect 88952 -43819 88968 -43805
rect 89070 -43805 89136 -43769
rect 89170 -43667 89204 -43625
rect 89170 -43735 89204 -43701
rect 89170 -43785 89204 -43769
rect 89238 -43667 89304 -43659
rect 89238 -43701 89254 -43667
rect 89288 -43701 89304 -43667
rect 89238 -43735 89304 -43701
rect 89238 -43769 89254 -43735
rect 89288 -43769 89304 -43735
rect 89070 -43819 89086 -43805
rect 88952 -43839 89086 -43819
rect 89120 -43819 89136 -43805
rect 89238 -43805 89304 -43769
rect 89338 -43667 89372 -43625
rect 89338 -43735 89372 -43701
rect 89338 -43785 89372 -43769
rect 89406 -43667 89472 -43659
rect 89406 -43701 89422 -43667
rect 89456 -43701 89472 -43667
rect 89406 -43735 89472 -43701
rect 89406 -43769 89422 -43735
rect 89456 -43769 89472 -43735
rect 89238 -43819 89254 -43805
rect 89120 -43839 89254 -43819
rect 89288 -43819 89304 -43805
rect 89406 -43805 89472 -43769
rect 89506 -43667 89540 -43625
rect 89506 -43735 89540 -43701
rect 89506 -43785 89540 -43769
rect 89574 -43667 89640 -43659
rect 89574 -43701 89590 -43667
rect 89624 -43701 89640 -43667
rect 89574 -43735 89640 -43701
rect 89574 -43769 89590 -43735
rect 89624 -43769 89640 -43735
rect 89406 -43819 89422 -43805
rect 89288 -43839 89422 -43819
rect 89456 -43819 89472 -43805
rect 89574 -43805 89640 -43769
rect 89674 -43667 89708 -43625
rect 89674 -43735 89708 -43701
rect 89674 -43785 89708 -43769
rect 89742 -43667 89808 -43659
rect 89742 -43701 89758 -43667
rect 89792 -43701 89808 -43667
rect 89742 -43735 89808 -43701
rect 89742 -43769 89758 -43735
rect 89792 -43769 89808 -43735
rect 89574 -43819 89590 -43805
rect 89456 -43839 89590 -43819
rect 89624 -43819 89640 -43805
rect 89742 -43805 89808 -43769
rect 89842 -43667 89884 -43625
rect 89876 -43701 89884 -43667
rect 89842 -43735 89884 -43701
rect 89876 -43769 89884 -43735
rect 89842 -43785 89884 -43769
rect 89962 -43667 90004 -43625
rect 89962 -43701 89970 -43667
rect 89962 -43735 90004 -43701
rect 89962 -43769 89970 -43735
rect 89742 -43810 89758 -43805
rect 89792 -43810 89808 -43805
rect 89742 -43819 89750 -43810
rect 89624 -43839 89750 -43819
rect 88566 -43853 89750 -43839
rect 88467 -43896 89555 -43889
rect 88467 -43903 88523 -43896
rect 89384 -43903 89555 -43896
rect 88467 -43937 88492 -43903
rect 89384 -43930 89505 -43903
rect 88526 -43937 88666 -43930
rect 88700 -43937 88834 -43930
rect 88868 -43937 89003 -43930
rect 89037 -43937 89170 -43930
rect 89204 -43937 89338 -43930
rect 89372 -43937 89505 -43930
rect 89539 -43937 89555 -43903
rect 89742 -43971 89750 -43853
rect 87094 -43991 88336 -43990
rect 87094 -44025 87110 -43991
rect 87144 -44009 87278 -43991
rect 87144 -44025 87160 -44009
rect 87094 -44059 87160 -44025
rect 87262 -44025 87278 -44009
rect 87312 -44009 87446 -43991
rect 87312 -44025 87328 -44009
rect 87094 -44093 87110 -44059
rect 87144 -44093 87160 -44059
rect 87094 -44101 87160 -44093
rect 87194 -44059 87228 -44043
rect 87194 -44135 87228 -44093
rect 87262 -44059 87328 -44025
rect 87430 -44025 87446 -44009
rect 87480 -44009 87614 -43991
rect 87480 -44025 87496 -44009
rect 87262 -44093 87278 -44059
rect 87312 -44093 87328 -44059
rect 87262 -44101 87328 -44093
rect 87362 -44059 87396 -44043
rect 87362 -44135 87396 -44093
rect 87430 -44059 87496 -44025
rect 87598 -44025 87614 -44009
rect 87648 -44009 87782 -43991
rect 87648 -44025 87664 -44009
rect 87430 -44093 87446 -44059
rect 87480 -44093 87496 -44059
rect 87430 -44101 87496 -44093
rect 87530 -44059 87564 -44043
rect 87530 -44135 87564 -44093
rect 87598 -44059 87664 -44025
rect 87766 -44025 87782 -44009
rect 87816 -44009 87950 -43991
rect 87816 -44025 87832 -44009
rect 87598 -44093 87614 -44059
rect 87648 -44093 87664 -44059
rect 87598 -44101 87664 -44093
rect 87698 -44059 87732 -44043
rect 87698 -44135 87732 -44093
rect 87766 -44059 87832 -44025
rect 87934 -44025 87950 -44009
rect 87984 -44009 88118 -43991
rect 87984 -44025 88000 -44009
rect 87766 -44093 87782 -44059
rect 87816 -44093 87832 -44059
rect 87766 -44101 87832 -44093
rect 87866 -44059 87900 -44043
rect 87866 -44135 87900 -44093
rect 87934 -44059 88000 -44025
rect 88102 -44025 88118 -44009
rect 88152 -44009 88286 -43991
rect 88152 -44025 88168 -44009
rect 87934 -44093 87950 -44059
rect 87984 -44093 88000 -44059
rect 87934 -44101 88000 -44093
rect 88034 -44059 88068 -44043
rect 88034 -44135 88068 -44093
rect 88102 -44059 88168 -44025
rect 88270 -44025 88286 -44009
rect 88320 -44025 88336 -43991
rect 88102 -44093 88118 -44059
rect 88152 -44093 88168 -44059
rect 88102 -44101 88168 -44093
rect 88202 -44059 88236 -44043
rect 88202 -44135 88236 -44093
rect 88270 -44059 88336 -44025
rect 88270 -44093 88286 -44059
rect 88320 -44093 88336 -44059
rect 88270 -44101 88336 -44093
rect 88370 -43991 88412 -43975
rect 88404 -44025 88412 -43991
rect 88370 -44059 88412 -44025
rect 88404 -44093 88412 -44059
rect 88370 -44135 88412 -44093
rect 88486 -43991 88532 -43975
rect 88486 -44025 88498 -43991
rect 88486 -44059 88532 -44025
rect 88486 -44093 88498 -44059
rect 88486 -44135 88532 -44093
rect 88566 -43991 89750 -43971
rect 88566 -44025 88582 -43991
rect 88616 -44009 88750 -43991
rect 88616 -44025 88632 -44009
rect 88566 -44059 88632 -44025
rect 88734 -44025 88750 -44009
rect 88784 -44009 88918 -43991
rect 88784 -44025 88800 -44009
rect 88566 -44093 88582 -44059
rect 88616 -44093 88632 -44059
rect 88566 -44101 88632 -44093
rect 88666 -44059 88700 -44043
rect 88666 -44135 88700 -44093
rect 88734 -44059 88800 -44025
rect 88902 -44025 88918 -44009
rect 88952 -44009 89086 -43991
rect 88952 -44025 88968 -44009
rect 88734 -44093 88750 -44059
rect 88784 -44093 88800 -44059
rect 88734 -44101 88800 -44093
rect 88834 -44059 88868 -44043
rect 88834 -44135 88868 -44093
rect 88902 -44059 88968 -44025
rect 89070 -44025 89086 -44009
rect 89120 -44009 89254 -43991
rect 89120 -44025 89136 -44009
rect 88902 -44093 88918 -44059
rect 88952 -44093 88968 -44059
rect 88902 -44101 88968 -44093
rect 89002 -44059 89036 -44043
rect 89002 -44135 89036 -44093
rect 89070 -44059 89136 -44025
rect 89238 -44025 89254 -44009
rect 89288 -44009 89422 -43991
rect 89288 -44025 89304 -44009
rect 89070 -44093 89086 -44059
rect 89120 -44093 89136 -44059
rect 89070 -44101 89136 -44093
rect 89170 -44059 89204 -44043
rect 89170 -44135 89204 -44093
rect 89238 -44059 89304 -44025
rect 89406 -44025 89422 -44009
rect 89456 -44009 89590 -43991
rect 89456 -44025 89472 -44009
rect 89238 -44093 89254 -44059
rect 89288 -44093 89304 -44059
rect 89238 -44101 89304 -44093
rect 89338 -44059 89372 -44043
rect 89338 -44135 89372 -44093
rect 89406 -44059 89472 -44025
rect 89574 -44025 89590 -44009
rect 89624 -44000 89750 -43991
rect 89800 -44000 89808 -43810
rect 89962 -43805 90004 -43769
rect 89962 -43839 89970 -43805
rect 89962 -43855 90004 -43839
rect 90038 -43667 90104 -43659
rect 90038 -43701 90054 -43667
rect 90088 -43701 90104 -43667
rect 90038 -43735 90104 -43701
rect 90038 -43769 90054 -43735
rect 90088 -43769 90104 -43735
rect 90038 -43805 90104 -43769
rect 90138 -43667 90172 -43625
rect 90138 -43735 90172 -43701
rect 90138 -43785 90172 -43769
rect 90206 -43667 90272 -43659
rect 90206 -43701 90222 -43667
rect 90256 -43701 90272 -43667
rect 90206 -43735 90272 -43701
rect 90206 -43769 90222 -43735
rect 90256 -43769 90272 -43735
rect 90038 -43839 90054 -43805
rect 90088 -43819 90104 -43805
rect 90206 -43805 90272 -43769
rect 90306 -43667 90340 -43625
rect 90306 -43735 90340 -43701
rect 90306 -43785 90340 -43769
rect 90374 -43667 90440 -43659
rect 90374 -43701 90390 -43667
rect 90424 -43701 90440 -43667
rect 90374 -43735 90440 -43701
rect 90374 -43769 90390 -43735
rect 90424 -43769 90440 -43735
rect 90206 -43819 90222 -43805
rect 90088 -43839 90222 -43819
rect 90256 -43819 90272 -43805
rect 90374 -43805 90440 -43769
rect 90474 -43667 90508 -43625
rect 90474 -43735 90508 -43701
rect 90474 -43785 90508 -43769
rect 90542 -43667 90608 -43659
rect 90542 -43701 90558 -43667
rect 90592 -43701 90608 -43667
rect 90542 -43735 90608 -43701
rect 90542 -43769 90558 -43735
rect 90592 -43769 90608 -43735
rect 90374 -43819 90390 -43805
rect 90256 -43839 90390 -43819
rect 90424 -43819 90440 -43805
rect 90542 -43805 90608 -43769
rect 90642 -43667 90676 -43625
rect 90642 -43735 90676 -43701
rect 90642 -43785 90676 -43769
rect 90710 -43667 90776 -43659
rect 90710 -43701 90726 -43667
rect 90760 -43701 90776 -43667
rect 90710 -43735 90776 -43701
rect 90710 -43769 90726 -43735
rect 90760 -43769 90776 -43735
rect 90542 -43819 90558 -43805
rect 90424 -43839 90558 -43819
rect 90592 -43819 90608 -43805
rect 90710 -43805 90776 -43769
rect 90810 -43667 90844 -43625
rect 90810 -43735 90844 -43701
rect 90810 -43785 90844 -43769
rect 90878 -43667 90944 -43659
rect 90878 -43701 90894 -43667
rect 90928 -43701 90944 -43667
rect 90878 -43735 90944 -43701
rect 90878 -43769 90894 -43735
rect 90928 -43769 90944 -43735
rect 90710 -43819 90726 -43805
rect 90592 -43839 90726 -43819
rect 90760 -43819 90776 -43805
rect 90878 -43805 90944 -43769
rect 90978 -43667 91012 -43625
rect 90978 -43735 91012 -43701
rect 90978 -43785 91012 -43769
rect 91046 -43667 91112 -43659
rect 91046 -43701 91062 -43667
rect 91096 -43701 91112 -43667
rect 91046 -43735 91112 -43701
rect 91046 -43769 91062 -43735
rect 91096 -43769 91112 -43735
rect 90878 -43819 90894 -43805
rect 90760 -43839 90894 -43819
rect 90928 -43819 90944 -43805
rect 91046 -43805 91112 -43769
rect 91146 -43667 91180 -43625
rect 91146 -43735 91180 -43701
rect 91146 -43785 91180 -43769
rect 91214 -43667 91280 -43659
rect 91214 -43701 91230 -43667
rect 91264 -43701 91280 -43667
rect 91214 -43735 91280 -43701
rect 91214 -43769 91230 -43735
rect 91264 -43769 91280 -43735
rect 91046 -43819 91062 -43805
rect 90928 -43839 91062 -43819
rect 91096 -43819 91112 -43805
rect 91214 -43805 91280 -43769
rect 91314 -43667 91356 -43625
rect 91348 -43701 91356 -43667
rect 91314 -43735 91356 -43701
rect 91348 -43769 91356 -43735
rect 91314 -43785 91356 -43769
rect 91214 -43810 91230 -43805
rect 91264 -43810 91280 -43805
rect 91214 -43819 91220 -43810
rect 91096 -43839 91220 -43819
rect 90038 -43853 91220 -43839
rect 89939 -43897 91027 -43889
rect 89939 -43899 89980 -43897
rect 90747 -43899 91027 -43897
rect 89939 -43903 89978 -43899
rect 90748 -43903 91027 -43899
rect 89939 -43937 89964 -43903
rect 90748 -43933 90810 -43903
rect 89998 -43937 90138 -43933
rect 90172 -43937 90306 -43933
rect 90340 -43937 90475 -43933
rect 90509 -43937 90642 -43933
rect 90676 -43937 90810 -43933
rect 90844 -43937 90977 -43903
rect 91011 -43937 91027 -43903
rect 91214 -43971 91220 -43853
rect 89624 -44009 89758 -44000
rect 89624 -44025 89640 -44009
rect 89406 -44093 89422 -44059
rect 89456 -44093 89472 -44059
rect 89406 -44101 89472 -44093
rect 89506 -44059 89540 -44043
rect 89506 -44135 89540 -44093
rect 89574 -44059 89640 -44025
rect 89742 -44025 89758 -44009
rect 89792 -44025 89808 -44000
rect 89574 -44093 89590 -44059
rect 89624 -44093 89640 -44059
rect 89574 -44101 89640 -44093
rect 89674 -44059 89708 -44043
rect 89674 -44135 89708 -44093
rect 89742 -44059 89808 -44025
rect 89742 -44093 89758 -44059
rect 89792 -44093 89808 -44059
rect 89742 -44101 89808 -44093
rect 89842 -43991 89884 -43975
rect 89876 -44025 89884 -43991
rect 89842 -44059 89884 -44025
rect 89876 -44093 89884 -44059
rect 89842 -44135 89884 -44093
rect 89958 -43991 90004 -43975
rect 89958 -44025 89970 -43991
rect 89958 -44059 90004 -44025
rect 89958 -44093 89970 -44059
rect 89958 -44135 90004 -44093
rect 90038 -43991 91220 -43971
rect 90038 -44025 90054 -43991
rect 90088 -44009 90222 -43991
rect 90088 -44025 90104 -44009
rect 90038 -44059 90104 -44025
rect 90206 -44025 90222 -44009
rect 90256 -44009 90390 -43991
rect 90256 -44025 90272 -44009
rect 90038 -44093 90054 -44059
rect 90088 -44093 90104 -44059
rect 90038 -44101 90104 -44093
rect 90138 -44059 90172 -44043
rect 90138 -44135 90172 -44093
rect 90206 -44059 90272 -44025
rect 90374 -44025 90390 -44009
rect 90424 -44009 90558 -43991
rect 90424 -44025 90440 -44009
rect 90206 -44093 90222 -44059
rect 90256 -44093 90272 -44059
rect 90206 -44101 90272 -44093
rect 90306 -44059 90340 -44043
rect 90306 -44135 90340 -44093
rect 90374 -44059 90440 -44025
rect 90542 -44025 90558 -44009
rect 90592 -44009 90726 -43991
rect 90592 -44025 90608 -44009
rect 90374 -44093 90390 -44059
rect 90424 -44093 90440 -44059
rect 90374 -44101 90440 -44093
rect 90474 -44059 90508 -44043
rect 90474 -44135 90508 -44093
rect 90542 -44059 90608 -44025
rect 90710 -44025 90726 -44009
rect 90760 -44009 90894 -43991
rect 90760 -44025 90776 -44009
rect 90542 -44093 90558 -44059
rect 90592 -44093 90608 -44059
rect 90542 -44101 90608 -44093
rect 90642 -44059 90676 -44043
rect 90642 -44135 90676 -44093
rect 90710 -44059 90776 -44025
rect 90878 -44025 90894 -44009
rect 90928 -44009 91062 -43991
rect 90928 -44025 90944 -44009
rect 90710 -44093 90726 -44059
rect 90760 -44093 90776 -44059
rect 90710 -44101 90776 -44093
rect 90810 -44059 90844 -44043
rect 90810 -44135 90844 -44093
rect 90878 -44059 90944 -44025
rect 91046 -44025 91062 -44009
rect 91096 -44000 91220 -43991
rect 91270 -44000 91280 -43810
rect 91096 -44009 91230 -44000
rect 91096 -44025 91112 -44009
rect 90878 -44093 90894 -44059
rect 90928 -44093 90944 -44059
rect 90878 -44101 90944 -44093
rect 90978 -44059 91012 -44043
rect 90978 -44135 91012 -44093
rect 91046 -44059 91112 -44025
rect 91214 -44025 91230 -44009
rect 91264 -44025 91280 -44000
rect 91046 -44093 91062 -44059
rect 91096 -44093 91112 -44059
rect 91046 -44101 91112 -44093
rect 91146 -44059 91180 -44043
rect 91146 -44135 91180 -44093
rect 91214 -44059 91280 -44025
rect 91214 -44093 91230 -44059
rect 91264 -44093 91280 -44059
rect 91214 -44101 91280 -44093
rect 91314 -43991 91356 -43975
rect 91348 -44025 91356 -43991
rect 91314 -44059 91356 -44025
rect 91348 -44093 91356 -44059
rect 91314 -44135 91356 -44093
rect 78153 -44157 78180 -44140
rect 78153 -44225 78180 -44191
rect 77595 -44359 77609 -44325
rect 77595 -44421 77643 -44359
rect 77677 -44275 78115 -44241
rect 77677 -44457 77711 -44275
rect 78052 -44309 78115 -44275
rect 77612 -44473 77711 -44457
rect 77612 -44507 77613 -44473
rect 77647 -44507 77711 -44473
rect 77755 -44325 77825 -44309
rect 77789 -44359 77825 -44325
rect 77755 -44440 77825 -44359
rect 77755 -44480 77770 -44440
rect 77810 -44480 77825 -44440
rect 77755 -44502 77825 -44480
rect 77861 -44320 77921 -44309
rect 77861 -44325 77870 -44320
rect 77861 -44360 77870 -44359
rect 77910 -44360 77921 -44320
rect 77861 -44410 77921 -44360
rect 77861 -44470 77870 -44410
rect 77910 -44470 77921 -44410
rect 77861 -44503 77921 -44470
rect 77957 -44325 78013 -44309
rect 77991 -44359 78013 -44325
rect 78052 -44325 78118 -44309
rect 78052 -44359 78068 -44325
rect 78102 -44359 78118 -44325
rect 77957 -44360 78013 -44359
rect 77957 -44460 77970 -44360
rect 78010 -44460 78013 -44360
rect 77957 -44503 78013 -44460
rect 78049 -44413 78103 -44397
rect 78153 -44413 78180 -44259
rect 78049 -44447 78054 -44413
rect 78088 -44447 78103 -44413
rect 78049 -44481 78103 -44447
rect 77612 -44523 77711 -44507
rect 78049 -44515 78054 -44481
rect 78088 -44515 78103 -44481
rect 78137 -44447 78153 -44413
rect 78137 -44460 78180 -44447
rect 78290 -44460 78310 -44140
rect 82838 -44169 82867 -44135
rect 82901 -44169 82959 -44135
rect 82993 -44169 83051 -44135
rect 83085 -44169 83143 -44135
rect 83177 -44169 83235 -44135
rect 83269 -44169 83327 -44135
rect 83361 -44169 83419 -44135
rect 83453 -44169 83511 -44135
rect 83545 -44169 83603 -44135
rect 83637 -44169 83695 -44135
rect 83729 -44169 83787 -44135
rect 83821 -44169 83879 -44135
rect 83913 -44169 83971 -44135
rect 84005 -44169 84063 -44135
rect 84097 -44169 84155 -44135
rect 84189 -44169 84247 -44135
rect 84281 -44169 84339 -44135
rect 84373 -44169 84431 -44135
rect 84465 -44169 84523 -44135
rect 84557 -44169 84615 -44135
rect 84649 -44169 84707 -44135
rect 84741 -44169 84799 -44135
rect 84833 -44169 84891 -44135
rect 84925 -44169 84983 -44135
rect 85017 -44169 85075 -44135
rect 85109 -44169 85167 -44135
rect 85201 -44169 85259 -44135
rect 85293 -44169 85351 -44135
rect 85385 -44169 85443 -44135
rect 85477 -44169 85535 -44135
rect 85569 -44169 85627 -44135
rect 85661 -44169 85719 -44135
rect 85753 -44169 85811 -44135
rect 85845 -44169 85903 -44135
rect 85937 -44169 85995 -44135
rect 86029 -44169 86087 -44135
rect 86121 -44169 86179 -44135
rect 86213 -44169 86271 -44135
rect 86305 -44169 86363 -44135
rect 86397 -44169 86455 -44135
rect 86489 -44169 86547 -44135
rect 86581 -44169 86639 -44135
rect 86673 -44169 86731 -44135
rect 86765 -44169 86823 -44135
rect 86857 -44169 86915 -44135
rect 86949 -44169 87007 -44135
rect 87041 -44169 87099 -44135
rect 87133 -44169 87191 -44135
rect 87225 -44169 87283 -44135
rect 87317 -44169 87375 -44135
rect 87409 -44169 87467 -44135
rect 87501 -44169 87559 -44135
rect 87593 -44169 87651 -44135
rect 87685 -44169 87743 -44135
rect 87777 -44169 87835 -44135
rect 87869 -44169 87927 -44135
rect 87961 -44169 88019 -44135
rect 88053 -44169 88111 -44135
rect 88145 -44169 88203 -44135
rect 88237 -44169 88295 -44135
rect 88329 -44169 88387 -44135
rect 88421 -44169 88479 -44135
rect 88513 -44169 88571 -44135
rect 88605 -44169 88663 -44135
rect 88697 -44169 88755 -44135
rect 88789 -44169 88847 -44135
rect 88881 -44169 88939 -44135
rect 88973 -44169 89031 -44135
rect 89065 -44169 89123 -44135
rect 89157 -44169 89215 -44135
rect 89249 -44169 89307 -44135
rect 89341 -44169 89399 -44135
rect 89433 -44169 89491 -44135
rect 89525 -44169 89583 -44135
rect 89617 -44169 89675 -44135
rect 89709 -44169 89767 -44135
rect 89801 -44169 89859 -44135
rect 89893 -44169 89951 -44135
rect 89985 -44169 90043 -44135
rect 90077 -44169 90135 -44135
rect 90169 -44169 90227 -44135
rect 90261 -44169 90319 -44135
rect 90353 -44169 90411 -44135
rect 90445 -44169 90503 -44135
rect 90537 -44169 90595 -44135
rect 90629 -44169 90687 -44135
rect 90721 -44169 90779 -44135
rect 90813 -44169 90871 -44135
rect 90905 -44169 90963 -44135
rect 90997 -44169 91055 -44135
rect 91089 -44169 91147 -44135
rect 91181 -44169 91239 -44135
rect 91273 -44169 91331 -44135
rect 91365 -44169 91394 -44135
rect 78137 -44481 78310 -44460
rect 78137 -44515 78153 -44481
rect 78187 -44510 78310 -44481
rect 78187 -44515 78205 -44510
rect 78049 -44557 78103 -44515
rect 77578 -44591 77607 -44557
rect 77641 -44591 77699 -44557
rect 77733 -44591 77791 -44557
rect 77825 -44591 77883 -44557
rect 77917 -44591 77975 -44557
rect 78009 -44591 78067 -44557
rect 78101 -44591 78159 -44557
rect 78193 -44591 78222 -44557
rect 77578 -44665 77607 -44631
rect 77641 -44665 77699 -44631
rect 77733 -44665 77791 -44631
rect 77825 -44665 77883 -44631
rect 77917 -44665 77975 -44631
rect 78009 -44665 78067 -44631
rect 78101 -44665 78159 -44631
rect 78193 -44665 78222 -44631
rect 77612 -44715 77711 -44699
rect 77612 -44749 77613 -44715
rect 77647 -44749 77711 -44715
rect 78049 -44707 78103 -44665
rect 53896 -44792 53992 -44758
rect 54966 -44792 55062 -44758
rect 77612 -44765 77711 -44749
rect 53896 -44854 53930 -44792
rect 55028 -44854 55062 -44792
rect 54075 -44906 54091 -44872
rect 54867 -44906 54883 -44872
rect 53998 -44934 54032 -44918
rect 53998 -44988 54032 -44972
rect 54926 -44934 54960 -44918
rect 54926 -44988 54960 -44972
rect 54075 -45034 54091 -45000
rect 54867 -45034 54883 -45000
rect 53896 -45114 53930 -45052
rect 77560 -44801 77640 -44800
rect 77560 -44863 77643 -44801
rect 77560 -44897 77609 -44863
rect 55028 -45114 55062 -45052
rect 77560 -44950 77643 -44897
rect 77560 -45040 77580 -44950
rect 77630 -45040 77643 -44950
rect 77677 -44947 77711 -44765
rect 77755 -44740 77825 -44720
rect 77755 -44780 77770 -44740
rect 77810 -44780 77825 -44740
rect 77755 -44863 77825 -44780
rect 77789 -44897 77825 -44863
rect 77755 -44913 77825 -44897
rect 77861 -44850 77921 -44719
rect 77861 -44863 77870 -44850
rect 77910 -44890 77921 -44850
rect 77895 -44897 77921 -44890
rect 77861 -44913 77921 -44897
rect 77957 -44860 78013 -44719
rect 78049 -44741 78054 -44707
rect 78088 -44741 78103 -44707
rect 78049 -44775 78103 -44741
rect 78049 -44809 78054 -44775
rect 78088 -44809 78103 -44775
rect 78137 -44741 78153 -44707
rect 78187 -44741 78205 -44707
rect 78137 -44775 78205 -44741
rect 78137 -44809 78153 -44775
rect 78187 -44809 78205 -44775
rect 78049 -44825 78103 -44809
rect 77957 -44863 77960 -44860
rect 77957 -44910 77960 -44897
rect 78010 -44910 78013 -44860
rect 77957 -44913 78013 -44910
rect 78052 -44897 78068 -44863
rect 78102 -44897 78118 -44863
rect 78052 -44913 78118 -44897
rect 78052 -44947 78115 -44913
rect 77677 -44981 78115 -44947
rect 78153 -44920 78205 -44809
rect 78153 -44950 78290 -44920
rect 78153 -44963 78190 -44950
rect 77560 -45060 77643 -45040
rect 77595 -45063 77643 -45060
rect 55960 -45108 56040 -45098
rect 53896 -45148 53992 -45114
rect 54966 -45148 55062 -45114
rect 35802 -45390 35836 -45328
rect 53350 -45238 53790 -45204
rect 53350 -45300 53384 -45238
rect 53510 -45340 53526 -45306
rect 53614 -45340 53630 -45306
rect 25780 -45428 35836 -45390
rect 35802 -45490 35836 -45428
rect 53464 -45390 53498 -45374
rect 53464 -46182 53498 -46166
rect 53642 -45390 53676 -45374
rect 53642 -46182 53676 -46166
rect 53756 -45864 53790 -45238
rect 53896 -45210 53930 -45148
rect 55028 -45210 55062 -45148
rect 55710 -45154 56040 -45108
rect 77697 -45091 77747 -44981
rect 54075 -45262 54091 -45228
rect 54867 -45262 54883 -45228
rect 53998 -45290 54032 -45274
rect 53998 -45344 54032 -45328
rect 54926 -45290 54960 -45274
rect 54926 -45344 54960 -45328
rect 54075 -45390 54091 -45356
rect 54867 -45390 54883 -45356
rect 53896 -45470 53930 -45408
rect 55706 -45188 55802 -45154
rect 56050 -45188 56146 -45154
rect 55706 -45250 55740 -45188
rect 55028 -45470 55062 -45408
rect 53896 -45504 53992 -45470
rect 54966 -45504 55062 -45470
rect 55176 -45300 55272 -45266
rect 55430 -45300 55526 -45266
rect 55176 -45362 55210 -45300
rect 55492 -45362 55526 -45300
rect 55318 -45402 55334 -45368
rect 55368 -45402 55384 -45368
rect 55290 -45452 55324 -45436
rect 55290 -45644 55324 -45628
rect 55378 -45452 55412 -45436
rect 55378 -45644 55412 -45628
rect 55176 -45718 55210 -45656
rect 55492 -45718 55526 -45656
rect 54870 -45752 55272 -45718
rect 55430 -45752 55706 -45718
rect 54870 -45758 55706 -45752
rect 54870 -45864 54904 -45758
rect 53756 -45898 53852 -45864
rect 54808 -45898 54904 -45864
rect 53756 -45960 53790 -45898
rect 54870 -45960 54904 -45898
rect 55126 -45908 55142 -45874
rect 55494 -45908 55510 -45874
rect 53926 -46012 53942 -45978
rect 54718 -46012 54734 -45978
rect 53858 -46040 53892 -46024
rect 53858 -46144 53892 -46128
rect 54768 -46040 54802 -46024
rect 54768 -46144 54802 -46128
rect 53926 -46190 53942 -46156
rect 54718 -46190 54734 -46156
rect 53510 -46250 53526 -46216
rect 53614 -46250 53630 -46216
rect 53756 -46270 53790 -46208
rect 55046 -45960 55080 -45944
rect 55046 -46010 55080 -45994
rect 55556 -45960 55590 -45944
rect 55556 -46010 55590 -45994
rect 55126 -46080 55142 -46046
rect 55494 -46080 55510 -46046
rect 54870 -46238 54904 -46208
rect 55700 -46206 55706 -45758
rect 56112 -45250 56146 -45188
rect 77596 -45133 77613 -45099
rect 77647 -45133 77663 -45099
rect 58930 -45167 59026 -45133
rect 59600 -45167 59696 -45133
rect 58930 -45210 58964 -45167
rect 58926 -45220 58966 -45210
rect 55866 -45290 55882 -45256
rect 55970 -45290 55986 -45256
rect 55820 -45340 55854 -45324
rect 55820 -46132 55854 -46116
rect 55998 -45340 56032 -45324
rect 55998 -46132 56032 -46116
rect 55866 -46200 55882 -46166
rect 55970 -46200 55986 -46166
rect 55700 -46238 55740 -46206
rect 57096 -45279 57125 -45245
rect 57159 -45279 57217 -45245
rect 57251 -45279 57309 -45245
rect 57343 -45279 57372 -45245
rect 57129 -45329 57165 -45313
rect 57129 -45363 57131 -45329
rect 57129 -45397 57165 -45363
rect 57129 -45431 57131 -45397
rect 57201 -45329 57267 -45279
rect 57201 -45363 57217 -45329
rect 57251 -45363 57267 -45329
rect 57201 -45397 57267 -45363
rect 57201 -45431 57217 -45397
rect 57251 -45431 57267 -45397
rect 57301 -45329 57355 -45313
rect 57301 -45363 57303 -45329
rect 57337 -45363 57355 -45329
rect 57301 -45410 57355 -45363
rect 57129 -45465 57165 -45431
rect 57301 -45444 57303 -45410
rect 57337 -45444 57355 -45410
rect 57129 -45499 57264 -45465
rect 57301 -45494 57355 -45444
rect 57230 -45528 57264 -45499
rect 57117 -45544 57185 -45535
rect 57117 -45594 57118 -45544
rect 57178 -45594 57185 -45544
rect 57117 -45609 57185 -45594
rect 57230 -45544 57285 -45528
rect 57230 -45578 57251 -45544
rect 57230 -45594 57285 -45578
rect 57319 -45540 57355 -45494
rect 59662 -45229 59696 -45167
rect 77596 -45175 77663 -45133
rect 77697 -45125 77705 -45091
rect 77739 -45125 77747 -45091
rect 77697 -45141 77747 -45125
rect 77791 -45099 77857 -45031
rect 77791 -45133 77807 -45099
rect 77841 -45133 77857 -45099
rect 77791 -45175 77857 -45133
rect 77894 -45091 77944 -44981
rect 78187 -44997 78190 -44963
rect 77894 -45125 77902 -45091
rect 77936 -45125 77944 -45091
rect 77894 -45141 77944 -45125
rect 78037 -45031 78103 -45015
rect 78037 -45065 78053 -45031
rect 78087 -45065 78103 -45031
rect 78037 -45099 78103 -45065
rect 78153 -45031 78190 -44997
rect 78187 -45065 78190 -45031
rect 78153 -45080 78190 -45065
rect 78260 -45080 78290 -44950
rect 78153 -45089 78290 -45080
rect 78037 -45133 78053 -45099
rect 78087 -45133 78103 -45099
rect 78037 -45175 78103 -45133
rect 78137 -45099 78290 -45089
rect 78137 -45133 78153 -45099
rect 78187 -45100 78290 -45099
rect 78187 -45133 78205 -45100
rect 78137 -45141 78205 -45133
rect 77578 -45209 77607 -45175
rect 77641 -45209 77699 -45175
rect 77733 -45209 77791 -45175
rect 77825 -45209 77883 -45175
rect 77917 -45209 77975 -45175
rect 78009 -45209 78067 -45175
rect 78101 -45209 78159 -45175
rect 78193 -45209 78222 -45175
rect 59109 -45281 59125 -45247
rect 59501 -45281 59517 -45247
rect 59560 -45301 59594 -45285
rect 59560 -45351 59594 -45335
rect 59109 -45389 59125 -45355
rect 59501 -45389 59517 -45355
rect 59032 -45409 59066 -45393
rect 59032 -45459 59066 -45443
rect 59109 -45497 59125 -45463
rect 59501 -45497 59517 -45463
rect 77578 -45285 77607 -45251
rect 77641 -45285 77699 -45251
rect 77733 -45285 77791 -45251
rect 77825 -45285 77883 -45251
rect 77917 -45285 77975 -45251
rect 78009 -45285 78067 -45251
rect 78101 -45285 78159 -45251
rect 78193 -45285 78251 -45251
rect 78285 -45285 78343 -45251
rect 78377 -45285 78435 -45251
rect 78469 -45285 78527 -45251
rect 78561 -45285 78619 -45251
rect 78653 -45285 78711 -45251
rect 78745 -45285 78803 -45251
rect 78837 -45285 78895 -45251
rect 78929 -45285 78987 -45251
rect 79021 -45285 79050 -45251
rect 77595 -45396 77716 -45285
rect 77751 -45336 77847 -45319
rect 77785 -45352 77847 -45336
rect 77751 -45387 77770 -45370
rect 77830 -45387 77847 -45352
rect 77881 -45327 77932 -45285
rect 77881 -45361 77885 -45327
rect 77919 -45361 77932 -45327
rect 77881 -45394 77932 -45361
rect 77966 -45341 78021 -45319
rect 77966 -45375 77969 -45341
rect 78003 -45375 78021 -45341
rect 77595 -45416 77718 -45396
rect 77681 -45421 77718 -45416
rect 77966 -45409 78021 -45375
rect 77681 -45436 77747 -45421
rect 58926 -45540 58966 -45520
rect 57319 -45580 57326 -45540
rect 58930 -45576 58964 -45540
rect 57230 -45645 57264 -45594
rect 57131 -45679 57264 -45645
rect 57319 -45654 57355 -45580
rect 57131 -45700 57165 -45679
rect 56316 -45718 56412 -45704
rect 54830 -46248 55830 -46238
rect 54830 -46270 55030 -46248
rect 53756 -46304 53852 -46270
rect 54808 -46304 55030 -46270
rect 53510 -46358 53526 -46324
rect 53614 -46358 53630 -46324
rect 53756 -46366 53790 -46304
rect 54830 -46328 55030 -46304
rect 55110 -46268 55740 -46248
rect 55810 -46268 55830 -46248
rect 56112 -46268 56146 -46206
rect 55110 -46308 55160 -46268
rect 55600 -46308 55740 -46268
rect 56050 -46302 56146 -46268
rect 55110 -46328 55740 -46308
rect 55810 -46328 55830 -46302
rect 54830 -46338 55830 -46328
rect 53464 -46408 53498 -46392
rect 35802 -46988 35836 -46926
rect 25780 -47022 35836 -46988
rect 35802 -47084 35836 -47022
rect 53464 -47200 53498 -47184
rect 53642 -46408 53676 -46392
rect 53642 -47200 53676 -47184
rect 54870 -46366 54904 -46338
rect 53926 -46418 53942 -46384
rect 54718 -46418 54734 -46384
rect 53858 -46446 53892 -46430
rect 53858 -46550 53892 -46534
rect 54768 -46446 54802 -46430
rect 54768 -46550 54802 -46534
rect 53926 -46596 53942 -46562
rect 54718 -46596 54734 -46562
rect 53756 -46676 53790 -46614
rect 55700 -46364 55740 -46338
rect 55126 -46530 55142 -46496
rect 55494 -46530 55510 -46496
rect 54870 -46676 54904 -46614
rect 55046 -46582 55080 -46566
rect 55046 -46632 55080 -46616
rect 55556 -46582 55590 -46566
rect 55556 -46632 55590 -46616
rect 53756 -46710 53852 -46676
rect 54808 -46710 54904 -46676
rect 55126 -46702 55142 -46668
rect 55494 -46702 55510 -46668
rect 53510 -47268 53526 -47234
rect 53614 -47268 53630 -47234
rect 53350 -47336 53384 -47274
rect 53756 -47336 53790 -46710
rect 54870 -46818 54904 -46710
rect 55700 -46818 55706 -46364
rect 54870 -46824 55706 -46818
rect 54870 -46858 55262 -46824
rect 55420 -46858 55706 -46824
rect 55166 -46920 55200 -46858
rect 53350 -47370 53446 -47336
rect 53694 -47370 53790 -47336
rect 53886 -47108 53982 -47074
rect 54956 -47108 55052 -47074
rect 53886 -47170 53920 -47108
rect 55018 -47170 55052 -47108
rect 54065 -47222 54081 -47188
rect 54857 -47222 54873 -47188
rect 53988 -47250 54022 -47234
rect 53988 -47304 54022 -47288
rect 54916 -47250 54950 -47234
rect 54916 -47304 54950 -47288
rect 54065 -47350 54081 -47316
rect 54857 -47350 54873 -47316
rect 53886 -47430 53920 -47368
rect 55482 -46920 55516 -46858
rect 55280 -46948 55314 -46932
rect 55280 -47140 55314 -47124
rect 55368 -46948 55402 -46932
rect 55368 -47140 55402 -47124
rect 55308 -47208 55324 -47174
rect 55358 -47208 55374 -47174
rect 55166 -47276 55200 -47214
rect 55482 -47276 55516 -47214
rect 55166 -47310 55262 -47276
rect 55420 -47310 55516 -47276
rect 55018 -47430 55052 -47368
rect 56112 -46364 56146 -46302
rect 56350 -45738 56412 -45718
rect 56610 -45738 56706 -45704
rect 56672 -45800 56706 -45738
rect 57303 -45683 57355 -45654
rect 57131 -45755 57165 -45734
rect 57201 -45747 57217 -45713
rect 57251 -45747 57267 -45713
rect 57201 -45789 57267 -45747
rect 57337 -45717 57355 -45683
rect 57303 -45755 57355 -45717
rect 58930 -45610 59026 -45576
rect 59214 -45577 59310 -45576
rect 59662 -45577 59696 -45520
rect 59772 -45494 59866 -45460
rect 60426 -45494 60520 -45460
rect 59772 -45550 59806 -45494
rect 59214 -45610 59696 -45577
rect 58930 -45611 59696 -45610
rect 58930 -45672 58964 -45611
rect 59276 -45672 59310 -45611
rect 59087 -45712 59103 -45678
rect 59137 -45712 59153 -45678
rect 56476 -45840 56492 -45806
rect 56530 -45840 56546 -45806
rect 55866 -46404 55882 -46370
rect 55970 -46404 55986 -46370
rect 55820 -46454 55854 -46438
rect 55820 -47246 55854 -47230
rect 55998 -46454 56032 -46438
rect 55998 -47246 56032 -47230
rect 55866 -47314 55882 -47280
rect 55970 -47314 55986 -47280
rect 55706 -47382 55740 -47320
rect 56430 -45899 56464 -45883
rect 56430 -46691 56464 -46675
rect 56558 -45899 56592 -45883
rect 56558 -46691 56592 -46675
rect 56476 -46768 56492 -46734
rect 56530 -46768 56546 -46734
rect 56316 -46836 56350 -46774
rect 57096 -45823 57125 -45789
rect 57159 -45823 57217 -45789
rect 57251 -45823 57309 -45789
rect 57343 -45823 57372 -45789
rect 59044 -45771 59078 -45755
rect 59044 -46163 59078 -46147
rect 59162 -45771 59196 -45755
rect 59162 -46163 59196 -46147
rect 59087 -46240 59103 -46206
rect 59137 -46240 59153 -46206
rect 60486 -45556 60520 -45494
rect 59942 -45608 59958 -45574
rect 60334 -45608 60350 -45574
rect 59874 -45628 59908 -45612
rect 59874 -45678 59908 -45662
rect 60384 -45628 60418 -45612
rect 60384 -45678 60418 -45662
rect 59942 -45716 59958 -45682
rect 60334 -45716 60350 -45682
rect 59772 -45796 59806 -45740
rect 77595 -45466 77647 -45450
rect 77595 -45500 77613 -45466
rect 77681 -45470 77697 -45436
rect 77731 -45470 77747 -45436
rect 77781 -45455 77932 -45435
rect 77781 -45485 77790 -45455
rect 77778 -45489 77790 -45485
rect 77824 -45489 77932 -45455
rect 77966 -45443 77969 -45409
rect 78003 -45443 78021 -45409
rect 78095 -45369 78151 -45285
rect 78285 -45327 78351 -45285
rect 78095 -45403 78109 -45369
rect 78143 -45403 78151 -45369
rect 78095 -45419 78151 -45403
rect 78185 -45369 78245 -45353
rect 78185 -45403 78193 -45369
rect 78227 -45403 78245 -45369
rect 77966 -45459 78021 -45443
rect 77778 -45492 77932 -45489
rect 77775 -45494 77932 -45492
rect 77774 -45497 77953 -45494
rect 77770 -45500 77953 -45497
rect 77595 -45540 77647 -45500
rect 77766 -45502 77953 -45500
rect 77761 -45504 77953 -45502
rect 77747 -45510 77953 -45504
rect 77743 -45516 77953 -45510
rect 77739 -45522 77953 -45516
rect 77733 -45527 77953 -45522
rect 77726 -45534 77953 -45527
rect 77720 -45535 77953 -45534
rect 77720 -45536 77798 -45535
rect 77720 -45538 77793 -45536
rect 77720 -45539 77790 -45538
rect 77720 -45540 77787 -45539
rect 77595 -45541 77787 -45540
rect 77595 -45543 77785 -45541
rect 77595 -45544 77783 -45543
rect 77595 -45546 77781 -45544
rect 77595 -45548 77780 -45546
rect 77595 -45549 77779 -45548
rect 77595 -45552 77777 -45549
rect 77595 -45555 77776 -45552
rect 77595 -45560 77774 -45555
rect 77595 -45574 77773 -45560
rect 77907 -45563 77953 -45535
rect 77595 -45609 77705 -45608
rect 60486 -45796 60520 -45734
rect 77595 -45643 77613 -45609
rect 77647 -45620 77705 -45609
rect 77595 -45670 77620 -45643
rect 77690 -45670 77705 -45620
rect 77595 -45685 77705 -45670
rect 77739 -45719 77773 -45574
rect 77595 -45753 77613 -45719
rect 77647 -45753 77773 -45719
rect 77807 -45590 77823 -45569
rect 77857 -45590 77873 -45569
rect 77807 -45640 77820 -45590
rect 77860 -45640 77873 -45590
rect 77907 -45597 77919 -45563
rect 77907 -45614 77953 -45597
rect 77807 -45654 77873 -45640
rect 77807 -45751 77851 -45654
rect 77987 -45665 78021 -45459
rect 78185 -45463 78245 -45403
rect 78285 -45361 78301 -45327
rect 78335 -45361 78351 -45327
rect 78285 -45395 78351 -45361
rect 78285 -45429 78301 -45395
rect 78335 -45429 78351 -45395
rect 78389 -45320 78481 -45319
rect 78389 -45327 78840 -45320
rect 78389 -45361 78405 -45327
rect 78439 -45329 78840 -45327
rect 78881 -45327 78937 -45285
rect 78439 -45339 78847 -45329
rect 78439 -45361 78755 -45339
rect 78389 -45373 78755 -45361
rect 78789 -45373 78847 -45339
rect 78389 -45380 78847 -45373
rect 78389 -45395 78481 -45380
rect 78516 -45387 78847 -45380
rect 78881 -45361 78894 -45327
rect 78928 -45361 78937 -45327
rect 78389 -45429 78405 -45395
rect 78439 -45429 78481 -45395
rect 78881 -45395 78937 -45361
rect 78060 -45475 78150 -45470
rect 78058 -45490 78150 -45475
rect 78058 -45580 78080 -45490
rect 78130 -45547 78150 -45490
rect 78185 -45497 78373 -45463
rect 78339 -45547 78373 -45497
rect 78130 -45563 78193 -45547
rect 78058 -45597 78112 -45580
rect 78146 -45597 78193 -45563
rect 78237 -45550 78305 -45547
rect 78237 -45590 78250 -45550
rect 78290 -45590 78305 -45550
rect 78237 -45597 78253 -45590
rect 78287 -45597 78305 -45590
rect 78339 -45563 78397 -45547
rect 78339 -45597 78361 -45563
rect 78395 -45597 78397 -45563
rect 78339 -45613 78397 -45597
rect 78339 -45631 78373 -45613
rect 77969 -45670 78021 -45665
rect 78095 -45669 78373 -45631
rect 77969 -45680 78050 -45670
rect 77885 -45703 77935 -45687
rect 77919 -45737 77935 -45703
rect 77885 -45795 77935 -45737
rect 77969 -45693 77990 -45680
rect 78030 -45720 78050 -45680
rect 78003 -45727 78050 -45720
rect 77969 -45760 78050 -45727
rect 78095 -45691 78161 -45669
rect 78095 -45725 78109 -45691
rect 78143 -45725 78161 -45691
rect 78431 -45703 78481 -45429
rect 78516 -45455 78834 -45421
rect 78881 -45429 78894 -45395
rect 78928 -45429 78937 -45395
rect 78881 -45445 78937 -45429
rect 78979 -45320 79033 -45319
rect 78979 -45358 79090 -45320
rect 79013 -45370 79090 -45358
rect 79013 -45392 79020 -45370
rect 78979 -45426 79020 -45392
rect 78516 -45458 78580 -45455
rect 78516 -45492 78533 -45458
rect 78567 -45492 78580 -45458
rect 78800 -45479 78834 -45455
rect 79013 -45460 79020 -45426
rect 78516 -45513 78580 -45492
rect 78620 -45520 78762 -45489
rect 78800 -45513 78945 -45479
rect 78979 -45513 79020 -45460
rect 78516 -45560 78586 -45547
rect 78516 -45640 78530 -45560
rect 78570 -45640 78586 -45560
rect 78620 -45590 78650 -45520
rect 78730 -45590 78762 -45520
rect 78911 -45547 78945 -45513
rect 78620 -45597 78659 -45590
rect 78693 -45597 78762 -45590
rect 78620 -45613 78762 -45597
rect 78796 -45560 78877 -45547
rect 78796 -45600 78820 -45560
rect 78860 -45563 78877 -45560
rect 78869 -45597 78877 -45563
rect 78860 -45600 78877 -45597
rect 78796 -45613 78877 -45600
rect 78911 -45563 78965 -45547
rect 78911 -45597 78931 -45563
rect 78911 -45613 78965 -45597
rect 78516 -45661 78586 -45640
rect 78911 -45647 78945 -45613
rect 78623 -45681 78945 -45647
rect 78999 -45660 79020 -45513
rect 78979 -45677 79020 -45660
rect 78095 -45741 78161 -45725
rect 78285 -45719 78335 -45703
rect 78285 -45753 78301 -45719
rect 77969 -45761 78021 -45760
rect 78285 -45795 78335 -45753
rect 78369 -45719 78481 -45703
rect 78369 -45753 78385 -45719
rect 78419 -45753 78481 -45719
rect 78369 -45761 78481 -45753
rect 78517 -45729 78533 -45695
rect 78567 -45729 78583 -45695
rect 78517 -45795 78583 -45729
rect 78623 -45701 78657 -45681
rect 78797 -45701 78831 -45681
rect 78623 -45751 78657 -45735
rect 78697 -45749 78713 -45715
rect 78747 -45749 78763 -45715
rect 78697 -45795 78763 -45749
rect 79013 -45680 79020 -45677
rect 79070 -45680 79090 -45370
rect 79013 -45711 79090 -45680
rect 78797 -45751 78831 -45735
rect 78865 -45749 78891 -45715
rect 78925 -45749 78941 -45715
rect 78979 -45729 79090 -45711
rect 79000 -45730 79090 -45729
rect 78865 -45795 78941 -45749
rect 59388 -45830 59476 -45796
rect 59656 -45830 59800 -45796
rect 59958 -45830 60520 -45796
rect 77578 -45829 77607 -45795
rect 77641 -45829 77699 -45795
rect 77733 -45829 77791 -45795
rect 77825 -45829 77883 -45795
rect 77917 -45829 77975 -45795
rect 78009 -45829 78067 -45795
rect 78101 -45829 78159 -45795
rect 78193 -45829 78251 -45795
rect 78285 -45829 78343 -45795
rect 78377 -45829 78435 -45795
rect 78469 -45829 78527 -45795
rect 78561 -45829 78619 -45795
rect 78653 -45829 78711 -45795
rect 78745 -45829 78803 -45795
rect 78837 -45829 78895 -45795
rect 78929 -45829 78987 -45795
rect 79021 -45829 79050 -45795
rect 59388 -45890 59422 -45830
rect 59276 -46306 59310 -46246
rect 59530 -45932 59546 -45898
rect 59580 -45932 59596 -45898
rect 59502 -45982 59536 -45966
rect 59502 -46174 59536 -46158
rect 59590 -45982 59624 -45966
rect 59590 -46174 59624 -46158
rect 59530 -46242 59546 -46208
rect 59580 -46242 59596 -46208
rect 58966 -46342 59310 -46306
rect 59388 -46309 59422 -46250
rect 59704 -46309 59738 -45830
rect 60020 -45892 60054 -45830
rect 59846 -45932 59862 -45898
rect 59896 -45932 59912 -45898
rect 59818 -45982 59852 -45966
rect 59818 -46174 59852 -46158
rect 59906 -45982 59940 -45966
rect 59906 -46174 59940 -46158
rect 59846 -46242 59862 -46208
rect 59896 -46242 59912 -46208
rect 61186 -46000 61286 -45990
rect 61186 -46080 61196 -46000
rect 61186 -46090 61286 -46080
rect 60020 -46309 60054 -46248
rect 56672 -46836 56706 -46774
rect 57096 -46799 57125 -46765
rect 57159 -46799 57217 -46765
rect 57251 -46799 57309 -46765
rect 57343 -46799 57372 -46765
rect 56316 -46870 56412 -46836
rect 56610 -46870 56706 -46836
rect 57131 -46854 57165 -46833
rect 57201 -46841 57267 -46799
rect 57201 -46875 57217 -46841
rect 57251 -46875 57267 -46841
rect 57303 -46871 57355 -46833
rect 57131 -46909 57165 -46888
rect 57337 -46905 57355 -46871
rect 59276 -46402 59310 -46342
rect 59387 -46344 60054 -46309
rect 60127 -46154 60161 -46128
rect 60127 -46157 60253 -46154
rect 60161 -46173 60253 -46157
rect 60161 -46191 60203 -46173
rect 60127 -46207 60203 -46191
rect 60237 -46207 60253 -46173
rect 60359 -46160 60409 -46149
rect 60671 -46154 60705 -46128
rect 60359 -46165 60366 -46160
rect 60359 -46200 60366 -46199
rect 60406 -46200 60409 -46160
rect 60127 -46249 60161 -46207
rect 60127 -46341 60161 -46283
rect 60195 -46257 60325 -46241
rect 60195 -46291 60211 -46257
rect 60245 -46291 60325 -46257
rect 60195 -46307 60325 -46291
rect 59387 -46400 59421 -46344
rect 59087 -46442 59103 -46408
rect 59137 -46442 59153 -46408
rect 59044 -46501 59078 -46485
rect 57131 -46943 57264 -46909
rect 57303 -46934 57355 -46905
rect 57117 -46994 57185 -46979
rect 57117 -47044 57118 -46994
rect 57168 -47044 57185 -46994
rect 57117 -47053 57185 -47044
rect 57230 -46994 57264 -46943
rect 57319 -46970 57355 -46934
rect 57230 -47010 57285 -46994
rect 57230 -47044 57251 -47010
rect 57230 -47060 57285 -47044
rect 57319 -47010 57326 -46970
rect 59044 -46893 59078 -46877
rect 59162 -46501 59196 -46485
rect 59162 -46893 59196 -46877
rect 59087 -46970 59103 -46936
rect 59137 -46970 59153 -46936
rect 57230 -47089 57264 -47060
rect 57129 -47123 57264 -47089
rect 57319 -47094 57355 -47010
rect 57129 -47157 57165 -47123
rect 57301 -47144 57355 -47094
rect 58930 -47038 58964 -46976
rect 59529 -46445 59545 -46411
rect 59579 -46445 59595 -46411
rect 59501 -46495 59535 -46479
rect 59501 -46687 59535 -46671
rect 59589 -46495 59623 -46479
rect 59589 -46687 59623 -46671
rect 59529 -46755 59545 -46721
rect 59579 -46755 59595 -46721
rect 59387 -46823 59421 -46770
rect 59703 -46823 59737 -46344
rect 60019 -46405 60053 -46344
rect 59845 -46445 59861 -46411
rect 59895 -46445 59911 -46411
rect 59817 -46495 59851 -46479
rect 59817 -46687 59851 -46671
rect 59905 -46495 59939 -46479
rect 59905 -46687 59939 -46671
rect 59845 -46755 59861 -46721
rect 59895 -46755 59911 -46721
rect 60161 -46375 60203 -46341
rect 60237 -46375 60253 -46341
rect 60127 -46433 60161 -46375
rect 60289 -46409 60325 -46307
rect 60127 -46509 60161 -46467
rect 60195 -46425 60325 -46409
rect 60195 -46459 60211 -46425
rect 60245 -46459 60325 -46425
rect 60195 -46475 60325 -46459
rect 60359 -46250 60409 -46200
rect 60443 -46157 60705 -46154
rect 60443 -46173 60671 -46157
rect 60443 -46207 60459 -46173
rect 60493 -46207 60527 -46173
rect 60561 -46207 60595 -46173
rect 60629 -46191 60671 -46173
rect 60629 -46207 60705 -46191
rect 60359 -46257 60366 -46250
rect 60406 -46290 60409 -46250
rect 60393 -46291 60409 -46290
rect 60359 -46340 60409 -46291
rect 60359 -46341 60366 -46340
rect 60359 -46380 60366 -46375
rect 60406 -46380 60409 -46340
rect 60359 -46420 60409 -46380
rect 60359 -46425 60366 -46420
rect 60359 -46460 60366 -46459
rect 60406 -46460 60409 -46420
rect 60359 -46475 60409 -46460
rect 60443 -46257 60637 -46241
rect 60443 -46291 60459 -46257
rect 60493 -46291 60527 -46257
rect 60561 -46291 60595 -46257
rect 60629 -46291 60637 -46257
rect 60443 -46307 60637 -46291
rect 60671 -46249 60705 -46207
rect 60443 -46409 60477 -46307
rect 60671 -46341 60705 -46283
rect 60511 -46375 60527 -46341
rect 60561 -46375 60595 -46341
rect 60629 -46375 60671 -46341
rect 60443 -46425 60637 -46409
rect 60443 -46459 60459 -46425
rect 60493 -46459 60527 -46425
rect 60561 -46459 60595 -46425
rect 60629 -46459 60637 -46425
rect 60443 -46475 60637 -46459
rect 60671 -46433 60705 -46375
rect 60289 -46509 60325 -46475
rect 60443 -46509 60481 -46475
rect 60671 -46509 60705 -46467
rect 60127 -46525 60204 -46509
rect 60161 -46543 60204 -46525
rect 60238 -46543 60254 -46509
rect 60161 -46559 60254 -46543
rect 60289 -46525 60481 -46509
rect 60289 -46559 60297 -46525
rect 60331 -46559 60369 -46525
rect 60405 -46559 60449 -46525
rect 60579 -46543 60595 -46509
rect 60629 -46525 60705 -46509
rect 60629 -46543 60671 -46525
rect 60579 -46551 60671 -46543
rect 60127 -46588 60161 -46559
rect 60289 -46562 60481 -46559
rect 60671 -46588 60705 -46559
rect 60747 -46154 60781 -46128
rect 60747 -46157 61009 -46154
rect 60781 -46173 61009 -46157
rect 60781 -46191 60823 -46173
rect 60747 -46207 60823 -46191
rect 60857 -46207 60891 -46173
rect 60925 -46207 60959 -46173
rect 60993 -46207 61009 -46173
rect 61043 -46160 61093 -46149
rect 61291 -46154 61325 -46128
rect 61043 -46200 61046 -46160
rect 61086 -46165 61093 -46160
rect 61086 -46200 61093 -46199
rect 60747 -46249 60781 -46207
rect 60747 -46341 60781 -46283
rect 60815 -46257 61009 -46241
rect 60815 -46291 60823 -46257
rect 60857 -46291 60891 -46257
rect 60925 -46291 60959 -46257
rect 60993 -46291 61009 -46257
rect 60815 -46307 61009 -46291
rect 60781 -46375 60823 -46341
rect 60857 -46375 60891 -46341
rect 60925 -46375 60941 -46341
rect 60747 -46433 60781 -46375
rect 60975 -46409 61009 -46307
rect 60747 -46509 60781 -46467
rect 60815 -46425 61009 -46409
rect 60815 -46459 60823 -46425
rect 60857 -46459 60891 -46425
rect 60925 -46459 60959 -46425
rect 60993 -46459 61009 -46425
rect 60815 -46475 61009 -46459
rect 61043 -46250 61093 -46200
rect 61199 -46157 61325 -46154
rect 61199 -46173 61291 -46157
rect 61199 -46207 61215 -46173
rect 61249 -46191 61291 -46173
rect 61249 -46207 61325 -46191
rect 61043 -46290 61046 -46250
rect 61086 -46257 61093 -46250
rect 61043 -46291 61059 -46290
rect 61043 -46340 61093 -46291
rect 61043 -46380 61046 -46340
rect 61086 -46341 61093 -46340
rect 61086 -46380 61093 -46375
rect 61043 -46420 61093 -46380
rect 61043 -46460 61046 -46420
rect 61086 -46425 61093 -46420
rect 61086 -46460 61093 -46459
rect 61043 -46475 61093 -46460
rect 61127 -46257 61257 -46241
rect 61127 -46291 61207 -46257
rect 61241 -46291 61257 -46257
rect 61127 -46307 61257 -46291
rect 61291 -46249 61325 -46207
rect 61127 -46409 61163 -46307
rect 61291 -46341 61325 -46283
rect 61199 -46375 61215 -46341
rect 61249 -46375 61291 -46341
rect 61127 -46425 61257 -46409
rect 61127 -46459 61207 -46425
rect 61241 -46459 61257 -46425
rect 61127 -46475 61257 -46459
rect 61291 -46433 61325 -46375
rect 75506 -46445 75535 -46411
rect 75569 -46445 75627 -46411
rect 75661 -46445 75719 -46411
rect 75753 -46445 75811 -46411
rect 75845 -46445 75903 -46411
rect 75937 -46445 75995 -46411
rect 76029 -46445 76085 -46411
rect 76119 -46445 76177 -46411
rect 76211 -46445 76269 -46411
rect 76303 -46445 76361 -46411
rect 76395 -46445 76453 -46411
rect 76487 -46445 76545 -46411
rect 76579 -46445 76637 -46411
rect 76671 -46445 76729 -46411
rect 76763 -46445 76821 -46411
rect 76855 -46445 76884 -46411
rect 60971 -46509 61009 -46475
rect 61127 -46509 61163 -46475
rect 61291 -46509 61325 -46467
rect 60747 -46525 60823 -46509
rect 60781 -46543 60823 -46525
rect 60857 -46543 60873 -46509
rect 60781 -46551 60873 -46543
rect 60971 -46524 61163 -46509
rect 60971 -46525 61129 -46524
rect 60747 -46588 60781 -46559
rect 60971 -46559 60980 -46525
rect 61015 -46559 61053 -46525
rect 61088 -46558 61129 -46525
rect 61198 -46543 61214 -46509
rect 61248 -46525 61325 -46509
rect 61248 -46543 61291 -46525
rect 61088 -46559 61163 -46558
rect 61198 -46559 61291 -46543
rect 60971 -46562 61163 -46559
rect 61291 -46588 61325 -46559
rect 75570 -46491 75616 -46445
rect 75570 -46525 75582 -46491
rect 75570 -46559 75616 -46525
rect 75570 -46593 75582 -46559
rect 75570 -46609 75616 -46593
rect 75650 -46491 75716 -46479
rect 75650 -46525 75666 -46491
rect 75700 -46525 75716 -46491
rect 75650 -46557 75716 -46525
rect 75650 -46559 75670 -46557
rect 75650 -46593 75666 -46559
rect 75704 -46591 75716 -46557
rect 75700 -46593 75716 -46591
rect 75650 -46605 75716 -46593
rect 60466 -46660 60546 -46640
rect 60466 -46700 60486 -46660
rect 60526 -46700 60546 -46660
rect 60466 -46720 60546 -46700
rect 60606 -46660 60686 -46640
rect 60606 -46700 60626 -46660
rect 60666 -46700 60686 -46660
rect 60606 -46720 60686 -46700
rect 60746 -46660 60826 -46640
rect 60746 -46700 60766 -46660
rect 60806 -46700 60826 -46660
rect 60746 -46720 60826 -46700
rect 60886 -46660 60966 -46640
rect 60886 -46700 60906 -46660
rect 60946 -46700 60966 -46660
rect 75570 -46650 75586 -46643
rect 75570 -46690 75580 -46650
rect 75620 -46690 75636 -46643
rect 75570 -46691 75636 -46690
rect 75670 -46649 75716 -46605
rect 75846 -46491 75892 -46445
rect 75846 -46525 75858 -46491
rect 75846 -46559 75892 -46525
rect 75846 -46593 75858 -46559
rect 75846 -46609 75892 -46593
rect 75926 -46491 75992 -46479
rect 75926 -46525 75942 -46491
rect 75976 -46525 75992 -46491
rect 75926 -46559 75992 -46525
rect 75926 -46594 75942 -46559
rect 75976 -46594 75992 -46559
rect 75926 -46605 75992 -46594
rect 75704 -46683 75716 -46649
rect 60886 -46720 60966 -46700
rect 75670 -46725 75716 -46683
rect 75846 -46677 75862 -46643
rect 75896 -46677 75912 -46643
rect 75846 -46691 75912 -46677
rect 75946 -46649 75992 -46605
rect 76120 -46491 76166 -46445
rect 76120 -46525 76132 -46491
rect 76120 -46559 76166 -46525
rect 76120 -46593 76132 -46559
rect 76120 -46609 76166 -46593
rect 76200 -46491 76266 -46479
rect 76200 -46525 76216 -46491
rect 76250 -46525 76266 -46491
rect 76200 -46559 76266 -46525
rect 76200 -46593 76216 -46559
rect 76251 -46593 76266 -46559
rect 76200 -46605 76266 -46593
rect 75946 -46683 75947 -46649
rect 75981 -46683 75992 -46649
rect 75946 -46725 75992 -46683
rect 76120 -46650 76136 -46643
rect 76120 -46684 76128 -46650
rect 76170 -46677 76186 -46643
rect 76162 -46684 76186 -46677
rect 76120 -46691 76186 -46684
rect 76220 -46650 76266 -46605
rect 76396 -46491 76442 -46445
rect 76396 -46525 76408 -46491
rect 76396 -46559 76442 -46525
rect 76396 -46593 76408 -46559
rect 76396 -46609 76442 -46593
rect 76476 -46491 76542 -46479
rect 76476 -46525 76492 -46491
rect 76526 -46525 76542 -46491
rect 76476 -46559 76542 -46525
rect 76476 -46593 76492 -46559
rect 76526 -46593 76542 -46559
rect 76476 -46605 76542 -46593
rect 76220 -46684 76224 -46650
rect 76258 -46684 76266 -46650
rect 76220 -46725 76266 -46684
rect 76396 -46649 76412 -46643
rect 76396 -46683 76404 -46649
rect 76446 -46677 76462 -46643
rect 76438 -46683 76462 -46677
rect 76396 -46691 76462 -46683
rect 76496 -46649 76542 -46605
rect 76672 -46491 76718 -46445
rect 76672 -46525 76684 -46491
rect 76672 -46559 76718 -46525
rect 76672 -46593 76684 -46559
rect 76672 -46609 76718 -46593
rect 76752 -46491 76818 -46479
rect 76752 -46525 76768 -46491
rect 76802 -46525 76818 -46491
rect 76752 -46559 76818 -46525
rect 76752 -46595 76768 -46559
rect 76802 -46595 76818 -46559
rect 76752 -46605 76818 -46595
rect 76496 -46683 76497 -46649
rect 76531 -46683 76542 -46649
rect 76496 -46725 76542 -46683
rect 76672 -46649 76688 -46643
rect 76672 -46683 76680 -46649
rect 76722 -46677 76738 -46643
rect 76714 -46683 76738 -46677
rect 76672 -46691 76738 -46683
rect 76772 -46650 76818 -46605
rect 76806 -46684 76818 -46650
rect 76772 -46725 76818 -46684
rect 60019 -46823 60053 -46761
rect 59387 -46857 59476 -46823
rect 59646 -46857 59799 -46823
rect 59957 -46826 60053 -46823
rect 75574 -46743 75616 -46727
rect 75574 -46777 75582 -46743
rect 75574 -46811 75616 -46777
rect 59957 -46857 60520 -46826
rect 59772 -46860 60520 -46857
rect 59772 -46920 59806 -46860
rect 59276 -47038 59310 -46976
rect 58930 -47072 59026 -47038
rect 59214 -47040 59310 -47038
rect 59214 -47072 59696 -47040
rect 58930 -47074 59696 -47072
rect 58930 -47110 58964 -47074
rect 57129 -47191 57131 -47157
rect 57129 -47225 57165 -47191
rect 57129 -47259 57131 -47225
rect 57129 -47275 57165 -47259
rect 57201 -47191 57217 -47157
rect 57251 -47191 57267 -47157
rect 57201 -47225 57267 -47191
rect 57201 -47259 57217 -47225
rect 57251 -47259 57267 -47225
rect 57201 -47309 57267 -47259
rect 57301 -47178 57303 -47144
rect 57337 -47178 57355 -47144
rect 57301 -47225 57355 -47178
rect 57301 -47259 57303 -47225
rect 57337 -47259 57355 -47225
rect 57301 -47275 57355 -47259
rect 59662 -47130 59696 -47074
rect 60486 -46922 60520 -46860
rect 59942 -46974 59958 -46940
rect 60334 -46974 60350 -46940
rect 59874 -46994 59908 -46978
rect 59874 -47044 59908 -47028
rect 60384 -46994 60418 -46978
rect 60384 -47044 60418 -47028
rect 59942 -47082 59958 -47048
rect 60334 -47082 60350 -47048
rect 56112 -47382 56146 -47320
rect 57096 -47343 57125 -47309
rect 57159 -47343 57217 -47309
rect 57251 -47343 57309 -47309
rect 57343 -47343 57372 -47309
rect 55706 -47416 55802 -47382
rect 56050 -47416 56146 -47382
rect 53886 -47464 53982 -47430
rect 54956 -47464 55052 -47430
rect 53886 -47526 53920 -47464
rect 55018 -47526 55052 -47464
rect 55720 -47458 56090 -47416
rect 55720 -47468 56020 -47458
rect 54065 -47578 54081 -47544
rect 54857 -47578 54873 -47544
rect 53988 -47606 54022 -47590
rect 53988 -47660 54022 -47644
rect 54916 -47606 54950 -47590
rect 54916 -47660 54950 -47644
rect 54065 -47706 54081 -47672
rect 54857 -47706 54873 -47672
rect 53886 -47786 53920 -47724
rect 56010 -47608 56020 -47468
rect 56080 -47608 56090 -47458
rect 59109 -47188 59125 -47154
rect 59501 -47188 59517 -47154
rect 59560 -47208 59594 -47192
rect 59560 -47258 59594 -47242
rect 59109 -47296 59125 -47262
rect 59501 -47296 59517 -47262
rect 59032 -47316 59066 -47300
rect 59032 -47366 59066 -47350
rect 59109 -47404 59125 -47370
rect 59501 -47404 59517 -47370
rect 56010 -47618 56090 -47608
rect 59772 -47162 59806 -47100
rect 75574 -46845 75582 -46811
rect 75574 -46879 75616 -46845
rect 75574 -46913 75582 -46879
rect 75574 -46955 75616 -46913
rect 75650 -46738 75716 -46725
rect 75650 -46743 75670 -46738
rect 75650 -46777 75666 -46743
rect 75704 -46772 75716 -46738
rect 75700 -46777 75716 -46772
rect 75650 -46811 75716 -46777
rect 75650 -46845 75666 -46811
rect 75700 -46845 75716 -46811
rect 75650 -46879 75716 -46845
rect 75650 -46913 75666 -46879
rect 75700 -46913 75716 -46879
rect 75650 -46921 75716 -46913
rect 75850 -46743 75892 -46727
rect 75850 -46777 75858 -46743
rect 75850 -46811 75892 -46777
rect 75850 -46845 75858 -46811
rect 75850 -46879 75892 -46845
rect 75850 -46913 75858 -46879
rect 75850 -46955 75892 -46913
rect 75926 -46743 75992 -46725
rect 75926 -46777 75942 -46743
rect 75977 -46777 75992 -46743
rect 75926 -46811 75992 -46777
rect 75926 -46845 75942 -46811
rect 75976 -46845 75992 -46811
rect 75926 -46879 75992 -46845
rect 75926 -46913 75942 -46879
rect 75976 -46913 75992 -46879
rect 75926 -46921 75992 -46913
rect 76124 -46743 76166 -46727
rect 76124 -46777 76132 -46743
rect 76124 -46811 76166 -46777
rect 76124 -46845 76132 -46811
rect 76124 -46879 76166 -46845
rect 76124 -46913 76132 -46879
rect 76124 -46955 76166 -46913
rect 76200 -46743 76266 -46725
rect 76200 -46744 76216 -46743
rect 76200 -46778 76215 -46744
rect 76250 -46777 76266 -46743
rect 76249 -46778 76266 -46777
rect 76200 -46811 76266 -46778
rect 76200 -46845 76216 -46811
rect 76250 -46816 76266 -46811
rect 76200 -46850 76218 -46845
rect 76252 -46850 76266 -46816
rect 76200 -46879 76266 -46850
rect 76200 -46913 76216 -46879
rect 76250 -46913 76266 -46879
rect 76200 -46921 76266 -46913
rect 76400 -46743 76442 -46727
rect 76400 -46777 76408 -46743
rect 76400 -46811 76442 -46777
rect 76400 -46845 76408 -46811
rect 76400 -46879 76442 -46845
rect 76400 -46913 76408 -46879
rect 76400 -46955 76442 -46913
rect 76476 -46743 76542 -46725
rect 76476 -46777 76492 -46743
rect 76526 -46777 76542 -46743
rect 76476 -46811 76542 -46777
rect 76476 -46845 76492 -46811
rect 76526 -46845 76542 -46811
rect 76476 -46879 76542 -46845
rect 76476 -46913 76492 -46879
rect 76526 -46913 76542 -46879
rect 76476 -46921 76542 -46913
rect 76676 -46743 76718 -46727
rect 76676 -46777 76684 -46743
rect 76676 -46811 76718 -46777
rect 76676 -46845 76684 -46811
rect 76676 -46879 76718 -46845
rect 76676 -46913 76684 -46879
rect 76676 -46955 76718 -46913
rect 76752 -46743 76818 -46725
rect 76752 -46777 76768 -46743
rect 76802 -46777 76818 -46743
rect 76752 -46811 76818 -46777
rect 76752 -46845 76768 -46811
rect 76802 -46845 76818 -46811
rect 76752 -46879 76818 -46845
rect 76752 -46913 76768 -46879
rect 76802 -46913 76818 -46879
rect 76752 -46921 76818 -46913
rect 75506 -46989 75535 -46955
rect 75569 -46989 75627 -46955
rect 75661 -46989 75719 -46955
rect 75753 -46989 75811 -46955
rect 75845 -46989 75903 -46955
rect 75937 -46989 75995 -46955
rect 76029 -46989 76085 -46955
rect 76119 -46989 76177 -46955
rect 76211 -46989 76269 -46955
rect 76303 -46989 76361 -46955
rect 76395 -46989 76453 -46955
rect 76487 -46989 76545 -46955
rect 76579 -46989 76637 -46955
rect 76671 -46989 76729 -46955
rect 76763 -46989 76821 -46955
rect 76855 -46989 76884 -46955
rect 60486 -47162 60520 -47100
rect 77578 -47115 77607 -47081
rect 77641 -47115 77699 -47081
rect 77733 -47115 77791 -47081
rect 77825 -47115 77883 -47081
rect 77917 -47115 77975 -47081
rect 78009 -47115 78067 -47081
rect 78101 -47115 78159 -47081
rect 78193 -47115 78251 -47081
rect 78285 -47115 78343 -47081
rect 78377 -47115 78435 -47081
rect 78469 -47115 78527 -47081
rect 78561 -47115 78619 -47081
rect 78653 -47115 78711 -47081
rect 78745 -47115 78803 -47081
rect 78837 -47115 78895 -47081
rect 78929 -47115 78987 -47081
rect 79021 -47115 79050 -47081
rect 77961 -47157 78017 -47115
rect 77596 -47160 77927 -47159
rect 59772 -47196 59866 -47162
rect 60426 -47196 60520 -47162
rect 77410 -47169 77927 -47160
rect 77410 -47170 77835 -47169
rect 77410 -47210 77430 -47170
rect 77520 -47203 77835 -47170
rect 77869 -47203 77927 -47169
rect 77520 -47210 77927 -47203
rect 77410 -47220 77540 -47210
rect 77596 -47217 77927 -47210
rect 77961 -47191 77974 -47157
rect 78008 -47191 78017 -47157
rect 77961 -47225 78017 -47191
rect 77596 -47285 77914 -47251
rect 77961 -47259 77974 -47225
rect 78008 -47259 78017 -47225
rect 77961 -47275 78017 -47259
rect 78059 -47160 78113 -47149
rect 78419 -47157 78475 -47115
rect 78147 -47160 78385 -47159
rect 78059 -47169 78385 -47160
rect 78059 -47188 78293 -47169
rect 78093 -47203 78293 -47188
rect 78327 -47203 78385 -47169
rect 78093 -47210 78385 -47203
rect 78093 -47222 78113 -47210
rect 78147 -47217 78385 -47210
rect 78419 -47191 78432 -47157
rect 78466 -47191 78475 -47157
rect 78059 -47256 78113 -47222
rect 78419 -47225 78475 -47191
rect 77596 -47288 77660 -47285
rect 77596 -47322 77613 -47288
rect 77647 -47322 77660 -47288
rect 77880 -47309 77914 -47285
rect 78093 -47290 78113 -47256
rect 77596 -47343 77660 -47322
rect 77700 -47320 77842 -47319
rect 77700 -47360 77780 -47320
rect 77820 -47360 77842 -47320
rect 77880 -47343 78025 -47309
rect 78059 -47343 78113 -47290
rect 78151 -47285 78385 -47251
rect 78419 -47259 78432 -47225
rect 78466 -47259 78475 -47225
rect 78419 -47275 78475 -47259
rect 78517 -47188 78572 -47149
rect 78551 -47222 78572 -47188
rect 78517 -47256 78572 -47222
rect 78647 -47199 78703 -47115
rect 78837 -47157 78903 -47115
rect 78647 -47233 78661 -47199
rect 78695 -47233 78703 -47199
rect 78647 -47249 78703 -47233
rect 78737 -47199 78797 -47183
rect 78737 -47233 78745 -47199
rect 78779 -47233 78797 -47199
rect 78151 -47288 78216 -47285
rect 78151 -47322 78167 -47288
rect 78201 -47322 78216 -47288
rect 78351 -47309 78385 -47285
rect 78551 -47290 78572 -47256
rect 78517 -47300 78572 -47290
rect 78737 -47293 78797 -47233
rect 78837 -47191 78853 -47157
rect 78887 -47191 78903 -47157
rect 78837 -47225 78903 -47191
rect 78837 -47259 78853 -47225
rect 78887 -47259 78903 -47225
rect 78941 -47150 79033 -47149
rect 78941 -47157 79170 -47150
rect 78941 -47191 78957 -47157
rect 78991 -47191 79170 -47157
rect 78941 -47225 79170 -47191
rect 78941 -47259 78957 -47225
rect 78991 -47259 79170 -47225
rect 78151 -47343 78216 -47322
rect 77596 -47380 77666 -47377
rect 77220 -47393 77666 -47380
rect 77220 -47427 77613 -47393
rect 77647 -47427 77666 -47393
rect 59662 -47484 59696 -47430
rect 58966 -47500 59026 -47484
rect 58930 -47518 59026 -47500
rect 59600 -47518 59696 -47484
rect 77220 -47450 77666 -47427
rect 77700 -47393 77842 -47360
rect 77991 -47377 78025 -47343
rect 77700 -47427 77739 -47393
rect 77773 -47427 77842 -47393
rect 77700 -47443 77842 -47427
rect 77876 -47390 77957 -47377
rect 77876 -47430 77900 -47390
rect 77940 -47393 77957 -47390
rect 77949 -47427 77957 -47393
rect 77940 -47430 77957 -47427
rect 77876 -47443 77957 -47430
rect 77991 -47393 78045 -47377
rect 77991 -47427 78011 -47393
rect 77991 -47443 78045 -47427
rect 77220 -47490 77320 -47450
rect 77220 -47530 77240 -47490
rect 77300 -47530 77320 -47490
rect 77596 -47491 77666 -47450
rect 77991 -47477 78025 -47443
rect 77220 -47560 77320 -47530
rect 77703 -47511 78025 -47477
rect 78079 -47490 78113 -47343
rect 78250 -47377 78289 -47319
rect 78351 -47343 78483 -47309
rect 78517 -47343 78670 -47300
rect 78737 -47327 78925 -47293
rect 78449 -47377 78483 -47343
rect 78538 -47370 78670 -47343
rect 78147 -47390 78216 -47377
rect 78147 -47430 78160 -47390
rect 78200 -47430 78216 -47390
rect 78147 -47443 78216 -47430
rect 78250 -47390 78415 -47377
rect 78250 -47430 78290 -47390
rect 78330 -47430 78370 -47390
rect 78410 -47430 78415 -47390
rect 78250 -47443 78415 -47430
rect 78449 -47393 78504 -47377
rect 78449 -47427 78470 -47393
rect 78449 -47443 78504 -47427
rect 78538 -47410 78590 -47370
rect 78630 -47377 78670 -47370
rect 78891 -47377 78925 -47327
rect 78630 -47393 78745 -47377
rect 78630 -47410 78664 -47393
rect 78538 -47427 78664 -47410
rect 78698 -47427 78745 -47393
rect 78789 -47380 78857 -47377
rect 78789 -47420 78800 -47380
rect 78850 -47420 78857 -47380
rect 78789 -47427 78805 -47420
rect 78839 -47427 78857 -47420
rect 78891 -47393 78949 -47377
rect 78891 -47427 78913 -47393
rect 78947 -47427 78949 -47393
rect 78538 -47430 78610 -47427
rect 78449 -47477 78483 -47443
rect 78059 -47507 78113 -47490
rect 77597 -47559 77613 -47525
rect 77647 -47559 77663 -47525
rect 77597 -47625 77663 -47559
rect 77703 -47531 77737 -47511
rect 77877 -47531 77911 -47511
rect 77703 -47581 77737 -47565
rect 77777 -47579 77793 -47545
rect 77827 -47579 77843 -47545
rect 77777 -47625 77843 -47579
rect 78093 -47541 78113 -47507
rect 77877 -47581 77911 -47565
rect 77945 -47579 77971 -47545
rect 78005 -47579 78021 -47545
rect 78059 -47559 78113 -47541
rect 78150 -47511 78483 -47477
rect 78538 -47490 78572 -47430
rect 78891 -47443 78949 -47427
rect 78983 -47380 79170 -47259
rect 78983 -47440 79080 -47380
rect 79140 -47440 79170 -47380
rect 78891 -47461 78925 -47443
rect 78517 -47507 78572 -47490
rect 78150 -47531 78201 -47511
rect 77945 -47625 78021 -47579
rect 78150 -47565 78167 -47531
rect 78335 -47531 78369 -47511
rect 78150 -47581 78201 -47565
rect 78235 -47579 78251 -47545
rect 78285 -47579 78301 -47545
rect 78235 -47625 78301 -47579
rect 78551 -47541 78572 -47507
rect 78335 -47581 78369 -47565
rect 78403 -47579 78429 -47545
rect 78463 -47579 78479 -47545
rect 78517 -47559 78572 -47541
rect 78647 -47499 78925 -47461
rect 78983 -47490 79170 -47440
rect 78647 -47521 78713 -47499
rect 78647 -47555 78661 -47521
rect 78695 -47555 78713 -47521
rect 78983 -47533 79080 -47490
rect 78647 -47571 78713 -47555
rect 78837 -47549 78887 -47533
rect 78403 -47625 78479 -47579
rect 78837 -47583 78853 -47549
rect 78837 -47625 78887 -47583
rect 78921 -47549 79080 -47533
rect 78921 -47583 78937 -47549
rect 78971 -47550 79080 -47549
rect 79140 -47550 79170 -47490
rect 78971 -47583 79170 -47550
rect 78921 -47590 79170 -47583
rect 78921 -47591 79033 -47590
rect 55018 -47786 55052 -47724
rect 53886 -47820 53982 -47786
rect 54956 -47820 55052 -47786
rect 55176 -47678 55272 -47644
rect 55566 -47678 55662 -47644
rect 77578 -47659 77607 -47625
rect 77641 -47659 77699 -47625
rect 77733 -47659 77791 -47625
rect 77825 -47659 77883 -47625
rect 77917 -47659 77975 -47625
rect 78009 -47659 78067 -47625
rect 78101 -47659 78159 -47625
rect 78193 -47659 78251 -47625
rect 78285 -47659 78343 -47625
rect 78377 -47659 78435 -47625
rect 78469 -47659 78527 -47625
rect 78561 -47659 78619 -47625
rect 78653 -47659 78711 -47625
rect 78745 -47659 78803 -47625
rect 78837 -47659 78895 -47625
rect 78929 -47659 78987 -47625
rect 79021 -47659 79050 -47625
rect 55176 -47740 55210 -47678
rect 55628 -47740 55662 -47678
rect 55284 -47792 55300 -47758
rect 55476 -47792 55492 -47758
rect 55526 -47802 55560 -47786
rect 55284 -47880 55300 -47846
rect 55476 -47880 55492 -47846
rect 55526 -47852 55560 -47836
rect 55176 -47960 55210 -47898
rect 77578 -47745 77607 -47711
rect 77641 -47745 77699 -47711
rect 77733 -47745 77791 -47711
rect 77825 -47745 77883 -47711
rect 77917 -47745 77975 -47711
rect 78009 -47745 78067 -47711
rect 78101 -47745 78130 -47711
rect 55628 -47960 55662 -47898
rect 55176 -47994 55272 -47960
rect 55566 -47994 55662 -47960
rect 77150 -47830 77280 -47800
rect 77597 -47811 77663 -47745
rect 77150 -47880 77170 -47830
rect 77260 -47880 77280 -47830
rect 77597 -47845 77613 -47811
rect 77647 -47845 77663 -47811
rect 77703 -47805 77737 -47789
rect 77777 -47791 77843 -47745
rect 77777 -47825 77793 -47791
rect 77827 -47825 77843 -47791
rect 77877 -47805 77911 -47789
rect 77703 -47859 77737 -47839
rect 77945 -47791 78021 -47745
rect 82838 -47765 82867 -47731
rect 82901 -47765 82959 -47731
rect 82993 -47765 83051 -47731
rect 83085 -47765 83143 -47731
rect 83177 -47765 83235 -47731
rect 83269 -47765 83327 -47731
rect 83361 -47765 83419 -47731
rect 83453 -47765 83511 -47731
rect 83545 -47765 83603 -47731
rect 83637 -47765 83695 -47731
rect 83729 -47765 83787 -47731
rect 83821 -47765 83879 -47731
rect 83913 -47765 83971 -47731
rect 84005 -47765 84063 -47731
rect 84097 -47765 84155 -47731
rect 84189 -47765 84247 -47731
rect 84281 -47765 84339 -47731
rect 84373 -47765 84431 -47731
rect 84465 -47765 84523 -47731
rect 84557 -47765 84615 -47731
rect 84649 -47765 84707 -47731
rect 84741 -47765 84799 -47731
rect 84833 -47765 84891 -47731
rect 84925 -47765 84983 -47731
rect 85017 -47765 85075 -47731
rect 85109 -47765 85167 -47731
rect 85201 -47765 85259 -47731
rect 85293 -47765 85351 -47731
rect 85385 -47765 85443 -47731
rect 85477 -47765 85535 -47731
rect 85569 -47765 85627 -47731
rect 85661 -47765 85719 -47731
rect 85753 -47765 85811 -47731
rect 85845 -47765 85903 -47731
rect 85937 -47765 85995 -47731
rect 86029 -47765 86087 -47731
rect 86121 -47765 86179 -47731
rect 86213 -47765 86271 -47731
rect 86305 -47765 86363 -47731
rect 86397 -47765 86455 -47731
rect 86489 -47765 86547 -47731
rect 86581 -47765 86639 -47731
rect 86673 -47765 86731 -47731
rect 86765 -47765 86823 -47731
rect 86857 -47765 86915 -47731
rect 86949 -47765 87007 -47731
rect 87041 -47765 87099 -47731
rect 87133 -47765 87191 -47731
rect 87225 -47765 87283 -47731
rect 87317 -47765 87375 -47731
rect 87409 -47765 87467 -47731
rect 87501 -47765 87559 -47731
rect 87593 -47765 87651 -47731
rect 87685 -47765 87743 -47731
rect 87777 -47765 87835 -47731
rect 87869 -47765 87927 -47731
rect 87961 -47765 88019 -47731
rect 88053 -47765 88111 -47731
rect 88145 -47765 88203 -47731
rect 88237 -47765 88295 -47731
rect 88329 -47765 88387 -47731
rect 88421 -47765 88479 -47731
rect 88513 -47765 88571 -47731
rect 88605 -47765 88663 -47731
rect 88697 -47765 88755 -47731
rect 88789 -47765 88847 -47731
rect 88881 -47765 88939 -47731
rect 88973 -47765 89031 -47731
rect 89065 -47765 89123 -47731
rect 89157 -47765 89215 -47731
rect 89249 -47765 89307 -47731
rect 89341 -47765 89399 -47731
rect 89433 -47765 89491 -47731
rect 89525 -47765 89583 -47731
rect 89617 -47765 89675 -47731
rect 89709 -47765 89767 -47731
rect 89801 -47765 89859 -47731
rect 89893 -47765 89951 -47731
rect 89985 -47765 90043 -47731
rect 90077 -47765 90135 -47731
rect 90169 -47765 90227 -47731
rect 90261 -47765 90319 -47731
rect 90353 -47765 90411 -47731
rect 90445 -47765 90503 -47731
rect 90537 -47765 90595 -47731
rect 90629 -47765 90687 -47731
rect 90721 -47765 90779 -47731
rect 90813 -47765 90871 -47731
rect 90905 -47765 90963 -47731
rect 90997 -47765 91055 -47731
rect 91089 -47765 91147 -47731
rect 91181 -47765 91239 -47731
rect 91273 -47765 91331 -47731
rect 91365 -47765 91394 -47731
rect 77945 -47825 77971 -47791
rect 78005 -47825 78021 -47791
rect 78080 -47811 78220 -47810
rect 77877 -47859 77911 -47839
rect 78059 -47829 78220 -47811
rect 77596 -47880 77666 -47879
rect 77150 -47943 77666 -47880
rect 77703 -47893 78025 -47859
rect 78093 -47830 78220 -47829
rect 78093 -47863 78160 -47830
rect 78059 -47870 78160 -47863
rect 78200 -47870 78220 -47830
rect 78059 -47880 78220 -47870
rect 77991 -47927 78025 -47893
rect 77150 -47977 77613 -47943
rect 77647 -47977 77666 -47943
rect 77150 -47990 77666 -47977
rect 77596 -47993 77666 -47990
rect 77700 -47943 77842 -47927
rect 77700 -47977 77739 -47943
rect 77773 -47977 77842 -47943
rect 77700 -48000 77842 -47977
rect 77876 -47940 77957 -47927
rect 77876 -47980 77900 -47940
rect 77940 -47943 77957 -47940
rect 77949 -47977 77957 -47943
rect 77940 -47980 77957 -47977
rect 77876 -47993 77957 -47980
rect 77991 -47943 78045 -47927
rect 77991 -47977 78011 -47943
rect 77991 -47993 78045 -47977
rect 78079 -47940 78220 -47880
rect 83067 -47823 83133 -47765
rect 83067 -47857 83083 -47823
rect 83117 -47857 83133 -47823
rect 83067 -47891 83133 -47857
rect 78079 -47980 78160 -47940
rect 78200 -47980 78220 -47940
rect 77596 -48048 77660 -48027
rect 77596 -48082 77613 -48048
rect 77647 -48082 77660 -48048
rect 77700 -48040 77770 -48000
rect 77810 -48040 77842 -48000
rect 77991 -48027 78025 -47993
rect 78079 -48027 78220 -47980
rect 82892 -47943 82970 -47924
rect 83067 -47925 83083 -47891
rect 83117 -47925 83133 -47891
rect 83167 -47807 83274 -47799
rect 83167 -47841 83183 -47807
rect 83217 -47841 83274 -47807
rect 83167 -47875 83274 -47841
rect 83167 -47909 83183 -47875
rect 83217 -47909 83274 -47875
rect 83167 -47923 83274 -47909
rect 82892 -47977 82914 -47943
rect 82948 -47959 82970 -47943
rect 82948 -47977 83177 -47959
rect 82892 -47993 83177 -47977
rect 77700 -48051 77842 -48040
rect 77596 -48085 77660 -48082
rect 77880 -48061 78025 -48027
rect 78059 -48060 78220 -48027
rect 77880 -48085 77914 -48061
rect 77596 -48119 77914 -48085
rect 78059 -48080 78160 -48060
rect 77961 -48111 78017 -48095
rect 77400 -48160 77490 -48140
rect 77961 -48145 77974 -48111
rect 78008 -48145 78017 -48111
rect 77596 -48160 77927 -48153
rect 77400 -48210 77420 -48160
rect 77470 -48167 77927 -48160
rect 77470 -48201 77835 -48167
rect 77869 -48201 77927 -48167
rect 77470 -48210 77927 -48201
rect 77400 -48230 77490 -48210
rect 77596 -48211 77927 -48210
rect 77961 -48179 78017 -48145
rect 77961 -48213 77974 -48179
rect 78008 -48213 78017 -48179
rect 77961 -48255 78017 -48213
rect 78093 -48100 78160 -48080
rect 78200 -48100 78220 -48060
rect 78093 -48114 78220 -48100
rect 78059 -48140 78220 -48114
rect 82867 -48040 82938 -48027
rect 82867 -48130 82870 -48040
rect 82930 -48043 82938 -48040
rect 82930 -48130 82938 -48077
rect 82867 -48139 82938 -48130
rect 78059 -48148 78113 -48140
rect 78093 -48182 78113 -48148
rect 82972 -48173 83006 -47993
rect 83040 -48040 83093 -48027
rect 83040 -48043 83050 -48040
rect 83040 -48130 83050 -48077
rect 83090 -48130 83093 -48040
rect 83143 -48043 83177 -47993
rect 83143 -48093 83177 -48077
rect 83211 -48000 83274 -47923
rect 83366 -47807 83408 -47765
rect 83366 -47841 83374 -47807
rect 83366 -47875 83408 -47841
rect 83366 -47909 83374 -47875
rect 83366 -47943 83408 -47909
rect 83366 -47977 83374 -47943
rect 83366 -47993 83408 -47977
rect 83442 -47807 83508 -47799
rect 83442 -47841 83458 -47807
rect 83492 -47841 83508 -47807
rect 83442 -47875 83508 -47841
rect 83442 -47909 83458 -47875
rect 83492 -47909 83508 -47875
rect 83442 -47943 83508 -47909
rect 83442 -47977 83458 -47943
rect 83492 -47977 83508 -47943
rect 83442 -47995 83508 -47977
rect 83600 -47807 83653 -47765
rect 83600 -47841 83619 -47807
rect 83600 -47875 83653 -47841
rect 83600 -47909 83619 -47875
rect 83600 -47943 83653 -47909
rect 83600 -47977 83619 -47943
rect 83600 -47993 83653 -47977
rect 83687 -47807 83753 -47799
rect 83687 -47841 83703 -47807
rect 83737 -47841 83753 -47807
rect 83687 -47875 83753 -47841
rect 83687 -47909 83703 -47875
rect 83737 -47909 83753 -47875
rect 83687 -47943 83753 -47909
rect 83787 -47807 83821 -47765
rect 83787 -47875 83821 -47841
rect 83787 -47925 83821 -47909
rect 83855 -47807 83921 -47799
rect 83855 -47841 83871 -47807
rect 83905 -47841 83921 -47807
rect 83855 -47875 83921 -47841
rect 83955 -47807 83997 -47765
rect 83989 -47841 83997 -47807
rect 83955 -47857 83997 -47841
rect 84074 -47807 84116 -47765
rect 84074 -47841 84082 -47807
rect 83855 -47909 83871 -47875
rect 83905 -47909 83921 -47875
rect 83687 -47977 83703 -47943
rect 83737 -47959 83753 -47943
rect 83855 -47943 83921 -47909
rect 83855 -47959 83871 -47943
rect 83737 -47977 83871 -47959
rect 83905 -47955 83921 -47943
rect 84074 -47875 84116 -47841
rect 84074 -47909 84082 -47875
rect 84074 -47945 84116 -47909
rect 83905 -47977 84008 -47955
rect 83687 -47993 84008 -47977
rect 83211 -48030 83320 -48000
rect 83362 -48030 83428 -48029
rect 83211 -48043 83428 -48030
rect 83211 -48070 83378 -48043
rect 83211 -48110 83320 -48070
rect 83362 -48077 83378 -48070
rect 83412 -48077 83428 -48043
rect 83462 -48030 83508 -47995
rect 83595 -48030 83921 -48027
rect 83462 -48043 83921 -48030
rect 83462 -48077 83611 -48043
rect 83645 -48077 83703 -48043
rect 83737 -48077 83787 -48043
rect 83821 -48077 83871 -48043
rect 83905 -48077 83921 -48043
rect 83955 -48030 84008 -47993
rect 84074 -47979 84082 -47945
rect 84074 -47995 84116 -47979
rect 84150 -47807 84216 -47799
rect 84150 -47841 84166 -47807
rect 84200 -47841 84216 -47807
rect 84150 -47875 84216 -47841
rect 84150 -47909 84166 -47875
rect 84200 -47909 84216 -47875
rect 84150 -47945 84216 -47909
rect 84250 -47807 84284 -47765
rect 84250 -47875 84284 -47841
rect 84250 -47925 84284 -47909
rect 84318 -47807 84384 -47799
rect 84318 -47841 84334 -47807
rect 84368 -47841 84384 -47807
rect 84318 -47875 84384 -47841
rect 84318 -47909 84334 -47875
rect 84368 -47909 84384 -47875
rect 84150 -47979 84166 -47945
rect 84200 -47959 84216 -47945
rect 84318 -47945 84384 -47909
rect 84418 -47807 84452 -47765
rect 84418 -47875 84452 -47841
rect 84418 -47925 84452 -47909
rect 84486 -47807 84552 -47799
rect 84486 -47841 84502 -47807
rect 84536 -47841 84552 -47807
rect 84486 -47875 84552 -47841
rect 84486 -47909 84502 -47875
rect 84536 -47909 84552 -47875
rect 84318 -47959 84334 -47945
rect 84200 -47979 84334 -47959
rect 84368 -47959 84384 -47945
rect 84486 -47945 84552 -47909
rect 84586 -47807 84620 -47765
rect 84586 -47875 84620 -47841
rect 84586 -47925 84620 -47909
rect 84654 -47807 84720 -47799
rect 84654 -47841 84670 -47807
rect 84704 -47841 84720 -47807
rect 84654 -47875 84720 -47841
rect 84654 -47909 84670 -47875
rect 84704 -47909 84720 -47875
rect 84486 -47959 84502 -47945
rect 84368 -47979 84502 -47959
rect 84536 -47959 84552 -47945
rect 84654 -47945 84720 -47909
rect 84754 -47807 84788 -47765
rect 84754 -47875 84788 -47841
rect 84754 -47925 84788 -47909
rect 84822 -47807 84888 -47799
rect 84822 -47841 84838 -47807
rect 84872 -47841 84888 -47807
rect 84822 -47875 84888 -47841
rect 84822 -47909 84838 -47875
rect 84872 -47909 84888 -47875
rect 84654 -47959 84670 -47945
rect 84536 -47979 84670 -47959
rect 84704 -47959 84720 -47945
rect 84822 -47945 84888 -47909
rect 84922 -47807 84956 -47765
rect 84922 -47875 84956 -47841
rect 84922 -47925 84956 -47909
rect 84990 -47807 85056 -47799
rect 84990 -47841 85006 -47807
rect 85040 -47841 85056 -47807
rect 84990 -47875 85056 -47841
rect 84990 -47909 85006 -47875
rect 85040 -47909 85056 -47875
rect 84822 -47959 84838 -47945
rect 84704 -47979 84838 -47959
rect 84872 -47959 84888 -47945
rect 84990 -47945 85056 -47909
rect 85090 -47807 85124 -47765
rect 85090 -47875 85124 -47841
rect 85090 -47925 85124 -47909
rect 85158 -47807 85224 -47799
rect 85158 -47841 85174 -47807
rect 85208 -47841 85224 -47807
rect 85158 -47875 85224 -47841
rect 85158 -47909 85174 -47875
rect 85208 -47909 85224 -47875
rect 84990 -47959 85006 -47945
rect 84872 -47979 85006 -47959
rect 85040 -47959 85056 -47945
rect 85158 -47945 85224 -47909
rect 85258 -47807 85292 -47765
rect 85258 -47875 85292 -47841
rect 85258 -47925 85292 -47909
rect 85326 -47807 85392 -47799
rect 85326 -47841 85342 -47807
rect 85376 -47841 85392 -47807
rect 85326 -47875 85392 -47841
rect 85326 -47909 85342 -47875
rect 85376 -47909 85392 -47875
rect 85158 -47959 85174 -47945
rect 85040 -47979 85174 -47959
rect 85208 -47959 85224 -47945
rect 85326 -47945 85392 -47909
rect 85426 -47807 85468 -47765
rect 85460 -47841 85468 -47807
rect 85426 -47875 85468 -47841
rect 85460 -47909 85468 -47875
rect 85426 -47925 85468 -47909
rect 85546 -47807 85588 -47765
rect 85546 -47841 85554 -47807
rect 85546 -47875 85588 -47841
rect 85546 -47909 85554 -47875
rect 85326 -47958 85342 -47945
rect 85376 -47958 85392 -47945
rect 85326 -47959 85334 -47958
rect 85208 -47979 85334 -47959
rect 84150 -47993 85334 -47979
rect 84051 -48030 85139 -48029
rect 83955 -48043 85139 -48030
rect 83955 -48077 84076 -48043
rect 84110 -48077 84250 -48043
rect 84284 -48077 84418 -48043
rect 84452 -48077 84587 -48043
rect 84621 -48077 84754 -48043
rect 84788 -48077 84922 -48043
rect 84956 -48077 85089 -48043
rect 85123 -48077 85139 -48043
rect 83462 -48080 83660 -48077
rect 83955 -48080 84120 -48077
rect 83211 -48127 83274 -48110
rect 83040 -48139 83093 -48130
rect 83151 -48129 83274 -48127
rect 83151 -48163 83167 -48129
rect 83201 -48163 83274 -48129
rect 78059 -48221 78113 -48182
rect 82888 -48189 82936 -48173
rect 82888 -48223 82902 -48189
rect 77578 -48289 77607 -48255
rect 77641 -48289 77699 -48255
rect 77733 -48289 77791 -48255
rect 77825 -48289 77883 -48255
rect 77917 -48289 77975 -48255
rect 78009 -48289 78067 -48255
rect 78101 -48289 78130 -48255
rect 77578 -48365 77607 -48331
rect 77641 -48365 77699 -48331
rect 77733 -48365 77791 -48331
rect 77825 -48365 77883 -48331
rect 77917 -48365 77975 -48331
rect 78009 -48365 78038 -48331
rect 77635 -48449 77691 -48365
rect 77825 -48407 77891 -48365
rect 82888 -48275 82936 -48223
rect 82972 -48189 83028 -48173
rect 82972 -48223 82986 -48189
rect 83020 -48223 83028 -48189
rect 82972 -48239 83028 -48223
rect 83074 -48189 83117 -48173
rect 83074 -48223 83082 -48189
rect 83116 -48223 83117 -48189
rect 83074 -48275 83117 -48223
rect 83151 -48197 83274 -48163
rect 83151 -48231 83167 -48197
rect 83201 -48231 83274 -48197
rect 83151 -48241 83274 -48231
rect 83362 -48127 83408 -48111
rect 83462 -48115 83508 -48080
rect 83955 -48111 84008 -48080
rect 85326 -48111 85334 -47993
rect 83362 -48161 83374 -48127
rect 83362 -48195 83408 -48161
rect 83362 -48229 83374 -48195
rect 83362 -48275 83408 -48229
rect 83442 -48127 83508 -48115
rect 83442 -48161 83458 -48127
rect 83492 -48161 83508 -48127
rect 83442 -48195 83508 -48161
rect 83687 -48147 84008 -48111
rect 84070 -48131 84116 -48115
rect 83442 -48229 83458 -48195
rect 83492 -48229 83508 -48195
rect 83442 -48241 83508 -48229
rect 83600 -48199 83653 -48183
rect 83600 -48233 83619 -48199
rect 83600 -48275 83653 -48233
rect 83687 -48191 83753 -48147
rect 83687 -48225 83703 -48191
rect 83737 -48225 83753 -48191
rect 83687 -48241 83753 -48225
rect 83787 -48199 83821 -48183
rect 83787 -48275 83821 -48233
rect 83855 -48191 83921 -48147
rect 84070 -48165 84082 -48131
rect 83855 -48225 83871 -48191
rect 83905 -48225 83921 -48191
rect 83855 -48241 83921 -48225
rect 83955 -48198 84005 -48182
rect 83989 -48232 84005 -48198
rect 83955 -48275 84005 -48232
rect 84070 -48199 84116 -48165
rect 84070 -48233 84082 -48199
rect 84070 -48275 84116 -48233
rect 84150 -48128 85334 -48111
rect 85384 -48128 85392 -47958
rect 85546 -47945 85588 -47909
rect 85546 -47979 85554 -47945
rect 85546 -47995 85588 -47979
rect 85622 -47807 85688 -47799
rect 85622 -47841 85638 -47807
rect 85672 -47841 85688 -47807
rect 85622 -47875 85688 -47841
rect 85622 -47909 85638 -47875
rect 85672 -47909 85688 -47875
rect 85622 -47945 85688 -47909
rect 85722 -47807 85756 -47765
rect 85722 -47875 85756 -47841
rect 85722 -47925 85756 -47909
rect 85790 -47807 85856 -47799
rect 85790 -47841 85806 -47807
rect 85840 -47841 85856 -47807
rect 85790 -47875 85856 -47841
rect 85790 -47909 85806 -47875
rect 85840 -47909 85856 -47875
rect 85622 -47979 85638 -47945
rect 85672 -47959 85688 -47945
rect 85790 -47945 85856 -47909
rect 85890 -47807 85924 -47765
rect 85890 -47875 85924 -47841
rect 85890 -47925 85924 -47909
rect 85958 -47807 86024 -47799
rect 85958 -47841 85974 -47807
rect 86008 -47841 86024 -47807
rect 85958 -47875 86024 -47841
rect 85958 -47909 85974 -47875
rect 86008 -47909 86024 -47875
rect 85790 -47959 85806 -47945
rect 85672 -47979 85806 -47959
rect 85840 -47959 85856 -47945
rect 85958 -47945 86024 -47909
rect 86058 -47807 86092 -47765
rect 86058 -47875 86092 -47841
rect 86058 -47925 86092 -47909
rect 86126 -47807 86192 -47799
rect 86126 -47841 86142 -47807
rect 86176 -47841 86192 -47807
rect 86126 -47875 86192 -47841
rect 86126 -47909 86142 -47875
rect 86176 -47909 86192 -47875
rect 85958 -47959 85974 -47945
rect 85840 -47979 85974 -47959
rect 86008 -47959 86024 -47945
rect 86126 -47945 86192 -47909
rect 86226 -47807 86260 -47765
rect 86226 -47875 86260 -47841
rect 86226 -47925 86260 -47909
rect 86294 -47807 86360 -47799
rect 86294 -47841 86310 -47807
rect 86344 -47841 86360 -47807
rect 86294 -47875 86360 -47841
rect 86294 -47909 86310 -47875
rect 86344 -47909 86360 -47875
rect 86126 -47959 86142 -47945
rect 86008 -47979 86142 -47959
rect 86176 -47959 86192 -47945
rect 86294 -47945 86360 -47909
rect 86394 -47807 86428 -47765
rect 86394 -47875 86428 -47841
rect 86394 -47925 86428 -47909
rect 86462 -47807 86528 -47799
rect 86462 -47841 86478 -47807
rect 86512 -47841 86528 -47807
rect 86462 -47875 86528 -47841
rect 86462 -47909 86478 -47875
rect 86512 -47909 86528 -47875
rect 86294 -47959 86310 -47945
rect 86176 -47979 86310 -47959
rect 86344 -47959 86360 -47945
rect 86462 -47945 86528 -47909
rect 86562 -47807 86596 -47765
rect 86562 -47875 86596 -47841
rect 86562 -47925 86596 -47909
rect 86630 -47807 86696 -47799
rect 86630 -47841 86646 -47807
rect 86680 -47841 86696 -47807
rect 86630 -47875 86696 -47841
rect 86630 -47909 86646 -47875
rect 86680 -47909 86696 -47875
rect 86462 -47959 86478 -47945
rect 86344 -47979 86478 -47959
rect 86512 -47959 86528 -47945
rect 86630 -47945 86696 -47909
rect 86730 -47807 86764 -47765
rect 86730 -47875 86764 -47841
rect 86730 -47925 86764 -47909
rect 86798 -47807 86864 -47799
rect 86798 -47841 86814 -47807
rect 86848 -47841 86864 -47807
rect 86798 -47875 86864 -47841
rect 86798 -47909 86814 -47875
rect 86848 -47909 86864 -47875
rect 86630 -47959 86646 -47945
rect 86512 -47979 86646 -47959
rect 86680 -47959 86696 -47945
rect 86798 -47938 86864 -47909
rect 86898 -47807 86940 -47765
rect 86932 -47841 86940 -47807
rect 86898 -47875 86940 -47841
rect 86932 -47909 86940 -47875
rect 86898 -47925 86940 -47909
rect 87018 -47807 87060 -47765
rect 87018 -47841 87026 -47807
rect 87018 -47875 87060 -47841
rect 87018 -47909 87026 -47875
rect 86798 -47959 86814 -47938
rect 86680 -47979 86814 -47959
rect 85622 -47993 86814 -47979
rect 85523 -48035 86611 -48029
rect 85523 -48043 85614 -48035
rect 86475 -48043 86611 -48035
rect 85523 -48077 85548 -48043
rect 85582 -48069 85614 -48043
rect 86475 -48069 86561 -48043
rect 85582 -48077 85722 -48069
rect 85756 -48077 85890 -48069
rect 85924 -48077 86059 -48069
rect 86093 -48077 86226 -48069
rect 86260 -48077 86394 -48069
rect 86428 -48077 86561 -48069
rect 86595 -48077 86611 -48043
rect 86798 -48111 86814 -47993
rect 84150 -48131 85392 -48128
rect 84150 -48165 84166 -48131
rect 84200 -48149 84334 -48131
rect 84200 -48165 84216 -48149
rect 84150 -48199 84216 -48165
rect 84318 -48165 84334 -48149
rect 84368 -48149 84502 -48131
rect 84368 -48165 84384 -48149
rect 84150 -48233 84166 -48199
rect 84200 -48233 84216 -48199
rect 84150 -48241 84216 -48233
rect 84250 -48199 84284 -48183
rect 84250 -48275 84284 -48233
rect 84318 -48199 84384 -48165
rect 84486 -48165 84502 -48149
rect 84536 -48149 84670 -48131
rect 84536 -48165 84552 -48149
rect 84318 -48233 84334 -48199
rect 84368 -48233 84384 -48199
rect 84318 -48241 84384 -48233
rect 84418 -48199 84452 -48183
rect 84418 -48275 84452 -48233
rect 84486 -48199 84552 -48165
rect 84654 -48165 84670 -48149
rect 84704 -48149 84838 -48131
rect 84704 -48165 84720 -48149
rect 84486 -48233 84502 -48199
rect 84536 -48233 84552 -48199
rect 84486 -48241 84552 -48233
rect 84586 -48199 84620 -48183
rect 84586 -48275 84620 -48233
rect 84654 -48199 84720 -48165
rect 84822 -48165 84838 -48149
rect 84872 -48149 85006 -48131
rect 84872 -48165 84888 -48149
rect 84654 -48233 84670 -48199
rect 84704 -48233 84720 -48199
rect 84654 -48241 84720 -48233
rect 84754 -48199 84788 -48183
rect 84754 -48275 84788 -48233
rect 84822 -48199 84888 -48165
rect 84990 -48165 85006 -48149
rect 85040 -48149 85174 -48131
rect 85040 -48165 85056 -48149
rect 84822 -48233 84838 -48199
rect 84872 -48233 84888 -48199
rect 84822 -48241 84888 -48233
rect 84922 -48199 84956 -48183
rect 84922 -48275 84956 -48233
rect 84990 -48199 85056 -48165
rect 85158 -48165 85174 -48149
rect 85208 -48149 85342 -48131
rect 85208 -48165 85224 -48149
rect 84990 -48233 85006 -48199
rect 85040 -48233 85056 -48199
rect 84990 -48241 85056 -48233
rect 85090 -48199 85124 -48183
rect 85090 -48275 85124 -48233
rect 85158 -48199 85224 -48165
rect 85326 -48165 85342 -48149
rect 85376 -48165 85392 -48131
rect 85158 -48233 85174 -48199
rect 85208 -48233 85224 -48199
rect 85158 -48241 85224 -48233
rect 85258 -48199 85292 -48183
rect 85258 -48275 85292 -48233
rect 85326 -48199 85392 -48165
rect 85326 -48233 85342 -48199
rect 85376 -48233 85392 -48199
rect 85326 -48241 85392 -48233
rect 85426 -48131 85468 -48115
rect 85460 -48165 85468 -48131
rect 85426 -48199 85468 -48165
rect 85460 -48233 85468 -48199
rect 85426 -48275 85468 -48233
rect 85542 -48131 85588 -48115
rect 85542 -48165 85554 -48131
rect 85542 -48199 85588 -48165
rect 85542 -48233 85554 -48199
rect 85542 -48275 85588 -48233
rect 85622 -48128 86814 -48111
rect 87018 -47945 87060 -47909
rect 87018 -47979 87026 -47945
rect 87018 -47995 87060 -47979
rect 87094 -47807 87160 -47799
rect 87094 -47841 87110 -47807
rect 87144 -47841 87160 -47807
rect 87094 -47875 87160 -47841
rect 87094 -47909 87110 -47875
rect 87144 -47909 87160 -47875
rect 87094 -47945 87160 -47909
rect 87194 -47807 87228 -47765
rect 87194 -47875 87228 -47841
rect 87194 -47925 87228 -47909
rect 87262 -47807 87328 -47799
rect 87262 -47841 87278 -47807
rect 87312 -47841 87328 -47807
rect 87262 -47875 87328 -47841
rect 87262 -47909 87278 -47875
rect 87312 -47909 87328 -47875
rect 87094 -47979 87110 -47945
rect 87144 -47959 87160 -47945
rect 87262 -47945 87328 -47909
rect 87362 -47807 87396 -47765
rect 87362 -47875 87396 -47841
rect 87362 -47925 87396 -47909
rect 87430 -47807 87496 -47799
rect 87430 -47841 87446 -47807
rect 87480 -47841 87496 -47807
rect 87430 -47875 87496 -47841
rect 87430 -47909 87446 -47875
rect 87480 -47909 87496 -47875
rect 87262 -47959 87278 -47945
rect 87144 -47979 87278 -47959
rect 87312 -47959 87328 -47945
rect 87430 -47945 87496 -47909
rect 87530 -47807 87564 -47765
rect 87530 -47875 87564 -47841
rect 87530 -47925 87564 -47909
rect 87598 -47807 87664 -47799
rect 87598 -47841 87614 -47807
rect 87648 -47841 87664 -47807
rect 87598 -47875 87664 -47841
rect 87598 -47909 87614 -47875
rect 87648 -47909 87664 -47875
rect 87430 -47959 87446 -47945
rect 87312 -47979 87446 -47959
rect 87480 -47959 87496 -47945
rect 87598 -47945 87664 -47909
rect 87698 -47807 87732 -47765
rect 87698 -47875 87732 -47841
rect 87698 -47925 87732 -47909
rect 87766 -47807 87832 -47799
rect 87766 -47841 87782 -47807
rect 87816 -47841 87832 -47807
rect 87766 -47875 87832 -47841
rect 87766 -47909 87782 -47875
rect 87816 -47909 87832 -47875
rect 87598 -47959 87614 -47945
rect 87480 -47979 87614 -47959
rect 87648 -47959 87664 -47945
rect 87766 -47945 87832 -47909
rect 87866 -47807 87900 -47765
rect 87866 -47875 87900 -47841
rect 87866 -47925 87900 -47909
rect 87934 -47807 88000 -47799
rect 87934 -47841 87950 -47807
rect 87984 -47841 88000 -47807
rect 87934 -47875 88000 -47841
rect 87934 -47909 87950 -47875
rect 87984 -47909 88000 -47875
rect 87766 -47959 87782 -47945
rect 87648 -47979 87782 -47959
rect 87816 -47959 87832 -47945
rect 87934 -47945 88000 -47909
rect 88034 -47807 88068 -47765
rect 88034 -47875 88068 -47841
rect 88034 -47925 88068 -47909
rect 88102 -47807 88168 -47799
rect 88102 -47841 88118 -47807
rect 88152 -47841 88168 -47807
rect 88102 -47875 88168 -47841
rect 88102 -47909 88118 -47875
rect 88152 -47909 88168 -47875
rect 87934 -47959 87950 -47945
rect 87816 -47979 87950 -47959
rect 87984 -47959 88000 -47945
rect 88102 -47945 88168 -47909
rect 88202 -47807 88236 -47765
rect 88202 -47875 88236 -47841
rect 88202 -47925 88236 -47909
rect 88270 -47807 88336 -47799
rect 88270 -47841 88286 -47807
rect 88320 -47841 88336 -47807
rect 88270 -47875 88336 -47841
rect 88270 -47909 88286 -47875
rect 88320 -47909 88336 -47875
rect 88102 -47959 88118 -47945
rect 87984 -47979 88118 -47959
rect 88152 -47959 88168 -47945
rect 88270 -47945 88336 -47909
rect 88370 -47807 88412 -47765
rect 88404 -47841 88412 -47807
rect 88370 -47875 88412 -47841
rect 88404 -47909 88412 -47875
rect 88370 -47925 88412 -47909
rect 88490 -47807 88532 -47765
rect 88490 -47841 88498 -47807
rect 88490 -47875 88532 -47841
rect 88490 -47909 88498 -47875
rect 88270 -47948 88286 -47945
rect 88320 -47948 88336 -47945
rect 88270 -47959 88284 -47948
rect 88152 -47979 88284 -47959
rect 87094 -47993 88284 -47979
rect 86995 -48034 88083 -48029
rect 86995 -48043 87048 -48034
rect 87909 -48043 88083 -48034
rect 86995 -48077 87020 -48043
rect 87909 -48068 88033 -48043
rect 87054 -48077 87194 -48068
rect 87228 -48077 87362 -48068
rect 87396 -48077 87531 -48068
rect 87565 -48077 87698 -48068
rect 87732 -48077 87866 -48068
rect 87900 -48077 88033 -48068
rect 88067 -48077 88083 -48043
rect 88270 -48111 88284 -47993
rect 85622 -48131 86864 -48128
rect 85622 -48165 85638 -48131
rect 85672 -48149 85806 -48131
rect 85672 -48165 85688 -48149
rect 85622 -48199 85688 -48165
rect 85790 -48165 85806 -48149
rect 85840 -48149 85974 -48131
rect 85840 -48165 85856 -48149
rect 85622 -48233 85638 -48199
rect 85672 -48233 85688 -48199
rect 85622 -48241 85688 -48233
rect 85722 -48199 85756 -48183
rect 85722 -48275 85756 -48233
rect 85790 -48199 85856 -48165
rect 85958 -48165 85974 -48149
rect 86008 -48149 86142 -48131
rect 86008 -48165 86024 -48149
rect 85790 -48233 85806 -48199
rect 85840 -48233 85856 -48199
rect 85790 -48241 85856 -48233
rect 85890 -48199 85924 -48183
rect 85890 -48275 85924 -48233
rect 85958 -48199 86024 -48165
rect 86126 -48165 86142 -48149
rect 86176 -48149 86310 -48131
rect 86176 -48165 86192 -48149
rect 85958 -48233 85974 -48199
rect 86008 -48233 86024 -48199
rect 85958 -48241 86024 -48233
rect 86058 -48199 86092 -48183
rect 86058 -48275 86092 -48233
rect 86126 -48199 86192 -48165
rect 86294 -48165 86310 -48149
rect 86344 -48149 86478 -48131
rect 86344 -48165 86360 -48149
rect 86126 -48233 86142 -48199
rect 86176 -48233 86192 -48199
rect 86126 -48241 86192 -48233
rect 86226 -48199 86260 -48183
rect 86226 -48275 86260 -48233
rect 86294 -48199 86360 -48165
rect 86462 -48165 86478 -48149
rect 86512 -48149 86646 -48131
rect 86512 -48165 86528 -48149
rect 86294 -48233 86310 -48199
rect 86344 -48233 86360 -48199
rect 86294 -48241 86360 -48233
rect 86394 -48199 86428 -48183
rect 86394 -48275 86428 -48233
rect 86462 -48199 86528 -48165
rect 86630 -48165 86646 -48149
rect 86680 -48149 86814 -48131
rect 86680 -48165 86696 -48149
rect 86462 -48233 86478 -48199
rect 86512 -48233 86528 -48199
rect 86462 -48241 86528 -48233
rect 86562 -48199 86596 -48183
rect 86562 -48275 86596 -48233
rect 86630 -48199 86696 -48165
rect 86798 -48165 86814 -48149
rect 86848 -48165 86864 -48131
rect 86630 -48233 86646 -48199
rect 86680 -48233 86696 -48199
rect 86630 -48241 86696 -48233
rect 86730 -48199 86764 -48183
rect 86730 -48275 86764 -48233
rect 86798 -48199 86864 -48165
rect 86798 -48233 86814 -48199
rect 86848 -48233 86864 -48199
rect 86798 -48241 86864 -48233
rect 86898 -48131 86940 -48115
rect 86932 -48165 86940 -48131
rect 86898 -48199 86940 -48165
rect 86932 -48233 86940 -48199
rect 86898 -48275 86940 -48233
rect 87014 -48131 87060 -48115
rect 87014 -48165 87026 -48131
rect 87014 -48199 87060 -48165
rect 87014 -48233 87026 -48199
rect 87014 -48275 87060 -48233
rect 87094 -48128 88284 -48111
rect 88334 -48128 88336 -47948
rect 88490 -47945 88532 -47909
rect 88490 -47979 88498 -47945
rect 88490 -47995 88532 -47979
rect 88566 -47807 88632 -47799
rect 88566 -47841 88582 -47807
rect 88616 -47841 88632 -47807
rect 88566 -47875 88632 -47841
rect 88566 -47909 88582 -47875
rect 88616 -47909 88632 -47875
rect 88566 -47945 88632 -47909
rect 88666 -47807 88700 -47765
rect 88666 -47875 88700 -47841
rect 88666 -47925 88700 -47909
rect 88734 -47807 88800 -47799
rect 88734 -47841 88750 -47807
rect 88784 -47841 88800 -47807
rect 88734 -47875 88800 -47841
rect 88734 -47909 88750 -47875
rect 88784 -47909 88800 -47875
rect 88566 -47979 88582 -47945
rect 88616 -47959 88632 -47945
rect 88734 -47945 88800 -47909
rect 88834 -47807 88868 -47765
rect 88834 -47875 88868 -47841
rect 88834 -47925 88868 -47909
rect 88902 -47807 88968 -47799
rect 88902 -47841 88918 -47807
rect 88952 -47841 88968 -47807
rect 88902 -47875 88968 -47841
rect 88902 -47909 88918 -47875
rect 88952 -47909 88968 -47875
rect 88734 -47959 88750 -47945
rect 88616 -47979 88750 -47959
rect 88784 -47959 88800 -47945
rect 88902 -47945 88968 -47909
rect 89002 -47807 89036 -47765
rect 89002 -47875 89036 -47841
rect 89002 -47925 89036 -47909
rect 89070 -47807 89136 -47799
rect 89070 -47841 89086 -47807
rect 89120 -47841 89136 -47807
rect 89070 -47875 89136 -47841
rect 89070 -47909 89086 -47875
rect 89120 -47909 89136 -47875
rect 88902 -47959 88918 -47945
rect 88784 -47979 88918 -47959
rect 88952 -47959 88968 -47945
rect 89070 -47945 89136 -47909
rect 89170 -47807 89204 -47765
rect 89170 -47875 89204 -47841
rect 89170 -47925 89204 -47909
rect 89238 -47807 89304 -47799
rect 89238 -47841 89254 -47807
rect 89288 -47841 89304 -47807
rect 89238 -47875 89304 -47841
rect 89238 -47909 89254 -47875
rect 89288 -47909 89304 -47875
rect 89070 -47959 89086 -47945
rect 88952 -47979 89086 -47959
rect 89120 -47959 89136 -47945
rect 89238 -47945 89304 -47909
rect 89338 -47807 89372 -47765
rect 89338 -47875 89372 -47841
rect 89338 -47925 89372 -47909
rect 89406 -47807 89472 -47799
rect 89406 -47841 89422 -47807
rect 89456 -47841 89472 -47807
rect 89406 -47875 89472 -47841
rect 89406 -47909 89422 -47875
rect 89456 -47909 89472 -47875
rect 89238 -47959 89254 -47945
rect 89120 -47979 89254 -47959
rect 89288 -47959 89304 -47945
rect 89406 -47945 89472 -47909
rect 89506 -47807 89540 -47765
rect 89506 -47875 89540 -47841
rect 89506 -47925 89540 -47909
rect 89574 -47807 89640 -47799
rect 89574 -47841 89590 -47807
rect 89624 -47841 89640 -47807
rect 89574 -47875 89640 -47841
rect 89574 -47909 89590 -47875
rect 89624 -47909 89640 -47875
rect 89406 -47959 89422 -47945
rect 89288 -47979 89422 -47959
rect 89456 -47959 89472 -47945
rect 89574 -47945 89640 -47909
rect 89674 -47807 89708 -47765
rect 89674 -47875 89708 -47841
rect 89674 -47925 89708 -47909
rect 89742 -47807 89808 -47799
rect 89742 -47841 89758 -47807
rect 89792 -47841 89808 -47807
rect 89742 -47875 89808 -47841
rect 89742 -47909 89758 -47875
rect 89792 -47909 89808 -47875
rect 89574 -47959 89590 -47945
rect 89456 -47979 89590 -47959
rect 89624 -47959 89640 -47945
rect 89742 -47945 89808 -47909
rect 89842 -47807 89884 -47765
rect 89876 -47841 89884 -47807
rect 89842 -47875 89884 -47841
rect 89876 -47909 89884 -47875
rect 89842 -47925 89884 -47909
rect 89962 -47807 90004 -47765
rect 89962 -47841 89970 -47807
rect 89962 -47875 90004 -47841
rect 89962 -47909 89970 -47875
rect 89742 -47948 89758 -47945
rect 89792 -47948 89808 -47945
rect 89742 -47959 89754 -47948
rect 89624 -47979 89754 -47959
rect 88566 -47993 89754 -47979
rect 88467 -48034 89555 -48029
rect 88467 -48043 88527 -48034
rect 89388 -48043 89555 -48034
rect 88467 -48077 88492 -48043
rect 88526 -48068 88527 -48043
rect 89388 -48068 89505 -48043
rect 88526 -48077 88666 -48068
rect 88700 -48077 88834 -48068
rect 88868 -48077 89003 -48068
rect 89037 -48077 89170 -48068
rect 89204 -48077 89338 -48068
rect 89372 -48077 89505 -48068
rect 89539 -48077 89555 -48043
rect 89742 -48111 89754 -47993
rect 87094 -48131 88336 -48128
rect 87094 -48165 87110 -48131
rect 87144 -48149 87278 -48131
rect 87144 -48165 87160 -48149
rect 87094 -48199 87160 -48165
rect 87262 -48165 87278 -48149
rect 87312 -48149 87446 -48131
rect 87312 -48165 87328 -48149
rect 87094 -48233 87110 -48199
rect 87144 -48233 87160 -48199
rect 87094 -48241 87160 -48233
rect 87194 -48199 87228 -48183
rect 87194 -48275 87228 -48233
rect 87262 -48199 87328 -48165
rect 87430 -48165 87446 -48149
rect 87480 -48149 87614 -48131
rect 87480 -48165 87496 -48149
rect 87262 -48233 87278 -48199
rect 87312 -48233 87328 -48199
rect 87262 -48241 87328 -48233
rect 87362 -48199 87396 -48183
rect 87362 -48275 87396 -48233
rect 87430 -48199 87496 -48165
rect 87598 -48165 87614 -48149
rect 87648 -48149 87782 -48131
rect 87648 -48165 87664 -48149
rect 87430 -48233 87446 -48199
rect 87480 -48233 87496 -48199
rect 87430 -48241 87496 -48233
rect 87530 -48199 87564 -48183
rect 87530 -48275 87564 -48233
rect 87598 -48199 87664 -48165
rect 87766 -48165 87782 -48149
rect 87816 -48149 87950 -48131
rect 87816 -48165 87832 -48149
rect 87598 -48233 87614 -48199
rect 87648 -48233 87664 -48199
rect 87598 -48241 87664 -48233
rect 87698 -48199 87732 -48183
rect 87698 -48275 87732 -48233
rect 87766 -48199 87832 -48165
rect 87934 -48165 87950 -48149
rect 87984 -48149 88118 -48131
rect 87984 -48165 88000 -48149
rect 87766 -48233 87782 -48199
rect 87816 -48233 87832 -48199
rect 87766 -48241 87832 -48233
rect 87866 -48199 87900 -48183
rect 87866 -48275 87900 -48233
rect 87934 -48199 88000 -48165
rect 88102 -48165 88118 -48149
rect 88152 -48149 88286 -48131
rect 88152 -48165 88168 -48149
rect 87934 -48233 87950 -48199
rect 87984 -48233 88000 -48199
rect 87934 -48241 88000 -48233
rect 88034 -48199 88068 -48183
rect 88034 -48275 88068 -48233
rect 88102 -48199 88168 -48165
rect 88270 -48165 88286 -48149
rect 88320 -48165 88336 -48131
rect 88102 -48233 88118 -48199
rect 88152 -48233 88168 -48199
rect 88102 -48241 88168 -48233
rect 88202 -48199 88236 -48183
rect 88202 -48275 88236 -48233
rect 88270 -48199 88336 -48165
rect 88270 -48233 88286 -48199
rect 88320 -48233 88336 -48199
rect 88270 -48241 88336 -48233
rect 88370 -48131 88412 -48115
rect 88404 -48165 88412 -48131
rect 88370 -48199 88412 -48165
rect 88404 -48233 88412 -48199
rect 88370 -48275 88412 -48233
rect 88486 -48131 88532 -48115
rect 88486 -48165 88498 -48131
rect 88486 -48199 88532 -48165
rect 88486 -48233 88498 -48199
rect 88486 -48275 88532 -48233
rect 88566 -48131 89754 -48111
rect 88566 -48165 88582 -48131
rect 88616 -48149 88750 -48131
rect 88616 -48165 88632 -48149
rect 88566 -48199 88632 -48165
rect 88734 -48165 88750 -48149
rect 88784 -48149 88918 -48131
rect 88784 -48165 88800 -48149
rect 88566 -48233 88582 -48199
rect 88616 -48233 88632 -48199
rect 88566 -48241 88632 -48233
rect 88666 -48199 88700 -48183
rect 88666 -48275 88700 -48233
rect 88734 -48199 88800 -48165
rect 88902 -48165 88918 -48149
rect 88952 -48149 89086 -48131
rect 88952 -48165 88968 -48149
rect 88734 -48233 88750 -48199
rect 88784 -48233 88800 -48199
rect 88734 -48241 88800 -48233
rect 88834 -48199 88868 -48183
rect 88834 -48275 88868 -48233
rect 88902 -48199 88968 -48165
rect 89070 -48165 89086 -48149
rect 89120 -48149 89254 -48131
rect 89120 -48165 89136 -48149
rect 88902 -48233 88918 -48199
rect 88952 -48233 88968 -48199
rect 88902 -48241 88968 -48233
rect 89002 -48199 89036 -48183
rect 89002 -48275 89036 -48233
rect 89070 -48199 89136 -48165
rect 89238 -48165 89254 -48149
rect 89288 -48149 89422 -48131
rect 89288 -48165 89304 -48149
rect 89070 -48233 89086 -48199
rect 89120 -48233 89136 -48199
rect 89070 -48241 89136 -48233
rect 89170 -48199 89204 -48183
rect 89170 -48275 89204 -48233
rect 89238 -48199 89304 -48165
rect 89406 -48165 89422 -48149
rect 89456 -48149 89590 -48131
rect 89456 -48165 89472 -48149
rect 89238 -48233 89254 -48199
rect 89288 -48233 89304 -48199
rect 89238 -48241 89304 -48233
rect 89338 -48199 89372 -48183
rect 89338 -48275 89372 -48233
rect 89406 -48199 89472 -48165
rect 89574 -48165 89590 -48149
rect 89624 -48138 89754 -48131
rect 89804 -48138 89808 -47948
rect 89962 -47945 90004 -47909
rect 89962 -47979 89970 -47945
rect 89962 -47995 90004 -47979
rect 90038 -47807 90104 -47799
rect 90038 -47841 90054 -47807
rect 90088 -47841 90104 -47807
rect 90038 -47875 90104 -47841
rect 90038 -47909 90054 -47875
rect 90088 -47909 90104 -47875
rect 90038 -47945 90104 -47909
rect 90138 -47807 90172 -47765
rect 90138 -47875 90172 -47841
rect 90138 -47925 90172 -47909
rect 90206 -47807 90272 -47799
rect 90206 -47841 90222 -47807
rect 90256 -47841 90272 -47807
rect 90206 -47875 90272 -47841
rect 90206 -47909 90222 -47875
rect 90256 -47909 90272 -47875
rect 90038 -47979 90054 -47945
rect 90088 -47959 90104 -47945
rect 90206 -47945 90272 -47909
rect 90306 -47807 90340 -47765
rect 90306 -47875 90340 -47841
rect 90306 -47925 90340 -47909
rect 90374 -47807 90440 -47799
rect 90374 -47841 90390 -47807
rect 90424 -47841 90440 -47807
rect 90374 -47875 90440 -47841
rect 90374 -47909 90390 -47875
rect 90424 -47909 90440 -47875
rect 90206 -47959 90222 -47945
rect 90088 -47979 90222 -47959
rect 90256 -47959 90272 -47945
rect 90374 -47945 90440 -47909
rect 90474 -47807 90508 -47765
rect 90474 -47875 90508 -47841
rect 90474 -47925 90508 -47909
rect 90542 -47807 90608 -47799
rect 90542 -47841 90558 -47807
rect 90592 -47841 90608 -47807
rect 90542 -47875 90608 -47841
rect 90542 -47909 90558 -47875
rect 90592 -47909 90608 -47875
rect 90374 -47959 90390 -47945
rect 90256 -47979 90390 -47959
rect 90424 -47959 90440 -47945
rect 90542 -47945 90608 -47909
rect 90642 -47807 90676 -47765
rect 90642 -47875 90676 -47841
rect 90642 -47925 90676 -47909
rect 90710 -47807 90776 -47799
rect 90710 -47841 90726 -47807
rect 90760 -47841 90776 -47807
rect 90710 -47875 90776 -47841
rect 90710 -47909 90726 -47875
rect 90760 -47909 90776 -47875
rect 90542 -47959 90558 -47945
rect 90424 -47979 90558 -47959
rect 90592 -47959 90608 -47945
rect 90710 -47945 90776 -47909
rect 90810 -47807 90844 -47765
rect 90810 -47875 90844 -47841
rect 90810 -47925 90844 -47909
rect 90878 -47807 90944 -47799
rect 90878 -47841 90894 -47807
rect 90928 -47841 90944 -47807
rect 90878 -47875 90944 -47841
rect 90878 -47909 90894 -47875
rect 90928 -47909 90944 -47875
rect 90710 -47959 90726 -47945
rect 90592 -47979 90726 -47959
rect 90760 -47959 90776 -47945
rect 90878 -47945 90944 -47909
rect 90978 -47807 91012 -47765
rect 90978 -47875 91012 -47841
rect 90978 -47925 91012 -47909
rect 91046 -47807 91112 -47799
rect 91046 -47841 91062 -47807
rect 91096 -47841 91112 -47807
rect 91046 -47875 91112 -47841
rect 91046 -47909 91062 -47875
rect 91096 -47909 91112 -47875
rect 90878 -47959 90894 -47945
rect 90760 -47979 90894 -47959
rect 90928 -47959 90944 -47945
rect 91046 -47945 91112 -47909
rect 91146 -47807 91180 -47765
rect 91146 -47875 91180 -47841
rect 91146 -47925 91180 -47909
rect 91214 -47807 91280 -47799
rect 91214 -47841 91230 -47807
rect 91264 -47841 91280 -47807
rect 91214 -47875 91280 -47841
rect 91214 -47909 91230 -47875
rect 91264 -47909 91280 -47875
rect 91046 -47959 91062 -47945
rect 90928 -47979 91062 -47959
rect 91096 -47959 91112 -47945
rect 91214 -47945 91280 -47909
rect 91314 -47807 91356 -47765
rect 91348 -47841 91356 -47807
rect 91314 -47875 91356 -47841
rect 91348 -47909 91356 -47875
rect 91314 -47925 91356 -47909
rect 91214 -47948 91230 -47945
rect 91264 -47948 91280 -47945
rect 91214 -47959 91224 -47948
rect 91096 -47979 91224 -47959
rect 90038 -47993 91224 -47979
rect 89939 -48035 91027 -48029
rect 89939 -48037 89984 -48035
rect 90751 -48037 91027 -48035
rect 89939 -48043 89982 -48037
rect 90752 -48043 91027 -48037
rect 89939 -48077 89964 -48043
rect 90752 -48071 90810 -48043
rect 89998 -48077 90138 -48071
rect 90172 -48077 90306 -48071
rect 90340 -48077 90475 -48071
rect 90509 -48077 90642 -48071
rect 90676 -48077 90810 -48071
rect 90844 -48077 90977 -48043
rect 91011 -48077 91027 -48043
rect 91214 -48111 91224 -47993
rect 89624 -48149 89758 -48138
rect 89624 -48165 89640 -48149
rect 89406 -48233 89422 -48199
rect 89456 -48233 89472 -48199
rect 89406 -48241 89472 -48233
rect 89506 -48199 89540 -48183
rect 89506 -48275 89540 -48233
rect 89574 -48199 89640 -48165
rect 89742 -48165 89758 -48149
rect 89792 -48165 89808 -48138
rect 89574 -48233 89590 -48199
rect 89624 -48233 89640 -48199
rect 89574 -48241 89640 -48233
rect 89674 -48199 89708 -48183
rect 89674 -48275 89708 -48233
rect 89742 -48199 89808 -48165
rect 89742 -48233 89758 -48199
rect 89792 -48233 89808 -48199
rect 89742 -48241 89808 -48233
rect 89842 -48131 89884 -48115
rect 89876 -48165 89884 -48131
rect 89842 -48199 89884 -48165
rect 89876 -48233 89884 -48199
rect 89842 -48275 89884 -48233
rect 89958 -48131 90004 -48115
rect 89958 -48165 89970 -48131
rect 89958 -48199 90004 -48165
rect 89958 -48233 89970 -48199
rect 89958 -48275 90004 -48233
rect 90038 -48131 91224 -48111
rect 90038 -48165 90054 -48131
rect 90088 -48149 90222 -48131
rect 90088 -48165 90104 -48149
rect 90038 -48199 90104 -48165
rect 90206 -48165 90222 -48149
rect 90256 -48149 90390 -48131
rect 90256 -48165 90272 -48149
rect 90038 -48233 90054 -48199
rect 90088 -48233 90104 -48199
rect 90038 -48241 90104 -48233
rect 90138 -48199 90172 -48183
rect 90138 -48275 90172 -48233
rect 90206 -48199 90272 -48165
rect 90374 -48165 90390 -48149
rect 90424 -48149 90558 -48131
rect 90424 -48165 90440 -48149
rect 90206 -48233 90222 -48199
rect 90256 -48233 90272 -48199
rect 90206 -48241 90272 -48233
rect 90306 -48199 90340 -48183
rect 90306 -48275 90340 -48233
rect 90374 -48199 90440 -48165
rect 90542 -48165 90558 -48149
rect 90592 -48149 90726 -48131
rect 90592 -48165 90608 -48149
rect 90374 -48233 90390 -48199
rect 90424 -48233 90440 -48199
rect 90374 -48241 90440 -48233
rect 90474 -48199 90508 -48183
rect 90474 -48275 90508 -48233
rect 90542 -48199 90608 -48165
rect 90710 -48165 90726 -48149
rect 90760 -48149 90894 -48131
rect 90760 -48165 90776 -48149
rect 90542 -48233 90558 -48199
rect 90592 -48233 90608 -48199
rect 90542 -48241 90608 -48233
rect 90642 -48199 90676 -48183
rect 90642 -48275 90676 -48233
rect 90710 -48199 90776 -48165
rect 90878 -48165 90894 -48149
rect 90928 -48149 91062 -48131
rect 90928 -48165 90944 -48149
rect 90710 -48233 90726 -48199
rect 90760 -48233 90776 -48199
rect 90710 -48241 90776 -48233
rect 90810 -48199 90844 -48183
rect 90810 -48275 90844 -48233
rect 90878 -48199 90944 -48165
rect 91046 -48165 91062 -48149
rect 91096 -48138 91224 -48131
rect 91274 -48138 91280 -47948
rect 91096 -48149 91230 -48138
rect 91096 -48165 91112 -48149
rect 90878 -48233 90894 -48199
rect 90928 -48233 90944 -48199
rect 90878 -48241 90944 -48233
rect 90978 -48199 91012 -48183
rect 90978 -48275 91012 -48233
rect 91046 -48199 91112 -48165
rect 91214 -48165 91230 -48149
rect 91264 -48165 91280 -48138
rect 91046 -48233 91062 -48199
rect 91096 -48233 91112 -48199
rect 91046 -48241 91112 -48233
rect 91146 -48199 91180 -48183
rect 91146 -48275 91180 -48233
rect 91214 -48199 91280 -48165
rect 91214 -48233 91230 -48199
rect 91264 -48233 91280 -48199
rect 91214 -48241 91280 -48233
rect 91314 -48131 91356 -48115
rect 91348 -48165 91356 -48131
rect 91314 -48199 91356 -48165
rect 91348 -48233 91356 -48199
rect 91314 -48275 91356 -48233
rect 82838 -48309 82867 -48275
rect 82901 -48309 82959 -48275
rect 82993 -48309 83051 -48275
rect 83085 -48309 83143 -48275
rect 83177 -48309 83235 -48275
rect 83269 -48309 83327 -48275
rect 83361 -48309 83419 -48275
rect 83453 -48309 83511 -48275
rect 83545 -48309 83603 -48275
rect 83637 -48309 83695 -48275
rect 83729 -48309 83787 -48275
rect 83821 -48309 83879 -48275
rect 83913 -48309 83971 -48275
rect 84005 -48309 84063 -48275
rect 84097 -48309 84155 -48275
rect 84189 -48309 84247 -48275
rect 84281 -48309 84339 -48275
rect 84373 -48309 84431 -48275
rect 84465 -48309 84523 -48275
rect 84557 -48309 84615 -48275
rect 84649 -48309 84707 -48275
rect 84741 -48309 84799 -48275
rect 84833 -48309 84891 -48275
rect 84925 -48309 84983 -48275
rect 85017 -48309 85075 -48275
rect 85109 -48309 85167 -48275
rect 85201 -48309 85259 -48275
rect 85293 -48309 85351 -48275
rect 85385 -48309 85443 -48275
rect 85477 -48309 85535 -48275
rect 85569 -48309 85627 -48275
rect 85661 -48309 85719 -48275
rect 85753 -48309 85811 -48275
rect 85845 -48309 85903 -48275
rect 85937 -48309 85995 -48275
rect 86029 -48309 86087 -48275
rect 86121 -48309 86179 -48275
rect 86213 -48309 86271 -48275
rect 86305 -48309 86363 -48275
rect 86397 -48309 86455 -48275
rect 86489 -48309 86547 -48275
rect 86581 -48309 86639 -48275
rect 86673 -48309 86731 -48275
rect 86765 -48309 86823 -48275
rect 86857 -48309 86915 -48275
rect 86949 -48309 87007 -48275
rect 87041 -48309 87099 -48275
rect 87133 -48309 87191 -48275
rect 87225 -48309 87283 -48275
rect 87317 -48309 87375 -48275
rect 87409 -48309 87467 -48275
rect 87501 -48309 87559 -48275
rect 87593 -48309 87651 -48275
rect 87685 -48309 87743 -48275
rect 87777 -48309 87835 -48275
rect 87869 -48309 87927 -48275
rect 87961 -48309 88019 -48275
rect 88053 -48309 88111 -48275
rect 88145 -48309 88203 -48275
rect 88237 -48309 88295 -48275
rect 88329 -48309 88387 -48275
rect 88421 -48309 88479 -48275
rect 88513 -48309 88571 -48275
rect 88605 -48309 88663 -48275
rect 88697 -48309 88755 -48275
rect 88789 -48309 88847 -48275
rect 88881 -48309 88939 -48275
rect 88973 -48309 89031 -48275
rect 89065 -48309 89123 -48275
rect 89157 -48309 89215 -48275
rect 89249 -48309 89307 -48275
rect 89341 -48309 89399 -48275
rect 89433 -48309 89491 -48275
rect 89525 -48309 89583 -48275
rect 89617 -48309 89675 -48275
rect 89709 -48309 89767 -48275
rect 89801 -48309 89859 -48275
rect 89893 -48309 89951 -48275
rect 89985 -48309 90043 -48275
rect 90077 -48309 90135 -48275
rect 90169 -48309 90227 -48275
rect 90261 -48309 90319 -48275
rect 90353 -48309 90411 -48275
rect 90445 -48309 90503 -48275
rect 90537 -48309 90595 -48275
rect 90629 -48309 90687 -48275
rect 90721 -48309 90779 -48275
rect 90813 -48309 90871 -48275
rect 90905 -48309 90963 -48275
rect 90997 -48309 91055 -48275
rect 91089 -48309 91147 -48275
rect 91181 -48309 91239 -48275
rect 91273 -48309 91331 -48275
rect 91365 -48309 91394 -48275
rect 77635 -48483 77649 -48449
rect 77683 -48483 77691 -48449
rect 77635 -48499 77691 -48483
rect 77725 -48449 77785 -48433
rect 77725 -48483 77733 -48449
rect 77767 -48483 77785 -48449
rect 35802 -48582 35836 -48520
rect 77725 -48543 77785 -48483
rect 77825 -48441 77841 -48407
rect 77875 -48441 77891 -48407
rect 77825 -48475 77891 -48441
rect 77825 -48509 77841 -48475
rect 77875 -48509 77891 -48475
rect 77929 -48407 78021 -48399
rect 77929 -48441 77945 -48407
rect 77979 -48410 78021 -48407
rect 77979 -48441 78060 -48410
rect 77929 -48475 78060 -48441
rect 77929 -48509 77945 -48475
rect 77979 -48509 78060 -48475
rect 77598 -48560 77651 -48555
rect 25780 -48586 35836 -48582
rect 25780 -48620 25832 -48586
rect 35740 -48620 35836 -48586
rect 35802 -48682 35836 -48620
rect 77410 -48590 77651 -48560
rect 77725 -48577 77913 -48543
rect 77410 -48640 77460 -48590
rect 77510 -48620 77651 -48590
rect 77510 -48640 77740 -48620
rect 77879 -48627 77913 -48577
rect 77971 -48570 78060 -48509
rect 77971 -48610 78000 -48570
rect 78040 -48610 78060 -48570
rect 77410 -48643 77740 -48640
rect 77410 -48670 77652 -48643
rect 77598 -48677 77652 -48670
rect 77686 -48670 77740 -48643
rect 77777 -48630 77845 -48627
rect 77777 -48670 77790 -48630
rect 77830 -48670 77845 -48630
rect 77686 -48677 77733 -48670
rect 77777 -48677 77793 -48670
rect 77827 -48677 77845 -48670
rect 77879 -48643 77937 -48627
rect 77879 -48677 77901 -48643
rect 77935 -48677 77937 -48643
rect 77879 -48693 77937 -48677
rect 77971 -48660 78060 -48610
rect 77879 -48711 77913 -48693
rect 77635 -48749 77913 -48711
rect 77971 -48700 78000 -48660
rect 78040 -48700 78060 -48660
rect 77971 -48740 78060 -48700
rect 77635 -48771 77701 -48749
rect 77635 -48805 77649 -48771
rect 77683 -48805 77701 -48771
rect 77971 -48780 78000 -48740
rect 78040 -48780 78060 -48740
rect 77971 -48783 78060 -48780
rect 77635 -48821 77701 -48805
rect 77825 -48799 77875 -48783
rect 77825 -48833 77841 -48799
rect 77825 -48875 77875 -48833
rect 77909 -48799 78060 -48783
rect 77909 -48833 77925 -48799
rect 77959 -48830 78060 -48799
rect 77959 -48833 78021 -48830
rect 77909 -48841 78021 -48833
rect 77578 -48909 77607 -48875
rect 77641 -48909 77699 -48875
rect 77733 -48909 77791 -48875
rect 77825 -48909 77883 -48875
rect 77917 -48909 77975 -48875
rect 78009 -48909 78038 -48875
rect 77578 -48985 77607 -48951
rect 77641 -48985 77699 -48951
rect 77733 -48985 77791 -48951
rect 77825 -48985 77883 -48951
rect 77917 -48985 77975 -48951
rect 78009 -48985 78067 -48951
rect 78101 -48985 78159 -48951
rect 78193 -48985 78251 -48951
rect 78285 -48985 78343 -48951
rect 78377 -48985 78435 -48951
rect 78469 -48985 78527 -48951
rect 78561 -48985 78590 -48951
rect 77825 -49027 77875 -48985
rect 77635 -49055 77701 -49039
rect 77635 -49089 77649 -49055
rect 77683 -49089 77701 -49055
rect 77825 -49061 77841 -49027
rect 77825 -49077 77875 -49061
rect 77909 -49027 78021 -49019
rect 77909 -49061 77925 -49027
rect 77959 -49061 78021 -49027
rect 77909 -49077 78021 -49061
rect 77635 -49111 77701 -49089
rect 77635 -49149 77913 -49111
rect 77879 -49167 77913 -49149
rect 77879 -49183 77937 -49167
rect 77598 -49190 77652 -49183
rect 77430 -49217 77652 -49190
rect 77686 -49217 77733 -49183
rect 77430 -49220 77733 -49217
rect 77430 -49260 77470 -49220
rect 77510 -49233 77733 -49220
rect 77777 -49190 77793 -49183
rect 77827 -49190 77845 -49183
rect 77777 -49230 77790 -49190
rect 77830 -49230 77845 -49190
rect 77777 -49233 77845 -49230
rect 77879 -49217 77901 -49183
rect 77935 -49217 77937 -49183
rect 77879 -49233 77937 -49217
rect 77510 -49260 77651 -49233
rect 77430 -49300 77651 -49260
rect 77879 -49283 77913 -49233
rect 77598 -49305 77651 -49300
rect 77725 -49317 77913 -49283
rect 77635 -49377 77691 -49361
rect 77635 -49411 77649 -49377
rect 77683 -49411 77691 -49377
rect 77635 -49495 77691 -49411
rect 77725 -49377 77785 -49317
rect 77971 -49351 78021 -49077
rect 78057 -49051 78123 -48985
rect 78057 -49085 78073 -49051
rect 78107 -49085 78123 -49051
rect 78163 -49045 78197 -49029
rect 78237 -49031 78303 -48985
rect 78237 -49065 78253 -49031
rect 78287 -49065 78303 -49031
rect 78337 -49045 78371 -49029
rect 78163 -49099 78197 -49079
rect 78405 -49031 78481 -48985
rect 78405 -49065 78431 -49031
rect 78465 -49065 78481 -49031
rect 78540 -49051 78660 -49050
rect 78337 -49099 78371 -49079
rect 78519 -49069 78660 -49051
rect 78056 -49130 78126 -49119
rect 78056 -49220 78070 -49130
rect 78110 -49220 78126 -49130
rect 78163 -49133 78485 -49099
rect 78553 -49070 78660 -49069
rect 78553 -49103 78570 -49070
rect 78519 -49120 78570 -49103
rect 78451 -49167 78485 -49133
rect 78539 -49140 78570 -49120
rect 78640 -49140 78660 -49070
rect 78056 -49233 78126 -49220
rect 78160 -49180 78302 -49167
rect 77725 -49411 77733 -49377
rect 77767 -49411 77785 -49377
rect 77725 -49427 77785 -49411
rect 77825 -49385 77841 -49351
rect 77875 -49385 77891 -49351
rect 77825 -49419 77891 -49385
rect 77825 -49453 77841 -49419
rect 77875 -49453 77891 -49419
rect 77825 -49495 77891 -49453
rect 77929 -49385 77945 -49351
rect 77979 -49385 78021 -49351
rect 78056 -49288 78120 -49267
rect 78056 -49322 78073 -49288
rect 78107 -49322 78120 -49288
rect 78160 -49270 78190 -49180
rect 78280 -49270 78302 -49180
rect 78336 -49180 78417 -49167
rect 78336 -49220 78360 -49180
rect 78400 -49183 78417 -49180
rect 78409 -49217 78417 -49183
rect 78400 -49220 78417 -49217
rect 78336 -49233 78417 -49220
rect 78451 -49183 78505 -49167
rect 78451 -49217 78471 -49183
rect 78451 -49233 78505 -49217
rect 78539 -49210 78660 -49140
rect 78451 -49267 78485 -49233
rect 78539 -49267 78570 -49210
rect 78160 -49291 78302 -49270
rect 78056 -49325 78120 -49322
rect 78340 -49301 78485 -49267
rect 78519 -49280 78570 -49267
rect 78640 -49280 78660 -49210
rect 78340 -49325 78374 -49301
rect 78056 -49359 78374 -49325
rect 78519 -49320 78660 -49280
rect 78421 -49351 78477 -49335
rect 77929 -49400 78021 -49385
rect 78421 -49385 78434 -49351
rect 78468 -49385 78477 -49351
rect 78056 -49400 78387 -49393
rect 77929 -49407 78387 -49400
rect 77929 -49419 78295 -49407
rect 77929 -49453 77945 -49419
rect 77979 -49441 78295 -49419
rect 78329 -49441 78387 -49407
rect 77979 -49451 78387 -49441
rect 78421 -49419 78477 -49385
rect 77979 -49453 78380 -49451
rect 77929 -49460 78380 -49453
rect 78421 -49453 78434 -49419
rect 78468 -49453 78477 -49419
rect 77929 -49461 78021 -49460
rect 78421 -49495 78477 -49453
rect 78553 -49350 78660 -49320
rect 78553 -49354 78570 -49350
rect 78519 -49388 78570 -49354
rect 78553 -49420 78570 -49388
rect 78640 -49420 78660 -49350
rect 78553 -49422 78660 -49420
rect 78519 -49460 78660 -49422
rect 78519 -49461 78573 -49460
rect 77578 -49529 77607 -49495
rect 77641 -49529 77699 -49495
rect 77733 -49529 77791 -49495
rect 77825 -49529 77883 -49495
rect 77917 -49529 77975 -49495
rect 78009 -49529 78067 -49495
rect 78101 -49529 78159 -49495
rect 78193 -49529 78251 -49495
rect 78285 -49529 78343 -49495
rect 78377 -49529 78435 -49495
rect 78469 -49529 78527 -49495
rect 78561 -49529 78590 -49495
rect 77578 -49605 77607 -49571
rect 77641 -49605 77699 -49571
rect 77733 -49605 77791 -49571
rect 77825 -49605 77883 -49571
rect 77917 -49605 77975 -49571
rect 78009 -49605 78038 -49571
rect 77635 -49689 77691 -49605
rect 77825 -49647 77891 -49605
rect 77635 -49723 77649 -49689
rect 77683 -49723 77691 -49689
rect 77635 -49739 77691 -49723
rect 77725 -49689 77785 -49673
rect 77725 -49723 77733 -49689
rect 77767 -49723 77785 -49689
rect 77725 -49783 77785 -49723
rect 77825 -49681 77841 -49647
rect 77875 -49681 77891 -49647
rect 77825 -49715 77891 -49681
rect 77825 -49749 77841 -49715
rect 77875 -49749 77891 -49715
rect 77929 -49647 78021 -49639
rect 77929 -49681 77945 -49647
rect 77979 -49681 78021 -49647
rect 77929 -49715 78021 -49681
rect 77929 -49749 77945 -49715
rect 77979 -49749 78021 -49715
rect 77971 -49780 78021 -49749
rect 77598 -49800 77651 -49795
rect 77470 -49830 77690 -49800
rect 77725 -49817 77913 -49783
rect 77470 -49880 77510 -49830
rect 77560 -49867 77690 -49830
rect 77879 -49867 77913 -49817
rect 77971 -49820 77980 -49780
rect 78020 -49820 78021 -49780
rect 77560 -49880 77733 -49867
rect 77470 -49883 77733 -49880
rect 77470 -49910 77652 -49883
rect 77598 -49917 77652 -49910
rect 77686 -49917 77733 -49883
rect 77777 -49870 77845 -49867
rect 77777 -49910 77790 -49870
rect 77830 -49910 77845 -49870
rect 77777 -49917 77793 -49910
rect 77827 -49917 77845 -49910
rect 77879 -49883 77937 -49867
rect 77879 -49917 77901 -49883
rect 77935 -49917 77937 -49883
rect 77879 -49933 77937 -49917
rect 77971 -49900 78021 -49820
rect 77879 -49951 77913 -49933
rect 77635 -49989 77913 -49951
rect 77971 -49940 77980 -49900
rect 78020 -49940 78021 -49900
rect 77635 -50011 77701 -49989
rect 77635 -50045 77649 -50011
rect 77683 -50045 77701 -50011
rect 77971 -50000 78021 -49940
rect 77971 -50023 77980 -50000
rect 77635 -50061 77701 -50045
rect 77825 -50039 77875 -50023
rect 35802 -50180 35836 -50118
rect 25780 -50214 25832 -50180
rect 35740 -50214 35836 -50180
rect 25780 -50222 35836 -50214
rect 35802 -50284 35836 -50222
rect 53896 -50192 53992 -50158
rect 54966 -50192 55062 -50158
rect 53896 -50254 53930 -50192
rect 55028 -50254 55062 -50192
rect 54075 -50306 54091 -50272
rect 54867 -50306 54883 -50272
rect 53998 -50334 54032 -50318
rect 53998 -50388 54032 -50372
rect 54926 -50334 54960 -50318
rect 54926 -50388 54960 -50372
rect 54075 -50434 54091 -50400
rect 54867 -50434 54883 -50400
rect 53896 -50514 53930 -50452
rect 77825 -50073 77841 -50039
rect 77825 -50115 77875 -50073
rect 77909 -50039 77980 -50023
rect 77909 -50073 77925 -50039
rect 77959 -50040 77980 -50039
rect 78020 -50040 78021 -50000
rect 77959 -50073 78021 -50040
rect 77909 -50081 78021 -50073
rect 77578 -50149 77607 -50115
rect 77641 -50149 77699 -50115
rect 77733 -50149 77791 -50115
rect 77825 -50149 77883 -50115
rect 77917 -50149 77975 -50115
rect 78009 -50149 78038 -50115
rect 77580 -50239 77609 -50205
rect 77643 -50239 77701 -50205
rect 77735 -50239 77793 -50205
rect 77827 -50239 77885 -50205
rect 77919 -50239 77977 -50205
rect 78011 -50239 78040 -50205
rect 77827 -50281 77877 -50239
rect 77637 -50309 77703 -50293
rect 55028 -50514 55062 -50452
rect 77637 -50343 77651 -50309
rect 77685 -50343 77703 -50309
rect 77827 -50315 77843 -50281
rect 77827 -50331 77877 -50315
rect 77911 -50281 78023 -50273
rect 77911 -50315 77927 -50281
rect 77961 -50315 78023 -50281
rect 77911 -50331 78023 -50315
rect 77637 -50365 77703 -50343
rect 77637 -50403 77915 -50365
rect 77881 -50421 77915 -50403
rect 77973 -50380 78023 -50331
rect 77973 -50420 77980 -50380
rect 78020 -50420 78023 -50380
rect 77881 -50437 77939 -50421
rect 77600 -50440 77654 -50437
rect 77440 -50470 77654 -50440
rect 55960 -50508 56040 -50498
rect 53896 -50548 53992 -50514
rect 54966 -50548 55062 -50514
rect 53350 -50638 53790 -50604
rect 53350 -50700 53384 -50638
rect 53510 -50740 53526 -50706
rect 53614 -50740 53630 -50706
rect 35802 -51782 35836 -51720
rect 25780 -51820 35836 -51782
rect 35802 -51882 35836 -51820
rect 53464 -50790 53498 -50774
rect 53464 -51582 53498 -51566
rect 53642 -50790 53676 -50774
rect 53642 -51582 53676 -51566
rect 53756 -51264 53790 -50638
rect 53896 -50610 53930 -50548
rect 55028 -50610 55062 -50548
rect 55710 -50554 56040 -50508
rect 54075 -50662 54091 -50628
rect 54867 -50662 54883 -50628
rect 53998 -50690 54032 -50674
rect 53998 -50744 54032 -50728
rect 54926 -50690 54960 -50674
rect 54926 -50744 54960 -50728
rect 54075 -50790 54091 -50756
rect 54867 -50790 54883 -50756
rect 53896 -50870 53930 -50808
rect 55706 -50588 55802 -50554
rect 56050 -50588 56146 -50554
rect 55706 -50650 55740 -50588
rect 55028 -50870 55062 -50808
rect 53896 -50904 53992 -50870
rect 54966 -50904 55062 -50870
rect 55176 -50700 55272 -50666
rect 55430 -50700 55526 -50666
rect 55176 -50762 55210 -50700
rect 55492 -50762 55526 -50700
rect 55318 -50802 55334 -50768
rect 55368 -50802 55384 -50768
rect 55290 -50852 55324 -50836
rect 55290 -51044 55324 -51028
rect 55378 -50852 55412 -50836
rect 55378 -51044 55412 -51028
rect 55176 -51118 55210 -51056
rect 55492 -51118 55526 -51056
rect 54870 -51152 55272 -51118
rect 55430 -51152 55706 -51118
rect 54870 -51158 55706 -51152
rect 54870 -51264 54904 -51158
rect 53756 -51298 53852 -51264
rect 54808 -51298 54904 -51264
rect 53756 -51360 53790 -51298
rect 54870 -51360 54904 -51298
rect 55126 -51308 55142 -51274
rect 55494 -51308 55510 -51274
rect 53926 -51412 53942 -51378
rect 54718 -51412 54734 -51378
rect 53858 -51440 53892 -51424
rect 53858 -51544 53892 -51528
rect 54768 -51440 54802 -51424
rect 54768 -51544 54802 -51528
rect 53926 -51590 53942 -51556
rect 54718 -51590 54734 -51556
rect 53510 -51650 53526 -51616
rect 53614 -51650 53630 -51616
rect 53756 -51670 53790 -51608
rect 55046 -51360 55080 -51344
rect 55046 -51410 55080 -51394
rect 55556 -51360 55590 -51344
rect 55556 -51410 55590 -51394
rect 55126 -51480 55142 -51446
rect 55494 -51480 55510 -51446
rect 54870 -51638 54904 -51608
rect 55700 -51606 55706 -51158
rect 56112 -50650 56146 -50588
rect 77440 -50520 77490 -50470
rect 77540 -50471 77654 -50470
rect 77688 -50471 77735 -50437
rect 77540 -50487 77735 -50471
rect 77779 -50440 77795 -50437
rect 77829 -50440 77847 -50437
rect 77779 -50480 77790 -50440
rect 77830 -50480 77847 -50440
rect 77779 -50487 77847 -50480
rect 77881 -50471 77903 -50437
rect 77937 -50471 77939 -50437
rect 77881 -50487 77939 -50471
rect 77973 -50460 78023 -50420
rect 77540 -50520 77690 -50487
rect 58930 -50567 59026 -50533
rect 59600 -50567 59696 -50533
rect 77440 -50550 77690 -50520
rect 77881 -50537 77915 -50487
rect 77600 -50559 77653 -50550
rect 58930 -50610 58964 -50567
rect 58926 -50620 58966 -50610
rect 55866 -50690 55882 -50656
rect 55970 -50690 55986 -50656
rect 55820 -50740 55854 -50724
rect 55820 -51532 55854 -51516
rect 55998 -50740 56032 -50724
rect 55998 -51532 56032 -51516
rect 55866 -51600 55882 -51566
rect 55970 -51600 55986 -51566
rect 55700 -51638 55740 -51606
rect 57096 -50679 57125 -50645
rect 57159 -50679 57217 -50645
rect 57251 -50679 57309 -50645
rect 57343 -50679 57372 -50645
rect 57129 -50729 57165 -50713
rect 57129 -50763 57131 -50729
rect 57129 -50797 57165 -50763
rect 57129 -50831 57131 -50797
rect 57201 -50729 57267 -50679
rect 57201 -50763 57217 -50729
rect 57251 -50763 57267 -50729
rect 57201 -50797 57267 -50763
rect 57201 -50831 57217 -50797
rect 57251 -50831 57267 -50797
rect 57301 -50729 57355 -50713
rect 57301 -50763 57303 -50729
rect 57337 -50763 57355 -50729
rect 57301 -50810 57355 -50763
rect 57129 -50865 57165 -50831
rect 57301 -50844 57303 -50810
rect 57337 -50844 57355 -50810
rect 57129 -50899 57264 -50865
rect 57301 -50894 57355 -50844
rect 57230 -50928 57264 -50899
rect 57117 -50944 57185 -50935
rect 57117 -50994 57118 -50944
rect 57178 -50994 57185 -50944
rect 57117 -51009 57185 -50994
rect 57230 -50944 57285 -50928
rect 57230 -50978 57251 -50944
rect 57230 -50994 57285 -50978
rect 57319 -50940 57355 -50894
rect 59662 -50629 59696 -50567
rect 77727 -50571 77915 -50537
rect 77973 -50500 77980 -50460
rect 78020 -50500 78023 -50460
rect 77973 -50560 78023 -50500
rect 59109 -50681 59125 -50647
rect 59501 -50681 59517 -50647
rect 59560 -50701 59594 -50685
rect 59560 -50751 59594 -50735
rect 59109 -50789 59125 -50755
rect 59501 -50789 59517 -50755
rect 59032 -50809 59066 -50793
rect 59032 -50859 59066 -50843
rect 59109 -50897 59125 -50863
rect 59501 -50897 59517 -50863
rect 77637 -50631 77693 -50615
rect 77637 -50665 77651 -50631
rect 77685 -50665 77693 -50631
rect 77637 -50749 77693 -50665
rect 77727 -50631 77787 -50571
rect 77973 -50600 77980 -50560
rect 78020 -50600 78023 -50560
rect 77973 -50605 78023 -50600
rect 77727 -50665 77735 -50631
rect 77769 -50665 77787 -50631
rect 77727 -50681 77787 -50665
rect 77827 -50639 77843 -50605
rect 77877 -50639 77893 -50605
rect 77827 -50673 77893 -50639
rect 77827 -50707 77843 -50673
rect 77877 -50707 77893 -50673
rect 77827 -50749 77893 -50707
rect 77931 -50639 77947 -50605
rect 77981 -50639 78023 -50605
rect 77931 -50640 78023 -50639
rect 77931 -50673 77980 -50640
rect 77931 -50707 77947 -50673
rect 78020 -50680 78023 -50640
rect 77981 -50707 78023 -50680
rect 77931 -50715 78023 -50707
rect 77580 -50783 77609 -50749
rect 77643 -50783 77701 -50749
rect 77735 -50783 77793 -50749
rect 77827 -50783 77885 -50749
rect 77919 -50783 77977 -50749
rect 78011 -50783 78040 -50749
rect 77578 -50855 77607 -50821
rect 77641 -50855 77699 -50821
rect 77733 -50855 77791 -50821
rect 77825 -50855 77883 -50821
rect 77917 -50855 77975 -50821
rect 78009 -50855 78067 -50821
rect 78101 -50855 78159 -50821
rect 78193 -50855 78222 -50821
rect 78322 -50855 78351 -50821
rect 78385 -50855 78443 -50821
rect 78477 -50855 78535 -50821
rect 78569 -50855 78627 -50821
rect 78661 -50855 78719 -50821
rect 78753 -50855 78811 -50821
rect 78845 -50855 78874 -50821
rect 58926 -50940 58966 -50920
rect 57319 -50980 57326 -50940
rect 58930 -50976 58964 -50940
rect 57230 -51045 57264 -50994
rect 57131 -51079 57264 -51045
rect 57319 -51054 57355 -50980
rect 57131 -51100 57165 -51079
rect 56316 -51118 56412 -51104
rect 54830 -51648 55830 -51638
rect 54830 -51670 55030 -51648
rect 53756 -51704 53852 -51670
rect 54808 -51704 55030 -51670
rect 53510 -51758 53526 -51724
rect 53614 -51758 53630 -51724
rect 53756 -51766 53790 -51704
rect 54830 -51728 55030 -51704
rect 55110 -51668 55740 -51648
rect 55810 -51668 55830 -51648
rect 56112 -51668 56146 -51606
rect 55110 -51708 55160 -51668
rect 55600 -51708 55740 -51668
rect 56050 -51702 56146 -51668
rect 55110 -51728 55740 -51708
rect 55810 -51728 55830 -51702
rect 54830 -51738 55830 -51728
rect 53464 -51808 53498 -51792
rect 53464 -52600 53498 -52584
rect 53642 -51808 53676 -51792
rect 53642 -52600 53676 -52584
rect 54870 -51766 54904 -51738
rect 53926 -51818 53942 -51784
rect 54718 -51818 54734 -51784
rect 53858 -51846 53892 -51830
rect 53858 -51950 53892 -51934
rect 54768 -51846 54802 -51830
rect 54768 -51950 54802 -51934
rect 53926 -51996 53942 -51962
rect 54718 -51996 54734 -51962
rect 53756 -52076 53790 -52014
rect 55700 -51764 55740 -51738
rect 55126 -51930 55142 -51896
rect 55494 -51930 55510 -51896
rect 54870 -52076 54904 -52014
rect 55046 -51982 55080 -51966
rect 55046 -52032 55080 -52016
rect 55556 -51982 55590 -51966
rect 55556 -52032 55590 -52016
rect 53756 -52110 53852 -52076
rect 54808 -52110 54904 -52076
rect 55126 -52102 55142 -52068
rect 55494 -52102 55510 -52068
rect 53510 -52668 53526 -52634
rect 53614 -52668 53630 -52634
rect 53350 -52736 53384 -52674
rect 53756 -52736 53790 -52110
rect 54870 -52218 54904 -52110
rect 55700 -52218 55706 -51764
rect 54870 -52224 55706 -52218
rect 54870 -52258 55262 -52224
rect 55420 -52258 55706 -52224
rect 55166 -52320 55200 -52258
rect 53350 -52770 53446 -52736
rect 53694 -52770 53790 -52736
rect 53886 -52508 53982 -52474
rect 54956 -52508 55052 -52474
rect 53886 -52570 53920 -52508
rect 55018 -52570 55052 -52508
rect 54065 -52622 54081 -52588
rect 54857 -52622 54873 -52588
rect 53988 -52650 54022 -52634
rect 53988 -52704 54022 -52688
rect 54916 -52650 54950 -52634
rect 54916 -52704 54950 -52688
rect 54065 -52750 54081 -52716
rect 54857 -52750 54873 -52716
rect 53886 -52830 53920 -52768
rect 55482 -52320 55516 -52258
rect 55280 -52348 55314 -52332
rect 55280 -52540 55314 -52524
rect 55368 -52348 55402 -52332
rect 55368 -52540 55402 -52524
rect 55308 -52608 55324 -52574
rect 55358 -52608 55374 -52574
rect 55166 -52676 55200 -52614
rect 55482 -52676 55516 -52614
rect 55166 -52710 55262 -52676
rect 55420 -52710 55516 -52676
rect 55018 -52830 55052 -52768
rect 56112 -51764 56146 -51702
rect 56350 -51138 56412 -51118
rect 56610 -51138 56706 -51104
rect 56672 -51200 56706 -51138
rect 57303 -51083 57355 -51054
rect 57131 -51155 57165 -51134
rect 57201 -51147 57217 -51113
rect 57251 -51147 57267 -51113
rect 57201 -51189 57267 -51147
rect 57337 -51117 57355 -51083
rect 57303 -51155 57355 -51117
rect 58930 -51010 59026 -50976
rect 59214 -50977 59310 -50976
rect 59662 -50977 59696 -50920
rect 59772 -50894 59866 -50860
rect 60426 -50894 60520 -50860
rect 59772 -50950 59806 -50894
rect 59214 -51010 59696 -50977
rect 58930 -51011 59696 -51010
rect 58930 -51072 58964 -51011
rect 59276 -51072 59310 -51011
rect 59087 -51112 59103 -51078
rect 59137 -51112 59153 -51078
rect 56476 -51240 56492 -51206
rect 56530 -51240 56546 -51206
rect 55866 -51804 55882 -51770
rect 55970 -51804 55986 -51770
rect 55820 -51854 55854 -51838
rect 55820 -52646 55854 -52630
rect 55998 -51854 56032 -51838
rect 55998 -52646 56032 -52630
rect 55866 -52714 55882 -52680
rect 55970 -52714 55986 -52680
rect 55706 -52782 55740 -52720
rect 56430 -51299 56464 -51283
rect 56430 -52091 56464 -52075
rect 56558 -51299 56592 -51283
rect 56558 -52091 56592 -52075
rect 56476 -52168 56492 -52134
rect 56530 -52168 56546 -52134
rect 56316 -52236 56350 -52174
rect 57096 -51223 57125 -51189
rect 57159 -51223 57217 -51189
rect 57251 -51223 57309 -51189
rect 57343 -51223 57372 -51189
rect 59044 -51171 59078 -51155
rect 59044 -51563 59078 -51547
rect 59162 -51171 59196 -51155
rect 59162 -51563 59196 -51547
rect 59087 -51640 59103 -51606
rect 59137 -51640 59153 -51606
rect 60486 -50956 60520 -50894
rect 77596 -50897 77663 -50855
rect 77596 -50931 77613 -50897
rect 77647 -50931 77663 -50897
rect 77697 -50905 77747 -50889
rect 59942 -51008 59958 -50974
rect 60334 -51008 60350 -50974
rect 59874 -51028 59908 -51012
rect 59874 -51078 59908 -51062
rect 60384 -51028 60418 -51012
rect 60384 -51078 60418 -51062
rect 59942 -51116 59958 -51082
rect 60334 -51116 60350 -51082
rect 59772 -51196 59806 -51140
rect 77697 -50939 77705 -50905
rect 77739 -50939 77747 -50905
rect 77595 -50970 77643 -50967
rect 60486 -51196 60520 -51134
rect 59388 -51230 59476 -51196
rect 59656 -51230 59800 -51196
rect 59958 -51230 60520 -51196
rect 77570 -50980 77643 -50970
rect 77570 -51030 77580 -50980
rect 77630 -51030 77643 -50980
rect 77570 -51133 77643 -51030
rect 77697 -51049 77747 -50939
rect 77791 -50897 77857 -50855
rect 77791 -50931 77807 -50897
rect 77841 -50931 77857 -50897
rect 77791 -50999 77857 -50931
rect 77894 -50905 77944 -50889
rect 77894 -50939 77902 -50905
rect 77936 -50939 77944 -50905
rect 77894 -51049 77944 -50939
rect 78037 -50897 78103 -50855
rect 78037 -50931 78053 -50897
rect 78087 -50931 78103 -50897
rect 78037 -50965 78103 -50931
rect 78137 -50897 78205 -50889
rect 78137 -50931 78153 -50897
rect 78187 -50931 78205 -50897
rect 78137 -50941 78205 -50931
rect 78037 -50999 78053 -50965
rect 78087 -50999 78103 -50965
rect 78037 -51015 78103 -50999
rect 78153 -50965 78205 -50941
rect 78187 -50999 78205 -50965
rect 78240 -50899 78340 -50890
rect 78705 -50897 78761 -50855
rect 78240 -50909 78671 -50899
rect 78240 -50929 78579 -50909
rect 78240 -50963 78250 -50929
rect 78290 -50943 78579 -50929
rect 78613 -50943 78671 -50909
rect 78290 -50957 78671 -50943
rect 78705 -50931 78718 -50897
rect 78752 -50931 78761 -50897
rect 78290 -50960 78310 -50957
rect 78290 -50963 78300 -50960
rect 78240 -50990 78300 -50963
rect 78705 -50965 78761 -50931
rect 78153 -51033 78205 -50999
rect 77570 -51167 77609 -51133
rect 77570 -51229 77643 -51167
rect 77677 -51083 78115 -51049
rect 77570 -51230 77640 -51229
rect 59388 -51290 59422 -51230
rect 59276 -51706 59310 -51646
rect 59530 -51332 59546 -51298
rect 59580 -51332 59596 -51298
rect 59502 -51382 59536 -51366
rect 59502 -51574 59536 -51558
rect 59590 -51382 59624 -51366
rect 59590 -51574 59624 -51558
rect 59530 -51642 59546 -51608
rect 59580 -51642 59596 -51608
rect 58966 -51742 59310 -51706
rect 59388 -51709 59422 -51650
rect 59704 -51709 59738 -51230
rect 60020 -51292 60054 -51230
rect 59846 -51332 59862 -51298
rect 59896 -51332 59912 -51298
rect 59818 -51382 59852 -51366
rect 59818 -51574 59852 -51558
rect 59906 -51382 59940 -51366
rect 59906 -51574 59940 -51558
rect 59846 -51642 59862 -51608
rect 59896 -51642 59912 -51608
rect 77677 -51265 77711 -51083
rect 78052 -51117 78115 -51083
rect 78187 -51050 78205 -51033
rect 78340 -51025 78658 -50991
rect 78705 -50999 78718 -50965
rect 78752 -50999 78761 -50965
rect 78705 -51015 78761 -50999
rect 78803 -50890 78857 -50889
rect 78803 -50928 78920 -50890
rect 78837 -50960 78920 -50928
rect 78837 -50962 78850 -50960
rect 78803 -50996 78850 -50962
rect 78340 -51028 78404 -51025
rect 77612 -51281 77711 -51265
rect 77612 -51315 77613 -51281
rect 77647 -51315 77711 -51281
rect 77755 -51130 77825 -51117
rect 77755 -51133 77770 -51130
rect 77755 -51170 77770 -51167
rect 77810 -51170 77825 -51130
rect 77755 -51310 77825 -51170
rect 77861 -51133 77921 -51117
rect 77895 -51160 77921 -51133
rect 77861 -51200 77870 -51167
rect 77910 -51200 77921 -51160
rect 77861 -51240 77921 -51200
rect 77861 -51280 77870 -51240
rect 77910 -51280 77921 -51240
rect 77861 -51311 77921 -51280
rect 77957 -51133 78013 -51117
rect 77991 -51167 78013 -51133
rect 78052 -51133 78118 -51117
rect 78052 -51167 78068 -51133
rect 78102 -51167 78118 -51133
rect 77957 -51250 78013 -51167
rect 77957 -51290 77970 -51250
rect 78010 -51290 78013 -51250
rect 77957 -51311 78013 -51290
rect 78049 -51221 78103 -51205
rect 78153 -51220 78170 -51067
rect 78340 -51062 78357 -51028
rect 78391 -51062 78404 -51028
rect 78624 -51049 78658 -51025
rect 78837 -51010 78850 -50996
rect 78900 -51010 78920 -50960
rect 78837 -51030 78920 -51010
rect 78340 -51083 78404 -51062
rect 78444 -51080 78586 -51059
rect 78153 -51221 78220 -51220
rect 78049 -51255 78054 -51221
rect 78088 -51255 78103 -51221
rect 78049 -51289 78103 -51255
rect 77612 -51331 77711 -51315
rect 78049 -51323 78054 -51289
rect 78088 -51323 78103 -51289
rect 78137 -51255 78153 -51221
rect 78187 -51240 78220 -51221
rect 78340 -51133 78410 -51117
rect 78340 -51167 78357 -51133
rect 78391 -51167 78410 -51133
rect 78340 -51180 78410 -51167
rect 78340 -51220 78350 -51180
rect 78400 -51220 78410 -51180
rect 78444 -51130 78470 -51080
rect 78560 -51130 78586 -51080
rect 78624 -51083 78769 -51049
rect 78803 -51080 78920 -51030
rect 78803 -51083 78850 -51080
rect 78735 -51117 78769 -51083
rect 78444 -51133 78586 -51130
rect 78444 -51167 78483 -51133
rect 78517 -51167 78586 -51133
rect 78444 -51183 78586 -51167
rect 78620 -51130 78701 -51117
rect 78620 -51170 78640 -51130
rect 78690 -51133 78701 -51130
rect 78693 -51167 78701 -51133
rect 78690 -51170 78701 -51167
rect 78620 -51183 78701 -51170
rect 78735 -51133 78789 -51117
rect 78735 -51167 78755 -51133
rect 78735 -51183 78789 -51167
rect 78823 -51130 78850 -51083
rect 78900 -51130 78920 -51080
rect 78735 -51217 78769 -51183
rect 78340 -51231 78410 -51220
rect 78187 -51255 78205 -51240
rect 78137 -51289 78205 -51255
rect 78447 -51251 78769 -51217
rect 78823 -51200 78920 -51130
rect 78823 -51230 78850 -51200
rect 78803 -51247 78850 -51230
rect 78137 -51323 78153 -51289
rect 78187 -51323 78205 -51289
rect 78341 -51299 78357 -51265
rect 78391 -51299 78407 -51265
rect 78049 -51365 78103 -51323
rect 78341 -51365 78407 -51299
rect 78447 -51271 78481 -51251
rect 78621 -51271 78655 -51251
rect 78447 -51321 78481 -51305
rect 78521 -51319 78537 -51285
rect 78571 -51319 78587 -51285
rect 78521 -51365 78587 -51319
rect 78837 -51250 78850 -51247
rect 78900 -51250 78920 -51200
rect 78837 -51281 78920 -51250
rect 78621 -51321 78655 -51305
rect 78689 -51319 78715 -51285
rect 78749 -51319 78765 -51285
rect 78803 -51299 78920 -51281
rect 78830 -51300 78920 -51299
rect 78689 -51365 78765 -51319
rect 61186 -51400 61286 -51390
rect 77578 -51399 77607 -51365
rect 77641 -51399 77699 -51365
rect 77733 -51399 77791 -51365
rect 77825 -51399 77883 -51365
rect 77917 -51399 77975 -51365
rect 78009 -51399 78067 -51365
rect 78101 -51399 78159 -51365
rect 78193 -51399 78222 -51365
rect 78322 -51399 78351 -51365
rect 78385 -51399 78443 -51365
rect 78477 -51399 78535 -51365
rect 78569 -51399 78627 -51365
rect 78661 -51399 78719 -51365
rect 78753 -51399 78811 -51365
rect 78845 -51399 78874 -51365
rect 61186 -51480 61196 -51400
rect 82838 -51415 82867 -51381
rect 82901 -51415 82959 -51381
rect 82993 -51415 83051 -51381
rect 83085 -51415 83143 -51381
rect 83177 -51415 83235 -51381
rect 83269 -51415 83327 -51381
rect 83361 -51415 83419 -51381
rect 83453 -51415 83511 -51381
rect 83545 -51415 83603 -51381
rect 83637 -51415 83695 -51381
rect 83729 -51415 83787 -51381
rect 83821 -51415 83879 -51381
rect 83913 -51415 83971 -51381
rect 84005 -51415 84063 -51381
rect 84097 -51415 84155 -51381
rect 84189 -51415 84247 -51381
rect 84281 -51415 84339 -51381
rect 84373 -51415 84431 -51381
rect 84465 -51415 84523 -51381
rect 84557 -51415 84615 -51381
rect 84649 -51415 84707 -51381
rect 84741 -51415 84799 -51381
rect 84833 -51415 84891 -51381
rect 84925 -51415 84983 -51381
rect 85017 -51415 85075 -51381
rect 85109 -51415 85167 -51381
rect 85201 -51415 85259 -51381
rect 85293 -51415 85351 -51381
rect 85385 -51415 85443 -51381
rect 85477 -51415 85535 -51381
rect 85569 -51415 85627 -51381
rect 85661 -51415 85719 -51381
rect 85753 -51415 85811 -51381
rect 85845 -51415 85903 -51381
rect 85937 -51415 85995 -51381
rect 86029 -51415 86087 -51381
rect 86121 -51415 86179 -51381
rect 86213 -51415 86271 -51381
rect 86305 -51415 86363 -51381
rect 86397 -51415 86455 -51381
rect 86489 -51415 86547 -51381
rect 86581 -51415 86639 -51381
rect 86673 -51415 86731 -51381
rect 86765 -51415 86823 -51381
rect 86857 -51415 86915 -51381
rect 86949 -51415 87007 -51381
rect 87041 -51415 87099 -51381
rect 87133 -51415 87191 -51381
rect 87225 -51415 87283 -51381
rect 87317 -51415 87375 -51381
rect 87409 -51415 87467 -51381
rect 87501 -51415 87559 -51381
rect 87593 -51415 87651 -51381
rect 87685 -51415 87743 -51381
rect 87777 -51415 87835 -51381
rect 87869 -51415 87927 -51381
rect 87961 -51415 88019 -51381
rect 88053 -51415 88111 -51381
rect 88145 -51415 88203 -51381
rect 88237 -51415 88295 -51381
rect 88329 -51415 88387 -51381
rect 88421 -51415 88479 -51381
rect 88513 -51415 88571 -51381
rect 88605 -51415 88663 -51381
rect 88697 -51415 88755 -51381
rect 88789 -51415 88847 -51381
rect 88881 -51415 88939 -51381
rect 88973 -51415 89031 -51381
rect 89065 -51415 89123 -51381
rect 89157 -51415 89215 -51381
rect 89249 -51415 89307 -51381
rect 89341 -51415 89399 -51381
rect 89433 -51415 89491 -51381
rect 89525 -51415 89583 -51381
rect 89617 -51415 89675 -51381
rect 89709 -51415 89767 -51381
rect 89801 -51415 89859 -51381
rect 89893 -51415 89951 -51381
rect 89985 -51415 90043 -51381
rect 90077 -51415 90135 -51381
rect 90169 -51415 90227 -51381
rect 90261 -51415 90319 -51381
rect 90353 -51415 90411 -51381
rect 90445 -51415 90503 -51381
rect 90537 -51415 90595 -51381
rect 90629 -51415 90687 -51381
rect 90721 -51415 90779 -51381
rect 90813 -51415 90871 -51381
rect 90905 -51415 90963 -51381
rect 90997 -51415 91055 -51381
rect 91089 -51415 91147 -51381
rect 91181 -51415 91239 -51381
rect 91273 -51415 91331 -51381
rect 91365 -51415 91394 -51381
rect 61186 -51490 61286 -51480
rect 77578 -51471 77607 -51437
rect 77641 -51471 77699 -51437
rect 77733 -51471 77791 -51437
rect 77825 -51471 77883 -51437
rect 77917 -51471 77975 -51437
rect 78009 -51471 78067 -51437
rect 78101 -51471 78159 -51437
rect 78193 -51471 78222 -51437
rect 60020 -51709 60054 -51648
rect 56672 -52236 56706 -52174
rect 57096 -52199 57125 -52165
rect 57159 -52199 57217 -52165
rect 57251 -52199 57309 -52165
rect 57343 -52199 57372 -52165
rect 56316 -52270 56412 -52236
rect 56610 -52270 56706 -52236
rect 57131 -52254 57165 -52233
rect 57201 -52241 57267 -52199
rect 57201 -52275 57217 -52241
rect 57251 -52275 57267 -52241
rect 57303 -52271 57355 -52233
rect 57131 -52309 57165 -52288
rect 57337 -52305 57355 -52271
rect 59276 -51802 59310 -51742
rect 59387 -51744 60054 -51709
rect 60127 -51554 60161 -51528
rect 60127 -51557 60253 -51554
rect 60161 -51573 60253 -51557
rect 60161 -51591 60203 -51573
rect 60127 -51607 60203 -51591
rect 60237 -51607 60253 -51573
rect 60359 -51560 60409 -51549
rect 60671 -51554 60705 -51528
rect 60359 -51565 60366 -51560
rect 60359 -51600 60366 -51599
rect 60406 -51600 60409 -51560
rect 60127 -51649 60161 -51607
rect 60127 -51741 60161 -51683
rect 60195 -51657 60325 -51641
rect 60195 -51691 60211 -51657
rect 60245 -51691 60325 -51657
rect 60195 -51707 60325 -51691
rect 59387 -51800 59421 -51744
rect 59087 -51842 59103 -51808
rect 59137 -51842 59153 -51808
rect 59044 -51901 59078 -51885
rect 57131 -52343 57264 -52309
rect 57303 -52334 57355 -52305
rect 57117 -52394 57185 -52379
rect 57117 -52444 57118 -52394
rect 57168 -52444 57185 -52394
rect 57117 -52453 57185 -52444
rect 57230 -52394 57264 -52343
rect 57319 -52370 57355 -52334
rect 57230 -52410 57285 -52394
rect 57230 -52444 57251 -52410
rect 57230 -52460 57285 -52444
rect 57319 -52410 57326 -52370
rect 59044 -52293 59078 -52277
rect 59162 -51901 59196 -51885
rect 59162 -52293 59196 -52277
rect 59087 -52370 59103 -52336
rect 59137 -52370 59153 -52336
rect 57230 -52489 57264 -52460
rect 57129 -52523 57264 -52489
rect 57319 -52494 57355 -52410
rect 57129 -52557 57165 -52523
rect 57301 -52544 57355 -52494
rect 58930 -52438 58964 -52376
rect 59529 -51845 59545 -51811
rect 59579 -51845 59595 -51811
rect 59501 -51895 59535 -51879
rect 59501 -52087 59535 -52071
rect 59589 -51895 59623 -51879
rect 59589 -52087 59623 -52071
rect 59529 -52155 59545 -52121
rect 59579 -52155 59595 -52121
rect 59387 -52223 59421 -52170
rect 59703 -52223 59737 -51744
rect 60019 -51805 60053 -51744
rect 59845 -51845 59861 -51811
rect 59895 -51845 59911 -51811
rect 59817 -51895 59851 -51879
rect 59817 -52087 59851 -52071
rect 59905 -51895 59939 -51879
rect 59905 -52087 59939 -52071
rect 59845 -52155 59861 -52121
rect 59895 -52155 59911 -52121
rect 60161 -51775 60203 -51741
rect 60237 -51775 60253 -51741
rect 60127 -51833 60161 -51775
rect 60289 -51809 60325 -51707
rect 60127 -51909 60161 -51867
rect 60195 -51825 60325 -51809
rect 60195 -51859 60211 -51825
rect 60245 -51859 60325 -51825
rect 60195 -51875 60325 -51859
rect 60359 -51650 60409 -51600
rect 60443 -51557 60705 -51554
rect 60443 -51573 60671 -51557
rect 60443 -51607 60459 -51573
rect 60493 -51607 60527 -51573
rect 60561 -51607 60595 -51573
rect 60629 -51591 60671 -51573
rect 60629 -51607 60705 -51591
rect 60359 -51657 60366 -51650
rect 60406 -51690 60409 -51650
rect 60393 -51691 60409 -51690
rect 60359 -51740 60409 -51691
rect 60359 -51741 60366 -51740
rect 60359 -51780 60366 -51775
rect 60406 -51780 60409 -51740
rect 60359 -51820 60409 -51780
rect 60359 -51825 60366 -51820
rect 60359 -51860 60366 -51859
rect 60406 -51860 60409 -51820
rect 60359 -51875 60409 -51860
rect 60443 -51657 60637 -51641
rect 60443 -51691 60459 -51657
rect 60493 -51691 60527 -51657
rect 60561 -51691 60595 -51657
rect 60629 -51691 60637 -51657
rect 60443 -51707 60637 -51691
rect 60671 -51649 60705 -51607
rect 60443 -51809 60477 -51707
rect 60671 -51741 60705 -51683
rect 60511 -51775 60527 -51741
rect 60561 -51775 60595 -51741
rect 60629 -51775 60671 -51741
rect 60443 -51825 60637 -51809
rect 60443 -51859 60459 -51825
rect 60493 -51859 60527 -51825
rect 60561 -51859 60595 -51825
rect 60629 -51859 60637 -51825
rect 60443 -51875 60637 -51859
rect 60671 -51833 60705 -51775
rect 60289 -51909 60325 -51875
rect 60443 -51909 60481 -51875
rect 60671 -51909 60705 -51867
rect 60127 -51925 60204 -51909
rect 60161 -51943 60204 -51925
rect 60238 -51943 60254 -51909
rect 60161 -51959 60254 -51943
rect 60289 -51925 60481 -51909
rect 60289 -51959 60297 -51925
rect 60331 -51959 60369 -51925
rect 60405 -51959 60449 -51925
rect 60579 -51943 60595 -51909
rect 60629 -51925 60705 -51909
rect 60629 -51943 60671 -51925
rect 60579 -51951 60671 -51943
rect 60127 -51988 60161 -51959
rect 60289 -51962 60481 -51959
rect 60671 -51988 60705 -51959
rect 60747 -51554 60781 -51528
rect 60747 -51557 61009 -51554
rect 60781 -51573 61009 -51557
rect 60781 -51591 60823 -51573
rect 60747 -51607 60823 -51591
rect 60857 -51607 60891 -51573
rect 60925 -51607 60959 -51573
rect 60993 -51607 61009 -51573
rect 61043 -51560 61093 -51549
rect 61291 -51554 61325 -51528
rect 77612 -51521 77711 -51505
rect 61043 -51600 61046 -51560
rect 61086 -51565 61093 -51560
rect 61086 -51600 61093 -51599
rect 60747 -51649 60781 -51607
rect 60747 -51741 60781 -51683
rect 60815 -51657 61009 -51641
rect 60815 -51691 60823 -51657
rect 60857 -51691 60891 -51657
rect 60925 -51691 60959 -51657
rect 60993 -51691 61009 -51657
rect 60815 -51707 61009 -51691
rect 60781 -51775 60823 -51741
rect 60857 -51775 60891 -51741
rect 60925 -51775 60941 -51741
rect 60747 -51833 60781 -51775
rect 60975 -51809 61009 -51707
rect 60747 -51909 60781 -51867
rect 60815 -51825 61009 -51809
rect 60815 -51859 60823 -51825
rect 60857 -51859 60891 -51825
rect 60925 -51859 60959 -51825
rect 60993 -51859 61009 -51825
rect 60815 -51875 61009 -51859
rect 61043 -51650 61093 -51600
rect 61199 -51557 61325 -51554
rect 61199 -51573 61291 -51557
rect 61199 -51607 61215 -51573
rect 61249 -51591 61291 -51573
rect 77612 -51555 77613 -51521
rect 77647 -51555 77711 -51521
rect 78049 -51513 78103 -51471
rect 83067 -51473 83133 -51415
rect 83067 -51507 83083 -51473
rect 83117 -51507 83133 -51473
rect 77612 -51571 77711 -51555
rect 61249 -51607 61325 -51591
rect 61043 -51690 61046 -51650
rect 61086 -51657 61093 -51650
rect 61043 -51691 61059 -51690
rect 61043 -51740 61093 -51691
rect 61043 -51780 61046 -51740
rect 61086 -51741 61093 -51740
rect 61086 -51780 61093 -51775
rect 61043 -51820 61093 -51780
rect 61043 -51860 61046 -51820
rect 61086 -51825 61093 -51820
rect 61086 -51860 61093 -51859
rect 61043 -51875 61093 -51860
rect 61127 -51657 61257 -51641
rect 61127 -51691 61207 -51657
rect 61241 -51691 61257 -51657
rect 61127 -51707 61257 -51691
rect 61291 -51649 61325 -51607
rect 61127 -51809 61163 -51707
rect 61291 -51741 61325 -51683
rect 77595 -51669 77643 -51607
rect 77595 -51703 77609 -51669
rect 77595 -51740 77643 -51703
rect 61199 -51775 61215 -51741
rect 61249 -51775 61291 -51741
rect 61127 -51825 61257 -51809
rect 61127 -51859 61207 -51825
rect 61241 -51859 61257 -51825
rect 61127 -51875 61257 -51859
rect 61291 -51833 61325 -51775
rect 60971 -51909 61009 -51875
rect 61127 -51909 61163 -51875
rect 61291 -51909 61325 -51867
rect 77420 -51810 77643 -51740
rect 77677 -51753 77711 -51571
rect 77755 -51560 77825 -51526
rect 77755 -51600 77770 -51560
rect 77810 -51600 77825 -51560
rect 77755 -51650 77825 -51600
rect 77755 -51669 77770 -51650
rect 77810 -51690 77825 -51650
rect 77789 -51703 77825 -51690
rect 77755 -51719 77825 -51703
rect 77861 -51580 77921 -51525
rect 77861 -51620 77870 -51580
rect 77910 -51620 77921 -51580
rect 77861 -51660 77921 -51620
rect 77861 -51669 77870 -51660
rect 77910 -51700 77921 -51660
rect 77895 -51703 77921 -51700
rect 77861 -51719 77921 -51703
rect 77957 -51669 78013 -51525
rect 78049 -51547 78054 -51513
rect 78088 -51547 78103 -51513
rect 78049 -51581 78103 -51547
rect 78049 -51615 78054 -51581
rect 78088 -51615 78103 -51581
rect 78137 -51547 78153 -51513
rect 78187 -51530 78205 -51513
rect 78187 -51547 78300 -51530
rect 78137 -51550 78300 -51547
rect 78137 -51581 78200 -51550
rect 78137 -51615 78153 -51581
rect 78187 -51600 78200 -51581
rect 78280 -51600 78300 -51550
rect 83067 -51541 83133 -51507
rect 78187 -51615 78300 -51600
rect 78049 -51631 78103 -51615
rect 77991 -51670 78013 -51669
rect 77957 -51710 77970 -51703
rect 78010 -51710 78013 -51670
rect 77957 -51719 78013 -51710
rect 78052 -51703 78068 -51669
rect 78102 -51703 78118 -51669
rect 78052 -51719 78118 -51703
rect 78153 -51690 78300 -51615
rect 82892 -51593 82970 -51574
rect 83067 -51575 83083 -51541
rect 83117 -51575 83133 -51541
rect 83167 -51457 83274 -51449
rect 83167 -51491 83183 -51457
rect 83217 -51491 83274 -51457
rect 83167 -51525 83274 -51491
rect 83167 -51559 83183 -51525
rect 83217 -51559 83274 -51525
rect 83167 -51573 83274 -51559
rect 82892 -51627 82914 -51593
rect 82948 -51609 82970 -51593
rect 82948 -51627 83177 -51609
rect 82892 -51643 83177 -51627
rect 78052 -51753 78115 -51719
rect 77677 -51787 78115 -51753
rect 78153 -51740 78200 -51690
rect 78280 -51740 78300 -51690
rect 78153 -51769 78300 -51740
rect 77420 -51860 77440 -51810
rect 77490 -51860 77643 -51810
rect 77420 -51880 77530 -51860
rect 77595 -51869 77643 -51860
rect 77697 -51897 77747 -51787
rect 60747 -51925 60823 -51909
rect 60781 -51943 60823 -51925
rect 60857 -51943 60873 -51909
rect 60781 -51951 60873 -51943
rect 60971 -51924 61163 -51909
rect 60971 -51925 61129 -51924
rect 60747 -51988 60781 -51959
rect 60971 -51959 60980 -51925
rect 61015 -51959 61053 -51925
rect 61088 -51958 61129 -51925
rect 61198 -51943 61214 -51909
rect 61248 -51925 61325 -51909
rect 61248 -51943 61291 -51925
rect 61088 -51959 61163 -51958
rect 61198 -51959 61291 -51943
rect 60971 -51962 61163 -51959
rect 61291 -51988 61325 -51959
rect 77596 -51939 77613 -51905
rect 77647 -51939 77663 -51905
rect 77596 -51981 77663 -51939
rect 77697 -51931 77705 -51897
rect 77739 -51931 77747 -51897
rect 77697 -51947 77747 -51931
rect 77791 -51905 77857 -51837
rect 77791 -51939 77807 -51905
rect 77841 -51939 77857 -51905
rect 77791 -51981 77857 -51939
rect 77894 -51897 77944 -51787
rect 78187 -51803 78300 -51769
rect 82867 -51690 82938 -51677
rect 82867 -51780 82870 -51690
rect 82930 -51693 82938 -51690
rect 82930 -51780 82938 -51727
rect 82867 -51789 82938 -51780
rect 77894 -51931 77902 -51897
rect 77936 -51931 77944 -51897
rect 77894 -51947 77944 -51931
rect 78037 -51837 78103 -51821
rect 78037 -51871 78053 -51837
rect 78087 -51871 78103 -51837
rect 78037 -51905 78103 -51871
rect 78153 -51830 78300 -51803
rect 82972 -51823 83006 -51643
rect 83040 -51690 83093 -51677
rect 83090 -51780 83093 -51690
rect 83143 -51693 83177 -51643
rect 83143 -51743 83177 -51727
rect 83211 -51630 83274 -51573
rect 83366 -51457 83408 -51415
rect 83366 -51491 83374 -51457
rect 83366 -51525 83408 -51491
rect 83366 -51559 83374 -51525
rect 83366 -51593 83408 -51559
rect 83366 -51627 83374 -51593
rect 83211 -51680 83320 -51630
rect 83366 -51643 83408 -51627
rect 83442 -51457 83508 -51449
rect 83442 -51491 83458 -51457
rect 83492 -51491 83508 -51457
rect 83442 -51525 83508 -51491
rect 83442 -51559 83458 -51525
rect 83492 -51559 83508 -51525
rect 83442 -51593 83508 -51559
rect 83442 -51627 83458 -51593
rect 83492 -51627 83508 -51593
rect 83442 -51645 83508 -51627
rect 83600 -51457 83653 -51415
rect 83600 -51491 83619 -51457
rect 83600 -51525 83653 -51491
rect 83600 -51559 83619 -51525
rect 83600 -51593 83653 -51559
rect 83600 -51627 83619 -51593
rect 83600 -51643 83653 -51627
rect 83687 -51457 83753 -51449
rect 83687 -51491 83703 -51457
rect 83737 -51491 83753 -51457
rect 83687 -51525 83753 -51491
rect 83687 -51559 83703 -51525
rect 83737 -51559 83753 -51525
rect 83687 -51593 83753 -51559
rect 83787 -51457 83821 -51415
rect 83787 -51525 83821 -51491
rect 83787 -51575 83821 -51559
rect 83855 -51457 83921 -51449
rect 83855 -51491 83871 -51457
rect 83905 -51491 83921 -51457
rect 83855 -51525 83921 -51491
rect 83955 -51457 83997 -51415
rect 83989 -51491 83997 -51457
rect 83955 -51507 83997 -51491
rect 84074 -51457 84116 -51415
rect 84074 -51491 84082 -51457
rect 83855 -51559 83871 -51525
rect 83905 -51559 83921 -51525
rect 83687 -51627 83703 -51593
rect 83737 -51609 83753 -51593
rect 83855 -51593 83921 -51559
rect 83855 -51609 83871 -51593
rect 83737 -51627 83871 -51609
rect 83905 -51605 83921 -51593
rect 84074 -51525 84116 -51491
rect 84074 -51559 84082 -51525
rect 84074 -51595 84116 -51559
rect 83905 -51627 84008 -51605
rect 83687 -51643 84008 -51627
rect 83362 -51680 83428 -51679
rect 83211 -51693 83428 -51680
rect 83211 -51720 83378 -51693
rect 83211 -51760 83320 -51720
rect 83362 -51727 83378 -51720
rect 83412 -51727 83428 -51693
rect 83462 -51680 83508 -51645
rect 83595 -51680 83921 -51677
rect 83462 -51693 83921 -51680
rect 83462 -51727 83611 -51693
rect 83645 -51727 83703 -51693
rect 83737 -51727 83787 -51693
rect 83821 -51727 83871 -51693
rect 83905 -51727 83921 -51693
rect 83955 -51680 84008 -51643
rect 84074 -51629 84082 -51595
rect 84074 -51645 84116 -51629
rect 84150 -51457 84216 -51449
rect 84150 -51491 84166 -51457
rect 84200 -51491 84216 -51457
rect 84150 -51525 84216 -51491
rect 84150 -51559 84166 -51525
rect 84200 -51559 84216 -51525
rect 84150 -51595 84216 -51559
rect 84250 -51457 84284 -51415
rect 84250 -51525 84284 -51491
rect 84250 -51575 84284 -51559
rect 84318 -51457 84384 -51449
rect 84318 -51491 84334 -51457
rect 84368 -51491 84384 -51457
rect 84318 -51525 84384 -51491
rect 84318 -51559 84334 -51525
rect 84368 -51559 84384 -51525
rect 84150 -51629 84166 -51595
rect 84200 -51609 84216 -51595
rect 84318 -51595 84384 -51559
rect 84418 -51457 84452 -51415
rect 84418 -51525 84452 -51491
rect 84418 -51575 84452 -51559
rect 84486 -51457 84552 -51449
rect 84486 -51491 84502 -51457
rect 84536 -51491 84552 -51457
rect 84486 -51525 84552 -51491
rect 84486 -51559 84502 -51525
rect 84536 -51559 84552 -51525
rect 84318 -51609 84334 -51595
rect 84200 -51629 84334 -51609
rect 84368 -51609 84384 -51595
rect 84486 -51595 84552 -51559
rect 84586 -51457 84620 -51415
rect 84586 -51525 84620 -51491
rect 84586 -51575 84620 -51559
rect 84654 -51457 84720 -51449
rect 84654 -51491 84670 -51457
rect 84704 -51491 84720 -51457
rect 84654 -51525 84720 -51491
rect 84654 -51559 84670 -51525
rect 84704 -51559 84720 -51525
rect 84486 -51609 84502 -51595
rect 84368 -51629 84502 -51609
rect 84536 -51609 84552 -51595
rect 84654 -51595 84720 -51559
rect 84754 -51457 84788 -51415
rect 84754 -51525 84788 -51491
rect 84754 -51575 84788 -51559
rect 84822 -51457 84888 -51449
rect 84822 -51491 84838 -51457
rect 84872 -51491 84888 -51457
rect 84822 -51525 84888 -51491
rect 84822 -51559 84838 -51525
rect 84872 -51559 84888 -51525
rect 84654 -51609 84670 -51595
rect 84536 -51629 84670 -51609
rect 84704 -51609 84720 -51595
rect 84822 -51595 84888 -51559
rect 84922 -51457 84956 -51415
rect 84922 -51525 84956 -51491
rect 84922 -51575 84956 -51559
rect 84990 -51457 85056 -51449
rect 84990 -51491 85006 -51457
rect 85040 -51491 85056 -51457
rect 84990 -51525 85056 -51491
rect 84990 -51559 85006 -51525
rect 85040 -51559 85056 -51525
rect 84822 -51609 84838 -51595
rect 84704 -51629 84838 -51609
rect 84872 -51609 84888 -51595
rect 84990 -51595 85056 -51559
rect 85090 -51457 85124 -51415
rect 85090 -51525 85124 -51491
rect 85090 -51575 85124 -51559
rect 85158 -51457 85224 -51449
rect 85158 -51491 85174 -51457
rect 85208 -51491 85224 -51457
rect 85158 -51525 85224 -51491
rect 85158 -51559 85174 -51525
rect 85208 -51559 85224 -51525
rect 84990 -51609 85006 -51595
rect 84872 -51629 85006 -51609
rect 85040 -51609 85056 -51595
rect 85158 -51595 85224 -51559
rect 85258 -51457 85292 -51415
rect 85258 -51525 85292 -51491
rect 85258 -51575 85292 -51559
rect 85326 -51457 85392 -51449
rect 85326 -51491 85342 -51457
rect 85376 -51491 85392 -51457
rect 85326 -51525 85392 -51491
rect 85326 -51559 85342 -51525
rect 85376 -51559 85392 -51525
rect 85158 -51609 85174 -51595
rect 85040 -51629 85174 -51609
rect 85208 -51609 85224 -51595
rect 85326 -51595 85392 -51559
rect 85426 -51457 85468 -51415
rect 85460 -51491 85468 -51457
rect 85426 -51525 85468 -51491
rect 85460 -51559 85468 -51525
rect 85426 -51575 85468 -51559
rect 85546 -51457 85588 -51415
rect 85546 -51491 85554 -51457
rect 85546 -51525 85588 -51491
rect 85546 -51559 85554 -51525
rect 85326 -51609 85342 -51595
rect 85208 -51610 85342 -51609
rect 85376 -51610 85392 -51595
rect 85208 -51629 85330 -51610
rect 84150 -51643 85330 -51629
rect 84051 -51680 85139 -51679
rect 83955 -51693 85139 -51680
rect 83955 -51727 84076 -51693
rect 84110 -51727 84250 -51693
rect 84284 -51727 84418 -51693
rect 84452 -51727 84587 -51693
rect 84621 -51727 84754 -51693
rect 84788 -51727 84922 -51693
rect 84956 -51727 85089 -51693
rect 85123 -51727 85139 -51693
rect 83462 -51730 83660 -51727
rect 83955 -51730 84110 -51727
rect 83211 -51777 83274 -51760
rect 83040 -51789 83093 -51780
rect 83151 -51779 83274 -51777
rect 83151 -51813 83167 -51779
rect 83201 -51813 83274 -51779
rect 78153 -51837 78200 -51830
rect 78187 -51871 78200 -51837
rect 78153 -51880 78200 -51871
rect 78280 -51880 78300 -51830
rect 78153 -51895 78300 -51880
rect 78037 -51939 78053 -51905
rect 78087 -51939 78103 -51905
rect 78037 -51981 78103 -51939
rect 78137 -51905 78300 -51895
rect 78137 -51939 78153 -51905
rect 78187 -51920 78300 -51905
rect 82888 -51839 82936 -51823
rect 82888 -51873 82902 -51839
rect 78187 -51939 78205 -51920
rect 82888 -51925 82936 -51873
rect 82972 -51839 83028 -51823
rect 82972 -51873 82986 -51839
rect 83020 -51873 83028 -51839
rect 82972 -51889 83028 -51873
rect 83074 -51839 83117 -51823
rect 83074 -51873 83082 -51839
rect 83116 -51873 83117 -51839
rect 83074 -51925 83117 -51873
rect 83151 -51847 83274 -51813
rect 83151 -51881 83167 -51847
rect 83201 -51881 83274 -51847
rect 83151 -51891 83274 -51881
rect 83362 -51777 83408 -51761
rect 83462 -51765 83508 -51730
rect 83955 -51761 84008 -51730
rect 85326 -51761 85330 -51643
rect 83362 -51811 83374 -51777
rect 83362 -51845 83408 -51811
rect 83362 -51879 83374 -51845
rect 83362 -51925 83408 -51879
rect 83442 -51777 83508 -51765
rect 83442 -51811 83458 -51777
rect 83492 -51811 83508 -51777
rect 83442 -51845 83508 -51811
rect 83687 -51797 84008 -51761
rect 84070 -51781 84116 -51765
rect 83442 -51879 83458 -51845
rect 83492 -51879 83508 -51845
rect 83442 -51891 83508 -51879
rect 83600 -51849 83653 -51833
rect 83600 -51883 83619 -51849
rect 83600 -51925 83653 -51883
rect 83687 -51841 83753 -51797
rect 83687 -51875 83703 -51841
rect 83737 -51875 83753 -51841
rect 83687 -51891 83753 -51875
rect 83787 -51849 83821 -51833
rect 83787 -51925 83821 -51883
rect 83855 -51841 83921 -51797
rect 84070 -51815 84082 -51781
rect 83855 -51875 83871 -51841
rect 83905 -51875 83921 -51841
rect 83855 -51891 83921 -51875
rect 83955 -51848 84005 -51832
rect 83989 -51882 84005 -51848
rect 83955 -51925 84005 -51882
rect 84070 -51849 84116 -51815
rect 84070 -51883 84082 -51849
rect 84070 -51925 84116 -51883
rect 84150 -51780 85330 -51761
rect 85380 -51780 85392 -51610
rect 85546 -51595 85588 -51559
rect 85546 -51629 85554 -51595
rect 85546 -51645 85588 -51629
rect 85622 -51457 85688 -51449
rect 85622 -51491 85638 -51457
rect 85672 -51491 85688 -51457
rect 85622 -51525 85688 -51491
rect 85622 -51559 85638 -51525
rect 85672 -51559 85688 -51525
rect 85622 -51595 85688 -51559
rect 85722 -51457 85756 -51415
rect 85722 -51525 85756 -51491
rect 85722 -51575 85756 -51559
rect 85790 -51457 85856 -51449
rect 85790 -51491 85806 -51457
rect 85840 -51491 85856 -51457
rect 85790 -51525 85856 -51491
rect 85790 -51559 85806 -51525
rect 85840 -51559 85856 -51525
rect 85622 -51629 85638 -51595
rect 85672 -51609 85688 -51595
rect 85790 -51595 85856 -51559
rect 85890 -51457 85924 -51415
rect 85890 -51525 85924 -51491
rect 85890 -51575 85924 -51559
rect 85958 -51457 86024 -51449
rect 85958 -51491 85974 -51457
rect 86008 -51491 86024 -51457
rect 85958 -51525 86024 -51491
rect 85958 -51559 85974 -51525
rect 86008 -51559 86024 -51525
rect 85790 -51609 85806 -51595
rect 85672 -51629 85806 -51609
rect 85840 -51609 85856 -51595
rect 85958 -51595 86024 -51559
rect 86058 -51457 86092 -51415
rect 86058 -51525 86092 -51491
rect 86058 -51575 86092 -51559
rect 86126 -51457 86192 -51449
rect 86126 -51491 86142 -51457
rect 86176 -51491 86192 -51457
rect 86126 -51525 86192 -51491
rect 86126 -51559 86142 -51525
rect 86176 -51559 86192 -51525
rect 85958 -51609 85974 -51595
rect 85840 -51629 85974 -51609
rect 86008 -51609 86024 -51595
rect 86126 -51595 86192 -51559
rect 86226 -51457 86260 -51415
rect 86226 -51525 86260 -51491
rect 86226 -51575 86260 -51559
rect 86294 -51457 86360 -51449
rect 86294 -51491 86310 -51457
rect 86344 -51491 86360 -51457
rect 86294 -51525 86360 -51491
rect 86294 -51559 86310 -51525
rect 86344 -51559 86360 -51525
rect 86126 -51609 86142 -51595
rect 86008 -51629 86142 -51609
rect 86176 -51609 86192 -51595
rect 86294 -51595 86360 -51559
rect 86394 -51457 86428 -51415
rect 86394 -51525 86428 -51491
rect 86394 -51575 86428 -51559
rect 86462 -51457 86528 -51449
rect 86462 -51491 86478 -51457
rect 86512 -51491 86528 -51457
rect 86462 -51525 86528 -51491
rect 86462 -51559 86478 -51525
rect 86512 -51559 86528 -51525
rect 86294 -51609 86310 -51595
rect 86176 -51629 86310 -51609
rect 86344 -51609 86360 -51595
rect 86462 -51595 86528 -51559
rect 86562 -51457 86596 -51415
rect 86562 -51525 86596 -51491
rect 86562 -51575 86596 -51559
rect 86630 -51457 86696 -51449
rect 86630 -51491 86646 -51457
rect 86680 -51491 86696 -51457
rect 86630 -51525 86696 -51491
rect 86630 -51559 86646 -51525
rect 86680 -51559 86696 -51525
rect 86462 -51609 86478 -51595
rect 86344 -51629 86478 -51609
rect 86512 -51609 86528 -51595
rect 86630 -51595 86696 -51559
rect 86730 -51457 86764 -51415
rect 86730 -51525 86764 -51491
rect 86730 -51575 86764 -51559
rect 86798 -51457 86864 -51449
rect 86798 -51491 86814 -51457
rect 86848 -51491 86864 -51457
rect 86798 -51525 86864 -51491
rect 86798 -51559 86814 -51525
rect 86848 -51559 86864 -51525
rect 86630 -51609 86646 -51595
rect 86512 -51629 86646 -51609
rect 86680 -51609 86696 -51595
rect 86798 -51590 86864 -51559
rect 86898 -51457 86940 -51415
rect 86932 -51491 86940 -51457
rect 86898 -51525 86940 -51491
rect 86932 -51559 86940 -51525
rect 86898 -51575 86940 -51559
rect 87018 -51457 87060 -51415
rect 87018 -51491 87026 -51457
rect 87018 -51525 87060 -51491
rect 87018 -51559 87026 -51525
rect 86798 -51609 86810 -51590
rect 86680 -51629 86810 -51609
rect 85622 -51643 86810 -51629
rect 85523 -51687 86611 -51679
rect 85523 -51693 85610 -51687
rect 86471 -51693 86611 -51687
rect 85523 -51727 85548 -51693
rect 85582 -51721 85610 -51693
rect 86471 -51721 86561 -51693
rect 85582 -51727 85722 -51721
rect 85756 -51727 85890 -51721
rect 85924 -51727 86059 -51721
rect 86093 -51727 86226 -51721
rect 86260 -51727 86394 -51721
rect 86428 -51727 86561 -51721
rect 86595 -51727 86611 -51693
rect 86798 -51761 86810 -51643
rect 84150 -51781 85392 -51780
rect 84150 -51815 84166 -51781
rect 84200 -51799 84334 -51781
rect 84200 -51815 84216 -51799
rect 84150 -51849 84216 -51815
rect 84318 -51815 84334 -51799
rect 84368 -51799 84502 -51781
rect 84368 -51815 84384 -51799
rect 84150 -51883 84166 -51849
rect 84200 -51883 84216 -51849
rect 84150 -51891 84216 -51883
rect 84250 -51849 84284 -51833
rect 84250 -51925 84284 -51883
rect 84318 -51849 84384 -51815
rect 84486 -51815 84502 -51799
rect 84536 -51799 84670 -51781
rect 84536 -51815 84552 -51799
rect 84318 -51883 84334 -51849
rect 84368 -51883 84384 -51849
rect 84318 -51891 84384 -51883
rect 84418 -51849 84452 -51833
rect 84418 -51925 84452 -51883
rect 84486 -51849 84552 -51815
rect 84654 -51815 84670 -51799
rect 84704 -51799 84838 -51781
rect 84704 -51815 84720 -51799
rect 84486 -51883 84502 -51849
rect 84536 -51883 84552 -51849
rect 84486 -51891 84552 -51883
rect 84586 -51849 84620 -51833
rect 84586 -51925 84620 -51883
rect 84654 -51849 84720 -51815
rect 84822 -51815 84838 -51799
rect 84872 -51799 85006 -51781
rect 84872 -51815 84888 -51799
rect 84654 -51883 84670 -51849
rect 84704 -51883 84720 -51849
rect 84654 -51891 84720 -51883
rect 84754 -51849 84788 -51833
rect 84754 -51925 84788 -51883
rect 84822 -51849 84888 -51815
rect 84990 -51815 85006 -51799
rect 85040 -51799 85174 -51781
rect 85040 -51815 85056 -51799
rect 84822 -51883 84838 -51849
rect 84872 -51883 84888 -51849
rect 84822 -51891 84888 -51883
rect 84922 -51849 84956 -51833
rect 84922 -51925 84956 -51883
rect 84990 -51849 85056 -51815
rect 85158 -51815 85174 -51799
rect 85208 -51799 85342 -51781
rect 85208 -51815 85224 -51799
rect 84990 -51883 85006 -51849
rect 85040 -51883 85056 -51849
rect 84990 -51891 85056 -51883
rect 85090 -51849 85124 -51833
rect 85090 -51925 85124 -51883
rect 85158 -51849 85224 -51815
rect 85326 -51815 85342 -51799
rect 85376 -51815 85392 -51781
rect 85158 -51883 85174 -51849
rect 85208 -51883 85224 -51849
rect 85158 -51891 85224 -51883
rect 85258 -51849 85292 -51833
rect 85258 -51925 85292 -51883
rect 85326 -51849 85392 -51815
rect 85326 -51883 85342 -51849
rect 85376 -51883 85392 -51849
rect 85326 -51891 85392 -51883
rect 85426 -51781 85468 -51765
rect 85460 -51815 85468 -51781
rect 85426 -51849 85468 -51815
rect 85460 -51883 85468 -51849
rect 85426 -51925 85468 -51883
rect 85542 -51781 85588 -51765
rect 85542 -51815 85554 -51781
rect 85542 -51849 85588 -51815
rect 85542 -51883 85554 -51849
rect 85542 -51925 85588 -51883
rect 85622 -51780 86810 -51761
rect 86860 -51780 86864 -51590
rect 87018 -51595 87060 -51559
rect 87018 -51629 87026 -51595
rect 87018 -51645 87060 -51629
rect 87094 -51457 87160 -51449
rect 87094 -51491 87110 -51457
rect 87144 -51491 87160 -51457
rect 87094 -51525 87160 -51491
rect 87094 -51559 87110 -51525
rect 87144 -51559 87160 -51525
rect 87094 -51595 87160 -51559
rect 87194 -51457 87228 -51415
rect 87194 -51525 87228 -51491
rect 87194 -51575 87228 -51559
rect 87262 -51457 87328 -51449
rect 87262 -51491 87278 -51457
rect 87312 -51491 87328 -51457
rect 87262 -51525 87328 -51491
rect 87262 -51559 87278 -51525
rect 87312 -51559 87328 -51525
rect 87094 -51629 87110 -51595
rect 87144 -51609 87160 -51595
rect 87262 -51595 87328 -51559
rect 87362 -51457 87396 -51415
rect 87362 -51525 87396 -51491
rect 87362 -51575 87396 -51559
rect 87430 -51457 87496 -51449
rect 87430 -51491 87446 -51457
rect 87480 -51491 87496 -51457
rect 87430 -51525 87496 -51491
rect 87430 -51559 87446 -51525
rect 87480 -51559 87496 -51525
rect 87262 -51609 87278 -51595
rect 87144 -51629 87278 -51609
rect 87312 -51609 87328 -51595
rect 87430 -51595 87496 -51559
rect 87530 -51457 87564 -51415
rect 87530 -51525 87564 -51491
rect 87530 -51575 87564 -51559
rect 87598 -51457 87664 -51449
rect 87598 -51491 87614 -51457
rect 87648 -51491 87664 -51457
rect 87598 -51525 87664 -51491
rect 87598 -51559 87614 -51525
rect 87648 -51559 87664 -51525
rect 87430 -51609 87446 -51595
rect 87312 -51629 87446 -51609
rect 87480 -51609 87496 -51595
rect 87598 -51595 87664 -51559
rect 87698 -51457 87732 -51415
rect 87698 -51525 87732 -51491
rect 87698 -51575 87732 -51559
rect 87766 -51457 87832 -51449
rect 87766 -51491 87782 -51457
rect 87816 -51491 87832 -51457
rect 87766 -51525 87832 -51491
rect 87766 -51559 87782 -51525
rect 87816 -51559 87832 -51525
rect 87598 -51609 87614 -51595
rect 87480 -51629 87614 -51609
rect 87648 -51609 87664 -51595
rect 87766 -51595 87832 -51559
rect 87866 -51457 87900 -51415
rect 87866 -51525 87900 -51491
rect 87866 -51575 87900 -51559
rect 87934 -51457 88000 -51449
rect 87934 -51491 87950 -51457
rect 87984 -51491 88000 -51457
rect 87934 -51525 88000 -51491
rect 87934 -51559 87950 -51525
rect 87984 -51559 88000 -51525
rect 87766 -51609 87782 -51595
rect 87648 -51629 87782 -51609
rect 87816 -51609 87832 -51595
rect 87934 -51595 88000 -51559
rect 88034 -51457 88068 -51415
rect 88034 -51525 88068 -51491
rect 88034 -51575 88068 -51559
rect 88102 -51457 88168 -51449
rect 88102 -51491 88118 -51457
rect 88152 -51491 88168 -51457
rect 88102 -51525 88168 -51491
rect 88102 -51559 88118 -51525
rect 88152 -51559 88168 -51525
rect 87934 -51609 87950 -51595
rect 87816 -51629 87950 -51609
rect 87984 -51609 88000 -51595
rect 88102 -51595 88168 -51559
rect 88202 -51457 88236 -51415
rect 88202 -51525 88236 -51491
rect 88202 -51575 88236 -51559
rect 88270 -51457 88336 -51449
rect 88270 -51491 88286 -51457
rect 88320 -51491 88336 -51457
rect 88270 -51525 88336 -51491
rect 88270 -51559 88286 -51525
rect 88320 -51559 88336 -51525
rect 88102 -51609 88118 -51595
rect 87984 -51629 88118 -51609
rect 88152 -51609 88168 -51595
rect 88270 -51595 88336 -51559
rect 88370 -51457 88412 -51415
rect 88404 -51491 88412 -51457
rect 88370 -51525 88412 -51491
rect 88404 -51559 88412 -51525
rect 88370 -51575 88412 -51559
rect 88490 -51457 88532 -51415
rect 88490 -51491 88498 -51457
rect 88490 -51525 88532 -51491
rect 88490 -51559 88498 -51525
rect 88270 -51600 88286 -51595
rect 88320 -51600 88336 -51595
rect 88270 -51609 88280 -51600
rect 88152 -51629 88280 -51609
rect 87094 -51643 88280 -51629
rect 86995 -51686 88083 -51679
rect 86995 -51693 87044 -51686
rect 87905 -51693 88083 -51686
rect 86995 -51727 87020 -51693
rect 87905 -51720 88033 -51693
rect 87054 -51727 87194 -51720
rect 87228 -51727 87362 -51720
rect 87396 -51727 87531 -51720
rect 87565 -51727 87698 -51720
rect 87732 -51727 87866 -51720
rect 87900 -51727 88033 -51720
rect 88067 -51727 88083 -51693
rect 88270 -51761 88280 -51643
rect 85622 -51781 86864 -51780
rect 85622 -51815 85638 -51781
rect 85672 -51799 85806 -51781
rect 85672 -51815 85688 -51799
rect 85622 -51849 85688 -51815
rect 85790 -51815 85806 -51799
rect 85840 -51799 85974 -51781
rect 85840 -51815 85856 -51799
rect 85622 -51883 85638 -51849
rect 85672 -51883 85688 -51849
rect 85622 -51891 85688 -51883
rect 85722 -51849 85756 -51833
rect 85722 -51925 85756 -51883
rect 85790 -51849 85856 -51815
rect 85958 -51815 85974 -51799
rect 86008 -51799 86142 -51781
rect 86008 -51815 86024 -51799
rect 85790 -51883 85806 -51849
rect 85840 -51883 85856 -51849
rect 85790 -51891 85856 -51883
rect 85890 -51849 85924 -51833
rect 85890 -51925 85924 -51883
rect 85958 -51849 86024 -51815
rect 86126 -51815 86142 -51799
rect 86176 -51799 86310 -51781
rect 86176 -51815 86192 -51799
rect 85958 -51883 85974 -51849
rect 86008 -51883 86024 -51849
rect 85958 -51891 86024 -51883
rect 86058 -51849 86092 -51833
rect 86058 -51925 86092 -51883
rect 86126 -51849 86192 -51815
rect 86294 -51815 86310 -51799
rect 86344 -51799 86478 -51781
rect 86344 -51815 86360 -51799
rect 86126 -51883 86142 -51849
rect 86176 -51883 86192 -51849
rect 86126 -51891 86192 -51883
rect 86226 -51849 86260 -51833
rect 86226 -51925 86260 -51883
rect 86294 -51849 86360 -51815
rect 86462 -51815 86478 -51799
rect 86512 -51799 86646 -51781
rect 86512 -51815 86528 -51799
rect 86294 -51883 86310 -51849
rect 86344 -51883 86360 -51849
rect 86294 -51891 86360 -51883
rect 86394 -51849 86428 -51833
rect 86394 -51925 86428 -51883
rect 86462 -51849 86528 -51815
rect 86630 -51815 86646 -51799
rect 86680 -51799 86814 -51781
rect 86680 -51815 86696 -51799
rect 86462 -51883 86478 -51849
rect 86512 -51883 86528 -51849
rect 86462 -51891 86528 -51883
rect 86562 -51849 86596 -51833
rect 86562 -51925 86596 -51883
rect 86630 -51849 86696 -51815
rect 86798 -51815 86814 -51799
rect 86848 -51815 86864 -51781
rect 86630 -51883 86646 -51849
rect 86680 -51883 86696 -51849
rect 86630 -51891 86696 -51883
rect 86730 -51849 86764 -51833
rect 86730 -51925 86764 -51883
rect 86798 -51849 86864 -51815
rect 86798 -51883 86814 -51849
rect 86848 -51883 86864 -51849
rect 86798 -51891 86864 -51883
rect 86898 -51781 86940 -51765
rect 86932 -51815 86940 -51781
rect 86898 -51849 86940 -51815
rect 86932 -51883 86940 -51849
rect 86898 -51925 86940 -51883
rect 87014 -51781 87060 -51765
rect 87014 -51815 87026 -51781
rect 87014 -51849 87060 -51815
rect 87014 -51883 87026 -51849
rect 87014 -51925 87060 -51883
rect 87094 -51780 88280 -51761
rect 88330 -51780 88336 -51600
rect 88490 -51595 88532 -51559
rect 88490 -51629 88498 -51595
rect 88490 -51645 88532 -51629
rect 88566 -51457 88632 -51449
rect 88566 -51491 88582 -51457
rect 88616 -51491 88632 -51457
rect 88566 -51525 88632 -51491
rect 88566 -51559 88582 -51525
rect 88616 -51559 88632 -51525
rect 88566 -51595 88632 -51559
rect 88666 -51457 88700 -51415
rect 88666 -51525 88700 -51491
rect 88666 -51575 88700 -51559
rect 88734 -51457 88800 -51449
rect 88734 -51491 88750 -51457
rect 88784 -51491 88800 -51457
rect 88734 -51525 88800 -51491
rect 88734 -51559 88750 -51525
rect 88784 -51559 88800 -51525
rect 88566 -51629 88582 -51595
rect 88616 -51609 88632 -51595
rect 88734 -51595 88800 -51559
rect 88834 -51457 88868 -51415
rect 88834 -51525 88868 -51491
rect 88834 -51575 88868 -51559
rect 88902 -51457 88968 -51449
rect 88902 -51491 88918 -51457
rect 88952 -51491 88968 -51457
rect 88902 -51525 88968 -51491
rect 88902 -51559 88918 -51525
rect 88952 -51559 88968 -51525
rect 88734 -51609 88750 -51595
rect 88616 -51629 88750 -51609
rect 88784 -51609 88800 -51595
rect 88902 -51595 88968 -51559
rect 89002 -51457 89036 -51415
rect 89002 -51525 89036 -51491
rect 89002 -51575 89036 -51559
rect 89070 -51457 89136 -51449
rect 89070 -51491 89086 -51457
rect 89120 -51491 89136 -51457
rect 89070 -51525 89136 -51491
rect 89070 -51559 89086 -51525
rect 89120 -51559 89136 -51525
rect 88902 -51609 88918 -51595
rect 88784 -51629 88918 -51609
rect 88952 -51609 88968 -51595
rect 89070 -51595 89136 -51559
rect 89170 -51457 89204 -51415
rect 89170 -51525 89204 -51491
rect 89170 -51575 89204 -51559
rect 89238 -51457 89304 -51449
rect 89238 -51491 89254 -51457
rect 89288 -51491 89304 -51457
rect 89238 -51525 89304 -51491
rect 89238 -51559 89254 -51525
rect 89288 -51559 89304 -51525
rect 89070 -51609 89086 -51595
rect 88952 -51629 89086 -51609
rect 89120 -51609 89136 -51595
rect 89238 -51595 89304 -51559
rect 89338 -51457 89372 -51415
rect 89338 -51525 89372 -51491
rect 89338 -51575 89372 -51559
rect 89406 -51457 89472 -51449
rect 89406 -51491 89422 -51457
rect 89456 -51491 89472 -51457
rect 89406 -51525 89472 -51491
rect 89406 -51559 89422 -51525
rect 89456 -51559 89472 -51525
rect 89238 -51609 89254 -51595
rect 89120 -51629 89254 -51609
rect 89288 -51609 89304 -51595
rect 89406 -51595 89472 -51559
rect 89506 -51457 89540 -51415
rect 89506 -51525 89540 -51491
rect 89506 -51575 89540 -51559
rect 89574 -51457 89640 -51449
rect 89574 -51491 89590 -51457
rect 89624 -51491 89640 -51457
rect 89574 -51525 89640 -51491
rect 89574 -51559 89590 -51525
rect 89624 -51559 89640 -51525
rect 89406 -51609 89422 -51595
rect 89288 -51629 89422 -51609
rect 89456 -51609 89472 -51595
rect 89574 -51595 89640 -51559
rect 89674 -51457 89708 -51415
rect 89674 -51525 89708 -51491
rect 89674 -51575 89708 -51559
rect 89742 -51457 89808 -51449
rect 89742 -51491 89758 -51457
rect 89792 -51491 89808 -51457
rect 89742 -51525 89808 -51491
rect 89742 -51559 89758 -51525
rect 89792 -51559 89808 -51525
rect 89574 -51609 89590 -51595
rect 89456 -51629 89590 -51609
rect 89624 -51609 89640 -51595
rect 89742 -51595 89808 -51559
rect 89842 -51457 89884 -51415
rect 89876 -51491 89884 -51457
rect 89842 -51525 89884 -51491
rect 89876 -51559 89884 -51525
rect 89842 -51575 89884 -51559
rect 89962 -51457 90004 -51415
rect 89962 -51491 89970 -51457
rect 89962 -51525 90004 -51491
rect 89962 -51559 89970 -51525
rect 89742 -51600 89758 -51595
rect 89792 -51600 89808 -51595
rect 89742 -51609 89750 -51600
rect 89624 -51629 89750 -51609
rect 88566 -51643 89750 -51629
rect 88467 -51686 89555 -51679
rect 88467 -51693 88523 -51686
rect 89384 -51693 89555 -51686
rect 88467 -51727 88492 -51693
rect 89384 -51720 89505 -51693
rect 88526 -51727 88666 -51720
rect 88700 -51727 88834 -51720
rect 88868 -51727 89003 -51720
rect 89037 -51727 89170 -51720
rect 89204 -51727 89338 -51720
rect 89372 -51727 89505 -51720
rect 89539 -51727 89555 -51693
rect 89742 -51761 89750 -51643
rect 87094 -51781 88336 -51780
rect 87094 -51815 87110 -51781
rect 87144 -51799 87278 -51781
rect 87144 -51815 87160 -51799
rect 87094 -51849 87160 -51815
rect 87262 -51815 87278 -51799
rect 87312 -51799 87446 -51781
rect 87312 -51815 87328 -51799
rect 87094 -51883 87110 -51849
rect 87144 -51883 87160 -51849
rect 87094 -51891 87160 -51883
rect 87194 -51849 87228 -51833
rect 87194 -51925 87228 -51883
rect 87262 -51849 87328 -51815
rect 87430 -51815 87446 -51799
rect 87480 -51799 87614 -51781
rect 87480 -51815 87496 -51799
rect 87262 -51883 87278 -51849
rect 87312 -51883 87328 -51849
rect 87262 -51891 87328 -51883
rect 87362 -51849 87396 -51833
rect 87362 -51925 87396 -51883
rect 87430 -51849 87496 -51815
rect 87598 -51815 87614 -51799
rect 87648 -51799 87782 -51781
rect 87648 -51815 87664 -51799
rect 87430 -51883 87446 -51849
rect 87480 -51883 87496 -51849
rect 87430 -51891 87496 -51883
rect 87530 -51849 87564 -51833
rect 87530 -51925 87564 -51883
rect 87598 -51849 87664 -51815
rect 87766 -51815 87782 -51799
rect 87816 -51799 87950 -51781
rect 87816 -51815 87832 -51799
rect 87598 -51883 87614 -51849
rect 87648 -51883 87664 -51849
rect 87598 -51891 87664 -51883
rect 87698 -51849 87732 -51833
rect 87698 -51925 87732 -51883
rect 87766 -51849 87832 -51815
rect 87934 -51815 87950 -51799
rect 87984 -51799 88118 -51781
rect 87984 -51815 88000 -51799
rect 87766 -51883 87782 -51849
rect 87816 -51883 87832 -51849
rect 87766 -51891 87832 -51883
rect 87866 -51849 87900 -51833
rect 87866 -51925 87900 -51883
rect 87934 -51849 88000 -51815
rect 88102 -51815 88118 -51799
rect 88152 -51799 88286 -51781
rect 88152 -51815 88168 -51799
rect 87934 -51883 87950 -51849
rect 87984 -51883 88000 -51849
rect 87934 -51891 88000 -51883
rect 88034 -51849 88068 -51833
rect 88034 -51925 88068 -51883
rect 88102 -51849 88168 -51815
rect 88270 -51815 88286 -51799
rect 88320 -51815 88336 -51781
rect 88102 -51883 88118 -51849
rect 88152 -51883 88168 -51849
rect 88102 -51891 88168 -51883
rect 88202 -51849 88236 -51833
rect 88202 -51925 88236 -51883
rect 88270 -51849 88336 -51815
rect 88270 -51883 88286 -51849
rect 88320 -51883 88336 -51849
rect 88270 -51891 88336 -51883
rect 88370 -51781 88412 -51765
rect 88404 -51815 88412 -51781
rect 88370 -51849 88412 -51815
rect 88404 -51883 88412 -51849
rect 88370 -51925 88412 -51883
rect 88486 -51781 88532 -51765
rect 88486 -51815 88498 -51781
rect 88486 -51849 88532 -51815
rect 88486 -51883 88498 -51849
rect 88486 -51925 88532 -51883
rect 88566 -51781 89750 -51761
rect 88566 -51815 88582 -51781
rect 88616 -51799 88750 -51781
rect 88616 -51815 88632 -51799
rect 88566 -51849 88632 -51815
rect 88734 -51815 88750 -51799
rect 88784 -51799 88918 -51781
rect 88784 -51815 88800 -51799
rect 88566 -51883 88582 -51849
rect 88616 -51883 88632 -51849
rect 88566 -51891 88632 -51883
rect 88666 -51849 88700 -51833
rect 88666 -51925 88700 -51883
rect 88734 -51849 88800 -51815
rect 88902 -51815 88918 -51799
rect 88952 -51799 89086 -51781
rect 88952 -51815 88968 -51799
rect 88734 -51883 88750 -51849
rect 88784 -51883 88800 -51849
rect 88734 -51891 88800 -51883
rect 88834 -51849 88868 -51833
rect 88834 -51925 88868 -51883
rect 88902 -51849 88968 -51815
rect 89070 -51815 89086 -51799
rect 89120 -51799 89254 -51781
rect 89120 -51815 89136 -51799
rect 88902 -51883 88918 -51849
rect 88952 -51883 88968 -51849
rect 88902 -51891 88968 -51883
rect 89002 -51849 89036 -51833
rect 89002 -51925 89036 -51883
rect 89070 -51849 89136 -51815
rect 89238 -51815 89254 -51799
rect 89288 -51799 89422 -51781
rect 89288 -51815 89304 -51799
rect 89070 -51883 89086 -51849
rect 89120 -51883 89136 -51849
rect 89070 -51891 89136 -51883
rect 89170 -51849 89204 -51833
rect 89170 -51925 89204 -51883
rect 89238 -51849 89304 -51815
rect 89406 -51815 89422 -51799
rect 89456 -51799 89590 -51781
rect 89456 -51815 89472 -51799
rect 89238 -51883 89254 -51849
rect 89288 -51883 89304 -51849
rect 89238 -51891 89304 -51883
rect 89338 -51849 89372 -51833
rect 89338 -51925 89372 -51883
rect 89406 -51849 89472 -51815
rect 89574 -51815 89590 -51799
rect 89624 -51790 89750 -51781
rect 89800 -51790 89808 -51600
rect 89962 -51595 90004 -51559
rect 89962 -51629 89970 -51595
rect 89962 -51645 90004 -51629
rect 90038 -51457 90104 -51449
rect 90038 -51491 90054 -51457
rect 90088 -51491 90104 -51457
rect 90038 -51525 90104 -51491
rect 90038 -51559 90054 -51525
rect 90088 -51559 90104 -51525
rect 90038 -51595 90104 -51559
rect 90138 -51457 90172 -51415
rect 90138 -51525 90172 -51491
rect 90138 -51575 90172 -51559
rect 90206 -51457 90272 -51449
rect 90206 -51491 90222 -51457
rect 90256 -51491 90272 -51457
rect 90206 -51525 90272 -51491
rect 90206 -51559 90222 -51525
rect 90256 -51559 90272 -51525
rect 90038 -51629 90054 -51595
rect 90088 -51609 90104 -51595
rect 90206 -51595 90272 -51559
rect 90306 -51457 90340 -51415
rect 90306 -51525 90340 -51491
rect 90306 -51575 90340 -51559
rect 90374 -51457 90440 -51449
rect 90374 -51491 90390 -51457
rect 90424 -51491 90440 -51457
rect 90374 -51525 90440 -51491
rect 90374 -51559 90390 -51525
rect 90424 -51559 90440 -51525
rect 90206 -51609 90222 -51595
rect 90088 -51629 90222 -51609
rect 90256 -51609 90272 -51595
rect 90374 -51595 90440 -51559
rect 90474 -51457 90508 -51415
rect 90474 -51525 90508 -51491
rect 90474 -51575 90508 -51559
rect 90542 -51457 90608 -51449
rect 90542 -51491 90558 -51457
rect 90592 -51491 90608 -51457
rect 90542 -51525 90608 -51491
rect 90542 -51559 90558 -51525
rect 90592 -51559 90608 -51525
rect 90374 -51609 90390 -51595
rect 90256 -51629 90390 -51609
rect 90424 -51609 90440 -51595
rect 90542 -51595 90608 -51559
rect 90642 -51457 90676 -51415
rect 90642 -51525 90676 -51491
rect 90642 -51575 90676 -51559
rect 90710 -51457 90776 -51449
rect 90710 -51491 90726 -51457
rect 90760 -51491 90776 -51457
rect 90710 -51525 90776 -51491
rect 90710 -51559 90726 -51525
rect 90760 -51559 90776 -51525
rect 90542 -51609 90558 -51595
rect 90424 -51629 90558 -51609
rect 90592 -51609 90608 -51595
rect 90710 -51595 90776 -51559
rect 90810 -51457 90844 -51415
rect 90810 -51525 90844 -51491
rect 90810 -51575 90844 -51559
rect 90878 -51457 90944 -51449
rect 90878 -51491 90894 -51457
rect 90928 -51491 90944 -51457
rect 90878 -51525 90944 -51491
rect 90878 -51559 90894 -51525
rect 90928 -51559 90944 -51525
rect 90710 -51609 90726 -51595
rect 90592 -51629 90726 -51609
rect 90760 -51609 90776 -51595
rect 90878 -51595 90944 -51559
rect 90978 -51457 91012 -51415
rect 90978 -51525 91012 -51491
rect 90978 -51575 91012 -51559
rect 91046 -51457 91112 -51449
rect 91046 -51491 91062 -51457
rect 91096 -51491 91112 -51457
rect 91046 -51525 91112 -51491
rect 91046 -51559 91062 -51525
rect 91096 -51559 91112 -51525
rect 90878 -51609 90894 -51595
rect 90760 -51629 90894 -51609
rect 90928 -51609 90944 -51595
rect 91046 -51595 91112 -51559
rect 91146 -51457 91180 -51415
rect 91146 -51525 91180 -51491
rect 91146 -51575 91180 -51559
rect 91214 -51457 91280 -51449
rect 91214 -51491 91230 -51457
rect 91264 -51491 91280 -51457
rect 91214 -51525 91280 -51491
rect 91214 -51559 91230 -51525
rect 91264 -51559 91280 -51525
rect 91046 -51609 91062 -51595
rect 90928 -51629 91062 -51609
rect 91096 -51609 91112 -51595
rect 91214 -51595 91280 -51559
rect 91314 -51457 91356 -51415
rect 91348 -51491 91356 -51457
rect 91314 -51525 91356 -51491
rect 91348 -51559 91356 -51525
rect 91314 -51575 91356 -51559
rect 91214 -51600 91230 -51595
rect 91264 -51600 91280 -51595
rect 91214 -51609 91220 -51600
rect 91096 -51629 91220 -51609
rect 90038 -51643 91220 -51629
rect 89939 -51687 91027 -51679
rect 89939 -51689 89980 -51687
rect 90747 -51689 91027 -51687
rect 89939 -51693 89978 -51689
rect 90748 -51693 91027 -51689
rect 89939 -51727 89964 -51693
rect 90748 -51723 90810 -51693
rect 89998 -51727 90138 -51723
rect 90172 -51727 90306 -51723
rect 90340 -51727 90475 -51723
rect 90509 -51727 90642 -51723
rect 90676 -51727 90810 -51723
rect 90844 -51727 90977 -51693
rect 91011 -51727 91027 -51693
rect 91214 -51761 91220 -51643
rect 89624 -51799 89758 -51790
rect 89624 -51815 89640 -51799
rect 89406 -51883 89422 -51849
rect 89456 -51883 89472 -51849
rect 89406 -51891 89472 -51883
rect 89506 -51849 89540 -51833
rect 89506 -51925 89540 -51883
rect 89574 -51849 89640 -51815
rect 89742 -51815 89758 -51799
rect 89792 -51815 89808 -51790
rect 89574 -51883 89590 -51849
rect 89624 -51883 89640 -51849
rect 89574 -51891 89640 -51883
rect 89674 -51849 89708 -51833
rect 89674 -51925 89708 -51883
rect 89742 -51849 89808 -51815
rect 89742 -51883 89758 -51849
rect 89792 -51883 89808 -51849
rect 89742 -51891 89808 -51883
rect 89842 -51781 89884 -51765
rect 89876 -51815 89884 -51781
rect 89842 -51849 89884 -51815
rect 89876 -51883 89884 -51849
rect 89842 -51925 89884 -51883
rect 89958 -51781 90004 -51765
rect 89958 -51815 89970 -51781
rect 89958 -51849 90004 -51815
rect 89958 -51883 89970 -51849
rect 89958 -51925 90004 -51883
rect 90038 -51781 91220 -51761
rect 90038 -51815 90054 -51781
rect 90088 -51799 90222 -51781
rect 90088 -51815 90104 -51799
rect 90038 -51849 90104 -51815
rect 90206 -51815 90222 -51799
rect 90256 -51799 90390 -51781
rect 90256 -51815 90272 -51799
rect 90038 -51883 90054 -51849
rect 90088 -51883 90104 -51849
rect 90038 -51891 90104 -51883
rect 90138 -51849 90172 -51833
rect 90138 -51925 90172 -51883
rect 90206 -51849 90272 -51815
rect 90374 -51815 90390 -51799
rect 90424 -51799 90558 -51781
rect 90424 -51815 90440 -51799
rect 90206 -51883 90222 -51849
rect 90256 -51883 90272 -51849
rect 90206 -51891 90272 -51883
rect 90306 -51849 90340 -51833
rect 90306 -51925 90340 -51883
rect 90374 -51849 90440 -51815
rect 90542 -51815 90558 -51799
rect 90592 -51799 90726 -51781
rect 90592 -51815 90608 -51799
rect 90374 -51883 90390 -51849
rect 90424 -51883 90440 -51849
rect 90374 -51891 90440 -51883
rect 90474 -51849 90508 -51833
rect 90474 -51925 90508 -51883
rect 90542 -51849 90608 -51815
rect 90710 -51815 90726 -51799
rect 90760 -51799 90894 -51781
rect 90760 -51815 90776 -51799
rect 90542 -51883 90558 -51849
rect 90592 -51883 90608 -51849
rect 90542 -51891 90608 -51883
rect 90642 -51849 90676 -51833
rect 90642 -51925 90676 -51883
rect 90710 -51849 90776 -51815
rect 90878 -51815 90894 -51799
rect 90928 -51799 91062 -51781
rect 90928 -51815 90944 -51799
rect 90710 -51883 90726 -51849
rect 90760 -51883 90776 -51849
rect 90710 -51891 90776 -51883
rect 90810 -51849 90844 -51833
rect 90810 -51925 90844 -51883
rect 90878 -51849 90944 -51815
rect 91046 -51815 91062 -51799
rect 91096 -51790 91220 -51781
rect 91270 -51790 91280 -51600
rect 91096 -51799 91230 -51790
rect 91096 -51815 91112 -51799
rect 90878 -51883 90894 -51849
rect 90928 -51883 90944 -51849
rect 90878 -51891 90944 -51883
rect 90978 -51849 91012 -51833
rect 90978 -51925 91012 -51883
rect 91046 -51849 91112 -51815
rect 91214 -51815 91230 -51799
rect 91264 -51815 91280 -51790
rect 91046 -51883 91062 -51849
rect 91096 -51883 91112 -51849
rect 91046 -51891 91112 -51883
rect 91146 -51849 91180 -51833
rect 91146 -51925 91180 -51883
rect 91214 -51849 91280 -51815
rect 91214 -51883 91230 -51849
rect 91264 -51883 91280 -51849
rect 91214 -51891 91280 -51883
rect 91314 -51781 91356 -51765
rect 91348 -51815 91356 -51781
rect 91314 -51849 91356 -51815
rect 91348 -51883 91356 -51849
rect 91314 -51925 91356 -51883
rect 78137 -51947 78205 -51939
rect 82838 -51959 82867 -51925
rect 82901 -51959 82959 -51925
rect 82993 -51959 83051 -51925
rect 83085 -51959 83143 -51925
rect 83177 -51959 83235 -51925
rect 83269 -51959 83327 -51925
rect 83361 -51959 83419 -51925
rect 83453 -51959 83511 -51925
rect 83545 -51959 83603 -51925
rect 83637 -51959 83695 -51925
rect 83729 -51959 83787 -51925
rect 83821 -51959 83879 -51925
rect 83913 -51959 83971 -51925
rect 84005 -51959 84063 -51925
rect 84097 -51959 84155 -51925
rect 84189 -51959 84247 -51925
rect 84281 -51959 84339 -51925
rect 84373 -51959 84431 -51925
rect 84465 -51959 84523 -51925
rect 84557 -51959 84615 -51925
rect 84649 -51959 84707 -51925
rect 84741 -51959 84799 -51925
rect 84833 -51959 84891 -51925
rect 84925 -51959 84983 -51925
rect 85017 -51959 85075 -51925
rect 85109 -51959 85167 -51925
rect 85201 -51959 85259 -51925
rect 85293 -51959 85351 -51925
rect 85385 -51959 85443 -51925
rect 85477 -51959 85535 -51925
rect 85569 -51959 85627 -51925
rect 85661 -51959 85719 -51925
rect 85753 -51959 85811 -51925
rect 85845 -51959 85903 -51925
rect 85937 -51959 85995 -51925
rect 86029 -51959 86087 -51925
rect 86121 -51959 86179 -51925
rect 86213 -51959 86271 -51925
rect 86305 -51959 86363 -51925
rect 86397 -51959 86455 -51925
rect 86489 -51959 86547 -51925
rect 86581 -51959 86639 -51925
rect 86673 -51959 86731 -51925
rect 86765 -51959 86823 -51925
rect 86857 -51959 86915 -51925
rect 86949 -51959 87007 -51925
rect 87041 -51959 87099 -51925
rect 87133 -51959 87191 -51925
rect 87225 -51959 87283 -51925
rect 87317 -51959 87375 -51925
rect 87409 -51959 87467 -51925
rect 87501 -51959 87559 -51925
rect 87593 -51959 87651 -51925
rect 87685 -51959 87743 -51925
rect 87777 -51959 87835 -51925
rect 87869 -51959 87927 -51925
rect 87961 -51959 88019 -51925
rect 88053 -51959 88111 -51925
rect 88145 -51959 88203 -51925
rect 88237 -51959 88295 -51925
rect 88329 -51959 88387 -51925
rect 88421 -51959 88479 -51925
rect 88513 -51959 88571 -51925
rect 88605 -51959 88663 -51925
rect 88697 -51959 88755 -51925
rect 88789 -51959 88847 -51925
rect 88881 -51959 88939 -51925
rect 88973 -51959 89031 -51925
rect 89065 -51959 89123 -51925
rect 89157 -51959 89215 -51925
rect 89249 -51959 89307 -51925
rect 89341 -51959 89399 -51925
rect 89433 -51959 89491 -51925
rect 89525 -51959 89583 -51925
rect 89617 -51959 89675 -51925
rect 89709 -51959 89767 -51925
rect 89801 -51959 89859 -51925
rect 89893 -51959 89951 -51925
rect 89985 -51959 90043 -51925
rect 90077 -51959 90135 -51925
rect 90169 -51959 90227 -51925
rect 90261 -51959 90319 -51925
rect 90353 -51959 90411 -51925
rect 90445 -51959 90503 -51925
rect 90537 -51959 90595 -51925
rect 90629 -51959 90687 -51925
rect 90721 -51959 90779 -51925
rect 90813 -51959 90871 -51925
rect 90905 -51959 90963 -51925
rect 90997 -51959 91055 -51925
rect 91089 -51959 91147 -51925
rect 91181 -51959 91239 -51925
rect 91273 -51959 91331 -51925
rect 91365 -51959 91394 -51925
rect 77578 -52015 77607 -51981
rect 77641 -52015 77699 -51981
rect 77733 -52015 77791 -51981
rect 77825 -52015 77883 -51981
rect 77917 -52015 77975 -51981
rect 78009 -52015 78067 -51981
rect 78101 -52015 78159 -51981
rect 78193 -52015 78222 -51981
rect 60466 -52060 60546 -52040
rect 60466 -52100 60486 -52060
rect 60526 -52100 60546 -52060
rect 60466 -52120 60546 -52100
rect 60606 -52060 60686 -52040
rect 60606 -52100 60626 -52060
rect 60666 -52100 60686 -52060
rect 60606 -52120 60686 -52100
rect 60746 -52060 60826 -52040
rect 60746 -52100 60766 -52060
rect 60806 -52100 60826 -52060
rect 60746 -52120 60826 -52100
rect 60886 -52060 60966 -52040
rect 60886 -52100 60906 -52060
rect 60946 -52100 60966 -52060
rect 77578 -52087 77607 -52053
rect 77641 -52087 77699 -52053
rect 77733 -52087 77791 -52053
rect 77825 -52087 77883 -52053
rect 77917 -52087 77975 -52053
rect 78009 -52087 78067 -52053
rect 78101 -52087 78159 -52053
rect 78193 -52087 78222 -52053
rect 60886 -52120 60966 -52100
rect 60019 -52223 60053 -52161
rect 77596 -52129 77663 -52087
rect 77596 -52163 77613 -52129
rect 77647 -52163 77663 -52129
rect 77697 -52137 77747 -52121
rect 77697 -52171 77705 -52137
rect 77739 -52171 77747 -52137
rect 59387 -52257 59476 -52223
rect 59646 -52257 59799 -52223
rect 59957 -52226 60053 -52223
rect 77450 -52200 77530 -52190
rect 77595 -52200 77643 -52199
rect 77450 -52210 77643 -52200
rect 59957 -52257 60520 -52226
rect 59772 -52260 60520 -52257
rect 59772 -52320 59806 -52260
rect 59276 -52438 59310 -52376
rect 58930 -52472 59026 -52438
rect 59214 -52440 59310 -52438
rect 59214 -52472 59696 -52440
rect 58930 -52474 59696 -52472
rect 58930 -52510 58964 -52474
rect 57129 -52591 57131 -52557
rect 57129 -52625 57165 -52591
rect 57129 -52659 57131 -52625
rect 57129 -52675 57165 -52659
rect 57201 -52591 57217 -52557
rect 57251 -52591 57267 -52557
rect 57201 -52625 57267 -52591
rect 57201 -52659 57217 -52625
rect 57251 -52659 57267 -52625
rect 57201 -52709 57267 -52659
rect 57301 -52578 57303 -52544
rect 57337 -52578 57355 -52544
rect 57301 -52625 57355 -52578
rect 57301 -52659 57303 -52625
rect 57337 -52659 57355 -52625
rect 57301 -52675 57355 -52659
rect 59662 -52530 59696 -52474
rect 60486 -52322 60520 -52260
rect 77450 -52260 77470 -52210
rect 77510 -52260 77643 -52210
rect 77450 -52270 77643 -52260
rect 77450 -52280 77530 -52270
rect 59942 -52374 59958 -52340
rect 60334 -52374 60350 -52340
rect 59874 -52394 59908 -52378
rect 59874 -52444 59908 -52428
rect 60384 -52394 60418 -52378
rect 60384 -52444 60418 -52428
rect 59942 -52482 59958 -52448
rect 60334 -52482 60350 -52448
rect 56112 -52782 56146 -52720
rect 57096 -52743 57125 -52709
rect 57159 -52743 57217 -52709
rect 57251 -52743 57309 -52709
rect 57343 -52743 57372 -52709
rect 55706 -52816 55802 -52782
rect 56050 -52816 56146 -52782
rect 53886 -52864 53982 -52830
rect 54956 -52864 55052 -52830
rect 53886 -52926 53920 -52864
rect 55018 -52926 55052 -52864
rect 55720 -52858 56090 -52816
rect 55720 -52868 56020 -52858
rect 54065 -52978 54081 -52944
rect 54857 -52978 54873 -52944
rect 53988 -53006 54022 -52990
rect 53988 -53060 54022 -53044
rect 54916 -53006 54950 -52990
rect 54916 -53060 54950 -53044
rect 54065 -53106 54081 -53072
rect 54857 -53106 54873 -53072
rect 53886 -53186 53920 -53124
rect 56010 -53008 56020 -52868
rect 56080 -53008 56090 -52858
rect 59109 -52588 59125 -52554
rect 59501 -52588 59517 -52554
rect 59560 -52608 59594 -52592
rect 59560 -52658 59594 -52642
rect 59109 -52696 59125 -52662
rect 59501 -52696 59517 -52662
rect 59032 -52716 59066 -52700
rect 59032 -52766 59066 -52750
rect 59109 -52804 59125 -52770
rect 59501 -52804 59517 -52770
rect 56010 -53018 56090 -53008
rect 59772 -52562 59806 -52500
rect 77595 -52365 77643 -52270
rect 77697 -52281 77747 -52171
rect 77791 -52129 77857 -52087
rect 77791 -52163 77807 -52129
rect 77841 -52163 77857 -52129
rect 77791 -52231 77857 -52163
rect 77894 -52137 77944 -52121
rect 77894 -52171 77902 -52137
rect 77936 -52171 77944 -52137
rect 77894 -52281 77944 -52171
rect 78037 -52129 78103 -52087
rect 78037 -52163 78053 -52129
rect 78087 -52163 78103 -52129
rect 78037 -52197 78103 -52163
rect 78137 -52129 78205 -52121
rect 78137 -52163 78153 -52129
rect 78187 -52130 78205 -52129
rect 78187 -52163 78310 -52130
rect 78137 -52173 78310 -52163
rect 78037 -52231 78053 -52197
rect 78087 -52231 78103 -52197
rect 78037 -52247 78103 -52231
rect 78153 -52180 78310 -52173
rect 78153 -52197 78180 -52180
rect 78153 -52265 78180 -52231
rect 77595 -52399 77609 -52365
rect 60486 -52562 60520 -52500
rect 77595 -52461 77643 -52399
rect 77677 -52315 78115 -52281
rect 77677 -52497 77711 -52315
rect 78052 -52349 78115 -52315
rect 77612 -52513 77711 -52497
rect 59772 -52596 59866 -52562
rect 60426 -52596 60520 -52562
rect 77612 -52547 77613 -52513
rect 77647 -52547 77711 -52513
rect 77755 -52365 77825 -52349
rect 77789 -52399 77825 -52365
rect 77755 -52480 77825 -52399
rect 77755 -52520 77770 -52480
rect 77810 -52520 77825 -52480
rect 77755 -52542 77825 -52520
rect 77861 -52360 77921 -52349
rect 77861 -52365 77870 -52360
rect 77861 -52400 77870 -52399
rect 77910 -52400 77921 -52360
rect 77861 -52450 77921 -52400
rect 77861 -52510 77870 -52450
rect 77910 -52510 77921 -52450
rect 77861 -52543 77921 -52510
rect 77957 -52365 78013 -52349
rect 77991 -52399 78013 -52365
rect 78052 -52365 78118 -52349
rect 78052 -52399 78068 -52365
rect 78102 -52399 78118 -52365
rect 77957 -52400 78013 -52399
rect 77957 -52500 77970 -52400
rect 78010 -52500 78013 -52400
rect 77957 -52543 78013 -52500
rect 78049 -52453 78103 -52437
rect 78153 -52453 78180 -52299
rect 78049 -52487 78054 -52453
rect 78088 -52487 78103 -52453
rect 78049 -52521 78103 -52487
rect 77612 -52563 77711 -52547
rect 78049 -52555 78054 -52521
rect 78088 -52555 78103 -52521
rect 78137 -52487 78153 -52453
rect 78137 -52500 78180 -52487
rect 78290 -52500 78310 -52180
rect 78137 -52521 78310 -52500
rect 78137 -52555 78153 -52521
rect 78187 -52550 78310 -52521
rect 78187 -52555 78205 -52550
rect 78049 -52597 78103 -52555
rect 77578 -52631 77607 -52597
rect 77641 -52631 77699 -52597
rect 77733 -52631 77791 -52597
rect 77825 -52631 77883 -52597
rect 77917 -52631 77975 -52597
rect 78009 -52631 78067 -52597
rect 78101 -52631 78159 -52597
rect 78193 -52631 78222 -52597
rect 77578 -52705 77607 -52671
rect 77641 -52705 77699 -52671
rect 77733 -52705 77791 -52671
rect 77825 -52705 77883 -52671
rect 77917 -52705 77975 -52671
rect 78009 -52705 78067 -52671
rect 78101 -52705 78159 -52671
rect 78193 -52705 78222 -52671
rect 77612 -52755 77711 -52739
rect 77612 -52789 77613 -52755
rect 77647 -52789 77711 -52755
rect 78049 -52747 78103 -52705
rect 77612 -52805 77711 -52789
rect 59662 -52884 59696 -52830
rect 58966 -52900 59026 -52884
rect 58930 -52918 59026 -52900
rect 59600 -52918 59696 -52884
rect 77560 -52841 77640 -52840
rect 77560 -52903 77643 -52841
rect 77560 -52937 77609 -52903
rect 77560 -52990 77643 -52937
rect 55018 -53186 55052 -53124
rect 53886 -53220 53982 -53186
rect 54956 -53220 55052 -53186
rect 55176 -53078 55272 -53044
rect 55566 -53078 55662 -53044
rect 55176 -53140 55210 -53078
rect 55628 -53140 55662 -53078
rect 77560 -53080 77580 -52990
rect 77630 -53080 77643 -52990
rect 77677 -52987 77711 -52805
rect 77755 -52780 77825 -52760
rect 77755 -52820 77770 -52780
rect 77810 -52820 77825 -52780
rect 77755 -52903 77825 -52820
rect 77789 -52937 77825 -52903
rect 77755 -52953 77825 -52937
rect 77861 -52890 77921 -52759
rect 77861 -52903 77870 -52890
rect 77910 -52930 77921 -52890
rect 77895 -52937 77921 -52930
rect 77861 -52953 77921 -52937
rect 77957 -52900 78013 -52759
rect 78049 -52781 78054 -52747
rect 78088 -52781 78103 -52747
rect 78049 -52815 78103 -52781
rect 78049 -52849 78054 -52815
rect 78088 -52849 78103 -52815
rect 78137 -52781 78153 -52747
rect 78187 -52781 78205 -52747
rect 78137 -52815 78205 -52781
rect 78137 -52849 78153 -52815
rect 78187 -52849 78205 -52815
rect 78049 -52865 78103 -52849
rect 77957 -52903 77960 -52900
rect 77957 -52950 77960 -52937
rect 78010 -52950 78013 -52900
rect 77957 -52953 78013 -52950
rect 78052 -52937 78068 -52903
rect 78102 -52937 78118 -52903
rect 78052 -52953 78118 -52937
rect 78052 -52987 78115 -52953
rect 77677 -53021 78115 -52987
rect 78153 -52960 78205 -52849
rect 78153 -52990 78290 -52960
rect 78153 -53003 78190 -52990
rect 77560 -53100 77643 -53080
rect 77595 -53103 77643 -53100
rect 77697 -53131 77747 -53021
rect 55284 -53192 55300 -53158
rect 55476 -53192 55492 -53158
rect 55526 -53202 55560 -53186
rect 55284 -53280 55300 -53246
rect 55476 -53280 55492 -53246
rect 55526 -53252 55560 -53236
rect 35802 -53380 35836 -53318
rect 25780 -53388 35836 -53380
rect 55176 -53360 55210 -53298
rect 77596 -53173 77613 -53139
rect 77647 -53173 77663 -53139
rect 77596 -53215 77663 -53173
rect 77697 -53165 77705 -53131
rect 77739 -53165 77747 -53131
rect 77697 -53181 77747 -53165
rect 77791 -53139 77857 -53071
rect 77791 -53173 77807 -53139
rect 77841 -53173 77857 -53139
rect 77791 -53215 77857 -53173
rect 77894 -53131 77944 -53021
rect 78187 -53037 78190 -53003
rect 77894 -53165 77902 -53131
rect 77936 -53165 77944 -53131
rect 77894 -53181 77944 -53165
rect 78037 -53071 78103 -53055
rect 78037 -53105 78053 -53071
rect 78087 -53105 78103 -53071
rect 78037 -53139 78103 -53105
rect 78153 -53071 78190 -53037
rect 78187 -53105 78190 -53071
rect 78153 -53120 78190 -53105
rect 78260 -53120 78290 -52990
rect 78153 -53129 78290 -53120
rect 78037 -53173 78053 -53139
rect 78087 -53173 78103 -53139
rect 78037 -53215 78103 -53173
rect 78137 -53139 78290 -53129
rect 78137 -53173 78153 -53139
rect 78187 -53140 78290 -53139
rect 78187 -53173 78205 -53140
rect 78137 -53181 78205 -53173
rect 77578 -53249 77607 -53215
rect 77641 -53249 77699 -53215
rect 77733 -53249 77791 -53215
rect 77825 -53249 77883 -53215
rect 77917 -53249 77975 -53215
rect 78009 -53249 78067 -53215
rect 78101 -53249 78159 -53215
rect 78193 -53249 78222 -53215
rect 55628 -53360 55662 -53298
rect 77578 -53325 77607 -53291
rect 77641 -53325 77699 -53291
rect 77733 -53325 77791 -53291
rect 77825 -53325 77883 -53291
rect 77917 -53325 77975 -53291
rect 78009 -53325 78067 -53291
rect 78101 -53325 78159 -53291
rect 78193 -53325 78251 -53291
rect 78285 -53325 78343 -53291
rect 78377 -53325 78435 -53291
rect 78469 -53325 78527 -53291
rect 78561 -53325 78619 -53291
rect 78653 -53325 78711 -53291
rect 78745 -53325 78803 -53291
rect 78837 -53325 78895 -53291
rect 78929 -53325 78987 -53291
rect 79021 -53325 79050 -53291
rect 25780 -53422 35838 -53388
rect 55176 -53394 55272 -53360
rect 55566 -53394 55662 -53360
rect 35804 -53484 35838 -53422
rect 77595 -53436 77716 -53325
rect 77751 -53376 77847 -53359
rect 77785 -53392 77847 -53376
rect 77751 -53427 77770 -53410
rect 77830 -53427 77847 -53392
rect 77881 -53367 77932 -53325
rect 77881 -53401 77885 -53367
rect 77919 -53401 77932 -53367
rect 77881 -53434 77932 -53401
rect 77966 -53381 78021 -53359
rect 77966 -53415 77969 -53381
rect 78003 -53415 78021 -53381
rect 77595 -53456 77718 -53436
rect 77681 -53461 77718 -53456
rect 77966 -53449 78021 -53415
rect 77681 -53476 77747 -53461
rect 77595 -53506 77647 -53490
rect 77595 -53540 77613 -53506
rect 77681 -53510 77697 -53476
rect 77731 -53510 77747 -53476
rect 77781 -53495 77932 -53475
rect 77781 -53525 77790 -53495
rect 77778 -53529 77790 -53525
rect 77824 -53529 77932 -53495
rect 77966 -53483 77969 -53449
rect 78003 -53483 78021 -53449
rect 78095 -53409 78151 -53325
rect 78285 -53367 78351 -53325
rect 78095 -53443 78109 -53409
rect 78143 -53443 78151 -53409
rect 78095 -53459 78151 -53443
rect 78185 -53409 78245 -53393
rect 78185 -53443 78193 -53409
rect 78227 -53443 78245 -53409
rect 77966 -53499 78021 -53483
rect 77778 -53532 77932 -53529
rect 77775 -53534 77932 -53532
rect 77774 -53537 77953 -53534
rect 77770 -53540 77953 -53537
rect 77595 -53580 77647 -53540
rect 77766 -53542 77953 -53540
rect 77761 -53544 77953 -53542
rect 77747 -53550 77953 -53544
rect 77743 -53556 77953 -53550
rect 77739 -53562 77953 -53556
rect 77733 -53567 77953 -53562
rect 77726 -53574 77953 -53567
rect 77720 -53575 77953 -53574
rect 77720 -53576 77798 -53575
rect 77720 -53578 77793 -53576
rect 77720 -53579 77790 -53578
rect 77720 -53580 77787 -53579
rect 77595 -53581 77787 -53580
rect 77595 -53583 77785 -53581
rect 77595 -53584 77783 -53583
rect 77595 -53586 77781 -53584
rect 77595 -53588 77780 -53586
rect 77595 -53589 77779 -53588
rect 77595 -53592 77777 -53589
rect 77595 -53595 77776 -53592
rect 77595 -53600 77774 -53595
rect 77595 -53614 77773 -53600
rect 77907 -53603 77953 -53575
rect 77595 -53649 77705 -53648
rect 77595 -53683 77613 -53649
rect 77647 -53660 77705 -53649
rect 77595 -53710 77620 -53683
rect 77690 -53710 77705 -53660
rect 77595 -53725 77705 -53710
rect 77739 -53759 77773 -53614
rect 77595 -53793 77613 -53759
rect 77647 -53793 77773 -53759
rect 77807 -53630 77823 -53609
rect 77857 -53630 77873 -53609
rect 77807 -53680 77820 -53630
rect 77860 -53680 77873 -53630
rect 77907 -53637 77919 -53603
rect 77907 -53654 77953 -53637
rect 77807 -53694 77873 -53680
rect 77807 -53791 77851 -53694
rect 77987 -53705 78021 -53499
rect 78185 -53503 78245 -53443
rect 78285 -53401 78301 -53367
rect 78335 -53401 78351 -53367
rect 78285 -53435 78351 -53401
rect 78285 -53469 78301 -53435
rect 78335 -53469 78351 -53435
rect 78389 -53360 78481 -53359
rect 78389 -53367 78840 -53360
rect 78389 -53401 78405 -53367
rect 78439 -53369 78840 -53367
rect 78881 -53367 78937 -53325
rect 78439 -53379 78847 -53369
rect 78439 -53401 78755 -53379
rect 78389 -53413 78755 -53401
rect 78789 -53413 78847 -53379
rect 78389 -53420 78847 -53413
rect 78389 -53435 78481 -53420
rect 78516 -53427 78847 -53420
rect 78881 -53401 78894 -53367
rect 78928 -53401 78937 -53367
rect 78389 -53469 78405 -53435
rect 78439 -53469 78481 -53435
rect 78881 -53435 78937 -53401
rect 78060 -53515 78150 -53510
rect 78058 -53530 78150 -53515
rect 78058 -53620 78080 -53530
rect 78130 -53587 78150 -53530
rect 78185 -53537 78373 -53503
rect 78339 -53587 78373 -53537
rect 78130 -53603 78193 -53587
rect 78058 -53637 78112 -53620
rect 78146 -53637 78193 -53603
rect 78237 -53590 78305 -53587
rect 78237 -53630 78250 -53590
rect 78290 -53630 78305 -53590
rect 78237 -53637 78253 -53630
rect 78287 -53637 78305 -53630
rect 78339 -53603 78397 -53587
rect 78339 -53637 78361 -53603
rect 78395 -53637 78397 -53603
rect 78339 -53653 78397 -53637
rect 78339 -53671 78373 -53653
rect 77969 -53710 78021 -53705
rect 78095 -53709 78373 -53671
rect 77969 -53720 78050 -53710
rect 77885 -53743 77935 -53727
rect 77919 -53777 77935 -53743
rect 77885 -53835 77935 -53777
rect 77969 -53733 77990 -53720
rect 78030 -53760 78050 -53720
rect 78003 -53767 78050 -53760
rect 77969 -53800 78050 -53767
rect 78095 -53731 78161 -53709
rect 78095 -53765 78109 -53731
rect 78143 -53765 78161 -53731
rect 78431 -53743 78481 -53469
rect 78516 -53495 78834 -53461
rect 78881 -53469 78894 -53435
rect 78928 -53469 78937 -53435
rect 78881 -53485 78937 -53469
rect 78979 -53360 79033 -53359
rect 78979 -53398 79090 -53360
rect 79013 -53410 79090 -53398
rect 79013 -53432 79020 -53410
rect 78979 -53466 79020 -53432
rect 78516 -53498 78580 -53495
rect 78516 -53532 78533 -53498
rect 78567 -53532 78580 -53498
rect 78800 -53519 78834 -53495
rect 79013 -53500 79020 -53466
rect 78516 -53553 78580 -53532
rect 78620 -53560 78762 -53529
rect 78800 -53553 78945 -53519
rect 78979 -53553 79020 -53500
rect 78516 -53600 78586 -53587
rect 78516 -53680 78530 -53600
rect 78570 -53680 78586 -53600
rect 78620 -53630 78650 -53560
rect 78730 -53630 78762 -53560
rect 78911 -53587 78945 -53553
rect 78620 -53637 78659 -53630
rect 78693 -53637 78762 -53630
rect 78620 -53653 78762 -53637
rect 78796 -53600 78877 -53587
rect 78796 -53640 78820 -53600
rect 78860 -53603 78877 -53600
rect 78869 -53637 78877 -53603
rect 78860 -53640 78877 -53637
rect 78796 -53653 78877 -53640
rect 78911 -53603 78965 -53587
rect 78911 -53637 78931 -53603
rect 78911 -53653 78965 -53637
rect 78516 -53701 78586 -53680
rect 78911 -53687 78945 -53653
rect 78623 -53721 78945 -53687
rect 78999 -53700 79020 -53553
rect 78979 -53717 79020 -53700
rect 78095 -53781 78161 -53765
rect 78285 -53759 78335 -53743
rect 78285 -53793 78301 -53759
rect 77969 -53801 78021 -53800
rect 78285 -53835 78335 -53793
rect 78369 -53759 78481 -53743
rect 78369 -53793 78385 -53759
rect 78419 -53793 78481 -53759
rect 78369 -53801 78481 -53793
rect 78517 -53769 78533 -53735
rect 78567 -53769 78583 -53735
rect 78517 -53835 78583 -53769
rect 78623 -53741 78657 -53721
rect 78797 -53741 78831 -53721
rect 78623 -53791 78657 -53775
rect 78697 -53789 78713 -53755
rect 78747 -53789 78763 -53755
rect 78697 -53835 78763 -53789
rect 79013 -53720 79020 -53717
rect 79070 -53720 79090 -53410
rect 79013 -53751 79090 -53720
rect 78797 -53791 78831 -53775
rect 78865 -53789 78891 -53755
rect 78925 -53789 78941 -53755
rect 78979 -53769 79090 -53751
rect 79000 -53770 79090 -53769
rect 78865 -53835 78941 -53789
rect 77578 -53869 77607 -53835
rect 77641 -53869 77699 -53835
rect 77733 -53869 77791 -53835
rect 77825 -53869 77883 -53835
rect 77917 -53869 77975 -53835
rect 78009 -53869 78067 -53835
rect 78101 -53869 78159 -53835
rect 78193 -53869 78251 -53835
rect 78285 -53869 78343 -53835
rect 78377 -53869 78435 -53835
rect 78469 -53869 78527 -53835
rect 78561 -53869 78619 -53835
rect 78653 -53869 78711 -53835
rect 78745 -53869 78803 -53835
rect 78837 -53869 78895 -53835
rect 78929 -53869 78987 -53835
rect 79021 -53869 79050 -53835
rect 35804 -54982 35838 -54920
rect 25780 -55016 35838 -54982
rect 25780 -55020 35836 -55016
rect 35802 -55082 35836 -55020
rect 53896 -55592 53992 -55558
rect 54966 -55592 55062 -55558
rect 53896 -55654 53930 -55592
rect 55028 -55654 55062 -55592
rect 54075 -55706 54091 -55672
rect 54867 -55706 54883 -55672
rect 53998 -55734 54032 -55718
rect 53998 -55788 54032 -55772
rect 54926 -55734 54960 -55718
rect 54926 -55788 54960 -55772
rect 54075 -55834 54091 -55800
rect 54867 -55834 54883 -55800
rect 53896 -55914 53930 -55852
rect 55028 -55914 55062 -55852
rect 55960 -55908 56040 -55898
rect 53896 -55948 53992 -55914
rect 54966 -55948 55062 -55914
rect 53350 -56038 53790 -56004
rect 53350 -56100 53384 -56038
rect 53510 -56140 53526 -56106
rect 53614 -56140 53630 -56106
rect 35802 -56580 35836 -56518
rect 25780 -56620 35836 -56580
rect 35802 -56682 35836 -56620
rect 25736 -58180 25770 -58118
rect 53464 -56190 53498 -56174
rect 53464 -56982 53498 -56966
rect 53642 -56190 53676 -56174
rect 53642 -56982 53676 -56966
rect 53756 -56664 53790 -56038
rect 53896 -56010 53930 -55948
rect 55028 -56010 55062 -55948
rect 55710 -55954 56040 -55908
rect 54075 -56062 54091 -56028
rect 54867 -56062 54883 -56028
rect 53998 -56090 54032 -56074
rect 53998 -56144 54032 -56128
rect 54926 -56090 54960 -56074
rect 54926 -56144 54960 -56128
rect 54075 -56190 54091 -56156
rect 54867 -56190 54883 -56156
rect 53896 -56270 53930 -56208
rect 55706 -55988 55802 -55954
rect 56050 -55988 56146 -55954
rect 55706 -56050 55740 -55988
rect 55028 -56270 55062 -56208
rect 53896 -56304 53992 -56270
rect 54966 -56304 55062 -56270
rect 55176 -56100 55272 -56066
rect 55430 -56100 55526 -56066
rect 55176 -56162 55210 -56100
rect 55492 -56162 55526 -56100
rect 55318 -56202 55334 -56168
rect 55368 -56202 55384 -56168
rect 55290 -56252 55324 -56236
rect 55290 -56444 55324 -56428
rect 55378 -56252 55412 -56236
rect 55378 -56444 55412 -56428
rect 55176 -56518 55210 -56456
rect 55492 -56518 55526 -56456
rect 54870 -56552 55272 -56518
rect 55430 -56552 55706 -56518
rect 54870 -56558 55706 -56552
rect 54870 -56664 54904 -56558
rect 53756 -56698 53852 -56664
rect 54808 -56698 54904 -56664
rect 53756 -56760 53790 -56698
rect 54870 -56760 54904 -56698
rect 55126 -56708 55142 -56674
rect 55494 -56708 55510 -56674
rect 53926 -56812 53942 -56778
rect 54718 -56812 54734 -56778
rect 53858 -56840 53892 -56824
rect 53858 -56944 53892 -56928
rect 54768 -56840 54802 -56824
rect 54768 -56944 54802 -56928
rect 53926 -56990 53942 -56956
rect 54718 -56990 54734 -56956
rect 53510 -57050 53526 -57016
rect 53614 -57050 53630 -57016
rect 53756 -57070 53790 -57008
rect 55046 -56760 55080 -56744
rect 55046 -56810 55080 -56794
rect 55556 -56760 55590 -56744
rect 55556 -56810 55590 -56794
rect 55126 -56880 55142 -56846
rect 55494 -56880 55510 -56846
rect 54870 -57038 54904 -57008
rect 55700 -57006 55706 -56558
rect 56112 -56050 56146 -55988
rect 58930 -55967 59026 -55933
rect 59600 -55967 59696 -55933
rect 58930 -56010 58964 -55967
rect 58926 -56020 58966 -56010
rect 55866 -56090 55882 -56056
rect 55970 -56090 55986 -56056
rect 55820 -56140 55854 -56124
rect 55820 -56932 55854 -56916
rect 55998 -56140 56032 -56124
rect 55998 -56932 56032 -56916
rect 55866 -57000 55882 -56966
rect 55970 -57000 55986 -56966
rect 55700 -57038 55740 -57006
rect 57096 -56079 57125 -56045
rect 57159 -56079 57217 -56045
rect 57251 -56079 57309 -56045
rect 57343 -56079 57372 -56045
rect 57129 -56129 57165 -56113
rect 57129 -56163 57131 -56129
rect 57129 -56197 57165 -56163
rect 57129 -56231 57131 -56197
rect 57201 -56129 57267 -56079
rect 57201 -56163 57217 -56129
rect 57251 -56163 57267 -56129
rect 57201 -56197 57267 -56163
rect 57201 -56231 57217 -56197
rect 57251 -56231 57267 -56197
rect 57301 -56129 57355 -56113
rect 57301 -56163 57303 -56129
rect 57337 -56163 57355 -56129
rect 57301 -56210 57355 -56163
rect 57129 -56265 57165 -56231
rect 57301 -56244 57303 -56210
rect 57337 -56244 57355 -56210
rect 57129 -56299 57264 -56265
rect 57301 -56294 57355 -56244
rect 57230 -56328 57264 -56299
rect 57117 -56344 57185 -56335
rect 57117 -56394 57118 -56344
rect 57178 -56394 57185 -56344
rect 57117 -56409 57185 -56394
rect 57230 -56344 57285 -56328
rect 57230 -56378 57251 -56344
rect 57230 -56394 57285 -56378
rect 57319 -56340 57355 -56294
rect 59662 -56029 59696 -55967
rect 59109 -56081 59125 -56047
rect 59501 -56081 59517 -56047
rect 59560 -56101 59594 -56085
rect 59560 -56151 59594 -56135
rect 59109 -56189 59125 -56155
rect 59501 -56189 59517 -56155
rect 59032 -56209 59066 -56193
rect 59032 -56259 59066 -56243
rect 59109 -56297 59125 -56263
rect 59501 -56297 59517 -56263
rect 58926 -56340 58966 -56320
rect 57319 -56380 57326 -56340
rect 58930 -56376 58964 -56340
rect 57230 -56445 57264 -56394
rect 57131 -56479 57264 -56445
rect 57319 -56454 57355 -56380
rect 57131 -56500 57165 -56479
rect 56316 -56518 56412 -56504
rect 54830 -57048 55830 -57038
rect 54830 -57070 55030 -57048
rect 53756 -57104 53852 -57070
rect 54808 -57104 55030 -57070
rect 53510 -57158 53526 -57124
rect 53614 -57158 53630 -57124
rect 53756 -57166 53790 -57104
rect 54830 -57128 55030 -57104
rect 55110 -57068 55740 -57048
rect 55810 -57068 55830 -57048
rect 56112 -57068 56146 -57006
rect 55110 -57108 55160 -57068
rect 55600 -57108 55740 -57068
rect 56050 -57102 56146 -57068
rect 55110 -57128 55740 -57108
rect 55810 -57128 55830 -57102
rect 54830 -57138 55830 -57128
rect 53464 -57208 53498 -57192
rect 35802 -58180 35836 -58118
rect 53464 -58000 53498 -57984
rect 53642 -57208 53676 -57192
rect 53642 -58000 53676 -57984
rect 54870 -57166 54904 -57138
rect 53926 -57218 53942 -57184
rect 54718 -57218 54734 -57184
rect 53858 -57246 53892 -57230
rect 53858 -57350 53892 -57334
rect 54768 -57246 54802 -57230
rect 54768 -57350 54802 -57334
rect 53926 -57396 53942 -57362
rect 54718 -57396 54734 -57362
rect 53756 -57476 53790 -57414
rect 55700 -57164 55740 -57138
rect 55126 -57330 55142 -57296
rect 55494 -57330 55510 -57296
rect 54870 -57476 54904 -57414
rect 55046 -57382 55080 -57366
rect 55046 -57432 55080 -57416
rect 55556 -57382 55590 -57366
rect 55556 -57432 55590 -57416
rect 53756 -57510 53852 -57476
rect 54808 -57510 54904 -57476
rect 55126 -57502 55142 -57468
rect 55494 -57502 55510 -57468
rect 53510 -58068 53526 -58034
rect 53614 -58068 53630 -58034
rect 53350 -58136 53384 -58074
rect 53756 -58136 53790 -57510
rect 54870 -57618 54904 -57510
rect 55700 -57618 55706 -57164
rect 54870 -57624 55706 -57618
rect 54870 -57658 55262 -57624
rect 55420 -57658 55706 -57624
rect 55166 -57720 55200 -57658
rect 53350 -58170 53446 -58136
rect 53694 -58170 53790 -58136
rect 53886 -57908 53982 -57874
rect 54956 -57908 55052 -57874
rect 53886 -57970 53920 -57908
rect 55018 -57970 55052 -57908
rect 54065 -58022 54081 -57988
rect 54857 -58022 54873 -57988
rect 53988 -58050 54022 -58034
rect 53988 -58104 54022 -58088
rect 54916 -58050 54950 -58034
rect 54916 -58104 54950 -58088
rect 54065 -58150 54081 -58116
rect 54857 -58150 54873 -58116
rect 25736 -58214 25832 -58180
rect 35740 -58214 35836 -58180
rect 53886 -58230 53920 -58168
rect 55482 -57720 55516 -57658
rect 55280 -57748 55314 -57732
rect 55280 -57940 55314 -57924
rect 55368 -57748 55402 -57732
rect 55368 -57940 55402 -57924
rect 55308 -58008 55324 -57974
rect 55358 -58008 55374 -57974
rect 55166 -58076 55200 -58014
rect 55482 -58076 55516 -58014
rect 55166 -58110 55262 -58076
rect 55420 -58110 55516 -58076
rect 55018 -58230 55052 -58168
rect 56112 -57164 56146 -57102
rect 56350 -56538 56412 -56518
rect 56610 -56538 56706 -56504
rect 56672 -56600 56706 -56538
rect 57303 -56483 57355 -56454
rect 57131 -56555 57165 -56534
rect 57201 -56547 57217 -56513
rect 57251 -56547 57267 -56513
rect 57201 -56589 57267 -56547
rect 57337 -56517 57355 -56483
rect 57303 -56555 57355 -56517
rect 58930 -56410 59026 -56376
rect 59214 -56377 59310 -56376
rect 59662 -56377 59696 -56320
rect 59772 -56294 59866 -56260
rect 60426 -56294 60520 -56260
rect 59772 -56350 59806 -56294
rect 59214 -56410 59696 -56377
rect 58930 -56411 59696 -56410
rect 58930 -56472 58964 -56411
rect 59276 -56472 59310 -56411
rect 59087 -56512 59103 -56478
rect 59137 -56512 59153 -56478
rect 56476 -56640 56492 -56606
rect 56530 -56640 56546 -56606
rect 55866 -57204 55882 -57170
rect 55970 -57204 55986 -57170
rect 55820 -57254 55854 -57238
rect 55820 -58046 55854 -58030
rect 55998 -57254 56032 -57238
rect 55998 -58046 56032 -58030
rect 55866 -58114 55882 -58080
rect 55970 -58114 55986 -58080
rect 55706 -58182 55740 -58120
rect 56430 -56699 56464 -56683
rect 56430 -57491 56464 -57475
rect 56558 -56699 56592 -56683
rect 56558 -57491 56592 -57475
rect 56476 -57568 56492 -57534
rect 56530 -57568 56546 -57534
rect 56316 -57636 56350 -57574
rect 57096 -56623 57125 -56589
rect 57159 -56623 57217 -56589
rect 57251 -56623 57309 -56589
rect 57343 -56623 57372 -56589
rect 59044 -56571 59078 -56555
rect 59044 -56963 59078 -56947
rect 59162 -56571 59196 -56555
rect 59162 -56963 59196 -56947
rect 59087 -57040 59103 -57006
rect 59137 -57040 59153 -57006
rect 60486 -56356 60520 -56294
rect 59942 -56408 59958 -56374
rect 60334 -56408 60350 -56374
rect 59874 -56428 59908 -56412
rect 59874 -56478 59908 -56462
rect 60384 -56428 60418 -56412
rect 60384 -56478 60418 -56462
rect 59942 -56516 59958 -56482
rect 60334 -56516 60350 -56482
rect 59772 -56596 59806 -56540
rect 60486 -56596 60520 -56534
rect 59388 -56630 59476 -56596
rect 59656 -56630 59800 -56596
rect 59958 -56630 60520 -56596
rect 59388 -56690 59422 -56630
rect 59276 -57106 59310 -57046
rect 59530 -56732 59546 -56698
rect 59580 -56732 59596 -56698
rect 59502 -56782 59536 -56766
rect 59502 -56974 59536 -56958
rect 59590 -56782 59624 -56766
rect 59590 -56974 59624 -56958
rect 59530 -57042 59546 -57008
rect 59580 -57042 59596 -57008
rect 58966 -57142 59310 -57106
rect 59388 -57109 59422 -57050
rect 59704 -57109 59738 -56630
rect 60020 -56692 60054 -56630
rect 59846 -56732 59862 -56698
rect 59896 -56732 59912 -56698
rect 59818 -56782 59852 -56766
rect 59818 -56974 59852 -56958
rect 59906 -56782 59940 -56766
rect 59906 -56974 59940 -56958
rect 59846 -57042 59862 -57008
rect 59896 -57042 59912 -57008
rect 61186 -56800 61286 -56790
rect 61186 -56880 61196 -56800
rect 61186 -56890 61286 -56880
rect 60020 -57109 60054 -57048
rect 56672 -57636 56706 -57574
rect 57096 -57599 57125 -57565
rect 57159 -57599 57217 -57565
rect 57251 -57599 57309 -57565
rect 57343 -57599 57372 -57565
rect 56316 -57670 56412 -57636
rect 56610 -57670 56706 -57636
rect 57131 -57654 57165 -57633
rect 57201 -57641 57267 -57599
rect 57201 -57675 57217 -57641
rect 57251 -57675 57267 -57641
rect 57303 -57671 57355 -57633
rect 57131 -57709 57165 -57688
rect 57337 -57705 57355 -57671
rect 59276 -57202 59310 -57142
rect 59387 -57144 60054 -57109
rect 60127 -56954 60161 -56928
rect 60127 -56957 60253 -56954
rect 60161 -56973 60253 -56957
rect 60161 -56991 60203 -56973
rect 60127 -57007 60203 -56991
rect 60237 -57007 60253 -56973
rect 60359 -56960 60409 -56949
rect 60671 -56954 60705 -56928
rect 60359 -56965 60366 -56960
rect 60359 -57000 60366 -56999
rect 60406 -57000 60409 -56960
rect 60127 -57049 60161 -57007
rect 60127 -57141 60161 -57083
rect 60195 -57057 60325 -57041
rect 60195 -57091 60211 -57057
rect 60245 -57091 60325 -57057
rect 60195 -57107 60325 -57091
rect 59387 -57200 59421 -57144
rect 59087 -57242 59103 -57208
rect 59137 -57242 59153 -57208
rect 59044 -57301 59078 -57285
rect 57131 -57743 57264 -57709
rect 57303 -57734 57355 -57705
rect 57117 -57794 57185 -57779
rect 57117 -57844 57118 -57794
rect 57168 -57844 57185 -57794
rect 57117 -57853 57185 -57844
rect 57230 -57794 57264 -57743
rect 57319 -57770 57355 -57734
rect 57230 -57810 57285 -57794
rect 57230 -57844 57251 -57810
rect 57230 -57860 57285 -57844
rect 57319 -57810 57326 -57770
rect 59044 -57693 59078 -57677
rect 59162 -57301 59196 -57285
rect 59162 -57693 59196 -57677
rect 59087 -57770 59103 -57736
rect 59137 -57770 59153 -57736
rect 57230 -57889 57264 -57860
rect 57129 -57923 57264 -57889
rect 57319 -57894 57355 -57810
rect 57129 -57957 57165 -57923
rect 57301 -57944 57355 -57894
rect 58930 -57838 58964 -57776
rect 59529 -57245 59545 -57211
rect 59579 -57245 59595 -57211
rect 59501 -57295 59535 -57279
rect 59501 -57487 59535 -57471
rect 59589 -57295 59623 -57279
rect 59589 -57487 59623 -57471
rect 59529 -57555 59545 -57521
rect 59579 -57555 59595 -57521
rect 59387 -57623 59421 -57570
rect 59703 -57623 59737 -57144
rect 60019 -57205 60053 -57144
rect 59845 -57245 59861 -57211
rect 59895 -57245 59911 -57211
rect 59817 -57295 59851 -57279
rect 59817 -57487 59851 -57471
rect 59905 -57295 59939 -57279
rect 59905 -57487 59939 -57471
rect 59845 -57555 59861 -57521
rect 59895 -57555 59911 -57521
rect 60161 -57175 60203 -57141
rect 60237 -57175 60253 -57141
rect 60127 -57233 60161 -57175
rect 60289 -57209 60325 -57107
rect 60127 -57309 60161 -57267
rect 60195 -57225 60325 -57209
rect 60195 -57259 60211 -57225
rect 60245 -57259 60325 -57225
rect 60195 -57275 60325 -57259
rect 60359 -57050 60409 -57000
rect 60443 -56957 60705 -56954
rect 60443 -56973 60671 -56957
rect 60443 -57007 60459 -56973
rect 60493 -57007 60527 -56973
rect 60561 -57007 60595 -56973
rect 60629 -56991 60671 -56973
rect 60629 -57007 60705 -56991
rect 60359 -57057 60366 -57050
rect 60406 -57090 60409 -57050
rect 60393 -57091 60409 -57090
rect 60359 -57140 60409 -57091
rect 60359 -57141 60366 -57140
rect 60359 -57180 60366 -57175
rect 60406 -57180 60409 -57140
rect 60359 -57220 60409 -57180
rect 60359 -57225 60366 -57220
rect 60359 -57260 60366 -57259
rect 60406 -57260 60409 -57220
rect 60359 -57275 60409 -57260
rect 60443 -57057 60637 -57041
rect 60443 -57091 60459 -57057
rect 60493 -57091 60527 -57057
rect 60561 -57091 60595 -57057
rect 60629 -57091 60637 -57057
rect 60443 -57107 60637 -57091
rect 60671 -57049 60705 -57007
rect 60443 -57209 60477 -57107
rect 60671 -57141 60705 -57083
rect 60511 -57175 60527 -57141
rect 60561 -57175 60595 -57141
rect 60629 -57175 60671 -57141
rect 60443 -57225 60637 -57209
rect 60443 -57259 60459 -57225
rect 60493 -57259 60527 -57225
rect 60561 -57259 60595 -57225
rect 60629 -57259 60637 -57225
rect 60443 -57275 60637 -57259
rect 60671 -57233 60705 -57175
rect 60289 -57309 60325 -57275
rect 60443 -57309 60481 -57275
rect 60671 -57309 60705 -57267
rect 60127 -57325 60204 -57309
rect 60161 -57343 60204 -57325
rect 60238 -57343 60254 -57309
rect 60161 -57359 60254 -57343
rect 60289 -57325 60481 -57309
rect 60289 -57359 60297 -57325
rect 60331 -57359 60369 -57325
rect 60405 -57359 60449 -57325
rect 60579 -57343 60595 -57309
rect 60629 -57325 60705 -57309
rect 60629 -57343 60671 -57325
rect 60579 -57351 60671 -57343
rect 60127 -57388 60161 -57359
rect 60289 -57362 60481 -57359
rect 60671 -57388 60705 -57359
rect 60747 -56954 60781 -56928
rect 60747 -56957 61009 -56954
rect 60781 -56973 61009 -56957
rect 60781 -56991 60823 -56973
rect 60747 -57007 60823 -56991
rect 60857 -57007 60891 -56973
rect 60925 -57007 60959 -56973
rect 60993 -57007 61009 -56973
rect 61043 -56960 61093 -56949
rect 61291 -56954 61325 -56928
rect 61043 -57000 61046 -56960
rect 61086 -56965 61093 -56960
rect 61086 -57000 61093 -56999
rect 60747 -57049 60781 -57007
rect 60747 -57141 60781 -57083
rect 60815 -57057 61009 -57041
rect 60815 -57091 60823 -57057
rect 60857 -57091 60891 -57057
rect 60925 -57091 60959 -57057
rect 60993 -57091 61009 -57057
rect 60815 -57107 61009 -57091
rect 60781 -57175 60823 -57141
rect 60857 -57175 60891 -57141
rect 60925 -57175 60941 -57141
rect 60747 -57233 60781 -57175
rect 60975 -57209 61009 -57107
rect 60747 -57309 60781 -57267
rect 60815 -57225 61009 -57209
rect 60815 -57259 60823 -57225
rect 60857 -57259 60891 -57225
rect 60925 -57259 60959 -57225
rect 60993 -57259 61009 -57225
rect 60815 -57275 61009 -57259
rect 61043 -57050 61093 -57000
rect 61199 -56957 61325 -56954
rect 61199 -56973 61291 -56957
rect 61199 -57007 61215 -56973
rect 61249 -56991 61291 -56973
rect 61249 -57007 61325 -56991
rect 61043 -57090 61046 -57050
rect 61086 -57057 61093 -57050
rect 61043 -57091 61059 -57090
rect 61043 -57140 61093 -57091
rect 61043 -57180 61046 -57140
rect 61086 -57141 61093 -57140
rect 61086 -57180 61093 -57175
rect 61043 -57220 61093 -57180
rect 61043 -57260 61046 -57220
rect 61086 -57225 61093 -57220
rect 61086 -57260 61093 -57259
rect 61043 -57275 61093 -57260
rect 61127 -57057 61257 -57041
rect 61127 -57091 61207 -57057
rect 61241 -57091 61257 -57057
rect 61127 -57107 61257 -57091
rect 61291 -57049 61325 -57007
rect 61127 -57209 61163 -57107
rect 61291 -57141 61325 -57083
rect 61199 -57175 61215 -57141
rect 61249 -57175 61291 -57141
rect 61127 -57225 61257 -57209
rect 61127 -57259 61207 -57225
rect 61241 -57259 61257 -57225
rect 61127 -57275 61257 -57259
rect 61291 -57233 61325 -57175
rect 60971 -57309 61009 -57275
rect 61127 -57309 61163 -57275
rect 61291 -57309 61325 -57267
rect 60747 -57325 60823 -57309
rect 60781 -57343 60823 -57325
rect 60857 -57343 60873 -57309
rect 60781 -57351 60873 -57343
rect 60971 -57324 61163 -57309
rect 60971 -57325 61129 -57324
rect 60747 -57388 60781 -57359
rect 60971 -57359 60980 -57325
rect 61015 -57359 61053 -57325
rect 61088 -57358 61129 -57325
rect 61198 -57343 61214 -57309
rect 61248 -57325 61325 -57309
rect 61248 -57343 61291 -57325
rect 61088 -57359 61163 -57358
rect 61198 -57359 61291 -57343
rect 60971 -57362 61163 -57359
rect 61291 -57388 61325 -57359
rect 60466 -57460 60546 -57440
rect 60466 -57500 60486 -57460
rect 60526 -57500 60546 -57460
rect 60466 -57520 60546 -57500
rect 60606 -57460 60686 -57440
rect 60606 -57500 60626 -57460
rect 60666 -57500 60686 -57460
rect 60606 -57520 60686 -57500
rect 60746 -57460 60826 -57440
rect 60746 -57500 60766 -57460
rect 60806 -57500 60826 -57460
rect 60746 -57520 60826 -57500
rect 60886 -57460 60966 -57440
rect 60886 -57500 60906 -57460
rect 60946 -57500 60966 -57460
rect 60886 -57520 60966 -57500
rect 60019 -57623 60053 -57561
rect 59387 -57657 59476 -57623
rect 59646 -57657 59799 -57623
rect 59957 -57626 60053 -57623
rect 59957 -57657 60520 -57626
rect 59772 -57660 60520 -57657
rect 59772 -57720 59806 -57660
rect 59276 -57838 59310 -57776
rect 58930 -57872 59026 -57838
rect 59214 -57840 59310 -57838
rect 59214 -57872 59696 -57840
rect 58930 -57874 59696 -57872
rect 58930 -57910 58964 -57874
rect 57129 -57991 57131 -57957
rect 57129 -58025 57165 -57991
rect 57129 -58059 57131 -58025
rect 57129 -58075 57165 -58059
rect 57201 -57991 57217 -57957
rect 57251 -57991 57267 -57957
rect 57201 -58025 57267 -57991
rect 57201 -58059 57217 -58025
rect 57251 -58059 57267 -58025
rect 57201 -58109 57267 -58059
rect 57301 -57978 57303 -57944
rect 57337 -57978 57355 -57944
rect 57301 -58025 57355 -57978
rect 57301 -58059 57303 -58025
rect 57337 -58059 57355 -58025
rect 57301 -58075 57355 -58059
rect 59662 -57930 59696 -57874
rect 60486 -57722 60520 -57660
rect 59942 -57774 59958 -57740
rect 60334 -57774 60350 -57740
rect 59874 -57794 59908 -57778
rect 59874 -57844 59908 -57828
rect 60384 -57794 60418 -57778
rect 60384 -57844 60418 -57828
rect 59942 -57882 59958 -57848
rect 60334 -57882 60350 -57848
rect 56112 -58182 56146 -58120
rect 57096 -58143 57125 -58109
rect 57159 -58143 57217 -58109
rect 57251 -58143 57309 -58109
rect 57343 -58143 57372 -58109
rect 55706 -58216 55802 -58182
rect 56050 -58216 56146 -58182
rect 53886 -58264 53982 -58230
rect 54956 -58264 55052 -58230
rect 53886 -58326 53920 -58264
rect 55018 -58326 55052 -58264
rect 55720 -58258 56090 -58216
rect 55720 -58268 56020 -58258
rect 54065 -58378 54081 -58344
rect 54857 -58378 54873 -58344
rect 53988 -58406 54022 -58390
rect 53988 -58460 54022 -58444
rect 54916 -58406 54950 -58390
rect 54916 -58460 54950 -58444
rect 54065 -58506 54081 -58472
rect 54857 -58506 54873 -58472
rect 53886 -58586 53920 -58524
rect 56010 -58408 56020 -58268
rect 56080 -58408 56090 -58258
rect 59109 -57988 59125 -57954
rect 59501 -57988 59517 -57954
rect 59560 -58008 59594 -57992
rect 59560 -58058 59594 -58042
rect 59109 -58096 59125 -58062
rect 59501 -58096 59517 -58062
rect 59032 -58116 59066 -58100
rect 59032 -58166 59066 -58150
rect 59109 -58204 59125 -58170
rect 59501 -58204 59517 -58170
rect 56010 -58418 56090 -58408
rect 59772 -57962 59806 -57900
rect 60486 -57962 60520 -57900
rect 59772 -57996 59866 -57962
rect 60426 -57996 60520 -57962
rect 59662 -58284 59696 -58230
rect 58966 -58300 59026 -58284
rect 58930 -58318 59026 -58300
rect 59600 -58318 59696 -58284
rect 55018 -58586 55052 -58524
rect 53886 -58620 53982 -58586
rect 54956 -58620 55052 -58586
rect 55176 -58478 55272 -58444
rect 55566 -58478 55662 -58444
rect 55176 -58540 55210 -58478
rect 55628 -58540 55662 -58478
rect 55284 -58592 55300 -58558
rect 55476 -58592 55492 -58558
rect 55526 -58602 55560 -58586
rect 55284 -58680 55300 -58646
rect 55476 -58680 55492 -58646
rect 55526 -58652 55560 -58636
rect 55176 -58760 55210 -58698
rect 55628 -58760 55662 -58698
rect 55176 -58794 55272 -58760
rect 55566 -58794 55662 -58760
rect 53896 -60992 53992 -60958
rect 54966 -60992 55062 -60958
rect 53896 -61054 53930 -60992
rect 55028 -61054 55062 -60992
rect 54075 -61106 54091 -61072
rect 54867 -61106 54883 -61072
rect 53998 -61134 54032 -61118
rect 53998 -61188 54032 -61172
rect 54926 -61134 54960 -61118
rect 54926 -61188 54960 -61172
rect 54075 -61234 54091 -61200
rect 54867 -61234 54883 -61200
rect 53896 -61314 53930 -61252
rect 55028 -61314 55062 -61252
rect 55960 -61308 56040 -61298
rect 53896 -61348 53992 -61314
rect 54966 -61348 55062 -61314
rect 53350 -61438 53790 -61404
rect 53350 -61500 53384 -61438
rect 53510 -61540 53526 -61506
rect 53614 -61540 53630 -61506
rect 53464 -61590 53498 -61574
rect 53464 -62382 53498 -62366
rect 53642 -61590 53676 -61574
rect 53642 -62382 53676 -62366
rect 53756 -62064 53790 -61438
rect 53896 -61410 53930 -61348
rect 55028 -61410 55062 -61348
rect 55710 -61354 56040 -61308
rect 54075 -61462 54091 -61428
rect 54867 -61462 54883 -61428
rect 53998 -61490 54032 -61474
rect 53998 -61544 54032 -61528
rect 54926 -61490 54960 -61474
rect 54926 -61544 54960 -61528
rect 54075 -61590 54091 -61556
rect 54867 -61590 54883 -61556
rect 53896 -61670 53930 -61608
rect 55706 -61388 55802 -61354
rect 56050 -61388 56146 -61354
rect 55706 -61450 55740 -61388
rect 55028 -61670 55062 -61608
rect 53896 -61704 53992 -61670
rect 54966 -61704 55062 -61670
rect 55176 -61500 55272 -61466
rect 55430 -61500 55526 -61466
rect 55176 -61562 55210 -61500
rect 55492 -61562 55526 -61500
rect 55318 -61602 55334 -61568
rect 55368 -61602 55384 -61568
rect 55290 -61652 55324 -61636
rect 55290 -61844 55324 -61828
rect 55378 -61652 55412 -61636
rect 55378 -61844 55412 -61828
rect 55176 -61918 55210 -61856
rect 55492 -61918 55526 -61856
rect 54870 -61952 55272 -61918
rect 55430 -61952 55706 -61918
rect 54870 -61958 55706 -61952
rect 54870 -62064 54904 -61958
rect 53756 -62098 53852 -62064
rect 54808 -62098 54904 -62064
rect 53756 -62160 53790 -62098
rect 54870 -62160 54904 -62098
rect 55126 -62108 55142 -62074
rect 55494 -62108 55510 -62074
rect 53926 -62212 53942 -62178
rect 54718 -62212 54734 -62178
rect 53858 -62240 53892 -62224
rect 53858 -62344 53892 -62328
rect 54768 -62240 54802 -62224
rect 54768 -62344 54802 -62328
rect 53926 -62390 53942 -62356
rect 54718 -62390 54734 -62356
rect 53510 -62450 53526 -62416
rect 53614 -62450 53630 -62416
rect 53756 -62470 53790 -62408
rect 55046 -62160 55080 -62144
rect 55046 -62210 55080 -62194
rect 55556 -62160 55590 -62144
rect 55556 -62210 55590 -62194
rect 55126 -62280 55142 -62246
rect 55494 -62280 55510 -62246
rect 54870 -62438 54904 -62408
rect 55700 -62406 55706 -61958
rect 56112 -61450 56146 -61388
rect 58930 -61367 59026 -61333
rect 59600 -61367 59696 -61333
rect 58930 -61410 58964 -61367
rect 58926 -61420 58966 -61410
rect 55866 -61490 55882 -61456
rect 55970 -61490 55986 -61456
rect 55820 -61540 55854 -61524
rect 55820 -62332 55854 -62316
rect 55998 -61540 56032 -61524
rect 55998 -62332 56032 -62316
rect 55866 -62400 55882 -62366
rect 55970 -62400 55986 -62366
rect 55700 -62438 55740 -62406
rect 57096 -61479 57125 -61445
rect 57159 -61479 57217 -61445
rect 57251 -61479 57309 -61445
rect 57343 -61479 57372 -61445
rect 57129 -61529 57165 -61513
rect 57129 -61563 57131 -61529
rect 57129 -61597 57165 -61563
rect 57129 -61631 57131 -61597
rect 57201 -61529 57267 -61479
rect 57201 -61563 57217 -61529
rect 57251 -61563 57267 -61529
rect 57201 -61597 57267 -61563
rect 57201 -61631 57217 -61597
rect 57251 -61631 57267 -61597
rect 57301 -61529 57355 -61513
rect 57301 -61563 57303 -61529
rect 57337 -61563 57355 -61529
rect 57301 -61610 57355 -61563
rect 57129 -61665 57165 -61631
rect 57301 -61644 57303 -61610
rect 57337 -61644 57355 -61610
rect 57129 -61699 57264 -61665
rect 57301 -61694 57355 -61644
rect 57230 -61728 57264 -61699
rect 57117 -61744 57185 -61735
rect 57117 -61794 57118 -61744
rect 57178 -61794 57185 -61744
rect 57117 -61809 57185 -61794
rect 57230 -61744 57285 -61728
rect 57230 -61778 57251 -61744
rect 57230 -61794 57285 -61778
rect 57319 -61740 57355 -61694
rect 59662 -61429 59696 -61367
rect 59109 -61481 59125 -61447
rect 59501 -61481 59517 -61447
rect 59560 -61501 59594 -61485
rect 59560 -61551 59594 -61535
rect 59109 -61589 59125 -61555
rect 59501 -61589 59517 -61555
rect 59032 -61609 59066 -61593
rect 59032 -61659 59066 -61643
rect 59109 -61697 59125 -61663
rect 59501 -61697 59517 -61663
rect 58926 -61740 58966 -61720
rect 57319 -61780 57326 -61740
rect 58930 -61776 58964 -61740
rect 57230 -61845 57264 -61794
rect 57131 -61879 57264 -61845
rect 57319 -61854 57355 -61780
rect 57131 -61900 57165 -61879
rect 56316 -61918 56412 -61904
rect 54830 -62448 55830 -62438
rect 54830 -62470 55030 -62448
rect 53756 -62504 53852 -62470
rect 54808 -62504 55030 -62470
rect 53510 -62558 53526 -62524
rect 53614 -62558 53630 -62524
rect 53756 -62566 53790 -62504
rect 54830 -62528 55030 -62504
rect 55110 -62468 55740 -62448
rect 55810 -62468 55830 -62448
rect 56112 -62468 56146 -62406
rect 55110 -62508 55160 -62468
rect 55600 -62508 55740 -62468
rect 56050 -62502 56146 -62468
rect 55110 -62528 55740 -62508
rect 55810 -62528 55830 -62502
rect 54830 -62538 55830 -62528
rect 53464 -62608 53498 -62592
rect 53464 -63400 53498 -63384
rect 53642 -62608 53676 -62592
rect 53642 -63400 53676 -63384
rect 54870 -62566 54904 -62538
rect 53926 -62618 53942 -62584
rect 54718 -62618 54734 -62584
rect 53858 -62646 53892 -62630
rect 53858 -62750 53892 -62734
rect 54768 -62646 54802 -62630
rect 54768 -62750 54802 -62734
rect 53926 -62796 53942 -62762
rect 54718 -62796 54734 -62762
rect 53756 -62876 53790 -62814
rect 55700 -62564 55740 -62538
rect 55126 -62730 55142 -62696
rect 55494 -62730 55510 -62696
rect 54870 -62876 54904 -62814
rect 55046 -62782 55080 -62766
rect 55046 -62832 55080 -62816
rect 55556 -62782 55590 -62766
rect 55556 -62832 55590 -62816
rect 53756 -62910 53852 -62876
rect 54808 -62910 54904 -62876
rect 55126 -62902 55142 -62868
rect 55494 -62902 55510 -62868
rect 53510 -63468 53526 -63434
rect 53614 -63468 53630 -63434
rect 53350 -63536 53384 -63474
rect 53756 -63536 53790 -62910
rect 54870 -63018 54904 -62910
rect 55700 -63018 55706 -62564
rect 54870 -63024 55706 -63018
rect 54870 -63058 55262 -63024
rect 55420 -63058 55706 -63024
rect 55166 -63120 55200 -63058
rect 53350 -63570 53446 -63536
rect 53694 -63570 53790 -63536
rect 53886 -63308 53982 -63274
rect 54956 -63308 55052 -63274
rect 53886 -63370 53920 -63308
rect 55018 -63370 55052 -63308
rect 54065 -63422 54081 -63388
rect 54857 -63422 54873 -63388
rect 53988 -63450 54022 -63434
rect 53988 -63504 54022 -63488
rect 54916 -63450 54950 -63434
rect 54916 -63504 54950 -63488
rect 54065 -63550 54081 -63516
rect 54857 -63550 54873 -63516
rect 53886 -63630 53920 -63568
rect 55482 -63120 55516 -63058
rect 55280 -63148 55314 -63132
rect 55280 -63340 55314 -63324
rect 55368 -63148 55402 -63132
rect 55368 -63340 55402 -63324
rect 55308 -63408 55324 -63374
rect 55358 -63408 55374 -63374
rect 55166 -63476 55200 -63414
rect 55482 -63476 55516 -63414
rect 55166 -63510 55262 -63476
rect 55420 -63510 55516 -63476
rect 55018 -63630 55052 -63568
rect 56112 -62564 56146 -62502
rect 56350 -61938 56412 -61918
rect 56610 -61938 56706 -61904
rect 56672 -62000 56706 -61938
rect 57303 -61883 57355 -61854
rect 57131 -61955 57165 -61934
rect 57201 -61947 57217 -61913
rect 57251 -61947 57267 -61913
rect 57201 -61989 57267 -61947
rect 57337 -61917 57355 -61883
rect 57303 -61955 57355 -61917
rect 58930 -61810 59026 -61776
rect 59214 -61777 59310 -61776
rect 59662 -61777 59696 -61720
rect 59772 -61694 59866 -61660
rect 60426 -61694 60520 -61660
rect 59772 -61750 59806 -61694
rect 59214 -61810 59696 -61777
rect 58930 -61811 59696 -61810
rect 58930 -61872 58964 -61811
rect 59276 -61872 59310 -61811
rect 59087 -61912 59103 -61878
rect 59137 -61912 59153 -61878
rect 56476 -62040 56492 -62006
rect 56530 -62040 56546 -62006
rect 55866 -62604 55882 -62570
rect 55970 -62604 55986 -62570
rect 55820 -62654 55854 -62638
rect 55820 -63446 55854 -63430
rect 55998 -62654 56032 -62638
rect 55998 -63446 56032 -63430
rect 55866 -63514 55882 -63480
rect 55970 -63514 55986 -63480
rect 55706 -63582 55740 -63520
rect 56430 -62099 56464 -62083
rect 56430 -62891 56464 -62875
rect 56558 -62099 56592 -62083
rect 56558 -62891 56592 -62875
rect 56476 -62968 56492 -62934
rect 56530 -62968 56546 -62934
rect 56316 -63036 56350 -62974
rect 57096 -62023 57125 -61989
rect 57159 -62023 57217 -61989
rect 57251 -62023 57309 -61989
rect 57343 -62023 57372 -61989
rect 59044 -61971 59078 -61955
rect 59044 -62363 59078 -62347
rect 59162 -61971 59196 -61955
rect 59162 -62363 59196 -62347
rect 59087 -62440 59103 -62406
rect 59137 -62440 59153 -62406
rect 60486 -61756 60520 -61694
rect 59942 -61808 59958 -61774
rect 60334 -61808 60350 -61774
rect 59874 -61828 59908 -61812
rect 59874 -61878 59908 -61862
rect 60384 -61828 60418 -61812
rect 60384 -61878 60418 -61862
rect 59942 -61916 59958 -61882
rect 60334 -61916 60350 -61882
rect 59772 -61996 59806 -61940
rect 60486 -61996 60520 -61934
rect 59388 -62030 59476 -61996
rect 59656 -62030 59800 -61996
rect 59958 -62030 60520 -61996
rect 59388 -62090 59422 -62030
rect 59276 -62506 59310 -62446
rect 59530 -62132 59546 -62098
rect 59580 -62132 59596 -62098
rect 59502 -62182 59536 -62166
rect 59502 -62374 59536 -62358
rect 59590 -62182 59624 -62166
rect 59590 -62374 59624 -62358
rect 59530 -62442 59546 -62408
rect 59580 -62442 59596 -62408
rect 58966 -62542 59310 -62506
rect 59388 -62509 59422 -62450
rect 59704 -62509 59738 -62030
rect 60020 -62092 60054 -62030
rect 59846 -62132 59862 -62098
rect 59896 -62132 59912 -62098
rect 59818 -62182 59852 -62166
rect 59818 -62374 59852 -62358
rect 59906 -62182 59940 -62166
rect 59906 -62374 59940 -62358
rect 59846 -62442 59862 -62408
rect 59896 -62442 59912 -62408
rect 61186 -62200 61286 -62190
rect 61186 -62280 61196 -62200
rect 61186 -62290 61286 -62280
rect 60020 -62509 60054 -62448
rect 56672 -63036 56706 -62974
rect 57096 -62999 57125 -62965
rect 57159 -62999 57217 -62965
rect 57251 -62999 57309 -62965
rect 57343 -62999 57372 -62965
rect 56316 -63070 56412 -63036
rect 56610 -63070 56706 -63036
rect 57131 -63054 57165 -63033
rect 57201 -63041 57267 -62999
rect 57201 -63075 57217 -63041
rect 57251 -63075 57267 -63041
rect 57303 -63071 57355 -63033
rect 57131 -63109 57165 -63088
rect 57337 -63105 57355 -63071
rect 59276 -62602 59310 -62542
rect 59387 -62544 60054 -62509
rect 60127 -62354 60161 -62328
rect 60127 -62357 60253 -62354
rect 60161 -62373 60253 -62357
rect 60161 -62391 60203 -62373
rect 60127 -62407 60203 -62391
rect 60237 -62407 60253 -62373
rect 60359 -62360 60409 -62349
rect 60671 -62354 60705 -62328
rect 60359 -62365 60366 -62360
rect 60359 -62400 60366 -62399
rect 60406 -62400 60409 -62360
rect 60127 -62449 60161 -62407
rect 60127 -62541 60161 -62483
rect 60195 -62457 60325 -62441
rect 60195 -62491 60211 -62457
rect 60245 -62491 60325 -62457
rect 60195 -62507 60325 -62491
rect 59387 -62600 59421 -62544
rect 59087 -62642 59103 -62608
rect 59137 -62642 59153 -62608
rect 59044 -62701 59078 -62685
rect 57131 -63143 57264 -63109
rect 57303 -63134 57355 -63105
rect 57117 -63194 57185 -63179
rect 57117 -63244 57118 -63194
rect 57168 -63244 57185 -63194
rect 57117 -63253 57185 -63244
rect 57230 -63194 57264 -63143
rect 57319 -63170 57355 -63134
rect 57230 -63210 57285 -63194
rect 57230 -63244 57251 -63210
rect 57230 -63260 57285 -63244
rect 57319 -63210 57326 -63170
rect 59044 -63093 59078 -63077
rect 59162 -62701 59196 -62685
rect 59162 -63093 59196 -63077
rect 59087 -63170 59103 -63136
rect 59137 -63170 59153 -63136
rect 57230 -63289 57264 -63260
rect 57129 -63323 57264 -63289
rect 57319 -63294 57355 -63210
rect 57129 -63357 57165 -63323
rect 57301 -63344 57355 -63294
rect 58930 -63238 58964 -63176
rect 59529 -62645 59545 -62611
rect 59579 -62645 59595 -62611
rect 59501 -62695 59535 -62679
rect 59501 -62887 59535 -62871
rect 59589 -62695 59623 -62679
rect 59589 -62887 59623 -62871
rect 59529 -62955 59545 -62921
rect 59579 -62955 59595 -62921
rect 59387 -63023 59421 -62970
rect 59703 -63023 59737 -62544
rect 60019 -62605 60053 -62544
rect 59845 -62645 59861 -62611
rect 59895 -62645 59911 -62611
rect 59817 -62695 59851 -62679
rect 59817 -62887 59851 -62871
rect 59905 -62695 59939 -62679
rect 59905 -62887 59939 -62871
rect 59845 -62955 59861 -62921
rect 59895 -62955 59911 -62921
rect 60161 -62575 60203 -62541
rect 60237 -62575 60253 -62541
rect 60127 -62633 60161 -62575
rect 60289 -62609 60325 -62507
rect 60127 -62709 60161 -62667
rect 60195 -62625 60325 -62609
rect 60195 -62659 60211 -62625
rect 60245 -62659 60325 -62625
rect 60195 -62675 60325 -62659
rect 60359 -62450 60409 -62400
rect 60443 -62357 60705 -62354
rect 60443 -62373 60671 -62357
rect 60443 -62407 60459 -62373
rect 60493 -62407 60527 -62373
rect 60561 -62407 60595 -62373
rect 60629 -62391 60671 -62373
rect 60629 -62407 60705 -62391
rect 60359 -62457 60366 -62450
rect 60406 -62490 60409 -62450
rect 60393 -62491 60409 -62490
rect 60359 -62540 60409 -62491
rect 60359 -62541 60366 -62540
rect 60359 -62580 60366 -62575
rect 60406 -62580 60409 -62540
rect 60359 -62620 60409 -62580
rect 60359 -62625 60366 -62620
rect 60359 -62660 60366 -62659
rect 60406 -62660 60409 -62620
rect 60359 -62675 60409 -62660
rect 60443 -62457 60637 -62441
rect 60443 -62491 60459 -62457
rect 60493 -62491 60527 -62457
rect 60561 -62491 60595 -62457
rect 60629 -62491 60637 -62457
rect 60443 -62507 60637 -62491
rect 60671 -62449 60705 -62407
rect 60443 -62609 60477 -62507
rect 60671 -62541 60705 -62483
rect 60511 -62575 60527 -62541
rect 60561 -62575 60595 -62541
rect 60629 -62575 60671 -62541
rect 60443 -62625 60637 -62609
rect 60443 -62659 60459 -62625
rect 60493 -62659 60527 -62625
rect 60561 -62659 60595 -62625
rect 60629 -62659 60637 -62625
rect 60443 -62675 60637 -62659
rect 60671 -62633 60705 -62575
rect 60289 -62709 60325 -62675
rect 60443 -62709 60481 -62675
rect 60671 -62709 60705 -62667
rect 60127 -62725 60204 -62709
rect 60161 -62743 60204 -62725
rect 60238 -62743 60254 -62709
rect 60161 -62759 60254 -62743
rect 60289 -62725 60481 -62709
rect 60289 -62759 60297 -62725
rect 60331 -62759 60369 -62725
rect 60405 -62759 60449 -62725
rect 60579 -62743 60595 -62709
rect 60629 -62725 60705 -62709
rect 60629 -62743 60671 -62725
rect 60579 -62751 60671 -62743
rect 60127 -62788 60161 -62759
rect 60289 -62762 60481 -62759
rect 60671 -62788 60705 -62759
rect 60747 -62354 60781 -62328
rect 60747 -62357 61009 -62354
rect 60781 -62373 61009 -62357
rect 60781 -62391 60823 -62373
rect 60747 -62407 60823 -62391
rect 60857 -62407 60891 -62373
rect 60925 -62407 60959 -62373
rect 60993 -62407 61009 -62373
rect 61043 -62360 61093 -62349
rect 61291 -62354 61325 -62328
rect 61043 -62400 61046 -62360
rect 61086 -62365 61093 -62360
rect 61086 -62400 61093 -62399
rect 60747 -62449 60781 -62407
rect 60747 -62541 60781 -62483
rect 60815 -62457 61009 -62441
rect 60815 -62491 60823 -62457
rect 60857 -62491 60891 -62457
rect 60925 -62491 60959 -62457
rect 60993 -62491 61009 -62457
rect 60815 -62507 61009 -62491
rect 60781 -62575 60823 -62541
rect 60857 -62575 60891 -62541
rect 60925 -62575 60941 -62541
rect 60747 -62633 60781 -62575
rect 60975 -62609 61009 -62507
rect 60747 -62709 60781 -62667
rect 60815 -62625 61009 -62609
rect 60815 -62659 60823 -62625
rect 60857 -62659 60891 -62625
rect 60925 -62659 60959 -62625
rect 60993 -62659 61009 -62625
rect 60815 -62675 61009 -62659
rect 61043 -62450 61093 -62400
rect 61199 -62357 61325 -62354
rect 61199 -62373 61291 -62357
rect 61199 -62407 61215 -62373
rect 61249 -62391 61291 -62373
rect 61249 -62407 61325 -62391
rect 61043 -62490 61046 -62450
rect 61086 -62457 61093 -62450
rect 61043 -62491 61059 -62490
rect 61043 -62540 61093 -62491
rect 61043 -62580 61046 -62540
rect 61086 -62541 61093 -62540
rect 61086 -62580 61093 -62575
rect 61043 -62620 61093 -62580
rect 61043 -62660 61046 -62620
rect 61086 -62625 61093 -62620
rect 61086 -62660 61093 -62659
rect 61043 -62675 61093 -62660
rect 61127 -62457 61257 -62441
rect 61127 -62491 61207 -62457
rect 61241 -62491 61257 -62457
rect 61127 -62507 61257 -62491
rect 61291 -62449 61325 -62407
rect 61127 -62609 61163 -62507
rect 61291 -62541 61325 -62483
rect 61199 -62575 61215 -62541
rect 61249 -62575 61291 -62541
rect 61127 -62625 61257 -62609
rect 61127 -62659 61207 -62625
rect 61241 -62659 61257 -62625
rect 61127 -62675 61257 -62659
rect 61291 -62633 61325 -62575
rect 60971 -62709 61009 -62675
rect 61127 -62709 61163 -62675
rect 61291 -62709 61325 -62667
rect 60747 -62725 60823 -62709
rect 60781 -62743 60823 -62725
rect 60857 -62743 60873 -62709
rect 60781 -62751 60873 -62743
rect 60971 -62724 61163 -62709
rect 60971 -62725 61129 -62724
rect 60747 -62788 60781 -62759
rect 60971 -62759 60980 -62725
rect 61015 -62759 61053 -62725
rect 61088 -62758 61129 -62725
rect 61198 -62743 61214 -62709
rect 61248 -62725 61325 -62709
rect 61248 -62743 61291 -62725
rect 61088 -62759 61163 -62758
rect 61198 -62759 61291 -62743
rect 60971 -62762 61163 -62759
rect 61291 -62788 61325 -62759
rect 60466 -62860 60546 -62840
rect 60466 -62900 60486 -62860
rect 60526 -62900 60546 -62860
rect 60466 -62920 60546 -62900
rect 60606 -62860 60686 -62840
rect 60606 -62900 60626 -62860
rect 60666 -62900 60686 -62860
rect 60606 -62920 60686 -62900
rect 60746 -62860 60826 -62840
rect 60746 -62900 60766 -62860
rect 60806 -62900 60826 -62860
rect 60746 -62920 60826 -62900
rect 60886 -62860 60966 -62840
rect 60886 -62900 60906 -62860
rect 60946 -62900 60966 -62860
rect 60886 -62920 60966 -62900
rect 60019 -63023 60053 -62961
rect 59387 -63057 59476 -63023
rect 59646 -63057 59799 -63023
rect 59957 -63026 60053 -63023
rect 59957 -63057 60520 -63026
rect 59772 -63060 60520 -63057
rect 59772 -63120 59806 -63060
rect 59276 -63238 59310 -63176
rect 58930 -63272 59026 -63238
rect 59214 -63240 59310 -63238
rect 59214 -63272 59696 -63240
rect 58930 -63274 59696 -63272
rect 58930 -63310 58964 -63274
rect 57129 -63391 57131 -63357
rect 57129 -63425 57165 -63391
rect 57129 -63459 57131 -63425
rect 57129 -63475 57165 -63459
rect 57201 -63391 57217 -63357
rect 57251 -63391 57267 -63357
rect 57201 -63425 57267 -63391
rect 57201 -63459 57217 -63425
rect 57251 -63459 57267 -63425
rect 57201 -63509 57267 -63459
rect 57301 -63378 57303 -63344
rect 57337 -63378 57355 -63344
rect 57301 -63425 57355 -63378
rect 57301 -63459 57303 -63425
rect 57337 -63459 57355 -63425
rect 57301 -63475 57355 -63459
rect 59662 -63330 59696 -63274
rect 60486 -63122 60520 -63060
rect 59942 -63174 59958 -63140
rect 60334 -63174 60350 -63140
rect 59874 -63194 59908 -63178
rect 59874 -63244 59908 -63228
rect 60384 -63194 60418 -63178
rect 60384 -63244 60418 -63228
rect 59942 -63282 59958 -63248
rect 60334 -63282 60350 -63248
rect 56112 -63582 56146 -63520
rect 57096 -63543 57125 -63509
rect 57159 -63543 57217 -63509
rect 57251 -63543 57309 -63509
rect 57343 -63543 57372 -63509
rect 55706 -63616 55802 -63582
rect 56050 -63616 56146 -63582
rect 53886 -63664 53982 -63630
rect 54956 -63664 55052 -63630
rect 53886 -63726 53920 -63664
rect 55018 -63726 55052 -63664
rect 55720 -63658 56090 -63616
rect 55720 -63668 56020 -63658
rect 54065 -63778 54081 -63744
rect 54857 -63778 54873 -63744
rect 53988 -63806 54022 -63790
rect 53988 -63860 54022 -63844
rect 54916 -63806 54950 -63790
rect 54916 -63860 54950 -63844
rect 54065 -63906 54081 -63872
rect 54857 -63906 54873 -63872
rect 53886 -63986 53920 -63924
rect 56010 -63808 56020 -63668
rect 56080 -63808 56090 -63658
rect 59109 -63388 59125 -63354
rect 59501 -63388 59517 -63354
rect 59560 -63408 59594 -63392
rect 59560 -63458 59594 -63442
rect 59109 -63496 59125 -63462
rect 59501 -63496 59517 -63462
rect 59032 -63516 59066 -63500
rect 59032 -63566 59066 -63550
rect 59109 -63604 59125 -63570
rect 59501 -63604 59517 -63570
rect 56010 -63818 56090 -63808
rect 59772 -63362 59806 -63300
rect 60486 -63362 60520 -63300
rect 59772 -63396 59866 -63362
rect 60426 -63396 60520 -63362
rect 59662 -63684 59696 -63630
rect 58966 -63700 59026 -63684
rect 58930 -63718 59026 -63700
rect 59600 -63718 59696 -63684
rect 55018 -63986 55052 -63924
rect 53886 -64020 53982 -63986
rect 54956 -64020 55052 -63986
rect 55176 -63878 55272 -63844
rect 55566 -63878 55662 -63844
rect 55176 -63940 55210 -63878
rect 55628 -63940 55662 -63878
rect 55284 -63992 55300 -63958
rect 55476 -63992 55492 -63958
rect 55526 -64002 55560 -63986
rect 55284 -64080 55300 -64046
rect 55476 -64080 55492 -64046
rect 55526 -64052 55560 -64036
rect 55176 -64160 55210 -64098
rect 55628 -64160 55662 -64098
rect 55176 -64194 55272 -64160
rect 55566 -64194 55662 -64160
rect 53896 -66392 53992 -66358
rect 54966 -66392 55062 -66358
rect 53896 -66454 53930 -66392
rect 55028 -66454 55062 -66392
rect 54075 -66506 54091 -66472
rect 54867 -66506 54883 -66472
rect 53998 -66534 54032 -66518
rect 53998 -66588 54032 -66572
rect 54926 -66534 54960 -66518
rect 54926 -66588 54960 -66572
rect 54075 -66634 54091 -66600
rect 54867 -66634 54883 -66600
rect 53896 -66714 53930 -66652
rect 55028 -66714 55062 -66652
rect 55960 -66708 56040 -66698
rect 53896 -66748 53992 -66714
rect 54966 -66748 55062 -66714
rect 53350 -66838 53790 -66804
rect 53350 -66900 53384 -66838
rect 53510 -66940 53526 -66906
rect 53614 -66940 53630 -66906
rect 53464 -66990 53498 -66974
rect 53464 -67782 53498 -67766
rect 53642 -66990 53676 -66974
rect 53642 -67782 53676 -67766
rect 53756 -67464 53790 -66838
rect 53896 -66810 53930 -66748
rect 55028 -66810 55062 -66748
rect 55710 -66754 56040 -66708
rect 54075 -66862 54091 -66828
rect 54867 -66862 54883 -66828
rect 53998 -66890 54032 -66874
rect 53998 -66944 54032 -66928
rect 54926 -66890 54960 -66874
rect 54926 -66944 54960 -66928
rect 54075 -66990 54091 -66956
rect 54867 -66990 54883 -66956
rect 53896 -67070 53930 -67008
rect 55706 -66788 55802 -66754
rect 56050 -66788 56146 -66754
rect 55706 -66850 55740 -66788
rect 55028 -67070 55062 -67008
rect 53896 -67104 53992 -67070
rect 54966 -67104 55062 -67070
rect 55176 -66900 55272 -66866
rect 55430 -66900 55526 -66866
rect 55176 -66962 55210 -66900
rect 55492 -66962 55526 -66900
rect 55318 -67002 55334 -66968
rect 55368 -67002 55384 -66968
rect 55290 -67052 55324 -67036
rect 55290 -67244 55324 -67228
rect 55378 -67052 55412 -67036
rect 55378 -67244 55412 -67228
rect 55176 -67318 55210 -67256
rect 55492 -67318 55526 -67256
rect 54870 -67352 55272 -67318
rect 55430 -67352 55706 -67318
rect 54870 -67358 55706 -67352
rect 54870 -67464 54904 -67358
rect 53756 -67498 53852 -67464
rect 54808 -67498 54904 -67464
rect 53756 -67560 53790 -67498
rect 54870 -67560 54904 -67498
rect 55126 -67508 55142 -67474
rect 55494 -67508 55510 -67474
rect 53926 -67612 53942 -67578
rect 54718 -67612 54734 -67578
rect 53858 -67640 53892 -67624
rect 53858 -67744 53892 -67728
rect 54768 -67640 54802 -67624
rect 54768 -67744 54802 -67728
rect 53926 -67790 53942 -67756
rect 54718 -67790 54734 -67756
rect 53510 -67850 53526 -67816
rect 53614 -67850 53630 -67816
rect 53756 -67870 53790 -67808
rect 55046 -67560 55080 -67544
rect 55046 -67610 55080 -67594
rect 55556 -67560 55590 -67544
rect 55556 -67610 55590 -67594
rect 55126 -67680 55142 -67646
rect 55494 -67680 55510 -67646
rect 54870 -67838 54904 -67808
rect 55700 -67806 55706 -67358
rect 56112 -66850 56146 -66788
rect 58930 -66767 59026 -66733
rect 59600 -66767 59696 -66733
rect 58930 -66810 58964 -66767
rect 58926 -66820 58966 -66810
rect 55866 -66890 55882 -66856
rect 55970 -66890 55986 -66856
rect 55820 -66940 55854 -66924
rect 55820 -67732 55854 -67716
rect 55998 -66940 56032 -66924
rect 55998 -67732 56032 -67716
rect 55866 -67800 55882 -67766
rect 55970 -67800 55986 -67766
rect 55700 -67838 55740 -67806
rect 57096 -66879 57125 -66845
rect 57159 -66879 57217 -66845
rect 57251 -66879 57309 -66845
rect 57343 -66879 57372 -66845
rect 57129 -66929 57165 -66913
rect 57129 -66963 57131 -66929
rect 57129 -66997 57165 -66963
rect 57129 -67031 57131 -66997
rect 57201 -66929 57267 -66879
rect 57201 -66963 57217 -66929
rect 57251 -66963 57267 -66929
rect 57201 -66997 57267 -66963
rect 57201 -67031 57217 -66997
rect 57251 -67031 57267 -66997
rect 57301 -66929 57355 -66913
rect 57301 -66963 57303 -66929
rect 57337 -66963 57355 -66929
rect 57301 -67010 57355 -66963
rect 57129 -67065 57165 -67031
rect 57301 -67044 57303 -67010
rect 57337 -67044 57355 -67010
rect 57129 -67099 57264 -67065
rect 57301 -67094 57355 -67044
rect 57230 -67128 57264 -67099
rect 57117 -67144 57185 -67135
rect 57117 -67194 57118 -67144
rect 57178 -67194 57185 -67144
rect 57117 -67209 57185 -67194
rect 57230 -67144 57285 -67128
rect 57230 -67178 57251 -67144
rect 57230 -67194 57285 -67178
rect 57319 -67140 57355 -67094
rect 59662 -66829 59696 -66767
rect 59109 -66881 59125 -66847
rect 59501 -66881 59517 -66847
rect 59560 -66901 59594 -66885
rect 59560 -66951 59594 -66935
rect 59109 -66989 59125 -66955
rect 59501 -66989 59517 -66955
rect 59032 -67009 59066 -66993
rect 59032 -67059 59066 -67043
rect 59109 -67097 59125 -67063
rect 59501 -67097 59517 -67063
rect 58926 -67140 58966 -67120
rect 57319 -67180 57326 -67140
rect 58930 -67176 58964 -67140
rect 57230 -67245 57264 -67194
rect 57131 -67279 57264 -67245
rect 57319 -67254 57355 -67180
rect 57131 -67300 57165 -67279
rect 56316 -67318 56412 -67304
rect 54830 -67848 55830 -67838
rect 54830 -67870 55030 -67848
rect 53756 -67904 53852 -67870
rect 54808 -67904 55030 -67870
rect 53510 -67958 53526 -67924
rect 53614 -67958 53630 -67924
rect 53756 -67966 53790 -67904
rect 54830 -67928 55030 -67904
rect 55110 -67868 55740 -67848
rect 55810 -67868 55830 -67848
rect 56112 -67868 56146 -67806
rect 55110 -67908 55160 -67868
rect 55600 -67908 55740 -67868
rect 56050 -67902 56146 -67868
rect 55110 -67928 55740 -67908
rect 55810 -67928 55830 -67902
rect 54830 -67938 55830 -67928
rect 53464 -68008 53498 -67992
rect 53464 -68800 53498 -68784
rect 53642 -68008 53676 -67992
rect 53642 -68800 53676 -68784
rect 54870 -67966 54904 -67938
rect 53926 -68018 53942 -67984
rect 54718 -68018 54734 -67984
rect 53858 -68046 53892 -68030
rect 53858 -68150 53892 -68134
rect 54768 -68046 54802 -68030
rect 54768 -68150 54802 -68134
rect 53926 -68196 53942 -68162
rect 54718 -68196 54734 -68162
rect 53756 -68276 53790 -68214
rect 55700 -67964 55740 -67938
rect 55126 -68130 55142 -68096
rect 55494 -68130 55510 -68096
rect 54870 -68276 54904 -68214
rect 55046 -68182 55080 -68166
rect 55046 -68232 55080 -68216
rect 55556 -68182 55590 -68166
rect 55556 -68232 55590 -68216
rect 53756 -68310 53852 -68276
rect 54808 -68310 54904 -68276
rect 55126 -68302 55142 -68268
rect 55494 -68302 55510 -68268
rect 53510 -68868 53526 -68834
rect 53614 -68868 53630 -68834
rect 53350 -68936 53384 -68874
rect 53756 -68936 53790 -68310
rect 54870 -68418 54904 -68310
rect 55700 -68418 55706 -67964
rect 54870 -68424 55706 -68418
rect 54870 -68458 55262 -68424
rect 55420 -68458 55706 -68424
rect 55166 -68520 55200 -68458
rect 53350 -68970 53446 -68936
rect 53694 -68970 53790 -68936
rect 53886 -68708 53982 -68674
rect 54956 -68708 55052 -68674
rect 53886 -68770 53920 -68708
rect 55018 -68770 55052 -68708
rect 54065 -68822 54081 -68788
rect 54857 -68822 54873 -68788
rect 53988 -68850 54022 -68834
rect 53988 -68904 54022 -68888
rect 54916 -68850 54950 -68834
rect 54916 -68904 54950 -68888
rect 54065 -68950 54081 -68916
rect 54857 -68950 54873 -68916
rect 53886 -69030 53920 -68968
rect 55482 -68520 55516 -68458
rect 55280 -68548 55314 -68532
rect 55280 -68740 55314 -68724
rect 55368 -68548 55402 -68532
rect 55368 -68740 55402 -68724
rect 55308 -68808 55324 -68774
rect 55358 -68808 55374 -68774
rect 55166 -68876 55200 -68814
rect 55482 -68876 55516 -68814
rect 55166 -68910 55262 -68876
rect 55420 -68910 55516 -68876
rect 55018 -69030 55052 -68968
rect 56112 -67964 56146 -67902
rect 56350 -67338 56412 -67318
rect 56610 -67338 56706 -67304
rect 56672 -67400 56706 -67338
rect 57303 -67283 57355 -67254
rect 57131 -67355 57165 -67334
rect 57201 -67347 57217 -67313
rect 57251 -67347 57267 -67313
rect 57201 -67389 57267 -67347
rect 57337 -67317 57355 -67283
rect 57303 -67355 57355 -67317
rect 58930 -67210 59026 -67176
rect 59214 -67177 59310 -67176
rect 59662 -67177 59696 -67120
rect 59772 -67094 59866 -67060
rect 60426 -67094 60520 -67060
rect 59772 -67150 59806 -67094
rect 59214 -67210 59696 -67177
rect 58930 -67211 59696 -67210
rect 58930 -67272 58964 -67211
rect 59276 -67272 59310 -67211
rect 59087 -67312 59103 -67278
rect 59137 -67312 59153 -67278
rect 56476 -67440 56492 -67406
rect 56530 -67440 56546 -67406
rect 55866 -68004 55882 -67970
rect 55970 -68004 55986 -67970
rect 55820 -68054 55854 -68038
rect 55820 -68846 55854 -68830
rect 55998 -68054 56032 -68038
rect 55998 -68846 56032 -68830
rect 55866 -68914 55882 -68880
rect 55970 -68914 55986 -68880
rect 55706 -68982 55740 -68920
rect 56430 -67499 56464 -67483
rect 56430 -68291 56464 -68275
rect 56558 -67499 56592 -67483
rect 56558 -68291 56592 -68275
rect 56476 -68368 56492 -68334
rect 56530 -68368 56546 -68334
rect 56316 -68436 56350 -68374
rect 57096 -67423 57125 -67389
rect 57159 -67423 57217 -67389
rect 57251 -67423 57309 -67389
rect 57343 -67423 57372 -67389
rect 59044 -67371 59078 -67355
rect 59044 -67763 59078 -67747
rect 59162 -67371 59196 -67355
rect 59162 -67763 59196 -67747
rect 59087 -67840 59103 -67806
rect 59137 -67840 59153 -67806
rect 60486 -67156 60520 -67094
rect 59942 -67208 59958 -67174
rect 60334 -67208 60350 -67174
rect 59874 -67228 59908 -67212
rect 59874 -67278 59908 -67262
rect 60384 -67228 60418 -67212
rect 60384 -67278 60418 -67262
rect 59942 -67316 59958 -67282
rect 60334 -67316 60350 -67282
rect 59772 -67396 59806 -67340
rect 60486 -67396 60520 -67334
rect 59388 -67430 59476 -67396
rect 59656 -67430 59800 -67396
rect 59958 -67430 60520 -67396
rect 59388 -67490 59422 -67430
rect 59276 -67906 59310 -67846
rect 59530 -67532 59546 -67498
rect 59580 -67532 59596 -67498
rect 59502 -67582 59536 -67566
rect 59502 -67774 59536 -67758
rect 59590 -67582 59624 -67566
rect 59590 -67774 59624 -67758
rect 59530 -67842 59546 -67808
rect 59580 -67842 59596 -67808
rect 58966 -67942 59310 -67906
rect 59388 -67909 59422 -67850
rect 59704 -67909 59738 -67430
rect 60020 -67492 60054 -67430
rect 59846 -67532 59862 -67498
rect 59896 -67532 59912 -67498
rect 59818 -67582 59852 -67566
rect 59818 -67774 59852 -67758
rect 59906 -67582 59940 -67566
rect 59906 -67774 59940 -67758
rect 59846 -67842 59862 -67808
rect 59896 -67842 59912 -67808
rect 61186 -67600 61286 -67590
rect 61186 -67680 61196 -67600
rect 61186 -67690 61286 -67680
rect 60020 -67909 60054 -67848
rect 56672 -68436 56706 -68374
rect 57096 -68399 57125 -68365
rect 57159 -68399 57217 -68365
rect 57251 -68399 57309 -68365
rect 57343 -68399 57372 -68365
rect 56316 -68470 56412 -68436
rect 56610 -68470 56706 -68436
rect 57131 -68454 57165 -68433
rect 57201 -68441 57267 -68399
rect 57201 -68475 57217 -68441
rect 57251 -68475 57267 -68441
rect 57303 -68471 57355 -68433
rect 57131 -68509 57165 -68488
rect 57337 -68505 57355 -68471
rect 59276 -68002 59310 -67942
rect 59387 -67944 60054 -67909
rect 60127 -67754 60161 -67728
rect 60127 -67757 60253 -67754
rect 60161 -67773 60253 -67757
rect 60161 -67791 60203 -67773
rect 60127 -67807 60203 -67791
rect 60237 -67807 60253 -67773
rect 60359 -67760 60409 -67749
rect 60671 -67754 60705 -67728
rect 60359 -67765 60366 -67760
rect 60359 -67800 60366 -67799
rect 60406 -67800 60409 -67760
rect 60127 -67849 60161 -67807
rect 60127 -67941 60161 -67883
rect 60195 -67857 60325 -67841
rect 60195 -67891 60211 -67857
rect 60245 -67891 60325 -67857
rect 60195 -67907 60325 -67891
rect 59387 -68000 59421 -67944
rect 59087 -68042 59103 -68008
rect 59137 -68042 59153 -68008
rect 59044 -68101 59078 -68085
rect 57131 -68543 57264 -68509
rect 57303 -68534 57355 -68505
rect 57117 -68594 57185 -68579
rect 57117 -68644 57118 -68594
rect 57168 -68644 57185 -68594
rect 57117 -68653 57185 -68644
rect 57230 -68594 57264 -68543
rect 57319 -68570 57355 -68534
rect 57230 -68610 57285 -68594
rect 57230 -68644 57251 -68610
rect 57230 -68660 57285 -68644
rect 57319 -68610 57326 -68570
rect 59044 -68493 59078 -68477
rect 59162 -68101 59196 -68085
rect 59162 -68493 59196 -68477
rect 59087 -68570 59103 -68536
rect 59137 -68570 59153 -68536
rect 57230 -68689 57264 -68660
rect 57129 -68723 57264 -68689
rect 57319 -68694 57355 -68610
rect 57129 -68757 57165 -68723
rect 57301 -68744 57355 -68694
rect 58930 -68638 58964 -68576
rect 59529 -68045 59545 -68011
rect 59579 -68045 59595 -68011
rect 59501 -68095 59535 -68079
rect 59501 -68287 59535 -68271
rect 59589 -68095 59623 -68079
rect 59589 -68287 59623 -68271
rect 59529 -68355 59545 -68321
rect 59579 -68355 59595 -68321
rect 59387 -68423 59421 -68370
rect 59703 -68423 59737 -67944
rect 60019 -68005 60053 -67944
rect 59845 -68045 59861 -68011
rect 59895 -68045 59911 -68011
rect 59817 -68095 59851 -68079
rect 59817 -68287 59851 -68271
rect 59905 -68095 59939 -68079
rect 59905 -68287 59939 -68271
rect 59845 -68355 59861 -68321
rect 59895 -68355 59911 -68321
rect 60161 -67975 60203 -67941
rect 60237 -67975 60253 -67941
rect 60127 -68033 60161 -67975
rect 60289 -68009 60325 -67907
rect 60127 -68109 60161 -68067
rect 60195 -68025 60325 -68009
rect 60195 -68059 60211 -68025
rect 60245 -68059 60325 -68025
rect 60195 -68075 60325 -68059
rect 60359 -67850 60409 -67800
rect 60443 -67757 60705 -67754
rect 60443 -67773 60671 -67757
rect 60443 -67807 60459 -67773
rect 60493 -67807 60527 -67773
rect 60561 -67807 60595 -67773
rect 60629 -67791 60671 -67773
rect 60629 -67807 60705 -67791
rect 60359 -67857 60366 -67850
rect 60406 -67890 60409 -67850
rect 60393 -67891 60409 -67890
rect 60359 -67940 60409 -67891
rect 60359 -67941 60366 -67940
rect 60359 -67980 60366 -67975
rect 60406 -67980 60409 -67940
rect 60359 -68020 60409 -67980
rect 60359 -68025 60366 -68020
rect 60359 -68060 60366 -68059
rect 60406 -68060 60409 -68020
rect 60359 -68075 60409 -68060
rect 60443 -67857 60637 -67841
rect 60443 -67891 60459 -67857
rect 60493 -67891 60527 -67857
rect 60561 -67891 60595 -67857
rect 60629 -67891 60637 -67857
rect 60443 -67907 60637 -67891
rect 60671 -67849 60705 -67807
rect 60443 -68009 60477 -67907
rect 60671 -67941 60705 -67883
rect 60511 -67975 60527 -67941
rect 60561 -67975 60595 -67941
rect 60629 -67975 60671 -67941
rect 60443 -68025 60637 -68009
rect 60443 -68059 60459 -68025
rect 60493 -68059 60527 -68025
rect 60561 -68059 60595 -68025
rect 60629 -68059 60637 -68025
rect 60443 -68075 60637 -68059
rect 60671 -68033 60705 -67975
rect 60289 -68109 60325 -68075
rect 60443 -68109 60481 -68075
rect 60671 -68109 60705 -68067
rect 60127 -68125 60204 -68109
rect 60161 -68143 60204 -68125
rect 60238 -68143 60254 -68109
rect 60161 -68159 60254 -68143
rect 60289 -68125 60481 -68109
rect 60289 -68159 60297 -68125
rect 60331 -68159 60369 -68125
rect 60405 -68159 60449 -68125
rect 60579 -68143 60595 -68109
rect 60629 -68125 60705 -68109
rect 60629 -68143 60671 -68125
rect 60579 -68151 60671 -68143
rect 60127 -68188 60161 -68159
rect 60289 -68162 60481 -68159
rect 60671 -68188 60705 -68159
rect 60747 -67754 60781 -67728
rect 60747 -67757 61009 -67754
rect 60781 -67773 61009 -67757
rect 60781 -67791 60823 -67773
rect 60747 -67807 60823 -67791
rect 60857 -67807 60891 -67773
rect 60925 -67807 60959 -67773
rect 60993 -67807 61009 -67773
rect 61043 -67760 61093 -67749
rect 61291 -67754 61325 -67728
rect 61043 -67800 61046 -67760
rect 61086 -67765 61093 -67760
rect 61086 -67800 61093 -67799
rect 60747 -67849 60781 -67807
rect 60747 -67941 60781 -67883
rect 60815 -67857 61009 -67841
rect 60815 -67891 60823 -67857
rect 60857 -67891 60891 -67857
rect 60925 -67891 60959 -67857
rect 60993 -67891 61009 -67857
rect 60815 -67907 61009 -67891
rect 60781 -67975 60823 -67941
rect 60857 -67975 60891 -67941
rect 60925 -67975 60941 -67941
rect 60747 -68033 60781 -67975
rect 60975 -68009 61009 -67907
rect 60747 -68109 60781 -68067
rect 60815 -68025 61009 -68009
rect 60815 -68059 60823 -68025
rect 60857 -68059 60891 -68025
rect 60925 -68059 60959 -68025
rect 60993 -68059 61009 -68025
rect 60815 -68075 61009 -68059
rect 61043 -67850 61093 -67800
rect 61199 -67757 61325 -67754
rect 61199 -67773 61291 -67757
rect 61199 -67807 61215 -67773
rect 61249 -67791 61291 -67773
rect 61249 -67807 61325 -67791
rect 61043 -67890 61046 -67850
rect 61086 -67857 61093 -67850
rect 61043 -67891 61059 -67890
rect 61043 -67940 61093 -67891
rect 61043 -67980 61046 -67940
rect 61086 -67941 61093 -67940
rect 61086 -67980 61093 -67975
rect 61043 -68020 61093 -67980
rect 61043 -68060 61046 -68020
rect 61086 -68025 61093 -68020
rect 61086 -68060 61093 -68059
rect 61043 -68075 61093 -68060
rect 61127 -67857 61257 -67841
rect 61127 -67891 61207 -67857
rect 61241 -67891 61257 -67857
rect 61127 -67907 61257 -67891
rect 61291 -67849 61325 -67807
rect 61127 -68009 61163 -67907
rect 61291 -67941 61325 -67883
rect 61199 -67975 61215 -67941
rect 61249 -67975 61291 -67941
rect 61127 -68025 61257 -68009
rect 61127 -68059 61207 -68025
rect 61241 -68059 61257 -68025
rect 61127 -68075 61257 -68059
rect 61291 -68033 61325 -67975
rect 60971 -68109 61009 -68075
rect 61127 -68109 61163 -68075
rect 61291 -68109 61325 -68067
rect 60747 -68125 60823 -68109
rect 60781 -68143 60823 -68125
rect 60857 -68143 60873 -68109
rect 60781 -68151 60873 -68143
rect 60971 -68124 61163 -68109
rect 60971 -68125 61129 -68124
rect 60747 -68188 60781 -68159
rect 60971 -68159 60980 -68125
rect 61015 -68159 61053 -68125
rect 61088 -68158 61129 -68125
rect 61198 -68143 61214 -68109
rect 61248 -68125 61325 -68109
rect 61248 -68143 61291 -68125
rect 61088 -68159 61163 -68158
rect 61198 -68159 61291 -68143
rect 60971 -68162 61163 -68159
rect 61291 -68188 61325 -68159
rect 60466 -68260 60546 -68240
rect 60466 -68300 60486 -68260
rect 60526 -68300 60546 -68260
rect 60466 -68320 60546 -68300
rect 60606 -68260 60686 -68240
rect 60606 -68300 60626 -68260
rect 60666 -68300 60686 -68260
rect 60606 -68320 60686 -68300
rect 60746 -68260 60826 -68240
rect 60746 -68300 60766 -68260
rect 60806 -68300 60826 -68260
rect 60746 -68320 60826 -68300
rect 60886 -68260 60966 -68240
rect 60886 -68300 60906 -68260
rect 60946 -68300 60966 -68260
rect 60886 -68320 60966 -68300
rect 60019 -68423 60053 -68361
rect 59387 -68457 59476 -68423
rect 59646 -68457 59799 -68423
rect 59957 -68426 60053 -68423
rect 59957 -68457 60520 -68426
rect 59772 -68460 60520 -68457
rect 59772 -68520 59806 -68460
rect 59276 -68638 59310 -68576
rect 58930 -68672 59026 -68638
rect 59214 -68640 59310 -68638
rect 59214 -68672 59696 -68640
rect 58930 -68674 59696 -68672
rect 58930 -68710 58964 -68674
rect 57129 -68791 57131 -68757
rect 57129 -68825 57165 -68791
rect 57129 -68859 57131 -68825
rect 57129 -68875 57165 -68859
rect 57201 -68791 57217 -68757
rect 57251 -68791 57267 -68757
rect 57201 -68825 57267 -68791
rect 57201 -68859 57217 -68825
rect 57251 -68859 57267 -68825
rect 57201 -68909 57267 -68859
rect 57301 -68778 57303 -68744
rect 57337 -68778 57355 -68744
rect 57301 -68825 57355 -68778
rect 57301 -68859 57303 -68825
rect 57337 -68859 57355 -68825
rect 57301 -68875 57355 -68859
rect 59662 -68730 59696 -68674
rect 60486 -68522 60520 -68460
rect 59942 -68574 59958 -68540
rect 60334 -68574 60350 -68540
rect 59874 -68594 59908 -68578
rect 59874 -68644 59908 -68628
rect 60384 -68594 60418 -68578
rect 60384 -68644 60418 -68628
rect 59942 -68682 59958 -68648
rect 60334 -68682 60350 -68648
rect 56112 -68982 56146 -68920
rect 57096 -68943 57125 -68909
rect 57159 -68943 57217 -68909
rect 57251 -68943 57309 -68909
rect 57343 -68943 57372 -68909
rect 55706 -69016 55802 -68982
rect 56050 -69016 56146 -68982
rect 53886 -69064 53982 -69030
rect 54956 -69064 55052 -69030
rect 53886 -69126 53920 -69064
rect 55018 -69126 55052 -69064
rect 55720 -69058 56090 -69016
rect 55720 -69068 56020 -69058
rect 54065 -69178 54081 -69144
rect 54857 -69178 54873 -69144
rect 53988 -69206 54022 -69190
rect 53988 -69260 54022 -69244
rect 54916 -69206 54950 -69190
rect 54916 -69260 54950 -69244
rect 54065 -69306 54081 -69272
rect 54857 -69306 54873 -69272
rect 53886 -69386 53920 -69324
rect 56010 -69208 56020 -69068
rect 56080 -69208 56090 -69058
rect 59109 -68788 59125 -68754
rect 59501 -68788 59517 -68754
rect 59560 -68808 59594 -68792
rect 59560 -68858 59594 -68842
rect 59109 -68896 59125 -68862
rect 59501 -68896 59517 -68862
rect 59032 -68916 59066 -68900
rect 59032 -68966 59066 -68950
rect 59109 -69004 59125 -68970
rect 59501 -69004 59517 -68970
rect 56010 -69218 56090 -69208
rect 59772 -68762 59806 -68700
rect 60486 -68762 60520 -68700
rect 59772 -68796 59866 -68762
rect 60426 -68796 60520 -68762
rect 59662 -69084 59696 -69030
rect 58966 -69100 59026 -69084
rect 58930 -69118 59026 -69100
rect 59600 -69118 59696 -69084
rect 55018 -69386 55052 -69324
rect 53886 -69420 53982 -69386
rect 54956 -69420 55052 -69386
rect 55176 -69278 55272 -69244
rect 55566 -69278 55662 -69244
rect 55176 -69340 55210 -69278
rect 55628 -69340 55662 -69278
rect 55284 -69392 55300 -69358
rect 55476 -69392 55492 -69358
rect 55526 -69402 55560 -69386
rect 55284 -69480 55300 -69446
rect 55476 -69480 55492 -69446
rect 55526 -69452 55560 -69436
rect 55176 -69560 55210 -69498
rect 55628 -69560 55662 -69498
rect 55176 -69594 55272 -69560
rect 55566 -69594 55662 -69560
rect 53896 -71792 53992 -71758
rect 54966 -71792 55062 -71758
rect 53896 -71854 53930 -71792
rect 55028 -71854 55062 -71792
rect 54075 -71906 54091 -71872
rect 54867 -71906 54883 -71872
rect 53998 -71934 54032 -71918
rect 53998 -71988 54032 -71972
rect 54926 -71934 54960 -71918
rect 54926 -71988 54960 -71972
rect 54075 -72034 54091 -72000
rect 54867 -72034 54883 -72000
rect 53896 -72114 53930 -72052
rect 55028 -72114 55062 -72052
rect 55960 -72108 56040 -72098
rect 53896 -72148 53992 -72114
rect 54966 -72148 55062 -72114
rect 53350 -72238 53790 -72204
rect 53350 -72300 53384 -72238
rect 53510 -72340 53526 -72306
rect 53614 -72340 53630 -72306
rect 53464 -72390 53498 -72374
rect 53464 -73182 53498 -73166
rect 53642 -72390 53676 -72374
rect 53642 -73182 53676 -73166
rect 53756 -72864 53790 -72238
rect 53896 -72210 53930 -72148
rect 55028 -72210 55062 -72148
rect 55710 -72154 56040 -72108
rect 54075 -72262 54091 -72228
rect 54867 -72262 54883 -72228
rect 53998 -72290 54032 -72274
rect 53998 -72344 54032 -72328
rect 54926 -72290 54960 -72274
rect 54926 -72344 54960 -72328
rect 54075 -72390 54091 -72356
rect 54867 -72390 54883 -72356
rect 53896 -72470 53930 -72408
rect 55706 -72188 55802 -72154
rect 56050 -72188 56146 -72154
rect 55706 -72250 55740 -72188
rect 55028 -72470 55062 -72408
rect 53896 -72504 53992 -72470
rect 54966 -72504 55062 -72470
rect 55176 -72300 55272 -72266
rect 55430 -72300 55526 -72266
rect 55176 -72362 55210 -72300
rect 55492 -72362 55526 -72300
rect 55318 -72402 55334 -72368
rect 55368 -72402 55384 -72368
rect 55290 -72452 55324 -72436
rect 55290 -72644 55324 -72628
rect 55378 -72452 55412 -72436
rect 55378 -72644 55412 -72628
rect 55176 -72718 55210 -72656
rect 55492 -72718 55526 -72656
rect 54870 -72752 55272 -72718
rect 55430 -72752 55706 -72718
rect 54870 -72758 55706 -72752
rect 54870 -72864 54904 -72758
rect 53756 -72898 53852 -72864
rect 54808 -72898 54904 -72864
rect 53756 -72960 53790 -72898
rect 54870 -72960 54904 -72898
rect 55126 -72908 55142 -72874
rect 55494 -72908 55510 -72874
rect 53926 -73012 53942 -72978
rect 54718 -73012 54734 -72978
rect 53858 -73040 53892 -73024
rect 53858 -73144 53892 -73128
rect 54768 -73040 54802 -73024
rect 54768 -73144 54802 -73128
rect 53926 -73190 53942 -73156
rect 54718 -73190 54734 -73156
rect 53510 -73250 53526 -73216
rect 53614 -73250 53630 -73216
rect 53756 -73270 53790 -73208
rect 55046 -72960 55080 -72944
rect 55046 -73010 55080 -72994
rect 55556 -72960 55590 -72944
rect 55556 -73010 55590 -72994
rect 55126 -73080 55142 -73046
rect 55494 -73080 55510 -73046
rect 54870 -73238 54904 -73208
rect 55700 -73206 55706 -72758
rect 56112 -72250 56146 -72188
rect 58930 -72167 59026 -72133
rect 59600 -72167 59696 -72133
rect 58930 -72210 58964 -72167
rect 58926 -72220 58966 -72210
rect 55866 -72290 55882 -72256
rect 55970 -72290 55986 -72256
rect 55820 -72340 55854 -72324
rect 55820 -73132 55854 -73116
rect 55998 -72340 56032 -72324
rect 55998 -73132 56032 -73116
rect 55866 -73200 55882 -73166
rect 55970 -73200 55986 -73166
rect 55700 -73238 55740 -73206
rect 57096 -72279 57125 -72245
rect 57159 -72279 57217 -72245
rect 57251 -72279 57309 -72245
rect 57343 -72279 57372 -72245
rect 57129 -72329 57165 -72313
rect 57129 -72363 57131 -72329
rect 57129 -72397 57165 -72363
rect 57129 -72431 57131 -72397
rect 57201 -72329 57267 -72279
rect 57201 -72363 57217 -72329
rect 57251 -72363 57267 -72329
rect 57201 -72397 57267 -72363
rect 57201 -72431 57217 -72397
rect 57251 -72431 57267 -72397
rect 57301 -72329 57355 -72313
rect 57301 -72363 57303 -72329
rect 57337 -72363 57355 -72329
rect 57301 -72410 57355 -72363
rect 57129 -72465 57165 -72431
rect 57301 -72444 57303 -72410
rect 57337 -72444 57355 -72410
rect 57129 -72499 57264 -72465
rect 57301 -72494 57355 -72444
rect 57230 -72528 57264 -72499
rect 57117 -72544 57185 -72535
rect 57117 -72594 57118 -72544
rect 57178 -72594 57185 -72544
rect 57117 -72609 57185 -72594
rect 57230 -72544 57285 -72528
rect 57230 -72578 57251 -72544
rect 57230 -72594 57285 -72578
rect 57319 -72540 57355 -72494
rect 59662 -72229 59696 -72167
rect 59109 -72281 59125 -72247
rect 59501 -72281 59517 -72247
rect 59560 -72301 59594 -72285
rect 59560 -72351 59594 -72335
rect 59109 -72389 59125 -72355
rect 59501 -72389 59517 -72355
rect 59032 -72409 59066 -72393
rect 59032 -72459 59066 -72443
rect 59109 -72497 59125 -72463
rect 59501 -72497 59517 -72463
rect 58926 -72540 58966 -72520
rect 57319 -72580 57326 -72540
rect 58930 -72576 58964 -72540
rect 57230 -72645 57264 -72594
rect 57131 -72679 57264 -72645
rect 57319 -72654 57355 -72580
rect 57131 -72700 57165 -72679
rect 56316 -72718 56412 -72704
rect 54830 -73248 55830 -73238
rect 54830 -73270 55030 -73248
rect 53756 -73304 53852 -73270
rect 54808 -73304 55030 -73270
rect 53510 -73358 53526 -73324
rect 53614 -73358 53630 -73324
rect 53756 -73366 53790 -73304
rect 54830 -73328 55030 -73304
rect 55110 -73268 55740 -73248
rect 55810 -73268 55830 -73248
rect 56112 -73268 56146 -73206
rect 55110 -73308 55160 -73268
rect 55600 -73308 55740 -73268
rect 56050 -73302 56146 -73268
rect 55110 -73328 55740 -73308
rect 55810 -73328 55830 -73302
rect 54830 -73338 55830 -73328
rect 53464 -73408 53498 -73392
rect 53464 -74200 53498 -74184
rect 53642 -73408 53676 -73392
rect 53642 -74200 53676 -74184
rect 54870 -73366 54904 -73338
rect 53926 -73418 53942 -73384
rect 54718 -73418 54734 -73384
rect 53858 -73446 53892 -73430
rect 53858 -73550 53892 -73534
rect 54768 -73446 54802 -73430
rect 54768 -73550 54802 -73534
rect 53926 -73596 53942 -73562
rect 54718 -73596 54734 -73562
rect 53756 -73676 53790 -73614
rect 55700 -73364 55740 -73338
rect 55126 -73530 55142 -73496
rect 55494 -73530 55510 -73496
rect 54870 -73676 54904 -73614
rect 55046 -73582 55080 -73566
rect 55046 -73632 55080 -73616
rect 55556 -73582 55590 -73566
rect 55556 -73632 55590 -73616
rect 53756 -73710 53852 -73676
rect 54808 -73710 54904 -73676
rect 55126 -73702 55142 -73668
rect 55494 -73702 55510 -73668
rect 53510 -74268 53526 -74234
rect 53614 -74268 53630 -74234
rect 53350 -74336 53384 -74274
rect 53756 -74336 53790 -73710
rect 54870 -73818 54904 -73710
rect 55700 -73818 55706 -73364
rect 54870 -73824 55706 -73818
rect 54870 -73858 55262 -73824
rect 55420 -73858 55706 -73824
rect 55166 -73920 55200 -73858
rect 53350 -74370 53446 -74336
rect 53694 -74370 53790 -74336
rect 53886 -74108 53982 -74074
rect 54956 -74108 55052 -74074
rect 53886 -74170 53920 -74108
rect 55018 -74170 55052 -74108
rect 54065 -74222 54081 -74188
rect 54857 -74222 54873 -74188
rect 53988 -74250 54022 -74234
rect 53988 -74304 54022 -74288
rect 54916 -74250 54950 -74234
rect 54916 -74304 54950 -74288
rect 54065 -74350 54081 -74316
rect 54857 -74350 54873 -74316
rect 53886 -74430 53920 -74368
rect 55482 -73920 55516 -73858
rect 55280 -73948 55314 -73932
rect 55280 -74140 55314 -74124
rect 55368 -73948 55402 -73932
rect 55368 -74140 55402 -74124
rect 55308 -74208 55324 -74174
rect 55358 -74208 55374 -74174
rect 55166 -74276 55200 -74214
rect 55482 -74276 55516 -74214
rect 55166 -74310 55262 -74276
rect 55420 -74310 55516 -74276
rect 55018 -74430 55052 -74368
rect 56112 -73364 56146 -73302
rect 56350 -72738 56412 -72718
rect 56610 -72738 56706 -72704
rect 56672 -72800 56706 -72738
rect 57303 -72683 57355 -72654
rect 57131 -72755 57165 -72734
rect 57201 -72747 57217 -72713
rect 57251 -72747 57267 -72713
rect 57201 -72789 57267 -72747
rect 57337 -72717 57355 -72683
rect 57303 -72755 57355 -72717
rect 58930 -72610 59026 -72576
rect 59214 -72577 59310 -72576
rect 59662 -72577 59696 -72520
rect 59772 -72494 59866 -72460
rect 60426 -72494 60520 -72460
rect 59772 -72550 59806 -72494
rect 59214 -72610 59696 -72577
rect 58930 -72611 59696 -72610
rect 58930 -72672 58964 -72611
rect 59276 -72672 59310 -72611
rect 59087 -72712 59103 -72678
rect 59137 -72712 59153 -72678
rect 56476 -72840 56492 -72806
rect 56530 -72840 56546 -72806
rect 55866 -73404 55882 -73370
rect 55970 -73404 55986 -73370
rect 55820 -73454 55854 -73438
rect 55820 -74246 55854 -74230
rect 55998 -73454 56032 -73438
rect 55998 -74246 56032 -74230
rect 55866 -74314 55882 -74280
rect 55970 -74314 55986 -74280
rect 55706 -74382 55740 -74320
rect 56430 -72899 56464 -72883
rect 56430 -73691 56464 -73675
rect 56558 -72899 56592 -72883
rect 56558 -73691 56592 -73675
rect 56476 -73768 56492 -73734
rect 56530 -73768 56546 -73734
rect 56316 -73836 56350 -73774
rect 57096 -72823 57125 -72789
rect 57159 -72823 57217 -72789
rect 57251 -72823 57309 -72789
rect 57343 -72823 57372 -72789
rect 59044 -72771 59078 -72755
rect 59044 -73163 59078 -73147
rect 59162 -72771 59196 -72755
rect 59162 -73163 59196 -73147
rect 59087 -73240 59103 -73206
rect 59137 -73240 59153 -73206
rect 60486 -72556 60520 -72494
rect 59942 -72608 59958 -72574
rect 60334 -72608 60350 -72574
rect 59874 -72628 59908 -72612
rect 59874 -72678 59908 -72662
rect 60384 -72628 60418 -72612
rect 60384 -72678 60418 -72662
rect 59942 -72716 59958 -72682
rect 60334 -72716 60350 -72682
rect 59772 -72796 59806 -72740
rect 60486 -72796 60520 -72734
rect 59388 -72830 59476 -72796
rect 59656 -72830 59800 -72796
rect 59958 -72830 60520 -72796
rect 59388 -72890 59422 -72830
rect 59276 -73306 59310 -73246
rect 59530 -72932 59546 -72898
rect 59580 -72932 59596 -72898
rect 59502 -72982 59536 -72966
rect 59502 -73174 59536 -73158
rect 59590 -72982 59624 -72966
rect 59590 -73174 59624 -73158
rect 59530 -73242 59546 -73208
rect 59580 -73242 59596 -73208
rect 58966 -73342 59310 -73306
rect 59388 -73309 59422 -73250
rect 59704 -73309 59738 -72830
rect 60020 -72892 60054 -72830
rect 59846 -72932 59862 -72898
rect 59896 -72932 59912 -72898
rect 59818 -72982 59852 -72966
rect 59818 -73174 59852 -73158
rect 59906 -72982 59940 -72966
rect 59906 -73174 59940 -73158
rect 59846 -73242 59862 -73208
rect 59896 -73242 59912 -73208
rect 61186 -73000 61286 -72990
rect 61186 -73080 61196 -73000
rect 61186 -73090 61286 -73080
rect 60020 -73309 60054 -73248
rect 56672 -73836 56706 -73774
rect 57096 -73799 57125 -73765
rect 57159 -73799 57217 -73765
rect 57251 -73799 57309 -73765
rect 57343 -73799 57372 -73765
rect 56316 -73870 56412 -73836
rect 56610 -73870 56706 -73836
rect 57131 -73854 57165 -73833
rect 57201 -73841 57267 -73799
rect 57201 -73875 57217 -73841
rect 57251 -73875 57267 -73841
rect 57303 -73871 57355 -73833
rect 57131 -73909 57165 -73888
rect 57337 -73905 57355 -73871
rect 59276 -73402 59310 -73342
rect 59387 -73344 60054 -73309
rect 60127 -73154 60161 -73128
rect 60127 -73157 60253 -73154
rect 60161 -73173 60253 -73157
rect 60161 -73191 60203 -73173
rect 60127 -73207 60203 -73191
rect 60237 -73207 60253 -73173
rect 60359 -73160 60409 -73149
rect 60671 -73154 60705 -73128
rect 60359 -73165 60366 -73160
rect 60359 -73200 60366 -73199
rect 60406 -73200 60409 -73160
rect 60127 -73249 60161 -73207
rect 60127 -73341 60161 -73283
rect 60195 -73257 60325 -73241
rect 60195 -73291 60211 -73257
rect 60245 -73291 60325 -73257
rect 60195 -73307 60325 -73291
rect 59387 -73400 59421 -73344
rect 59087 -73442 59103 -73408
rect 59137 -73442 59153 -73408
rect 59044 -73501 59078 -73485
rect 57131 -73943 57264 -73909
rect 57303 -73934 57355 -73905
rect 57117 -73994 57185 -73979
rect 57117 -74044 57118 -73994
rect 57168 -74044 57185 -73994
rect 57117 -74053 57185 -74044
rect 57230 -73994 57264 -73943
rect 57319 -73970 57355 -73934
rect 57230 -74010 57285 -73994
rect 57230 -74044 57251 -74010
rect 57230 -74060 57285 -74044
rect 57319 -74010 57326 -73970
rect 59044 -73893 59078 -73877
rect 59162 -73501 59196 -73485
rect 59162 -73893 59196 -73877
rect 59087 -73970 59103 -73936
rect 59137 -73970 59153 -73936
rect 57230 -74089 57264 -74060
rect 57129 -74123 57264 -74089
rect 57319 -74094 57355 -74010
rect 57129 -74157 57165 -74123
rect 57301 -74144 57355 -74094
rect 58930 -74038 58964 -73976
rect 59529 -73445 59545 -73411
rect 59579 -73445 59595 -73411
rect 59501 -73495 59535 -73479
rect 59501 -73687 59535 -73671
rect 59589 -73495 59623 -73479
rect 59589 -73687 59623 -73671
rect 59529 -73755 59545 -73721
rect 59579 -73755 59595 -73721
rect 59387 -73823 59421 -73770
rect 59703 -73823 59737 -73344
rect 60019 -73405 60053 -73344
rect 59845 -73445 59861 -73411
rect 59895 -73445 59911 -73411
rect 59817 -73495 59851 -73479
rect 59817 -73687 59851 -73671
rect 59905 -73495 59939 -73479
rect 59905 -73687 59939 -73671
rect 59845 -73755 59861 -73721
rect 59895 -73755 59911 -73721
rect 60161 -73375 60203 -73341
rect 60237 -73375 60253 -73341
rect 60127 -73433 60161 -73375
rect 60289 -73409 60325 -73307
rect 60127 -73509 60161 -73467
rect 60195 -73425 60325 -73409
rect 60195 -73459 60211 -73425
rect 60245 -73459 60325 -73425
rect 60195 -73475 60325 -73459
rect 60359 -73250 60409 -73200
rect 60443 -73157 60705 -73154
rect 60443 -73173 60671 -73157
rect 60443 -73207 60459 -73173
rect 60493 -73207 60527 -73173
rect 60561 -73207 60595 -73173
rect 60629 -73191 60671 -73173
rect 60629 -73207 60705 -73191
rect 60359 -73257 60366 -73250
rect 60406 -73290 60409 -73250
rect 60393 -73291 60409 -73290
rect 60359 -73340 60409 -73291
rect 60359 -73341 60366 -73340
rect 60359 -73380 60366 -73375
rect 60406 -73380 60409 -73340
rect 60359 -73420 60409 -73380
rect 60359 -73425 60366 -73420
rect 60359 -73460 60366 -73459
rect 60406 -73460 60409 -73420
rect 60359 -73475 60409 -73460
rect 60443 -73257 60637 -73241
rect 60443 -73291 60459 -73257
rect 60493 -73291 60527 -73257
rect 60561 -73291 60595 -73257
rect 60629 -73291 60637 -73257
rect 60443 -73307 60637 -73291
rect 60671 -73249 60705 -73207
rect 60443 -73409 60477 -73307
rect 60671 -73341 60705 -73283
rect 60511 -73375 60527 -73341
rect 60561 -73375 60595 -73341
rect 60629 -73375 60671 -73341
rect 60443 -73425 60637 -73409
rect 60443 -73459 60459 -73425
rect 60493 -73459 60527 -73425
rect 60561 -73459 60595 -73425
rect 60629 -73459 60637 -73425
rect 60443 -73475 60637 -73459
rect 60671 -73433 60705 -73375
rect 60289 -73509 60325 -73475
rect 60443 -73509 60481 -73475
rect 60671 -73509 60705 -73467
rect 60127 -73525 60204 -73509
rect 60161 -73543 60204 -73525
rect 60238 -73543 60254 -73509
rect 60161 -73559 60254 -73543
rect 60289 -73525 60481 -73509
rect 60289 -73559 60297 -73525
rect 60331 -73559 60369 -73525
rect 60405 -73559 60449 -73525
rect 60579 -73543 60595 -73509
rect 60629 -73525 60705 -73509
rect 60629 -73543 60671 -73525
rect 60579 -73551 60671 -73543
rect 60127 -73588 60161 -73559
rect 60289 -73562 60481 -73559
rect 60671 -73588 60705 -73559
rect 60747 -73154 60781 -73128
rect 60747 -73157 61009 -73154
rect 60781 -73173 61009 -73157
rect 60781 -73191 60823 -73173
rect 60747 -73207 60823 -73191
rect 60857 -73207 60891 -73173
rect 60925 -73207 60959 -73173
rect 60993 -73207 61009 -73173
rect 61043 -73160 61093 -73149
rect 61291 -73154 61325 -73128
rect 61043 -73200 61046 -73160
rect 61086 -73165 61093 -73160
rect 61086 -73200 61093 -73199
rect 60747 -73249 60781 -73207
rect 60747 -73341 60781 -73283
rect 60815 -73257 61009 -73241
rect 60815 -73291 60823 -73257
rect 60857 -73291 60891 -73257
rect 60925 -73291 60959 -73257
rect 60993 -73291 61009 -73257
rect 60815 -73307 61009 -73291
rect 60781 -73375 60823 -73341
rect 60857 -73375 60891 -73341
rect 60925 -73375 60941 -73341
rect 60747 -73433 60781 -73375
rect 60975 -73409 61009 -73307
rect 60747 -73509 60781 -73467
rect 60815 -73425 61009 -73409
rect 60815 -73459 60823 -73425
rect 60857 -73459 60891 -73425
rect 60925 -73459 60959 -73425
rect 60993 -73459 61009 -73425
rect 60815 -73475 61009 -73459
rect 61043 -73250 61093 -73200
rect 61199 -73157 61325 -73154
rect 61199 -73173 61291 -73157
rect 61199 -73207 61215 -73173
rect 61249 -73191 61291 -73173
rect 61249 -73207 61325 -73191
rect 61043 -73290 61046 -73250
rect 61086 -73257 61093 -73250
rect 61043 -73291 61059 -73290
rect 61043 -73340 61093 -73291
rect 61043 -73380 61046 -73340
rect 61086 -73341 61093 -73340
rect 61086 -73380 61093 -73375
rect 61043 -73420 61093 -73380
rect 61043 -73460 61046 -73420
rect 61086 -73425 61093 -73420
rect 61086 -73460 61093 -73459
rect 61043 -73475 61093 -73460
rect 61127 -73257 61257 -73241
rect 61127 -73291 61207 -73257
rect 61241 -73291 61257 -73257
rect 61127 -73307 61257 -73291
rect 61291 -73249 61325 -73207
rect 61127 -73409 61163 -73307
rect 61291 -73341 61325 -73283
rect 61199 -73375 61215 -73341
rect 61249 -73375 61291 -73341
rect 61127 -73425 61257 -73409
rect 61127 -73459 61207 -73425
rect 61241 -73459 61257 -73425
rect 61127 -73475 61257 -73459
rect 61291 -73433 61325 -73375
rect 60971 -73509 61009 -73475
rect 61127 -73509 61163 -73475
rect 61291 -73509 61325 -73467
rect 60747 -73525 60823 -73509
rect 60781 -73543 60823 -73525
rect 60857 -73543 60873 -73509
rect 60781 -73551 60873 -73543
rect 60971 -73524 61163 -73509
rect 60971 -73525 61129 -73524
rect 60747 -73588 60781 -73559
rect 60971 -73559 60980 -73525
rect 61015 -73559 61053 -73525
rect 61088 -73558 61129 -73525
rect 61198 -73543 61214 -73509
rect 61248 -73525 61325 -73509
rect 61248 -73543 61291 -73525
rect 61088 -73559 61163 -73558
rect 61198 -73559 61291 -73543
rect 60971 -73562 61163 -73559
rect 61291 -73588 61325 -73559
rect 60466 -73660 60546 -73640
rect 60466 -73700 60486 -73660
rect 60526 -73700 60546 -73660
rect 60466 -73720 60546 -73700
rect 60606 -73660 60686 -73640
rect 60606 -73700 60626 -73660
rect 60666 -73700 60686 -73660
rect 60606 -73720 60686 -73700
rect 60746 -73660 60826 -73640
rect 60746 -73700 60766 -73660
rect 60806 -73700 60826 -73660
rect 60746 -73720 60826 -73700
rect 60886 -73660 60966 -73640
rect 60886 -73700 60906 -73660
rect 60946 -73700 60966 -73660
rect 60886 -73720 60966 -73700
rect 60019 -73823 60053 -73761
rect 59387 -73857 59476 -73823
rect 59646 -73857 59799 -73823
rect 59957 -73826 60053 -73823
rect 59957 -73857 60520 -73826
rect 59772 -73860 60520 -73857
rect 59772 -73920 59806 -73860
rect 59276 -74038 59310 -73976
rect 58930 -74072 59026 -74038
rect 59214 -74040 59310 -74038
rect 59214 -74072 59696 -74040
rect 58930 -74074 59696 -74072
rect 58930 -74110 58964 -74074
rect 57129 -74191 57131 -74157
rect 57129 -74225 57165 -74191
rect 57129 -74259 57131 -74225
rect 57129 -74275 57165 -74259
rect 57201 -74191 57217 -74157
rect 57251 -74191 57267 -74157
rect 57201 -74225 57267 -74191
rect 57201 -74259 57217 -74225
rect 57251 -74259 57267 -74225
rect 57201 -74309 57267 -74259
rect 57301 -74178 57303 -74144
rect 57337 -74178 57355 -74144
rect 57301 -74225 57355 -74178
rect 57301 -74259 57303 -74225
rect 57337 -74259 57355 -74225
rect 57301 -74275 57355 -74259
rect 59662 -74130 59696 -74074
rect 60486 -73922 60520 -73860
rect 59942 -73974 59958 -73940
rect 60334 -73974 60350 -73940
rect 59874 -73994 59908 -73978
rect 59874 -74044 59908 -74028
rect 60384 -73994 60418 -73978
rect 60384 -74044 60418 -74028
rect 59942 -74082 59958 -74048
rect 60334 -74082 60350 -74048
rect 56112 -74382 56146 -74320
rect 57096 -74343 57125 -74309
rect 57159 -74343 57217 -74309
rect 57251 -74343 57309 -74309
rect 57343 -74343 57372 -74309
rect 55706 -74416 55802 -74382
rect 56050 -74416 56146 -74382
rect 53886 -74464 53982 -74430
rect 54956 -74464 55052 -74430
rect 53886 -74526 53920 -74464
rect 55018 -74526 55052 -74464
rect 55720 -74458 56090 -74416
rect 55720 -74468 56020 -74458
rect 54065 -74578 54081 -74544
rect 54857 -74578 54873 -74544
rect 53988 -74606 54022 -74590
rect 53988 -74660 54022 -74644
rect 54916 -74606 54950 -74590
rect 54916 -74660 54950 -74644
rect 54065 -74706 54081 -74672
rect 54857 -74706 54873 -74672
rect 53886 -74786 53920 -74724
rect 56010 -74608 56020 -74468
rect 56080 -74608 56090 -74458
rect 59109 -74188 59125 -74154
rect 59501 -74188 59517 -74154
rect 59560 -74208 59594 -74192
rect 59560 -74258 59594 -74242
rect 59109 -74296 59125 -74262
rect 59501 -74296 59517 -74262
rect 59032 -74316 59066 -74300
rect 59032 -74366 59066 -74350
rect 59109 -74404 59125 -74370
rect 59501 -74404 59517 -74370
rect 56010 -74618 56090 -74608
rect 59772 -74162 59806 -74100
rect 60486 -74162 60520 -74100
rect 59772 -74196 59866 -74162
rect 60426 -74196 60520 -74162
rect 59662 -74484 59696 -74430
rect 58966 -74500 59026 -74484
rect 58930 -74518 59026 -74500
rect 59600 -74518 59696 -74484
rect 55018 -74786 55052 -74724
rect 53886 -74820 53982 -74786
rect 54956 -74820 55052 -74786
rect 55176 -74678 55272 -74644
rect 55566 -74678 55662 -74644
rect 55176 -74740 55210 -74678
rect 55628 -74740 55662 -74678
rect 55284 -74792 55300 -74758
rect 55476 -74792 55492 -74758
rect 55526 -74802 55560 -74786
rect 55284 -74880 55300 -74846
rect 55476 -74880 55492 -74846
rect 55526 -74852 55560 -74836
rect 55176 -74960 55210 -74898
rect 55628 -74960 55662 -74898
rect 55176 -74994 55272 -74960
rect 55566 -74994 55662 -74960
rect 53896 -77192 53992 -77158
rect 54966 -77192 55062 -77158
rect 53896 -77254 53930 -77192
rect 55028 -77254 55062 -77192
rect 54075 -77306 54091 -77272
rect 54867 -77306 54883 -77272
rect 53998 -77334 54032 -77318
rect 53998 -77388 54032 -77372
rect 54926 -77334 54960 -77318
rect 54926 -77388 54960 -77372
rect 54075 -77434 54091 -77400
rect 54867 -77434 54883 -77400
rect 53896 -77514 53930 -77452
rect 55028 -77514 55062 -77452
rect 55960 -77508 56040 -77498
rect 53896 -77548 53992 -77514
rect 54966 -77548 55062 -77514
rect 53350 -77638 53790 -77604
rect 53350 -77700 53384 -77638
rect 53510 -77740 53526 -77706
rect 53614 -77740 53630 -77706
rect 53464 -77790 53498 -77774
rect 53464 -78582 53498 -78566
rect 53642 -77790 53676 -77774
rect 53642 -78582 53676 -78566
rect 53756 -78264 53790 -77638
rect 53896 -77610 53930 -77548
rect 55028 -77610 55062 -77548
rect 55710 -77554 56040 -77508
rect 54075 -77662 54091 -77628
rect 54867 -77662 54883 -77628
rect 53998 -77690 54032 -77674
rect 53998 -77744 54032 -77728
rect 54926 -77690 54960 -77674
rect 54926 -77744 54960 -77728
rect 54075 -77790 54091 -77756
rect 54867 -77790 54883 -77756
rect 53896 -77870 53930 -77808
rect 55706 -77588 55802 -77554
rect 56050 -77588 56146 -77554
rect 55706 -77650 55740 -77588
rect 55028 -77870 55062 -77808
rect 53896 -77904 53992 -77870
rect 54966 -77904 55062 -77870
rect 55176 -77700 55272 -77666
rect 55430 -77700 55526 -77666
rect 55176 -77762 55210 -77700
rect 55492 -77762 55526 -77700
rect 55318 -77802 55334 -77768
rect 55368 -77802 55384 -77768
rect 55290 -77852 55324 -77836
rect 55290 -78044 55324 -78028
rect 55378 -77852 55412 -77836
rect 55378 -78044 55412 -78028
rect 55176 -78118 55210 -78056
rect 55492 -78118 55526 -78056
rect 54870 -78152 55272 -78118
rect 55430 -78152 55706 -78118
rect 54870 -78158 55706 -78152
rect 54870 -78264 54904 -78158
rect 53756 -78298 53852 -78264
rect 54808 -78298 54904 -78264
rect 53756 -78360 53790 -78298
rect 54870 -78360 54904 -78298
rect 55126 -78308 55142 -78274
rect 55494 -78308 55510 -78274
rect 53926 -78412 53942 -78378
rect 54718 -78412 54734 -78378
rect 53858 -78440 53892 -78424
rect 53858 -78544 53892 -78528
rect 54768 -78440 54802 -78424
rect 54768 -78544 54802 -78528
rect 53926 -78590 53942 -78556
rect 54718 -78590 54734 -78556
rect 53510 -78650 53526 -78616
rect 53614 -78650 53630 -78616
rect 53756 -78670 53790 -78608
rect 55046 -78360 55080 -78344
rect 55046 -78410 55080 -78394
rect 55556 -78360 55590 -78344
rect 55556 -78410 55590 -78394
rect 55126 -78480 55142 -78446
rect 55494 -78480 55510 -78446
rect 54870 -78638 54904 -78608
rect 55700 -78606 55706 -78158
rect 56112 -77650 56146 -77588
rect 58930 -77567 59026 -77533
rect 59600 -77567 59696 -77533
rect 58930 -77610 58964 -77567
rect 58926 -77620 58966 -77610
rect 55866 -77690 55882 -77656
rect 55970 -77690 55986 -77656
rect 55820 -77740 55854 -77724
rect 55820 -78532 55854 -78516
rect 55998 -77740 56032 -77724
rect 55998 -78532 56032 -78516
rect 55866 -78600 55882 -78566
rect 55970 -78600 55986 -78566
rect 55700 -78638 55740 -78606
rect 57096 -77679 57125 -77645
rect 57159 -77679 57217 -77645
rect 57251 -77679 57309 -77645
rect 57343 -77679 57372 -77645
rect 57129 -77729 57165 -77713
rect 57129 -77763 57131 -77729
rect 57129 -77797 57165 -77763
rect 57129 -77831 57131 -77797
rect 57201 -77729 57267 -77679
rect 57201 -77763 57217 -77729
rect 57251 -77763 57267 -77729
rect 57201 -77797 57267 -77763
rect 57201 -77831 57217 -77797
rect 57251 -77831 57267 -77797
rect 57301 -77729 57355 -77713
rect 57301 -77763 57303 -77729
rect 57337 -77763 57355 -77729
rect 57301 -77810 57355 -77763
rect 57129 -77865 57165 -77831
rect 57301 -77844 57303 -77810
rect 57337 -77844 57355 -77810
rect 57129 -77899 57264 -77865
rect 57301 -77894 57355 -77844
rect 57230 -77928 57264 -77899
rect 57117 -77944 57185 -77935
rect 57117 -77994 57118 -77944
rect 57178 -77994 57185 -77944
rect 57117 -78009 57185 -77994
rect 57230 -77944 57285 -77928
rect 57230 -77978 57251 -77944
rect 57230 -77994 57285 -77978
rect 57319 -77940 57355 -77894
rect 59662 -77629 59696 -77567
rect 59109 -77681 59125 -77647
rect 59501 -77681 59517 -77647
rect 59560 -77701 59594 -77685
rect 59560 -77751 59594 -77735
rect 59109 -77789 59125 -77755
rect 59501 -77789 59517 -77755
rect 59032 -77809 59066 -77793
rect 59032 -77859 59066 -77843
rect 59109 -77897 59125 -77863
rect 59501 -77897 59517 -77863
rect 58926 -77940 58966 -77920
rect 57319 -77980 57326 -77940
rect 58930 -77976 58964 -77940
rect 57230 -78045 57264 -77994
rect 57131 -78079 57264 -78045
rect 57319 -78054 57355 -77980
rect 57131 -78100 57165 -78079
rect 56316 -78118 56412 -78104
rect 54830 -78648 55830 -78638
rect 54830 -78670 55030 -78648
rect 53756 -78704 53852 -78670
rect 54808 -78704 55030 -78670
rect 53510 -78758 53526 -78724
rect 53614 -78758 53630 -78724
rect 53756 -78766 53790 -78704
rect 54830 -78728 55030 -78704
rect 55110 -78668 55740 -78648
rect 55810 -78668 55830 -78648
rect 56112 -78668 56146 -78606
rect 55110 -78708 55160 -78668
rect 55600 -78708 55740 -78668
rect 56050 -78702 56146 -78668
rect 55110 -78728 55740 -78708
rect 55810 -78728 55830 -78702
rect 54830 -78738 55830 -78728
rect 53464 -78808 53498 -78792
rect 53464 -79600 53498 -79584
rect 53642 -78808 53676 -78792
rect 53642 -79600 53676 -79584
rect 54870 -78766 54904 -78738
rect 53926 -78818 53942 -78784
rect 54718 -78818 54734 -78784
rect 53858 -78846 53892 -78830
rect 53858 -78950 53892 -78934
rect 54768 -78846 54802 -78830
rect 54768 -78950 54802 -78934
rect 53926 -78996 53942 -78962
rect 54718 -78996 54734 -78962
rect 53756 -79076 53790 -79014
rect 55700 -78764 55740 -78738
rect 55126 -78930 55142 -78896
rect 55494 -78930 55510 -78896
rect 54870 -79076 54904 -79014
rect 55046 -78982 55080 -78966
rect 55046 -79032 55080 -79016
rect 55556 -78982 55590 -78966
rect 55556 -79032 55590 -79016
rect 53756 -79110 53852 -79076
rect 54808 -79110 54904 -79076
rect 55126 -79102 55142 -79068
rect 55494 -79102 55510 -79068
rect 53510 -79668 53526 -79634
rect 53614 -79668 53630 -79634
rect 53350 -79736 53384 -79674
rect 53756 -79736 53790 -79110
rect 54870 -79218 54904 -79110
rect 55700 -79218 55706 -78764
rect 54870 -79224 55706 -79218
rect 54870 -79258 55262 -79224
rect 55420 -79258 55706 -79224
rect 55166 -79320 55200 -79258
rect 53350 -79770 53446 -79736
rect 53694 -79770 53790 -79736
rect 53886 -79508 53982 -79474
rect 54956 -79508 55052 -79474
rect 53886 -79570 53920 -79508
rect 55018 -79570 55052 -79508
rect 54065 -79622 54081 -79588
rect 54857 -79622 54873 -79588
rect 53988 -79650 54022 -79634
rect 53988 -79704 54022 -79688
rect 54916 -79650 54950 -79634
rect 54916 -79704 54950 -79688
rect 54065 -79750 54081 -79716
rect 54857 -79750 54873 -79716
rect 53886 -79830 53920 -79768
rect 55482 -79320 55516 -79258
rect 55280 -79348 55314 -79332
rect 55280 -79540 55314 -79524
rect 55368 -79348 55402 -79332
rect 55368 -79540 55402 -79524
rect 55308 -79608 55324 -79574
rect 55358 -79608 55374 -79574
rect 55166 -79676 55200 -79614
rect 55482 -79676 55516 -79614
rect 55166 -79710 55262 -79676
rect 55420 -79710 55516 -79676
rect 55018 -79830 55052 -79768
rect 56112 -78764 56146 -78702
rect 56350 -78138 56412 -78118
rect 56610 -78138 56706 -78104
rect 56672 -78200 56706 -78138
rect 57303 -78083 57355 -78054
rect 57131 -78155 57165 -78134
rect 57201 -78147 57217 -78113
rect 57251 -78147 57267 -78113
rect 57201 -78189 57267 -78147
rect 57337 -78117 57355 -78083
rect 57303 -78155 57355 -78117
rect 58930 -78010 59026 -77976
rect 59214 -77977 59310 -77976
rect 59662 -77977 59696 -77920
rect 59772 -77894 59866 -77860
rect 60426 -77894 60520 -77860
rect 59772 -77950 59806 -77894
rect 59214 -78010 59696 -77977
rect 58930 -78011 59696 -78010
rect 58930 -78072 58964 -78011
rect 59276 -78072 59310 -78011
rect 59087 -78112 59103 -78078
rect 59137 -78112 59153 -78078
rect 56476 -78240 56492 -78206
rect 56530 -78240 56546 -78206
rect 55866 -78804 55882 -78770
rect 55970 -78804 55986 -78770
rect 55820 -78854 55854 -78838
rect 55820 -79646 55854 -79630
rect 55998 -78854 56032 -78838
rect 55998 -79646 56032 -79630
rect 55866 -79714 55882 -79680
rect 55970 -79714 55986 -79680
rect 55706 -79782 55740 -79720
rect 56430 -78299 56464 -78283
rect 56430 -79091 56464 -79075
rect 56558 -78299 56592 -78283
rect 56558 -79091 56592 -79075
rect 56476 -79168 56492 -79134
rect 56530 -79168 56546 -79134
rect 56316 -79236 56350 -79174
rect 57096 -78223 57125 -78189
rect 57159 -78223 57217 -78189
rect 57251 -78223 57309 -78189
rect 57343 -78223 57372 -78189
rect 59044 -78171 59078 -78155
rect 59044 -78563 59078 -78547
rect 59162 -78171 59196 -78155
rect 59162 -78563 59196 -78547
rect 59087 -78640 59103 -78606
rect 59137 -78640 59153 -78606
rect 60486 -77956 60520 -77894
rect 59942 -78008 59958 -77974
rect 60334 -78008 60350 -77974
rect 59874 -78028 59908 -78012
rect 59874 -78078 59908 -78062
rect 60384 -78028 60418 -78012
rect 60384 -78078 60418 -78062
rect 59942 -78116 59958 -78082
rect 60334 -78116 60350 -78082
rect 59772 -78196 59806 -78140
rect 60486 -78196 60520 -78134
rect 59388 -78230 59476 -78196
rect 59656 -78230 59800 -78196
rect 59958 -78230 60520 -78196
rect 59388 -78290 59422 -78230
rect 59276 -78706 59310 -78646
rect 59530 -78332 59546 -78298
rect 59580 -78332 59596 -78298
rect 59502 -78382 59536 -78366
rect 59502 -78574 59536 -78558
rect 59590 -78382 59624 -78366
rect 59590 -78574 59624 -78558
rect 59530 -78642 59546 -78608
rect 59580 -78642 59596 -78608
rect 58966 -78742 59310 -78706
rect 59388 -78709 59422 -78650
rect 59704 -78709 59738 -78230
rect 60020 -78292 60054 -78230
rect 59846 -78332 59862 -78298
rect 59896 -78332 59912 -78298
rect 59818 -78382 59852 -78366
rect 59818 -78574 59852 -78558
rect 59906 -78382 59940 -78366
rect 59906 -78574 59940 -78558
rect 59846 -78642 59862 -78608
rect 59896 -78642 59912 -78608
rect 61186 -78400 61286 -78390
rect 61186 -78480 61196 -78400
rect 61186 -78490 61286 -78480
rect 60020 -78709 60054 -78648
rect 56672 -79236 56706 -79174
rect 57096 -79199 57125 -79165
rect 57159 -79199 57217 -79165
rect 57251 -79199 57309 -79165
rect 57343 -79199 57372 -79165
rect 56316 -79270 56412 -79236
rect 56610 -79270 56706 -79236
rect 57131 -79254 57165 -79233
rect 57201 -79241 57267 -79199
rect 57201 -79275 57217 -79241
rect 57251 -79275 57267 -79241
rect 57303 -79271 57355 -79233
rect 57131 -79309 57165 -79288
rect 57337 -79305 57355 -79271
rect 59276 -78802 59310 -78742
rect 59387 -78744 60054 -78709
rect 60127 -78554 60161 -78528
rect 60127 -78557 60253 -78554
rect 60161 -78573 60253 -78557
rect 60161 -78591 60203 -78573
rect 60127 -78607 60203 -78591
rect 60237 -78607 60253 -78573
rect 60359 -78560 60409 -78549
rect 60671 -78554 60705 -78528
rect 60359 -78565 60366 -78560
rect 60359 -78600 60366 -78599
rect 60406 -78600 60409 -78560
rect 60127 -78649 60161 -78607
rect 60127 -78741 60161 -78683
rect 60195 -78657 60325 -78641
rect 60195 -78691 60211 -78657
rect 60245 -78691 60325 -78657
rect 60195 -78707 60325 -78691
rect 59387 -78800 59421 -78744
rect 59087 -78842 59103 -78808
rect 59137 -78842 59153 -78808
rect 59044 -78901 59078 -78885
rect 57131 -79343 57264 -79309
rect 57303 -79334 57355 -79305
rect 57117 -79394 57185 -79379
rect 57117 -79444 57118 -79394
rect 57168 -79444 57185 -79394
rect 57117 -79453 57185 -79444
rect 57230 -79394 57264 -79343
rect 57319 -79370 57355 -79334
rect 57230 -79410 57285 -79394
rect 57230 -79444 57251 -79410
rect 57230 -79460 57285 -79444
rect 57319 -79410 57326 -79370
rect 59044 -79293 59078 -79277
rect 59162 -78901 59196 -78885
rect 59162 -79293 59196 -79277
rect 59087 -79370 59103 -79336
rect 59137 -79370 59153 -79336
rect 57230 -79489 57264 -79460
rect 57129 -79523 57264 -79489
rect 57319 -79494 57355 -79410
rect 57129 -79557 57165 -79523
rect 57301 -79544 57355 -79494
rect 58930 -79438 58964 -79376
rect 59529 -78845 59545 -78811
rect 59579 -78845 59595 -78811
rect 59501 -78895 59535 -78879
rect 59501 -79087 59535 -79071
rect 59589 -78895 59623 -78879
rect 59589 -79087 59623 -79071
rect 59529 -79155 59545 -79121
rect 59579 -79155 59595 -79121
rect 59387 -79223 59421 -79170
rect 59703 -79223 59737 -78744
rect 60019 -78805 60053 -78744
rect 59845 -78845 59861 -78811
rect 59895 -78845 59911 -78811
rect 59817 -78895 59851 -78879
rect 59817 -79087 59851 -79071
rect 59905 -78895 59939 -78879
rect 59905 -79087 59939 -79071
rect 59845 -79155 59861 -79121
rect 59895 -79155 59911 -79121
rect 60161 -78775 60203 -78741
rect 60237 -78775 60253 -78741
rect 60127 -78833 60161 -78775
rect 60289 -78809 60325 -78707
rect 60127 -78909 60161 -78867
rect 60195 -78825 60325 -78809
rect 60195 -78859 60211 -78825
rect 60245 -78859 60325 -78825
rect 60195 -78875 60325 -78859
rect 60359 -78650 60409 -78600
rect 60443 -78557 60705 -78554
rect 60443 -78573 60671 -78557
rect 60443 -78607 60459 -78573
rect 60493 -78607 60527 -78573
rect 60561 -78607 60595 -78573
rect 60629 -78591 60671 -78573
rect 60629 -78607 60705 -78591
rect 60359 -78657 60366 -78650
rect 60406 -78690 60409 -78650
rect 60393 -78691 60409 -78690
rect 60359 -78740 60409 -78691
rect 60359 -78741 60366 -78740
rect 60359 -78780 60366 -78775
rect 60406 -78780 60409 -78740
rect 60359 -78820 60409 -78780
rect 60359 -78825 60366 -78820
rect 60359 -78860 60366 -78859
rect 60406 -78860 60409 -78820
rect 60359 -78875 60409 -78860
rect 60443 -78657 60637 -78641
rect 60443 -78691 60459 -78657
rect 60493 -78691 60527 -78657
rect 60561 -78691 60595 -78657
rect 60629 -78691 60637 -78657
rect 60443 -78707 60637 -78691
rect 60671 -78649 60705 -78607
rect 60443 -78809 60477 -78707
rect 60671 -78741 60705 -78683
rect 60511 -78775 60527 -78741
rect 60561 -78775 60595 -78741
rect 60629 -78775 60671 -78741
rect 60443 -78825 60637 -78809
rect 60443 -78859 60459 -78825
rect 60493 -78859 60527 -78825
rect 60561 -78859 60595 -78825
rect 60629 -78859 60637 -78825
rect 60443 -78875 60637 -78859
rect 60671 -78833 60705 -78775
rect 60289 -78909 60325 -78875
rect 60443 -78909 60481 -78875
rect 60671 -78909 60705 -78867
rect 60127 -78925 60204 -78909
rect 60161 -78943 60204 -78925
rect 60238 -78943 60254 -78909
rect 60161 -78959 60254 -78943
rect 60289 -78925 60481 -78909
rect 60289 -78959 60297 -78925
rect 60331 -78959 60369 -78925
rect 60405 -78959 60449 -78925
rect 60579 -78943 60595 -78909
rect 60629 -78925 60705 -78909
rect 60629 -78943 60671 -78925
rect 60579 -78951 60671 -78943
rect 60127 -78988 60161 -78959
rect 60289 -78962 60481 -78959
rect 60671 -78988 60705 -78959
rect 60747 -78554 60781 -78528
rect 60747 -78557 61009 -78554
rect 60781 -78573 61009 -78557
rect 60781 -78591 60823 -78573
rect 60747 -78607 60823 -78591
rect 60857 -78607 60891 -78573
rect 60925 -78607 60959 -78573
rect 60993 -78607 61009 -78573
rect 61043 -78560 61093 -78549
rect 61291 -78554 61325 -78528
rect 61043 -78600 61046 -78560
rect 61086 -78565 61093 -78560
rect 61086 -78600 61093 -78599
rect 60747 -78649 60781 -78607
rect 60747 -78741 60781 -78683
rect 60815 -78657 61009 -78641
rect 60815 -78691 60823 -78657
rect 60857 -78691 60891 -78657
rect 60925 -78691 60959 -78657
rect 60993 -78691 61009 -78657
rect 60815 -78707 61009 -78691
rect 60781 -78775 60823 -78741
rect 60857 -78775 60891 -78741
rect 60925 -78775 60941 -78741
rect 60747 -78833 60781 -78775
rect 60975 -78809 61009 -78707
rect 60747 -78909 60781 -78867
rect 60815 -78825 61009 -78809
rect 60815 -78859 60823 -78825
rect 60857 -78859 60891 -78825
rect 60925 -78859 60959 -78825
rect 60993 -78859 61009 -78825
rect 60815 -78875 61009 -78859
rect 61043 -78650 61093 -78600
rect 61199 -78557 61325 -78554
rect 61199 -78573 61291 -78557
rect 61199 -78607 61215 -78573
rect 61249 -78591 61291 -78573
rect 61249 -78607 61325 -78591
rect 61043 -78690 61046 -78650
rect 61086 -78657 61093 -78650
rect 61043 -78691 61059 -78690
rect 61043 -78740 61093 -78691
rect 61043 -78780 61046 -78740
rect 61086 -78741 61093 -78740
rect 61086 -78780 61093 -78775
rect 61043 -78820 61093 -78780
rect 61043 -78860 61046 -78820
rect 61086 -78825 61093 -78820
rect 61086 -78860 61093 -78859
rect 61043 -78875 61093 -78860
rect 61127 -78657 61257 -78641
rect 61127 -78691 61207 -78657
rect 61241 -78691 61257 -78657
rect 61127 -78707 61257 -78691
rect 61291 -78649 61325 -78607
rect 61127 -78809 61163 -78707
rect 61291 -78741 61325 -78683
rect 61199 -78775 61215 -78741
rect 61249 -78775 61291 -78741
rect 61127 -78825 61257 -78809
rect 61127 -78859 61207 -78825
rect 61241 -78859 61257 -78825
rect 61127 -78875 61257 -78859
rect 61291 -78833 61325 -78775
rect 60971 -78909 61009 -78875
rect 61127 -78909 61163 -78875
rect 61291 -78909 61325 -78867
rect 60747 -78925 60823 -78909
rect 60781 -78943 60823 -78925
rect 60857 -78943 60873 -78909
rect 60781 -78951 60873 -78943
rect 60971 -78924 61163 -78909
rect 60971 -78925 61129 -78924
rect 60747 -78988 60781 -78959
rect 60971 -78959 60980 -78925
rect 61015 -78959 61053 -78925
rect 61088 -78958 61129 -78925
rect 61198 -78943 61214 -78909
rect 61248 -78925 61325 -78909
rect 61248 -78943 61291 -78925
rect 61088 -78959 61163 -78958
rect 61198 -78959 61291 -78943
rect 60971 -78962 61163 -78959
rect 61291 -78988 61325 -78959
rect 60466 -79060 60546 -79040
rect 60466 -79100 60486 -79060
rect 60526 -79100 60546 -79060
rect 60466 -79120 60546 -79100
rect 60606 -79060 60686 -79040
rect 60606 -79100 60626 -79060
rect 60666 -79100 60686 -79060
rect 60606 -79120 60686 -79100
rect 60746 -79060 60826 -79040
rect 60746 -79100 60766 -79060
rect 60806 -79100 60826 -79060
rect 60746 -79120 60826 -79100
rect 60886 -79060 60966 -79040
rect 60886 -79100 60906 -79060
rect 60946 -79100 60966 -79060
rect 60886 -79120 60966 -79100
rect 60019 -79223 60053 -79161
rect 59387 -79257 59476 -79223
rect 59646 -79257 59799 -79223
rect 59957 -79226 60053 -79223
rect 59957 -79257 60520 -79226
rect 59772 -79260 60520 -79257
rect 59772 -79320 59806 -79260
rect 59276 -79438 59310 -79376
rect 58930 -79472 59026 -79438
rect 59214 -79440 59310 -79438
rect 59214 -79472 59696 -79440
rect 58930 -79474 59696 -79472
rect 58930 -79510 58964 -79474
rect 57129 -79591 57131 -79557
rect 57129 -79625 57165 -79591
rect 57129 -79659 57131 -79625
rect 57129 -79675 57165 -79659
rect 57201 -79591 57217 -79557
rect 57251 -79591 57267 -79557
rect 57201 -79625 57267 -79591
rect 57201 -79659 57217 -79625
rect 57251 -79659 57267 -79625
rect 57201 -79709 57267 -79659
rect 57301 -79578 57303 -79544
rect 57337 -79578 57355 -79544
rect 57301 -79625 57355 -79578
rect 57301 -79659 57303 -79625
rect 57337 -79659 57355 -79625
rect 57301 -79675 57355 -79659
rect 59662 -79530 59696 -79474
rect 60486 -79322 60520 -79260
rect 59942 -79374 59958 -79340
rect 60334 -79374 60350 -79340
rect 59874 -79394 59908 -79378
rect 59874 -79444 59908 -79428
rect 60384 -79394 60418 -79378
rect 60384 -79444 60418 -79428
rect 59942 -79482 59958 -79448
rect 60334 -79482 60350 -79448
rect 56112 -79782 56146 -79720
rect 57096 -79743 57125 -79709
rect 57159 -79743 57217 -79709
rect 57251 -79743 57309 -79709
rect 57343 -79743 57372 -79709
rect 55706 -79816 55802 -79782
rect 56050 -79816 56146 -79782
rect 53886 -79864 53982 -79830
rect 54956 -79864 55052 -79830
rect 53886 -79926 53920 -79864
rect 55018 -79926 55052 -79864
rect 55720 -79858 56090 -79816
rect 55720 -79868 56020 -79858
rect 54065 -79978 54081 -79944
rect 54857 -79978 54873 -79944
rect 53988 -80006 54022 -79990
rect 53988 -80060 54022 -80044
rect 54916 -80006 54950 -79990
rect 54916 -80060 54950 -80044
rect 54065 -80106 54081 -80072
rect 54857 -80106 54873 -80072
rect 53886 -80186 53920 -80124
rect 56010 -80008 56020 -79868
rect 56080 -80008 56090 -79858
rect 59109 -79588 59125 -79554
rect 59501 -79588 59517 -79554
rect 59560 -79608 59594 -79592
rect 59560 -79658 59594 -79642
rect 59109 -79696 59125 -79662
rect 59501 -79696 59517 -79662
rect 59032 -79716 59066 -79700
rect 59032 -79766 59066 -79750
rect 59109 -79804 59125 -79770
rect 59501 -79804 59517 -79770
rect 56010 -80018 56090 -80008
rect 59772 -79562 59806 -79500
rect 60486 -79562 60520 -79500
rect 59772 -79596 59866 -79562
rect 60426 -79596 60520 -79562
rect 59662 -79884 59696 -79830
rect 58966 -79900 59026 -79884
rect 58930 -79918 59026 -79900
rect 59600 -79918 59696 -79884
rect 55018 -80186 55052 -80124
rect 53886 -80220 53982 -80186
rect 54956 -80220 55052 -80186
rect 55176 -80078 55272 -80044
rect 55566 -80078 55662 -80044
rect 55176 -80140 55210 -80078
rect 55628 -80140 55662 -80078
rect 55284 -80192 55300 -80158
rect 55476 -80192 55492 -80158
rect 55526 -80202 55560 -80186
rect 55284 -80280 55300 -80246
rect 55476 -80280 55492 -80246
rect 55526 -80252 55560 -80236
rect 55176 -80360 55210 -80298
rect 55628 -80360 55662 -80298
rect 55176 -80394 55272 -80360
rect 55566 -80394 55662 -80360
rect 53896 -82592 53992 -82558
rect 54966 -82592 55062 -82558
rect 53896 -82654 53930 -82592
rect 55028 -82654 55062 -82592
rect 54075 -82706 54091 -82672
rect 54867 -82706 54883 -82672
rect 53998 -82734 54032 -82718
rect 53998 -82788 54032 -82772
rect 54926 -82734 54960 -82718
rect 54926 -82788 54960 -82772
rect 54075 -82834 54091 -82800
rect 54867 -82834 54883 -82800
rect 53896 -82914 53930 -82852
rect 55028 -82914 55062 -82852
rect 55960 -82908 56040 -82898
rect 53896 -82948 53992 -82914
rect 54966 -82948 55062 -82914
rect 53350 -83038 53790 -83004
rect 53350 -83100 53384 -83038
rect 53510 -83140 53526 -83106
rect 53614 -83140 53630 -83106
rect 53464 -83190 53498 -83174
rect 53464 -83982 53498 -83966
rect 53642 -83190 53676 -83174
rect 53642 -83982 53676 -83966
rect 53756 -83664 53790 -83038
rect 53896 -83010 53930 -82948
rect 55028 -83010 55062 -82948
rect 55710 -82954 56040 -82908
rect 54075 -83062 54091 -83028
rect 54867 -83062 54883 -83028
rect 53998 -83090 54032 -83074
rect 53998 -83144 54032 -83128
rect 54926 -83090 54960 -83074
rect 54926 -83144 54960 -83128
rect 54075 -83190 54091 -83156
rect 54867 -83190 54883 -83156
rect 53896 -83270 53930 -83208
rect 55706 -82988 55802 -82954
rect 56050 -82988 56146 -82954
rect 55706 -83050 55740 -82988
rect 55028 -83270 55062 -83208
rect 53896 -83304 53992 -83270
rect 54966 -83304 55062 -83270
rect 55176 -83100 55272 -83066
rect 55430 -83100 55526 -83066
rect 55176 -83162 55210 -83100
rect 55492 -83162 55526 -83100
rect 55318 -83202 55334 -83168
rect 55368 -83202 55384 -83168
rect 55290 -83252 55324 -83236
rect 55290 -83444 55324 -83428
rect 55378 -83252 55412 -83236
rect 55378 -83444 55412 -83428
rect 55176 -83518 55210 -83456
rect 55492 -83518 55526 -83456
rect 54870 -83552 55272 -83518
rect 55430 -83552 55706 -83518
rect 54870 -83558 55706 -83552
rect 54870 -83664 54904 -83558
rect 53756 -83698 53852 -83664
rect 54808 -83698 54904 -83664
rect 53756 -83760 53790 -83698
rect 54870 -83760 54904 -83698
rect 55126 -83708 55142 -83674
rect 55494 -83708 55510 -83674
rect 53926 -83812 53942 -83778
rect 54718 -83812 54734 -83778
rect 53858 -83840 53892 -83824
rect 53858 -83944 53892 -83928
rect 54768 -83840 54802 -83824
rect 54768 -83944 54802 -83928
rect 53926 -83990 53942 -83956
rect 54718 -83990 54734 -83956
rect 53510 -84050 53526 -84016
rect 53614 -84050 53630 -84016
rect 53756 -84070 53790 -84008
rect 55046 -83760 55080 -83744
rect 55046 -83810 55080 -83794
rect 55556 -83760 55590 -83744
rect 55556 -83810 55590 -83794
rect 55126 -83880 55142 -83846
rect 55494 -83880 55510 -83846
rect 54870 -84038 54904 -84008
rect 55700 -84006 55706 -83558
rect 56112 -83050 56146 -82988
rect 58930 -82967 59026 -82933
rect 59600 -82967 59696 -82933
rect 58930 -83010 58964 -82967
rect 58926 -83020 58966 -83010
rect 55866 -83090 55882 -83056
rect 55970 -83090 55986 -83056
rect 55820 -83140 55854 -83124
rect 55820 -83932 55854 -83916
rect 55998 -83140 56032 -83124
rect 55998 -83932 56032 -83916
rect 55866 -84000 55882 -83966
rect 55970 -84000 55986 -83966
rect 55700 -84038 55740 -84006
rect 57096 -83079 57125 -83045
rect 57159 -83079 57217 -83045
rect 57251 -83079 57309 -83045
rect 57343 -83079 57372 -83045
rect 57129 -83129 57165 -83113
rect 57129 -83163 57131 -83129
rect 57129 -83197 57165 -83163
rect 57129 -83231 57131 -83197
rect 57201 -83129 57267 -83079
rect 57201 -83163 57217 -83129
rect 57251 -83163 57267 -83129
rect 57201 -83197 57267 -83163
rect 57201 -83231 57217 -83197
rect 57251 -83231 57267 -83197
rect 57301 -83129 57355 -83113
rect 57301 -83163 57303 -83129
rect 57337 -83163 57355 -83129
rect 57301 -83210 57355 -83163
rect 57129 -83265 57165 -83231
rect 57301 -83244 57303 -83210
rect 57337 -83244 57355 -83210
rect 57129 -83299 57264 -83265
rect 57301 -83294 57355 -83244
rect 57230 -83328 57264 -83299
rect 57117 -83344 57185 -83335
rect 57117 -83394 57118 -83344
rect 57178 -83394 57185 -83344
rect 57117 -83409 57185 -83394
rect 57230 -83344 57285 -83328
rect 57230 -83378 57251 -83344
rect 57230 -83394 57285 -83378
rect 57319 -83340 57355 -83294
rect 59662 -83029 59696 -82967
rect 59109 -83081 59125 -83047
rect 59501 -83081 59517 -83047
rect 59560 -83101 59594 -83085
rect 59560 -83151 59594 -83135
rect 59109 -83189 59125 -83155
rect 59501 -83189 59517 -83155
rect 59032 -83209 59066 -83193
rect 59032 -83259 59066 -83243
rect 59109 -83297 59125 -83263
rect 59501 -83297 59517 -83263
rect 58926 -83340 58966 -83320
rect 57319 -83380 57326 -83340
rect 58930 -83376 58964 -83340
rect 57230 -83445 57264 -83394
rect 57131 -83479 57264 -83445
rect 57319 -83454 57355 -83380
rect 57131 -83500 57165 -83479
rect 56316 -83518 56412 -83504
rect 54830 -84048 55830 -84038
rect 54830 -84070 55030 -84048
rect 53756 -84104 53852 -84070
rect 54808 -84104 55030 -84070
rect 53510 -84158 53526 -84124
rect 53614 -84158 53630 -84124
rect 53756 -84166 53790 -84104
rect 54830 -84128 55030 -84104
rect 55110 -84068 55740 -84048
rect 55810 -84068 55830 -84048
rect 56112 -84068 56146 -84006
rect 55110 -84108 55160 -84068
rect 55600 -84108 55740 -84068
rect 56050 -84102 56146 -84068
rect 55110 -84128 55740 -84108
rect 55810 -84128 55830 -84102
rect 54830 -84138 55830 -84128
rect 53464 -84208 53498 -84192
rect 53464 -85000 53498 -84984
rect 53642 -84208 53676 -84192
rect 53642 -85000 53676 -84984
rect 54870 -84166 54904 -84138
rect 53926 -84218 53942 -84184
rect 54718 -84218 54734 -84184
rect 53858 -84246 53892 -84230
rect 53858 -84350 53892 -84334
rect 54768 -84246 54802 -84230
rect 54768 -84350 54802 -84334
rect 53926 -84396 53942 -84362
rect 54718 -84396 54734 -84362
rect 53756 -84476 53790 -84414
rect 55700 -84164 55740 -84138
rect 55126 -84330 55142 -84296
rect 55494 -84330 55510 -84296
rect 54870 -84476 54904 -84414
rect 55046 -84382 55080 -84366
rect 55046 -84432 55080 -84416
rect 55556 -84382 55590 -84366
rect 55556 -84432 55590 -84416
rect 53756 -84510 53852 -84476
rect 54808 -84510 54904 -84476
rect 55126 -84502 55142 -84468
rect 55494 -84502 55510 -84468
rect 53510 -85068 53526 -85034
rect 53614 -85068 53630 -85034
rect 53350 -85136 53384 -85074
rect 53756 -85136 53790 -84510
rect 54870 -84618 54904 -84510
rect 55700 -84618 55706 -84164
rect 54870 -84624 55706 -84618
rect 54870 -84658 55262 -84624
rect 55420 -84658 55706 -84624
rect 55166 -84720 55200 -84658
rect 53350 -85170 53446 -85136
rect 53694 -85170 53790 -85136
rect 53886 -84908 53982 -84874
rect 54956 -84908 55052 -84874
rect 53886 -84970 53920 -84908
rect 55018 -84970 55052 -84908
rect 54065 -85022 54081 -84988
rect 54857 -85022 54873 -84988
rect 53988 -85050 54022 -85034
rect 53988 -85104 54022 -85088
rect 54916 -85050 54950 -85034
rect 54916 -85104 54950 -85088
rect 54065 -85150 54081 -85116
rect 54857 -85150 54873 -85116
rect 53886 -85230 53920 -85168
rect 55482 -84720 55516 -84658
rect 55280 -84748 55314 -84732
rect 55280 -84940 55314 -84924
rect 55368 -84748 55402 -84732
rect 55368 -84940 55402 -84924
rect 55308 -85008 55324 -84974
rect 55358 -85008 55374 -84974
rect 55166 -85076 55200 -85014
rect 55482 -85076 55516 -85014
rect 55166 -85110 55262 -85076
rect 55420 -85110 55516 -85076
rect 55018 -85230 55052 -85168
rect 56112 -84164 56146 -84102
rect 56350 -83538 56412 -83518
rect 56610 -83538 56706 -83504
rect 56672 -83600 56706 -83538
rect 57303 -83483 57355 -83454
rect 57131 -83555 57165 -83534
rect 57201 -83547 57217 -83513
rect 57251 -83547 57267 -83513
rect 57201 -83589 57267 -83547
rect 57337 -83517 57355 -83483
rect 57303 -83555 57355 -83517
rect 58930 -83410 59026 -83376
rect 59214 -83377 59310 -83376
rect 59662 -83377 59696 -83320
rect 59772 -83294 59866 -83260
rect 60426 -83294 60520 -83260
rect 59772 -83350 59806 -83294
rect 59214 -83410 59696 -83377
rect 58930 -83411 59696 -83410
rect 58930 -83472 58964 -83411
rect 59276 -83472 59310 -83411
rect 59087 -83512 59103 -83478
rect 59137 -83512 59153 -83478
rect 56476 -83640 56492 -83606
rect 56530 -83640 56546 -83606
rect 55866 -84204 55882 -84170
rect 55970 -84204 55986 -84170
rect 55820 -84254 55854 -84238
rect 55820 -85046 55854 -85030
rect 55998 -84254 56032 -84238
rect 55998 -85046 56032 -85030
rect 55866 -85114 55882 -85080
rect 55970 -85114 55986 -85080
rect 55706 -85182 55740 -85120
rect 56430 -83699 56464 -83683
rect 56430 -84491 56464 -84475
rect 56558 -83699 56592 -83683
rect 56558 -84491 56592 -84475
rect 56476 -84568 56492 -84534
rect 56530 -84568 56546 -84534
rect 56316 -84636 56350 -84574
rect 57096 -83623 57125 -83589
rect 57159 -83623 57217 -83589
rect 57251 -83623 57309 -83589
rect 57343 -83623 57372 -83589
rect 59044 -83571 59078 -83555
rect 59044 -83963 59078 -83947
rect 59162 -83571 59196 -83555
rect 59162 -83963 59196 -83947
rect 59087 -84040 59103 -84006
rect 59137 -84040 59153 -84006
rect 60486 -83356 60520 -83294
rect 59942 -83408 59958 -83374
rect 60334 -83408 60350 -83374
rect 59874 -83428 59908 -83412
rect 59874 -83478 59908 -83462
rect 60384 -83428 60418 -83412
rect 60384 -83478 60418 -83462
rect 59942 -83516 59958 -83482
rect 60334 -83516 60350 -83482
rect 59772 -83596 59806 -83540
rect 60486 -83596 60520 -83534
rect 59388 -83630 59476 -83596
rect 59656 -83630 59800 -83596
rect 59958 -83630 60520 -83596
rect 59388 -83690 59422 -83630
rect 59276 -84106 59310 -84046
rect 59530 -83732 59546 -83698
rect 59580 -83732 59596 -83698
rect 59502 -83782 59536 -83766
rect 59502 -83974 59536 -83958
rect 59590 -83782 59624 -83766
rect 59590 -83974 59624 -83958
rect 59530 -84042 59546 -84008
rect 59580 -84042 59596 -84008
rect 58966 -84142 59310 -84106
rect 59388 -84109 59422 -84050
rect 59704 -84109 59738 -83630
rect 60020 -83692 60054 -83630
rect 59846 -83732 59862 -83698
rect 59896 -83732 59912 -83698
rect 59818 -83782 59852 -83766
rect 59818 -83974 59852 -83958
rect 59906 -83782 59940 -83766
rect 59906 -83974 59940 -83958
rect 59846 -84042 59862 -84008
rect 59896 -84042 59912 -84008
rect 61186 -83800 61286 -83790
rect 61186 -83880 61196 -83800
rect 61186 -83890 61286 -83880
rect 60020 -84109 60054 -84048
rect 56672 -84636 56706 -84574
rect 57096 -84599 57125 -84565
rect 57159 -84599 57217 -84565
rect 57251 -84599 57309 -84565
rect 57343 -84599 57372 -84565
rect 56316 -84670 56412 -84636
rect 56610 -84670 56706 -84636
rect 57131 -84654 57165 -84633
rect 57201 -84641 57267 -84599
rect 57201 -84675 57217 -84641
rect 57251 -84675 57267 -84641
rect 57303 -84671 57355 -84633
rect 57131 -84709 57165 -84688
rect 57337 -84705 57355 -84671
rect 59276 -84202 59310 -84142
rect 59387 -84144 60054 -84109
rect 60127 -83954 60161 -83928
rect 60127 -83957 60253 -83954
rect 60161 -83973 60253 -83957
rect 60161 -83991 60203 -83973
rect 60127 -84007 60203 -83991
rect 60237 -84007 60253 -83973
rect 60359 -83960 60409 -83949
rect 60671 -83954 60705 -83928
rect 60359 -83965 60366 -83960
rect 60359 -84000 60366 -83999
rect 60406 -84000 60409 -83960
rect 60127 -84049 60161 -84007
rect 60127 -84141 60161 -84083
rect 60195 -84057 60325 -84041
rect 60195 -84091 60211 -84057
rect 60245 -84091 60325 -84057
rect 60195 -84107 60325 -84091
rect 59387 -84200 59421 -84144
rect 59087 -84242 59103 -84208
rect 59137 -84242 59153 -84208
rect 59044 -84301 59078 -84285
rect 57131 -84743 57264 -84709
rect 57303 -84734 57355 -84705
rect 57117 -84794 57185 -84779
rect 57117 -84844 57118 -84794
rect 57168 -84844 57185 -84794
rect 57117 -84853 57185 -84844
rect 57230 -84794 57264 -84743
rect 57319 -84770 57355 -84734
rect 57230 -84810 57285 -84794
rect 57230 -84844 57251 -84810
rect 57230 -84860 57285 -84844
rect 57319 -84810 57326 -84770
rect 59044 -84693 59078 -84677
rect 59162 -84301 59196 -84285
rect 59162 -84693 59196 -84677
rect 59087 -84770 59103 -84736
rect 59137 -84770 59153 -84736
rect 57230 -84889 57264 -84860
rect 57129 -84923 57264 -84889
rect 57319 -84894 57355 -84810
rect 57129 -84957 57165 -84923
rect 57301 -84944 57355 -84894
rect 58930 -84838 58964 -84776
rect 59529 -84245 59545 -84211
rect 59579 -84245 59595 -84211
rect 59501 -84295 59535 -84279
rect 59501 -84487 59535 -84471
rect 59589 -84295 59623 -84279
rect 59589 -84487 59623 -84471
rect 59529 -84555 59545 -84521
rect 59579 -84555 59595 -84521
rect 59387 -84623 59421 -84570
rect 59703 -84623 59737 -84144
rect 60019 -84205 60053 -84144
rect 59845 -84245 59861 -84211
rect 59895 -84245 59911 -84211
rect 59817 -84295 59851 -84279
rect 59817 -84487 59851 -84471
rect 59905 -84295 59939 -84279
rect 59905 -84487 59939 -84471
rect 59845 -84555 59861 -84521
rect 59895 -84555 59911 -84521
rect 60161 -84175 60203 -84141
rect 60237 -84175 60253 -84141
rect 60127 -84233 60161 -84175
rect 60289 -84209 60325 -84107
rect 60127 -84309 60161 -84267
rect 60195 -84225 60325 -84209
rect 60195 -84259 60211 -84225
rect 60245 -84259 60325 -84225
rect 60195 -84275 60325 -84259
rect 60359 -84050 60409 -84000
rect 60443 -83957 60705 -83954
rect 60443 -83973 60671 -83957
rect 60443 -84007 60459 -83973
rect 60493 -84007 60527 -83973
rect 60561 -84007 60595 -83973
rect 60629 -83991 60671 -83973
rect 60629 -84007 60705 -83991
rect 60359 -84057 60366 -84050
rect 60406 -84090 60409 -84050
rect 60393 -84091 60409 -84090
rect 60359 -84140 60409 -84091
rect 60359 -84141 60366 -84140
rect 60359 -84180 60366 -84175
rect 60406 -84180 60409 -84140
rect 60359 -84220 60409 -84180
rect 60359 -84225 60366 -84220
rect 60359 -84260 60366 -84259
rect 60406 -84260 60409 -84220
rect 60359 -84275 60409 -84260
rect 60443 -84057 60637 -84041
rect 60443 -84091 60459 -84057
rect 60493 -84091 60527 -84057
rect 60561 -84091 60595 -84057
rect 60629 -84091 60637 -84057
rect 60443 -84107 60637 -84091
rect 60671 -84049 60705 -84007
rect 60443 -84209 60477 -84107
rect 60671 -84141 60705 -84083
rect 60511 -84175 60527 -84141
rect 60561 -84175 60595 -84141
rect 60629 -84175 60671 -84141
rect 60443 -84225 60637 -84209
rect 60443 -84259 60459 -84225
rect 60493 -84259 60527 -84225
rect 60561 -84259 60595 -84225
rect 60629 -84259 60637 -84225
rect 60443 -84275 60637 -84259
rect 60671 -84233 60705 -84175
rect 60289 -84309 60325 -84275
rect 60443 -84309 60481 -84275
rect 60671 -84309 60705 -84267
rect 60127 -84325 60204 -84309
rect 60161 -84343 60204 -84325
rect 60238 -84343 60254 -84309
rect 60161 -84359 60254 -84343
rect 60289 -84325 60481 -84309
rect 60289 -84359 60297 -84325
rect 60331 -84359 60369 -84325
rect 60405 -84359 60449 -84325
rect 60579 -84343 60595 -84309
rect 60629 -84325 60705 -84309
rect 60629 -84343 60671 -84325
rect 60579 -84351 60671 -84343
rect 60127 -84388 60161 -84359
rect 60289 -84362 60481 -84359
rect 60671 -84388 60705 -84359
rect 60747 -83954 60781 -83928
rect 60747 -83957 61009 -83954
rect 60781 -83973 61009 -83957
rect 60781 -83991 60823 -83973
rect 60747 -84007 60823 -83991
rect 60857 -84007 60891 -83973
rect 60925 -84007 60959 -83973
rect 60993 -84007 61009 -83973
rect 61043 -83960 61093 -83949
rect 61291 -83954 61325 -83928
rect 61043 -84000 61046 -83960
rect 61086 -83965 61093 -83960
rect 61086 -84000 61093 -83999
rect 60747 -84049 60781 -84007
rect 60747 -84141 60781 -84083
rect 60815 -84057 61009 -84041
rect 60815 -84091 60823 -84057
rect 60857 -84091 60891 -84057
rect 60925 -84091 60959 -84057
rect 60993 -84091 61009 -84057
rect 60815 -84107 61009 -84091
rect 60781 -84175 60823 -84141
rect 60857 -84175 60891 -84141
rect 60925 -84175 60941 -84141
rect 60747 -84233 60781 -84175
rect 60975 -84209 61009 -84107
rect 60747 -84309 60781 -84267
rect 60815 -84225 61009 -84209
rect 60815 -84259 60823 -84225
rect 60857 -84259 60891 -84225
rect 60925 -84259 60959 -84225
rect 60993 -84259 61009 -84225
rect 60815 -84275 61009 -84259
rect 61043 -84050 61093 -84000
rect 61199 -83957 61325 -83954
rect 61199 -83973 61291 -83957
rect 61199 -84007 61215 -83973
rect 61249 -83991 61291 -83973
rect 61249 -84007 61325 -83991
rect 61043 -84090 61046 -84050
rect 61086 -84057 61093 -84050
rect 61043 -84091 61059 -84090
rect 61043 -84140 61093 -84091
rect 61043 -84180 61046 -84140
rect 61086 -84141 61093 -84140
rect 61086 -84180 61093 -84175
rect 61043 -84220 61093 -84180
rect 61043 -84260 61046 -84220
rect 61086 -84225 61093 -84220
rect 61086 -84260 61093 -84259
rect 61043 -84275 61093 -84260
rect 61127 -84057 61257 -84041
rect 61127 -84091 61207 -84057
rect 61241 -84091 61257 -84057
rect 61127 -84107 61257 -84091
rect 61291 -84049 61325 -84007
rect 61127 -84209 61163 -84107
rect 61291 -84141 61325 -84083
rect 61199 -84175 61215 -84141
rect 61249 -84175 61291 -84141
rect 61127 -84225 61257 -84209
rect 61127 -84259 61207 -84225
rect 61241 -84259 61257 -84225
rect 61127 -84275 61257 -84259
rect 61291 -84233 61325 -84175
rect 60971 -84309 61009 -84275
rect 61127 -84309 61163 -84275
rect 61291 -84309 61325 -84267
rect 60747 -84325 60823 -84309
rect 60781 -84343 60823 -84325
rect 60857 -84343 60873 -84309
rect 60781 -84351 60873 -84343
rect 60971 -84324 61163 -84309
rect 60971 -84325 61129 -84324
rect 60747 -84388 60781 -84359
rect 60971 -84359 60980 -84325
rect 61015 -84359 61053 -84325
rect 61088 -84358 61129 -84325
rect 61198 -84343 61214 -84309
rect 61248 -84325 61325 -84309
rect 61248 -84343 61291 -84325
rect 61088 -84359 61163 -84358
rect 61198 -84359 61291 -84343
rect 60971 -84362 61163 -84359
rect 61291 -84388 61325 -84359
rect 60466 -84460 60546 -84440
rect 60466 -84500 60486 -84460
rect 60526 -84500 60546 -84460
rect 60466 -84520 60546 -84500
rect 60606 -84460 60686 -84440
rect 60606 -84500 60626 -84460
rect 60666 -84500 60686 -84460
rect 60606 -84520 60686 -84500
rect 60746 -84460 60826 -84440
rect 60746 -84500 60766 -84460
rect 60806 -84500 60826 -84460
rect 60746 -84520 60826 -84500
rect 60886 -84460 60966 -84440
rect 60886 -84500 60906 -84460
rect 60946 -84500 60966 -84460
rect 60886 -84520 60966 -84500
rect 60019 -84623 60053 -84561
rect 59387 -84657 59476 -84623
rect 59646 -84657 59799 -84623
rect 59957 -84626 60053 -84623
rect 59957 -84657 60520 -84626
rect 59772 -84660 60520 -84657
rect 59772 -84720 59806 -84660
rect 59276 -84838 59310 -84776
rect 58930 -84872 59026 -84838
rect 59214 -84840 59310 -84838
rect 59214 -84872 59696 -84840
rect 58930 -84874 59696 -84872
rect 58930 -84910 58964 -84874
rect 57129 -84991 57131 -84957
rect 57129 -85025 57165 -84991
rect 57129 -85059 57131 -85025
rect 57129 -85075 57165 -85059
rect 57201 -84991 57217 -84957
rect 57251 -84991 57267 -84957
rect 57201 -85025 57267 -84991
rect 57201 -85059 57217 -85025
rect 57251 -85059 57267 -85025
rect 57201 -85109 57267 -85059
rect 57301 -84978 57303 -84944
rect 57337 -84978 57355 -84944
rect 57301 -85025 57355 -84978
rect 57301 -85059 57303 -85025
rect 57337 -85059 57355 -85025
rect 57301 -85075 57355 -85059
rect 59662 -84930 59696 -84874
rect 60486 -84722 60520 -84660
rect 59942 -84774 59958 -84740
rect 60334 -84774 60350 -84740
rect 59874 -84794 59908 -84778
rect 59874 -84844 59908 -84828
rect 60384 -84794 60418 -84778
rect 60384 -84844 60418 -84828
rect 59942 -84882 59958 -84848
rect 60334 -84882 60350 -84848
rect 56112 -85182 56146 -85120
rect 57096 -85143 57125 -85109
rect 57159 -85143 57217 -85109
rect 57251 -85143 57309 -85109
rect 57343 -85143 57372 -85109
rect 55706 -85216 55802 -85182
rect 56050 -85216 56146 -85182
rect 53886 -85264 53982 -85230
rect 54956 -85264 55052 -85230
rect 53886 -85326 53920 -85264
rect 55018 -85326 55052 -85264
rect 55720 -85258 56090 -85216
rect 55720 -85268 56020 -85258
rect 54065 -85378 54081 -85344
rect 54857 -85378 54873 -85344
rect 53988 -85406 54022 -85390
rect 53988 -85460 54022 -85444
rect 54916 -85406 54950 -85390
rect 54916 -85460 54950 -85444
rect 54065 -85506 54081 -85472
rect 54857 -85506 54873 -85472
rect 53886 -85586 53920 -85524
rect 56010 -85408 56020 -85268
rect 56080 -85408 56090 -85258
rect 59109 -84988 59125 -84954
rect 59501 -84988 59517 -84954
rect 59560 -85008 59594 -84992
rect 59560 -85058 59594 -85042
rect 59109 -85096 59125 -85062
rect 59501 -85096 59517 -85062
rect 59032 -85116 59066 -85100
rect 59032 -85166 59066 -85150
rect 59109 -85204 59125 -85170
rect 59501 -85204 59517 -85170
rect 56010 -85418 56090 -85408
rect 59772 -84962 59806 -84900
rect 60486 -84962 60520 -84900
rect 59772 -84996 59866 -84962
rect 60426 -84996 60520 -84962
rect 59662 -85284 59696 -85230
rect 58966 -85300 59026 -85284
rect 58930 -85318 59026 -85300
rect 59600 -85318 59696 -85284
rect 55018 -85586 55052 -85524
rect 53886 -85620 53982 -85586
rect 54956 -85620 55052 -85586
rect 55176 -85478 55272 -85444
rect 55566 -85478 55662 -85444
rect 55176 -85540 55210 -85478
rect 55628 -85540 55662 -85478
rect 55284 -85592 55300 -85558
rect 55476 -85592 55492 -85558
rect 55526 -85602 55560 -85586
rect 55284 -85680 55300 -85646
rect 55476 -85680 55492 -85646
rect 55526 -85652 55560 -85636
rect 55176 -85760 55210 -85698
rect 55628 -85760 55662 -85698
rect 55176 -85794 55272 -85760
rect 55566 -85794 55662 -85760
<< viali >>
rect 54150 -1558 54850 -1508
rect 54150 -1592 54850 -1558
rect 54150 -1598 54850 -1592
rect 54091 -1706 54867 -1672
rect 53998 -1772 54032 -1734
rect 54926 -1772 54960 -1734
rect 54091 -1834 54867 -1800
rect 55960 -1898 56040 -1728
rect 53526 -2140 53614 -2106
rect 53330 -3518 53350 -2168
rect 53350 -3518 53384 -2168
rect 53384 -3518 53400 -2168
rect 53464 -2966 53498 -2190
rect 53642 -2966 53676 -2190
rect 57126 -1900 57356 -1870
rect 54091 -2062 54867 -2028
rect 53998 -2128 54032 -2090
rect 54926 -2128 54960 -2090
rect 54091 -2190 54867 -2156
rect 55334 -2202 55368 -2168
rect 55290 -2428 55324 -2252
rect 55378 -2428 55412 -2252
rect 55142 -2708 55494 -2674
rect 53942 -2812 54718 -2778
rect 53858 -2928 53892 -2840
rect 54768 -2928 54802 -2840
rect 53942 -2990 54718 -2956
rect 53526 -3050 53614 -3016
rect 55046 -2794 55080 -2760
rect 55556 -2794 55590 -2760
rect 55142 -2880 55494 -2846
rect 57126 -1970 57156 -1900
rect 57156 -1970 57316 -1900
rect 57316 -1970 57356 -1900
rect 57126 -2000 57356 -1970
rect 58926 -2029 58966 -2020
rect 55882 -2090 55970 -2056
rect 55820 -2916 55854 -2140
rect 55998 -2916 56032 -2140
rect 55882 -3000 55970 -2966
rect 57125 -2079 57159 -2045
rect 57217 -2079 57251 -2045
rect 57309 -2079 57343 -2045
rect 57118 -2357 57178 -2344
rect 57118 -2391 57133 -2357
rect 57133 -2391 57167 -2357
rect 57167 -2391 57178 -2357
rect 57118 -2394 57178 -2391
rect 58926 -2315 58930 -2029
rect 58930 -2315 58964 -2029
rect 58964 -2315 58966 -2029
rect 59125 -2081 59501 -2047
rect 59560 -2135 59594 -2101
rect 59125 -2189 59501 -2155
rect 59032 -2243 59066 -2209
rect 59125 -2297 59501 -2263
rect 58926 -2320 58966 -2315
rect 59656 -2315 59662 -2030
rect 59662 -2315 59696 -2030
rect 59656 -2320 59696 -2315
rect 57326 -2380 57366 -2340
rect 53526 -3158 53614 -3124
rect 55030 -3128 55110 -3048
rect 55740 -3068 55810 -3048
rect 55740 -3102 55802 -3068
rect 55802 -3102 55810 -3068
rect 55740 -3128 55810 -3102
rect 53464 -3984 53498 -3208
rect 53642 -3984 53676 -3208
rect 53942 -3218 54718 -3184
rect 53858 -3334 53892 -3246
rect 54768 -3334 54802 -3246
rect 53942 -3396 54718 -3362
rect 55142 -3330 55494 -3296
rect 55046 -3416 55080 -3382
rect 55556 -3416 55590 -3382
rect 55142 -3502 55494 -3468
rect 53526 -4068 53614 -4034
rect 54081 -4022 54857 -3988
rect 53988 -4088 54022 -4050
rect 54916 -4088 54950 -4050
rect 54081 -4150 54857 -4116
rect 55280 -3924 55314 -3748
rect 55368 -3924 55402 -3748
rect 55324 -4008 55358 -3974
rect 56280 -2600 56350 -2518
rect 56280 -3148 56316 -2600
rect 56316 -3148 56350 -2600
rect 59866 -2294 59868 -2260
rect 59868 -2294 60424 -2260
rect 60424 -2294 60426 -2260
rect 59866 -2300 60426 -2294
rect 59766 -2356 59806 -2350
rect 59103 -2512 59137 -2478
rect 56492 -2640 56530 -2606
rect 55882 -3204 55970 -3170
rect 55820 -4030 55854 -3254
rect 55998 -4030 56032 -3254
rect 55882 -4114 55970 -4080
rect 56430 -3475 56464 -2699
rect 56558 -3475 56592 -2699
rect 56492 -3568 56530 -3534
rect 57125 -2623 57159 -2589
rect 57217 -2623 57251 -2589
rect 57309 -2623 57343 -2589
rect 57086 -2710 57376 -2680
rect 57086 -2780 57116 -2710
rect 57116 -2780 57346 -2710
rect 57346 -2780 57376 -2710
rect 57086 -2810 57376 -2780
rect 58926 -3046 58930 -2560
rect 58930 -3046 58964 -2560
rect 58964 -3046 58966 -2560
rect 59044 -2947 59078 -2571
rect 59162 -2947 59196 -2571
rect 59103 -3040 59137 -3006
rect 58926 -3202 58966 -3046
rect 59766 -2534 59772 -2356
rect 59772 -2534 59806 -2356
rect 59958 -2408 60334 -2374
rect 59874 -2462 59908 -2428
rect 60384 -2462 60418 -2428
rect 59958 -2516 60334 -2482
rect 59766 -2540 59806 -2534
rect 59476 -2596 59656 -2590
rect 59476 -2630 59484 -2596
rect 59484 -2630 59642 -2596
rect 59642 -2630 59656 -2596
rect 59386 -2692 59426 -2690
rect 59386 -3048 59388 -2692
rect 59388 -3048 59422 -2692
rect 59422 -3048 59426 -2692
rect 59546 -2732 59580 -2698
rect 59502 -2958 59536 -2782
rect 59590 -2958 59624 -2782
rect 59546 -3042 59580 -3008
rect 59386 -3050 59426 -3048
rect 59862 -2732 59896 -2698
rect 59818 -2958 59852 -2782
rect 59906 -2958 59940 -2782
rect 59862 -3042 59896 -3008
rect 61196 -2820 61366 -2800
rect 61196 -2860 61216 -2820
rect 61216 -2860 61336 -2820
rect 61336 -2860 61366 -2820
rect 61196 -2880 61366 -2860
rect 57056 -3370 57416 -3340
rect 57056 -3450 57096 -3370
rect 57096 -3450 57376 -3370
rect 57376 -3450 57416 -3370
rect 57056 -3480 57416 -3450
rect 57125 -3599 57159 -3565
rect 57217 -3599 57251 -3565
rect 57309 -3599 57343 -3565
rect 58926 -3690 58930 -3202
rect 58930 -3690 58964 -3202
rect 58964 -3690 58966 -3202
rect 60127 -2991 60161 -2957
rect 60366 -2965 60406 -2960
rect 60366 -2999 60393 -2965
rect 60393 -2999 60406 -2965
rect 60366 -3000 60406 -2999
rect 60127 -3083 60161 -3049
rect 59103 -3242 59137 -3208
rect 59044 -3677 59078 -3301
rect 57118 -3797 57168 -3794
rect 57118 -3831 57133 -3797
rect 57133 -3831 57167 -3797
rect 57167 -3831 57168 -3797
rect 57118 -3844 57168 -3831
rect 57326 -3810 57376 -3770
rect 59162 -3677 59196 -3301
rect 59103 -3770 59137 -3736
rect 59386 -3205 59426 -3200
rect 59386 -3561 59387 -3205
rect 59387 -3561 59421 -3205
rect 59421 -3561 59426 -3205
rect 59545 -3245 59579 -3211
rect 59501 -3471 59535 -3295
rect 59589 -3471 59623 -3295
rect 59545 -3555 59579 -3521
rect 59386 -3570 59426 -3561
rect 59476 -3623 59646 -3620
rect 59861 -3245 59895 -3211
rect 59817 -3471 59851 -3295
rect 59905 -3471 59939 -3295
rect 59861 -3555 59895 -3521
rect 60127 -3175 60161 -3141
rect 60127 -3267 60161 -3233
rect 60671 -2991 60705 -2957
rect 60366 -3057 60406 -3050
rect 60366 -3090 60393 -3057
rect 60393 -3090 60406 -3057
rect 60366 -3141 60406 -3140
rect 60366 -3175 60393 -3141
rect 60393 -3175 60406 -3141
rect 60366 -3180 60406 -3175
rect 60366 -3225 60406 -3220
rect 60366 -3259 60393 -3225
rect 60393 -3259 60406 -3225
rect 60366 -3260 60406 -3259
rect 60671 -3083 60705 -3049
rect 60671 -3175 60705 -3141
rect 60671 -3267 60705 -3233
rect 60127 -3359 60161 -3325
rect 60297 -3359 60331 -3325
rect 60369 -3359 60405 -3325
rect 60449 -3359 60484 -3325
rect 60671 -3359 60705 -3325
rect 60747 -2991 60781 -2957
rect 61046 -2965 61086 -2960
rect 61046 -2999 61059 -2965
rect 61059 -2999 61086 -2965
rect 61046 -3000 61086 -2999
rect 60747 -3083 60781 -3049
rect 60747 -3175 60781 -3141
rect 60747 -3267 60781 -3233
rect 61291 -2991 61325 -2957
rect 61046 -3057 61086 -3050
rect 61046 -3090 61059 -3057
rect 61059 -3090 61086 -3057
rect 61046 -3141 61086 -3140
rect 61046 -3175 61059 -3141
rect 61059 -3175 61086 -3141
rect 61046 -3180 61086 -3175
rect 61046 -3225 61086 -3220
rect 61046 -3259 61059 -3225
rect 61059 -3259 61086 -3225
rect 61046 -3260 61086 -3259
rect 61291 -3083 61325 -3049
rect 61291 -3175 61325 -3141
rect 61291 -3267 61325 -3233
rect 60747 -3359 60781 -3325
rect 60980 -3359 61015 -3325
rect 61053 -3359 61088 -3325
rect 61129 -3358 61164 -3324
rect 61291 -3359 61325 -3325
rect 60486 -3500 60526 -3460
rect 60626 -3500 60666 -3460
rect 60766 -3500 60806 -3460
rect 60906 -3500 60946 -3460
rect 59476 -3657 59483 -3623
rect 59483 -3657 59641 -3623
rect 59641 -3657 59646 -3623
rect 59476 -3660 59646 -3657
rect 59766 -3722 59806 -3720
rect 58926 -3936 58966 -3910
rect 59766 -3900 59772 -3722
rect 59772 -3900 59806 -3722
rect 59958 -3774 60334 -3740
rect 59874 -3828 59908 -3794
rect 60384 -3828 60418 -3794
rect 59958 -3882 60334 -3848
rect 57125 -4143 57159 -4109
rect 57217 -4143 57251 -4109
rect 57309 -4143 57343 -4109
rect 54081 -4378 54857 -4344
rect 53988 -4444 54022 -4406
rect 54916 -4444 54950 -4406
rect 54081 -4506 54857 -4472
rect 56020 -4408 56080 -4258
rect 58926 -4222 58930 -3936
rect 58930 -4222 58964 -3936
rect 58964 -4222 58966 -3936
rect 59656 -3936 59706 -3930
rect 59125 -3988 59501 -3954
rect 59560 -4042 59594 -4008
rect 59125 -4096 59501 -4062
rect 59032 -4150 59066 -4116
rect 59125 -4204 59501 -4170
rect 57156 -4290 57316 -4260
rect 57156 -4390 57186 -4290
rect 57186 -4390 57286 -4290
rect 57286 -4390 57316 -4290
rect 58926 -4300 58966 -4222
rect 59656 -4222 59662 -3936
rect 59662 -4222 59696 -3936
rect 59696 -4222 59706 -3936
rect 59866 -3962 60426 -3960
rect 59866 -3996 59868 -3962
rect 59868 -3996 60424 -3962
rect 60424 -3996 60426 -3962
rect 59866 -4000 60426 -3996
rect 59656 -4230 59706 -4222
rect 57156 -4420 57316 -4390
rect 54150 -4620 54840 -4588
rect 54150 -4708 54840 -4620
rect 55300 -4592 55476 -4558
rect 55526 -4636 55560 -4602
rect 55300 -4680 55476 -4646
rect 55320 -4760 55470 -4748
rect 55320 -4794 55470 -4760
rect 55320 -4808 55470 -4794
rect 54150 -6958 54850 -6908
rect 54150 -6992 54850 -6958
rect 54150 -6998 54850 -6992
rect 54091 -7106 54867 -7072
rect 53998 -7172 54032 -7134
rect 54926 -7172 54960 -7134
rect 54091 -7234 54867 -7200
rect 55960 -7298 56040 -7128
rect 53526 -7540 53614 -7506
rect 20908 -7809 21076 -7775
rect 20846 -11644 20880 -7868
rect 21104 -11644 21138 -7868
rect 21394 -7809 21562 -7775
rect 21206 -11619 21218 -7889
rect 21218 -11619 21252 -7889
rect 21252 -11619 21256 -7889
rect 20908 -11737 21076 -11703
rect 21332 -11644 21366 -7868
rect 21590 -11644 21624 -7868
rect 21880 -7809 22048 -7775
rect 21706 -11629 21738 -7889
rect 21738 -11629 21756 -7889
rect 21394 -11737 21562 -11703
rect 21818 -11644 21852 -7868
rect 22076 -11644 22110 -7868
rect 21880 -11737 22048 -11703
rect 53330 -8918 53350 -7568
rect 53350 -8918 53384 -7568
rect 53384 -8918 53400 -7568
rect 53464 -8366 53498 -7590
rect 53642 -8366 53676 -7590
rect 57126 -7300 57356 -7270
rect 54091 -7462 54867 -7428
rect 53998 -7528 54032 -7490
rect 54926 -7528 54960 -7490
rect 54091 -7590 54867 -7556
rect 55334 -7602 55368 -7568
rect 55290 -7828 55324 -7652
rect 55378 -7828 55412 -7652
rect 55142 -8108 55494 -8074
rect 53942 -8212 54718 -8178
rect 53858 -8328 53892 -8240
rect 54768 -8328 54802 -8240
rect 53942 -8390 54718 -8356
rect 53526 -8450 53614 -8416
rect 55046 -8194 55080 -8160
rect 55556 -8194 55590 -8160
rect 55142 -8280 55494 -8246
rect 57126 -7370 57156 -7300
rect 57156 -7370 57316 -7300
rect 57316 -7370 57356 -7300
rect 57126 -7400 57356 -7370
rect 58926 -7429 58966 -7420
rect 55882 -7490 55970 -7456
rect 55820 -8316 55854 -7540
rect 55998 -8316 56032 -7540
rect 55882 -8400 55970 -8366
rect 57125 -7479 57159 -7445
rect 57217 -7479 57251 -7445
rect 57309 -7479 57343 -7445
rect 57118 -7757 57178 -7744
rect 57118 -7791 57133 -7757
rect 57133 -7791 57167 -7757
rect 57167 -7791 57178 -7757
rect 57118 -7794 57178 -7791
rect 58926 -7715 58930 -7429
rect 58930 -7715 58964 -7429
rect 58964 -7715 58966 -7429
rect 59125 -7481 59501 -7447
rect 59560 -7535 59594 -7501
rect 59125 -7589 59501 -7555
rect 59032 -7643 59066 -7609
rect 59125 -7697 59501 -7663
rect 58926 -7720 58966 -7715
rect 59656 -7715 59662 -7430
rect 59662 -7715 59696 -7430
rect 59656 -7720 59696 -7715
rect 57326 -7780 57366 -7740
rect 53526 -8558 53614 -8524
rect 55030 -8528 55110 -8448
rect 55740 -8468 55810 -8448
rect 55740 -8502 55802 -8468
rect 55802 -8502 55810 -8468
rect 55740 -8528 55810 -8502
rect 53464 -9384 53498 -8608
rect 53642 -9384 53676 -8608
rect 53942 -8618 54718 -8584
rect 53858 -8734 53892 -8646
rect 54768 -8734 54802 -8646
rect 53942 -8796 54718 -8762
rect 55142 -8730 55494 -8696
rect 55046 -8816 55080 -8782
rect 55556 -8816 55590 -8782
rect 55142 -8902 55494 -8868
rect 53526 -9468 53614 -9434
rect 54081 -9422 54857 -9388
rect 53988 -9488 54022 -9450
rect 54916 -9488 54950 -9450
rect 54081 -9550 54857 -9516
rect 55280 -9324 55314 -9148
rect 55368 -9324 55402 -9148
rect 55324 -9408 55358 -9374
rect 56280 -8000 56350 -7918
rect 56280 -8548 56316 -8000
rect 56316 -8548 56350 -8000
rect 59866 -7694 59868 -7660
rect 59868 -7694 60424 -7660
rect 60424 -7694 60426 -7660
rect 59866 -7700 60426 -7694
rect 59766 -7756 59806 -7750
rect 59103 -7912 59137 -7878
rect 56492 -8040 56530 -8006
rect 55882 -8604 55970 -8570
rect 55820 -9430 55854 -8654
rect 55998 -9430 56032 -8654
rect 55882 -9514 55970 -9480
rect 56430 -8875 56464 -8099
rect 56558 -8875 56592 -8099
rect 56492 -8968 56530 -8934
rect 57125 -8023 57159 -7989
rect 57217 -8023 57251 -7989
rect 57309 -8023 57343 -7989
rect 57086 -8110 57376 -8080
rect 57086 -8180 57116 -8110
rect 57116 -8180 57346 -8110
rect 57346 -8180 57376 -8110
rect 57086 -8210 57376 -8180
rect 58926 -8446 58930 -7960
rect 58930 -8446 58964 -7960
rect 58964 -8446 58966 -7960
rect 59044 -8347 59078 -7971
rect 59162 -8347 59196 -7971
rect 59103 -8440 59137 -8406
rect 58926 -8602 58966 -8446
rect 59766 -7934 59772 -7756
rect 59772 -7934 59806 -7756
rect 59958 -7808 60334 -7774
rect 59874 -7862 59908 -7828
rect 60384 -7862 60418 -7828
rect 59958 -7916 60334 -7882
rect 59766 -7940 59806 -7934
rect 59476 -7996 59656 -7990
rect 59476 -8030 59484 -7996
rect 59484 -8030 59642 -7996
rect 59642 -8030 59656 -7996
rect 59386 -8092 59426 -8090
rect 59386 -8448 59388 -8092
rect 59388 -8448 59422 -8092
rect 59422 -8448 59426 -8092
rect 59546 -8132 59580 -8098
rect 59502 -8358 59536 -8182
rect 59590 -8358 59624 -8182
rect 59546 -8442 59580 -8408
rect 59386 -8450 59426 -8448
rect 59862 -8132 59896 -8098
rect 59818 -8358 59852 -8182
rect 59906 -8358 59940 -8182
rect 59862 -8442 59896 -8408
rect 61196 -8220 61366 -8200
rect 61196 -8260 61216 -8220
rect 61216 -8260 61336 -8220
rect 61336 -8260 61366 -8220
rect 61196 -8280 61366 -8260
rect 57056 -8770 57416 -8740
rect 57056 -8850 57096 -8770
rect 57096 -8850 57376 -8770
rect 57376 -8850 57416 -8770
rect 57056 -8880 57416 -8850
rect 57125 -8999 57159 -8965
rect 57217 -8999 57251 -8965
rect 57309 -8999 57343 -8965
rect 58926 -9090 58930 -8602
rect 58930 -9090 58964 -8602
rect 58964 -9090 58966 -8602
rect 60127 -8391 60161 -8357
rect 60366 -8365 60406 -8360
rect 60366 -8399 60393 -8365
rect 60393 -8399 60406 -8365
rect 60366 -8400 60406 -8399
rect 60127 -8483 60161 -8449
rect 59103 -8642 59137 -8608
rect 59044 -9077 59078 -8701
rect 57118 -9197 57168 -9194
rect 57118 -9231 57133 -9197
rect 57133 -9231 57167 -9197
rect 57167 -9231 57168 -9197
rect 57118 -9244 57168 -9231
rect 57326 -9210 57376 -9170
rect 59162 -9077 59196 -8701
rect 59103 -9170 59137 -9136
rect 59386 -8605 59426 -8600
rect 59386 -8961 59387 -8605
rect 59387 -8961 59421 -8605
rect 59421 -8961 59426 -8605
rect 59545 -8645 59579 -8611
rect 59501 -8871 59535 -8695
rect 59589 -8871 59623 -8695
rect 59545 -8955 59579 -8921
rect 59386 -8970 59426 -8961
rect 59476 -9023 59646 -9020
rect 59861 -8645 59895 -8611
rect 59817 -8871 59851 -8695
rect 59905 -8871 59939 -8695
rect 59861 -8955 59895 -8921
rect 60127 -8575 60161 -8541
rect 60127 -8667 60161 -8633
rect 60671 -8391 60705 -8357
rect 60366 -8457 60406 -8450
rect 60366 -8490 60393 -8457
rect 60393 -8490 60406 -8457
rect 60366 -8541 60406 -8540
rect 60366 -8575 60393 -8541
rect 60393 -8575 60406 -8541
rect 60366 -8580 60406 -8575
rect 60366 -8625 60406 -8620
rect 60366 -8659 60393 -8625
rect 60393 -8659 60406 -8625
rect 60366 -8660 60406 -8659
rect 60671 -8483 60705 -8449
rect 60671 -8575 60705 -8541
rect 60671 -8667 60705 -8633
rect 60127 -8759 60161 -8725
rect 60297 -8759 60331 -8725
rect 60369 -8759 60405 -8725
rect 60449 -8759 60484 -8725
rect 60671 -8759 60705 -8725
rect 60747 -8391 60781 -8357
rect 61046 -8365 61086 -8360
rect 61046 -8399 61059 -8365
rect 61059 -8399 61086 -8365
rect 61046 -8400 61086 -8399
rect 60747 -8483 60781 -8449
rect 60747 -8575 60781 -8541
rect 60747 -8667 60781 -8633
rect 61291 -8391 61325 -8357
rect 61046 -8457 61086 -8450
rect 61046 -8490 61059 -8457
rect 61059 -8490 61086 -8457
rect 61046 -8541 61086 -8540
rect 61046 -8575 61059 -8541
rect 61059 -8575 61086 -8541
rect 61046 -8580 61086 -8575
rect 61046 -8625 61086 -8620
rect 61046 -8659 61059 -8625
rect 61059 -8659 61086 -8625
rect 61046 -8660 61086 -8659
rect 61291 -8483 61325 -8449
rect 61291 -8575 61325 -8541
rect 61291 -8667 61325 -8633
rect 60747 -8759 60781 -8725
rect 60980 -8759 61015 -8725
rect 61053 -8759 61088 -8725
rect 61129 -8758 61164 -8724
rect 61291 -8759 61325 -8725
rect 60486 -8900 60526 -8860
rect 60626 -8900 60666 -8860
rect 60766 -8900 60806 -8860
rect 60906 -8900 60946 -8860
rect 59476 -9057 59483 -9023
rect 59483 -9057 59641 -9023
rect 59641 -9057 59646 -9023
rect 59476 -9060 59646 -9057
rect 59766 -9122 59806 -9120
rect 58926 -9336 58966 -9310
rect 59766 -9300 59772 -9122
rect 59772 -9300 59806 -9122
rect 59958 -9174 60334 -9140
rect 59874 -9228 59908 -9194
rect 60384 -9228 60418 -9194
rect 59958 -9282 60334 -9248
rect 57125 -9543 57159 -9509
rect 57217 -9543 57251 -9509
rect 57309 -9543 57343 -9509
rect 54081 -9778 54857 -9744
rect 53988 -9844 54022 -9806
rect 54916 -9844 54950 -9806
rect 54081 -9906 54857 -9872
rect 56020 -9808 56080 -9658
rect 58926 -9622 58930 -9336
rect 58930 -9622 58964 -9336
rect 58964 -9622 58966 -9336
rect 59656 -9336 59706 -9330
rect 59125 -9388 59501 -9354
rect 59560 -9442 59594 -9408
rect 59125 -9496 59501 -9462
rect 59032 -9550 59066 -9516
rect 59125 -9604 59501 -9570
rect 57156 -9690 57316 -9660
rect 57156 -9790 57186 -9690
rect 57186 -9790 57286 -9690
rect 57286 -9790 57316 -9690
rect 58926 -9700 58966 -9622
rect 59656 -9622 59662 -9336
rect 59662 -9622 59696 -9336
rect 59696 -9622 59706 -9336
rect 59866 -9362 60426 -9360
rect 59866 -9396 59868 -9362
rect 59868 -9396 60424 -9362
rect 60424 -9396 60426 -9362
rect 59866 -9400 60426 -9396
rect 59656 -9630 59706 -9622
rect 57156 -9820 57316 -9790
rect 54150 -10020 54840 -9988
rect 54150 -10108 54840 -10020
rect 55300 -9992 55476 -9958
rect 55526 -10036 55560 -10002
rect 55300 -10080 55476 -10046
rect 55320 -10160 55470 -10148
rect 55320 -10194 55470 -10160
rect 55320 -10208 55470 -10194
rect 20280 -11964 20340 -11930
rect 20390 -12008 20424 -11974
rect 20280 -12052 20340 -12018
rect 16440 -12143 25410 -12122
rect 16440 -12177 16535 -12143
rect 16535 -12177 16783 -12143
rect 16783 -12177 16941 -12143
rect 16941 -12177 17189 -12143
rect 17189 -12177 17347 -12143
rect 17347 -12177 17595 -12143
rect 17595 -12177 17753 -12143
rect 17753 -12177 18001 -12143
rect 18001 -12177 18159 -12143
rect 18159 -12177 18407 -12143
rect 18407 -12177 18565 -12143
rect 18565 -12177 18813 -12143
rect 18813 -12177 18971 -12143
rect 18971 -12177 19219 -12143
rect 19219 -12177 19377 -12143
rect 19377 -12177 19625 -12143
rect 19625 -12177 19783 -12143
rect 19783 -12177 20031 -12143
rect 20031 -12177 20189 -12143
rect 20189 -12177 20437 -12143
rect 20437 -12177 20595 -12143
rect 20595 -12177 20843 -12143
rect 20843 -12177 21001 -12143
rect 21001 -12177 21249 -12143
rect 21249 -12177 21407 -12143
rect 21407 -12177 21655 -12143
rect 21655 -12177 21813 -12143
rect 21813 -12177 22061 -12143
rect 22061 -12177 22219 -12143
rect 22219 -12177 22467 -12143
rect 22467 -12177 22625 -12143
rect 22625 -12177 22873 -12143
rect 22873 -12177 23031 -12143
rect 23031 -12177 23279 -12143
rect 23279 -12177 23437 -12143
rect 23437 -12177 23685 -12143
rect 23685 -12177 23843 -12143
rect 23843 -12177 24091 -12143
rect 24091 -12177 24249 -12143
rect 24249 -12177 24497 -12143
rect 24497 -12177 24655 -12143
rect 24655 -12177 24903 -12143
rect 24903 -12177 25061 -12143
rect 25061 -12177 25309 -12143
rect 25309 -12177 25410 -12143
rect 16440 -12182 25410 -12177
rect 16615 -12279 16703 -12245
rect 16553 -13105 16587 -12329
rect 16731 -13105 16765 -12329
rect 16615 -13189 16703 -13155
rect 17021 -12279 17109 -12245
rect 16959 -13105 16993 -12329
rect 17137 -13105 17171 -12329
rect 17021 -13189 17109 -13155
rect 17427 -12279 17515 -12245
rect 17365 -13105 17399 -12329
rect 17543 -13105 17577 -12329
rect 17427 -13189 17515 -13155
rect 17833 -12279 17921 -12245
rect 17771 -13105 17805 -12329
rect 17949 -13105 17983 -12329
rect 17833 -13189 17921 -13155
rect 18239 -12279 18327 -12245
rect 18177 -13105 18211 -12329
rect 18355 -13105 18389 -12329
rect 18239 -13189 18327 -13155
rect 18645 -12279 18733 -12245
rect 18583 -13105 18617 -12329
rect 18761 -13105 18795 -12329
rect 18645 -13189 18733 -13155
rect 19051 -12279 19139 -12245
rect 18989 -13105 19023 -12329
rect 19167 -13105 19201 -12329
rect 19051 -13189 19139 -13155
rect 19457 -12279 19545 -12245
rect 19395 -13105 19429 -12329
rect 19573 -13105 19607 -12329
rect 19457 -13189 19545 -13155
rect 19863 -12279 19951 -12245
rect 19801 -13105 19835 -12329
rect 19979 -13105 20013 -12329
rect 19863 -13189 19951 -13155
rect 20269 -12279 20357 -12245
rect 20207 -13105 20241 -12329
rect 20385 -13105 20419 -12329
rect 20269 -13189 20357 -13155
rect 20675 -12279 20763 -12245
rect 20613 -13105 20647 -12329
rect 20791 -13105 20825 -12329
rect 20675 -13189 20763 -13155
rect 21081 -12279 21169 -12245
rect 21019 -13105 21053 -12329
rect 21197 -13105 21231 -12329
rect 21081 -13189 21169 -13155
rect 21487 -12279 21575 -12245
rect 21425 -13105 21459 -12329
rect 21603 -13105 21637 -12329
rect 21487 -13189 21575 -13155
rect 21893 -12279 21981 -12245
rect 21831 -13105 21865 -12329
rect 22009 -13105 22043 -12329
rect 21893 -13189 21981 -13155
rect 22299 -12279 22387 -12245
rect 22237 -13105 22271 -12329
rect 22415 -13105 22449 -12329
rect 22299 -13189 22387 -13155
rect 22705 -12279 22793 -12245
rect 22643 -13105 22677 -12329
rect 22821 -13105 22855 -12329
rect 22705 -13189 22793 -13155
rect 23111 -12279 23199 -12245
rect 23049 -13105 23083 -12329
rect 23227 -13105 23261 -12329
rect 23111 -13189 23199 -13155
rect 23517 -12279 23605 -12245
rect 23455 -13105 23489 -12329
rect 23633 -13105 23667 -12329
rect 23517 -13189 23605 -13155
rect 23923 -12279 24011 -12245
rect 23861 -13105 23895 -12329
rect 24039 -13105 24073 -12329
rect 23923 -13189 24011 -13155
rect 24329 -12279 24417 -12245
rect 24267 -13105 24301 -12329
rect 24445 -13105 24479 -12329
rect 24329 -13189 24417 -13155
rect 24735 -12279 24823 -12245
rect 24673 -13105 24707 -12329
rect 24851 -13105 24885 -12329
rect 24735 -13189 24823 -13155
rect 25360 -12239 25410 -12182
rect 25141 -12279 25229 -12245
rect 25360 -12276 25371 -12239
rect 25079 -13105 25113 -12329
rect 25257 -13105 25291 -12329
rect 25362 -13149 25371 -12276
rect 25141 -13189 25229 -13155
rect 25361 -13195 25371 -13149
rect 25371 -13195 25405 -12239
rect 25405 -13195 25410 -12239
rect 54150 -12358 54850 -12308
rect 54150 -12392 54850 -12358
rect 54150 -12398 54850 -12392
rect 54091 -12506 54867 -12472
rect 53998 -12572 54032 -12534
rect 54926 -12572 54960 -12534
rect 54091 -12634 54867 -12600
rect 55960 -12698 56040 -12528
rect 53526 -12940 53614 -12906
rect 25361 -13219 25410 -13195
rect 25360 -13254 25410 -13219
rect 16448 -13257 25410 -13254
rect 16448 -13291 16535 -13257
rect 16535 -13291 16783 -13257
rect 16783 -13291 16941 -13257
rect 16941 -13291 17189 -13257
rect 17189 -13291 17347 -13257
rect 17347 -13291 17595 -13257
rect 17595 -13291 17753 -13257
rect 17753 -13291 18001 -13257
rect 18001 -13291 18159 -13257
rect 18159 -13291 18407 -13257
rect 18407 -13291 18565 -13257
rect 18565 -13291 18813 -13257
rect 18813 -13291 18971 -13257
rect 18971 -13291 19219 -13257
rect 19219 -13291 19377 -13257
rect 19377 -13291 19625 -13257
rect 19625 -13291 19783 -13257
rect 19783 -13291 20031 -13257
rect 20031 -13291 20189 -13257
rect 20189 -13291 20437 -13257
rect 20437 -13291 20595 -13257
rect 20595 -13291 20843 -13257
rect 20843 -13291 21001 -13257
rect 21001 -13291 21249 -13257
rect 21249 -13291 21407 -13257
rect 21407 -13291 21655 -13257
rect 21655 -13291 21813 -13257
rect 21813 -13291 22061 -13257
rect 22061 -13291 22219 -13257
rect 22219 -13291 22467 -13257
rect 22467 -13291 22625 -13257
rect 22625 -13291 22873 -13257
rect 22873 -13291 23031 -13257
rect 23031 -13291 23279 -13257
rect 23279 -13291 23437 -13257
rect 23437 -13291 23685 -13257
rect 23685 -13291 23843 -13257
rect 23843 -13291 24091 -13257
rect 24091 -13291 24249 -13257
rect 24249 -13291 24497 -13257
rect 24497 -13291 24655 -13257
rect 24655 -13291 24903 -13257
rect 24903 -13291 25061 -13257
rect 25061 -13291 25309 -13257
rect 25309 -13291 25410 -13257
rect 16448 -13302 25410 -13291
rect 16448 -13314 25400 -13302
rect 16420 -13386 34720 -13362
rect 16420 -13420 16532 -13386
rect 16532 -13420 34620 -13386
rect 34620 -13420 34720 -13386
rect 16420 -13422 34720 -13420
rect 16420 -13482 16490 -13422
rect 16420 -14696 16436 -13482
rect 16436 -14696 16470 -13482
rect 16470 -14696 16490 -13482
rect 34630 -13482 34720 -13422
rect 16584 -14646 16981 -13532
rect 34171 -14646 34568 -13532
rect 16420 -14742 16490 -14696
rect 34630 -14696 34682 -13482
rect 34682 -14696 34716 -13482
rect 34716 -14696 34720 -13482
rect 53330 -14318 53350 -12968
rect 53350 -14318 53384 -12968
rect 53384 -14318 53400 -12968
rect 53464 -13766 53498 -12990
rect 53642 -13766 53676 -12990
rect 57126 -12700 57356 -12670
rect 54091 -12862 54867 -12828
rect 53998 -12928 54032 -12890
rect 54926 -12928 54960 -12890
rect 54091 -12990 54867 -12956
rect 55334 -13002 55368 -12968
rect 55290 -13228 55324 -13052
rect 55378 -13228 55412 -13052
rect 55142 -13508 55494 -13474
rect 53942 -13612 54718 -13578
rect 53858 -13728 53892 -13640
rect 54768 -13728 54802 -13640
rect 53942 -13790 54718 -13756
rect 53526 -13850 53614 -13816
rect 55046 -13594 55080 -13560
rect 55556 -13594 55590 -13560
rect 55142 -13680 55494 -13646
rect 57126 -12770 57156 -12700
rect 57156 -12770 57316 -12700
rect 57316 -12770 57356 -12700
rect 57126 -12800 57356 -12770
rect 58926 -12829 58966 -12820
rect 55882 -12890 55970 -12856
rect 55820 -13716 55854 -12940
rect 55998 -13716 56032 -12940
rect 55882 -13800 55970 -13766
rect 57125 -12879 57159 -12845
rect 57217 -12879 57251 -12845
rect 57309 -12879 57343 -12845
rect 57118 -13157 57178 -13144
rect 57118 -13191 57133 -13157
rect 57133 -13191 57167 -13157
rect 57167 -13191 57178 -13157
rect 57118 -13194 57178 -13191
rect 58926 -13115 58930 -12829
rect 58930 -13115 58964 -12829
rect 58964 -13115 58966 -12829
rect 59125 -12881 59501 -12847
rect 59560 -12935 59594 -12901
rect 59125 -12989 59501 -12955
rect 59032 -13043 59066 -13009
rect 59125 -13097 59501 -13063
rect 58926 -13120 58966 -13115
rect 59656 -13115 59662 -12830
rect 59662 -13115 59696 -12830
rect 59656 -13120 59696 -13115
rect 57326 -13180 57366 -13140
rect 53526 -13958 53614 -13924
rect 55030 -13928 55110 -13848
rect 55740 -13868 55810 -13848
rect 55740 -13902 55802 -13868
rect 55802 -13902 55810 -13868
rect 55740 -13928 55810 -13902
rect 34630 -14742 34720 -14696
rect 16420 -14758 34724 -14742
rect 16420 -14792 16532 -14758
rect 16532 -14792 34620 -14758
rect 34620 -14792 34724 -14758
rect 16420 -14802 34724 -14792
rect 16420 -14854 16490 -14802
rect 16420 -16068 16436 -14854
rect 16436 -16068 16470 -14854
rect 16470 -16068 16490 -14854
rect 34630 -14854 34720 -14802
rect 16584 -16018 16981 -14904
rect 34171 -16018 34568 -14904
rect 16420 -16092 16490 -16068
rect 34630 -16068 34682 -14854
rect 34682 -16068 34716 -14854
rect 34716 -16068 34720 -14854
rect 53464 -14784 53498 -14008
rect 53642 -14784 53676 -14008
rect 53942 -14018 54718 -13984
rect 53858 -14134 53892 -14046
rect 54768 -14134 54802 -14046
rect 53942 -14196 54718 -14162
rect 55142 -14130 55494 -14096
rect 55046 -14216 55080 -14182
rect 55556 -14216 55590 -14182
rect 55142 -14302 55494 -14268
rect 53526 -14868 53614 -14834
rect 54081 -14822 54857 -14788
rect 53988 -14888 54022 -14850
rect 54916 -14888 54950 -14850
rect 54081 -14950 54857 -14916
rect 55280 -14724 55314 -14548
rect 55368 -14724 55402 -14548
rect 55324 -14808 55358 -14774
rect 56280 -13400 56350 -13318
rect 56280 -13948 56316 -13400
rect 56316 -13948 56350 -13400
rect 59866 -13094 59868 -13060
rect 59868 -13094 60424 -13060
rect 60424 -13094 60426 -13060
rect 59866 -13100 60426 -13094
rect 59766 -13156 59806 -13150
rect 59103 -13312 59137 -13278
rect 56492 -13440 56530 -13406
rect 55882 -14004 55970 -13970
rect 55820 -14830 55854 -14054
rect 55998 -14830 56032 -14054
rect 55882 -14914 55970 -14880
rect 56430 -14275 56464 -13499
rect 56558 -14275 56592 -13499
rect 56492 -14368 56530 -14334
rect 57125 -13423 57159 -13389
rect 57217 -13423 57251 -13389
rect 57309 -13423 57343 -13389
rect 57086 -13510 57376 -13480
rect 57086 -13580 57116 -13510
rect 57116 -13580 57346 -13510
rect 57346 -13580 57376 -13510
rect 57086 -13610 57376 -13580
rect 58926 -13846 58930 -13360
rect 58930 -13846 58964 -13360
rect 58964 -13846 58966 -13360
rect 59044 -13747 59078 -13371
rect 59162 -13747 59196 -13371
rect 59103 -13840 59137 -13806
rect 58926 -14002 58966 -13846
rect 59766 -13334 59772 -13156
rect 59772 -13334 59806 -13156
rect 59958 -13208 60334 -13174
rect 59874 -13262 59908 -13228
rect 60384 -13262 60418 -13228
rect 59958 -13316 60334 -13282
rect 59766 -13340 59806 -13334
rect 59476 -13396 59656 -13390
rect 59476 -13430 59484 -13396
rect 59484 -13430 59642 -13396
rect 59642 -13430 59656 -13396
rect 59386 -13492 59426 -13490
rect 59386 -13848 59388 -13492
rect 59388 -13848 59422 -13492
rect 59422 -13848 59426 -13492
rect 59546 -13532 59580 -13498
rect 59502 -13758 59536 -13582
rect 59590 -13758 59624 -13582
rect 59546 -13842 59580 -13808
rect 59386 -13850 59426 -13848
rect 59862 -13532 59896 -13498
rect 59818 -13758 59852 -13582
rect 59906 -13758 59940 -13582
rect 59862 -13842 59896 -13808
rect 61196 -13620 61366 -13600
rect 61196 -13660 61216 -13620
rect 61216 -13660 61336 -13620
rect 61336 -13660 61366 -13620
rect 61196 -13680 61366 -13660
rect 57056 -14170 57416 -14140
rect 57056 -14250 57096 -14170
rect 57096 -14250 57376 -14170
rect 57376 -14250 57416 -14170
rect 57056 -14280 57416 -14250
rect 57125 -14399 57159 -14365
rect 57217 -14399 57251 -14365
rect 57309 -14399 57343 -14365
rect 58926 -14490 58930 -14002
rect 58930 -14490 58964 -14002
rect 58964 -14490 58966 -14002
rect 60127 -13791 60161 -13757
rect 60366 -13765 60406 -13760
rect 60366 -13799 60393 -13765
rect 60393 -13799 60406 -13765
rect 60366 -13800 60406 -13799
rect 60127 -13883 60161 -13849
rect 59103 -14042 59137 -14008
rect 59044 -14477 59078 -14101
rect 57118 -14597 57168 -14594
rect 57118 -14631 57133 -14597
rect 57133 -14631 57167 -14597
rect 57167 -14631 57168 -14597
rect 57118 -14644 57168 -14631
rect 57326 -14610 57376 -14570
rect 59162 -14477 59196 -14101
rect 59103 -14570 59137 -14536
rect 59386 -14005 59426 -14000
rect 59386 -14361 59387 -14005
rect 59387 -14361 59421 -14005
rect 59421 -14361 59426 -14005
rect 59545 -14045 59579 -14011
rect 59501 -14271 59535 -14095
rect 59589 -14271 59623 -14095
rect 59545 -14355 59579 -14321
rect 59386 -14370 59426 -14361
rect 59476 -14423 59646 -14420
rect 59861 -14045 59895 -14011
rect 59817 -14271 59851 -14095
rect 59905 -14271 59939 -14095
rect 59861 -14355 59895 -14321
rect 60127 -13975 60161 -13941
rect 60127 -14067 60161 -14033
rect 60671 -13791 60705 -13757
rect 60366 -13857 60406 -13850
rect 60366 -13890 60393 -13857
rect 60393 -13890 60406 -13857
rect 60366 -13941 60406 -13940
rect 60366 -13975 60393 -13941
rect 60393 -13975 60406 -13941
rect 60366 -13980 60406 -13975
rect 60366 -14025 60406 -14020
rect 60366 -14059 60393 -14025
rect 60393 -14059 60406 -14025
rect 60366 -14060 60406 -14059
rect 60671 -13883 60705 -13849
rect 60671 -13975 60705 -13941
rect 60671 -14067 60705 -14033
rect 60127 -14159 60161 -14125
rect 60297 -14159 60331 -14125
rect 60369 -14159 60405 -14125
rect 60449 -14159 60484 -14125
rect 60671 -14159 60705 -14125
rect 60747 -13791 60781 -13757
rect 61046 -13765 61086 -13760
rect 61046 -13799 61059 -13765
rect 61059 -13799 61086 -13765
rect 61046 -13800 61086 -13799
rect 60747 -13883 60781 -13849
rect 60747 -13975 60781 -13941
rect 60747 -14067 60781 -14033
rect 61291 -13791 61325 -13757
rect 61046 -13857 61086 -13850
rect 61046 -13890 61059 -13857
rect 61059 -13890 61086 -13857
rect 61046 -13941 61086 -13940
rect 61046 -13975 61059 -13941
rect 61059 -13975 61086 -13941
rect 61046 -13980 61086 -13975
rect 61046 -14025 61086 -14020
rect 61046 -14059 61059 -14025
rect 61059 -14059 61086 -14025
rect 61046 -14060 61086 -14059
rect 61291 -13883 61325 -13849
rect 61291 -13975 61325 -13941
rect 61291 -14067 61325 -14033
rect 60747 -14159 60781 -14125
rect 60980 -14159 61015 -14125
rect 61053 -14159 61088 -14125
rect 61129 -14158 61164 -14124
rect 61291 -14159 61325 -14125
rect 60486 -14300 60526 -14260
rect 60626 -14300 60666 -14260
rect 60766 -14300 60806 -14260
rect 60906 -14300 60946 -14260
rect 59476 -14457 59483 -14423
rect 59483 -14457 59641 -14423
rect 59641 -14457 59646 -14423
rect 59476 -14460 59646 -14457
rect 59766 -14522 59806 -14520
rect 58926 -14736 58966 -14710
rect 59766 -14700 59772 -14522
rect 59772 -14700 59806 -14522
rect 59958 -14574 60334 -14540
rect 59874 -14628 59908 -14594
rect 60384 -14628 60418 -14594
rect 59958 -14682 60334 -14648
rect 57125 -14943 57159 -14909
rect 57217 -14943 57251 -14909
rect 57309 -14943 57343 -14909
rect 54081 -15178 54857 -15144
rect 53988 -15244 54022 -15206
rect 54916 -15244 54950 -15206
rect 54081 -15306 54857 -15272
rect 56020 -15208 56080 -15058
rect 58926 -15022 58930 -14736
rect 58930 -15022 58964 -14736
rect 58964 -15022 58966 -14736
rect 59656 -14736 59706 -14730
rect 59125 -14788 59501 -14754
rect 59560 -14842 59594 -14808
rect 59125 -14896 59501 -14862
rect 59032 -14950 59066 -14916
rect 59125 -15004 59501 -14970
rect 57156 -15090 57316 -15060
rect 57156 -15190 57186 -15090
rect 57186 -15190 57286 -15090
rect 57286 -15190 57316 -15090
rect 58926 -15100 58966 -15022
rect 59656 -15022 59662 -14736
rect 59662 -15022 59696 -14736
rect 59696 -15022 59706 -14736
rect 59866 -14762 60426 -14760
rect 59866 -14796 59868 -14762
rect 59868 -14796 60424 -14762
rect 60424 -14796 60426 -14762
rect 59866 -14800 60426 -14796
rect 59656 -15030 59706 -15022
rect 57156 -15220 57316 -15190
rect 54150 -15420 54840 -15388
rect 54150 -15508 54840 -15420
rect 55300 -15392 55476 -15358
rect 55526 -15436 55560 -15402
rect 55300 -15480 55476 -15446
rect 55320 -15560 55470 -15548
rect 55320 -15594 55470 -15560
rect 55320 -15608 55470 -15594
rect 34630 -16092 34720 -16068
rect 16420 -16130 34730 -16092
rect 16420 -16164 16532 -16130
rect 16532 -16164 34620 -16130
rect 34620 -16164 34730 -16130
rect 16420 -16182 34730 -16164
rect 54150 -17758 54850 -17708
rect 54150 -17792 54850 -17758
rect 54150 -17798 54850 -17792
rect 54091 -17906 54867 -17872
rect 53998 -17972 54032 -17934
rect 54926 -17972 54960 -17934
rect 54091 -18034 54867 -18000
rect 55960 -18098 56040 -17928
rect 53526 -18340 53614 -18306
rect 53330 -19718 53350 -18368
rect 53350 -19718 53384 -18368
rect 53384 -19718 53400 -18368
rect 53464 -19166 53498 -18390
rect 53642 -19166 53676 -18390
rect 57126 -18100 57356 -18070
rect 54091 -18262 54867 -18228
rect 53998 -18328 54032 -18290
rect 54926 -18328 54960 -18290
rect 54091 -18390 54867 -18356
rect 55334 -18402 55368 -18368
rect 55290 -18628 55324 -18452
rect 55378 -18628 55412 -18452
rect 55142 -18908 55494 -18874
rect 53942 -19012 54718 -18978
rect 53858 -19128 53892 -19040
rect 54768 -19128 54802 -19040
rect 53942 -19190 54718 -19156
rect 53526 -19250 53614 -19216
rect 55046 -18994 55080 -18960
rect 55556 -18994 55590 -18960
rect 55142 -19080 55494 -19046
rect 57126 -18170 57156 -18100
rect 57156 -18170 57316 -18100
rect 57316 -18170 57356 -18100
rect 57126 -18200 57356 -18170
rect 58926 -18229 58966 -18220
rect 55882 -18290 55970 -18256
rect 55820 -19116 55854 -18340
rect 55998 -19116 56032 -18340
rect 55882 -19200 55970 -19166
rect 57125 -18279 57159 -18245
rect 57217 -18279 57251 -18245
rect 57309 -18279 57343 -18245
rect 57118 -18557 57178 -18544
rect 57118 -18591 57133 -18557
rect 57133 -18591 57167 -18557
rect 57167 -18591 57178 -18557
rect 57118 -18594 57178 -18591
rect 58926 -18515 58930 -18229
rect 58930 -18515 58964 -18229
rect 58964 -18515 58966 -18229
rect 59125 -18281 59501 -18247
rect 59560 -18335 59594 -18301
rect 59125 -18389 59501 -18355
rect 59032 -18443 59066 -18409
rect 59125 -18497 59501 -18463
rect 58926 -18520 58966 -18515
rect 59656 -18515 59662 -18230
rect 59662 -18515 59696 -18230
rect 59656 -18520 59696 -18515
rect 57326 -18580 57366 -18540
rect 53526 -19358 53614 -19324
rect 55030 -19328 55110 -19248
rect 55740 -19268 55810 -19248
rect 55740 -19302 55802 -19268
rect 55802 -19302 55810 -19268
rect 55740 -19328 55810 -19302
rect 53464 -20184 53498 -19408
rect 53642 -20184 53676 -19408
rect 53942 -19418 54718 -19384
rect 53858 -19534 53892 -19446
rect 54768 -19534 54802 -19446
rect 53942 -19596 54718 -19562
rect 55142 -19530 55494 -19496
rect 55046 -19616 55080 -19582
rect 55556 -19616 55590 -19582
rect 55142 -19702 55494 -19668
rect 53526 -20268 53614 -20234
rect 54081 -20222 54857 -20188
rect 53988 -20288 54022 -20250
rect 54916 -20288 54950 -20250
rect 54081 -20350 54857 -20316
rect 55280 -20124 55314 -19948
rect 55368 -20124 55402 -19948
rect 55324 -20208 55358 -20174
rect 56280 -18800 56350 -18718
rect 56280 -19348 56316 -18800
rect 56316 -19348 56350 -18800
rect 59866 -18494 59868 -18460
rect 59868 -18494 60424 -18460
rect 60424 -18494 60426 -18460
rect 59866 -18500 60426 -18494
rect 59766 -18556 59806 -18550
rect 59103 -18712 59137 -18678
rect 56492 -18840 56530 -18806
rect 55882 -19404 55970 -19370
rect 55820 -20230 55854 -19454
rect 55998 -20230 56032 -19454
rect 55882 -20314 55970 -20280
rect 56430 -19675 56464 -18899
rect 56558 -19675 56592 -18899
rect 56492 -19768 56530 -19734
rect 57125 -18823 57159 -18789
rect 57217 -18823 57251 -18789
rect 57309 -18823 57343 -18789
rect 57086 -18910 57376 -18880
rect 57086 -18980 57116 -18910
rect 57116 -18980 57346 -18910
rect 57346 -18980 57376 -18910
rect 57086 -19010 57376 -18980
rect 58926 -19246 58930 -18760
rect 58930 -19246 58964 -18760
rect 58964 -19246 58966 -18760
rect 59044 -19147 59078 -18771
rect 59162 -19147 59196 -18771
rect 59103 -19240 59137 -19206
rect 58926 -19402 58966 -19246
rect 59766 -18734 59772 -18556
rect 59772 -18734 59806 -18556
rect 59958 -18608 60334 -18574
rect 59874 -18662 59908 -18628
rect 60384 -18662 60418 -18628
rect 59958 -18716 60334 -18682
rect 59766 -18740 59806 -18734
rect 59476 -18796 59656 -18790
rect 59476 -18830 59484 -18796
rect 59484 -18830 59642 -18796
rect 59642 -18830 59656 -18796
rect 59386 -18892 59426 -18890
rect 59386 -19248 59388 -18892
rect 59388 -19248 59422 -18892
rect 59422 -19248 59426 -18892
rect 59546 -18932 59580 -18898
rect 59502 -19158 59536 -18982
rect 59590 -19158 59624 -18982
rect 59546 -19242 59580 -19208
rect 59386 -19250 59426 -19248
rect 59862 -18932 59896 -18898
rect 59818 -19158 59852 -18982
rect 59906 -19158 59940 -18982
rect 59862 -19242 59896 -19208
rect 61196 -19020 61366 -19000
rect 61196 -19060 61216 -19020
rect 61216 -19060 61336 -19020
rect 61336 -19060 61366 -19020
rect 61196 -19080 61366 -19060
rect 57056 -19570 57416 -19540
rect 57056 -19650 57096 -19570
rect 57096 -19650 57376 -19570
rect 57376 -19650 57416 -19570
rect 57056 -19680 57416 -19650
rect 57125 -19799 57159 -19765
rect 57217 -19799 57251 -19765
rect 57309 -19799 57343 -19765
rect 58926 -19890 58930 -19402
rect 58930 -19890 58964 -19402
rect 58964 -19890 58966 -19402
rect 60127 -19191 60161 -19157
rect 60366 -19165 60406 -19160
rect 60366 -19199 60393 -19165
rect 60393 -19199 60406 -19165
rect 60366 -19200 60406 -19199
rect 60127 -19283 60161 -19249
rect 59103 -19442 59137 -19408
rect 59044 -19877 59078 -19501
rect 57118 -19997 57168 -19994
rect 57118 -20031 57133 -19997
rect 57133 -20031 57167 -19997
rect 57167 -20031 57168 -19997
rect 57118 -20044 57168 -20031
rect 57326 -20010 57376 -19970
rect 59162 -19877 59196 -19501
rect 59103 -19970 59137 -19936
rect 59386 -19405 59426 -19400
rect 59386 -19761 59387 -19405
rect 59387 -19761 59421 -19405
rect 59421 -19761 59426 -19405
rect 59545 -19445 59579 -19411
rect 59501 -19671 59535 -19495
rect 59589 -19671 59623 -19495
rect 59545 -19755 59579 -19721
rect 59386 -19770 59426 -19761
rect 59476 -19823 59646 -19820
rect 59861 -19445 59895 -19411
rect 59817 -19671 59851 -19495
rect 59905 -19671 59939 -19495
rect 59861 -19755 59895 -19721
rect 60127 -19375 60161 -19341
rect 60127 -19467 60161 -19433
rect 60671 -19191 60705 -19157
rect 60366 -19257 60406 -19250
rect 60366 -19290 60393 -19257
rect 60393 -19290 60406 -19257
rect 60366 -19341 60406 -19340
rect 60366 -19375 60393 -19341
rect 60393 -19375 60406 -19341
rect 60366 -19380 60406 -19375
rect 60366 -19425 60406 -19420
rect 60366 -19459 60393 -19425
rect 60393 -19459 60406 -19425
rect 60366 -19460 60406 -19459
rect 60671 -19283 60705 -19249
rect 60671 -19375 60705 -19341
rect 60671 -19467 60705 -19433
rect 60127 -19559 60161 -19525
rect 60297 -19559 60331 -19525
rect 60369 -19559 60405 -19525
rect 60449 -19559 60484 -19525
rect 60671 -19559 60705 -19525
rect 60747 -19191 60781 -19157
rect 61046 -19165 61086 -19160
rect 61046 -19199 61059 -19165
rect 61059 -19199 61086 -19165
rect 61046 -19200 61086 -19199
rect 60747 -19283 60781 -19249
rect 60747 -19375 60781 -19341
rect 60747 -19467 60781 -19433
rect 61291 -19191 61325 -19157
rect 61046 -19257 61086 -19250
rect 61046 -19290 61059 -19257
rect 61059 -19290 61086 -19257
rect 61046 -19341 61086 -19340
rect 61046 -19375 61059 -19341
rect 61059 -19375 61086 -19341
rect 61046 -19380 61086 -19375
rect 61046 -19425 61086 -19420
rect 61046 -19459 61059 -19425
rect 61059 -19459 61086 -19425
rect 61046 -19460 61086 -19459
rect 61291 -19283 61325 -19249
rect 61291 -19375 61325 -19341
rect 61291 -19467 61325 -19433
rect 60747 -19559 60781 -19525
rect 60980 -19559 61015 -19525
rect 61053 -19559 61088 -19525
rect 61129 -19558 61164 -19524
rect 61291 -19559 61325 -19525
rect 60486 -19700 60526 -19660
rect 60626 -19700 60666 -19660
rect 60766 -19700 60806 -19660
rect 60906 -19700 60946 -19660
rect 59476 -19857 59483 -19823
rect 59483 -19857 59641 -19823
rect 59641 -19857 59646 -19823
rect 59476 -19860 59646 -19857
rect 59766 -19922 59806 -19920
rect 58926 -20136 58966 -20110
rect 59766 -20100 59772 -19922
rect 59772 -20100 59806 -19922
rect 59958 -19974 60334 -19940
rect 59874 -20028 59908 -19994
rect 60384 -20028 60418 -19994
rect 59958 -20082 60334 -20048
rect 57125 -20343 57159 -20309
rect 57217 -20343 57251 -20309
rect 57309 -20343 57343 -20309
rect 54081 -20578 54857 -20544
rect 53988 -20644 54022 -20606
rect 54916 -20644 54950 -20606
rect 54081 -20706 54857 -20672
rect 56020 -20608 56080 -20458
rect 58926 -20422 58930 -20136
rect 58930 -20422 58964 -20136
rect 58964 -20422 58966 -20136
rect 59656 -20136 59706 -20130
rect 59125 -20188 59501 -20154
rect 59560 -20242 59594 -20208
rect 59125 -20296 59501 -20262
rect 59032 -20350 59066 -20316
rect 59125 -20404 59501 -20370
rect 57156 -20490 57316 -20460
rect 57156 -20590 57186 -20490
rect 57186 -20590 57286 -20490
rect 57286 -20590 57316 -20490
rect 58926 -20500 58966 -20422
rect 59656 -20422 59662 -20136
rect 59662 -20422 59696 -20136
rect 59696 -20422 59706 -20136
rect 59866 -20162 60426 -20160
rect 59866 -20196 59868 -20162
rect 59868 -20196 60424 -20162
rect 60424 -20196 60426 -20162
rect 59866 -20200 60426 -20196
rect 59656 -20430 59706 -20422
rect 57156 -20620 57316 -20590
rect 54150 -20820 54840 -20788
rect 54150 -20908 54840 -20820
rect 55300 -20792 55476 -20758
rect 55526 -20836 55560 -20802
rect 55300 -20880 55476 -20846
rect 55320 -20960 55470 -20948
rect 55320 -20994 55470 -20960
rect 55320 -21008 55470 -20994
rect 54150 -23158 54850 -23108
rect 54150 -23192 54850 -23158
rect 54150 -23198 54850 -23192
rect 54091 -23306 54867 -23272
rect 53998 -23372 54032 -23334
rect 54926 -23372 54960 -23334
rect 54091 -23434 54867 -23400
rect 55960 -23498 56040 -23328
rect 53526 -23740 53614 -23706
rect 53330 -25118 53350 -23768
rect 53350 -25118 53384 -23768
rect 53384 -25118 53400 -23768
rect 53464 -24566 53498 -23790
rect 53642 -24566 53676 -23790
rect 57126 -23500 57356 -23470
rect 54091 -23662 54867 -23628
rect 53998 -23728 54032 -23690
rect 54926 -23728 54960 -23690
rect 54091 -23790 54867 -23756
rect 55334 -23802 55368 -23768
rect 55290 -24028 55324 -23852
rect 55378 -24028 55412 -23852
rect 55142 -24308 55494 -24274
rect 53942 -24412 54718 -24378
rect 53858 -24528 53892 -24440
rect 54768 -24528 54802 -24440
rect 53942 -24590 54718 -24556
rect 53526 -24650 53614 -24616
rect 55046 -24394 55080 -24360
rect 55556 -24394 55590 -24360
rect 55142 -24480 55494 -24446
rect 57126 -23570 57156 -23500
rect 57156 -23570 57316 -23500
rect 57316 -23570 57356 -23500
rect 57126 -23600 57356 -23570
rect 58926 -23629 58966 -23620
rect 55882 -23690 55970 -23656
rect 55820 -24516 55854 -23740
rect 55998 -24516 56032 -23740
rect 55882 -24600 55970 -24566
rect 57125 -23679 57159 -23645
rect 57217 -23679 57251 -23645
rect 57309 -23679 57343 -23645
rect 57118 -23957 57178 -23944
rect 57118 -23991 57133 -23957
rect 57133 -23991 57167 -23957
rect 57167 -23991 57178 -23957
rect 57118 -23994 57178 -23991
rect 58926 -23915 58930 -23629
rect 58930 -23915 58964 -23629
rect 58964 -23915 58966 -23629
rect 59125 -23681 59501 -23647
rect 59560 -23735 59594 -23701
rect 59125 -23789 59501 -23755
rect 59032 -23843 59066 -23809
rect 59125 -23897 59501 -23863
rect 58926 -23920 58966 -23915
rect 59656 -23915 59662 -23630
rect 59662 -23915 59696 -23630
rect 59656 -23920 59696 -23915
rect 57326 -23980 57366 -23940
rect 53526 -24758 53614 -24724
rect 55030 -24728 55110 -24648
rect 55740 -24668 55810 -24648
rect 55740 -24702 55802 -24668
rect 55802 -24702 55810 -24668
rect 55740 -24728 55810 -24702
rect 53464 -25584 53498 -24808
rect 53642 -25584 53676 -24808
rect 53942 -24818 54718 -24784
rect 53858 -24934 53892 -24846
rect 54768 -24934 54802 -24846
rect 53942 -24996 54718 -24962
rect 55142 -24930 55494 -24896
rect 55046 -25016 55080 -24982
rect 55556 -25016 55590 -24982
rect 55142 -25102 55494 -25068
rect 53526 -25668 53614 -25634
rect 54081 -25622 54857 -25588
rect 53988 -25688 54022 -25650
rect 54916 -25688 54950 -25650
rect 54081 -25750 54857 -25716
rect 55280 -25524 55314 -25348
rect 55368 -25524 55402 -25348
rect 55324 -25608 55358 -25574
rect 56280 -24200 56350 -24118
rect 56280 -24748 56316 -24200
rect 56316 -24748 56350 -24200
rect 59866 -23894 59868 -23860
rect 59868 -23894 60424 -23860
rect 60424 -23894 60426 -23860
rect 59866 -23900 60426 -23894
rect 59766 -23956 59806 -23950
rect 59103 -24112 59137 -24078
rect 56492 -24240 56530 -24206
rect 55882 -24804 55970 -24770
rect 55820 -25630 55854 -24854
rect 55998 -25630 56032 -24854
rect 55882 -25714 55970 -25680
rect 56430 -25075 56464 -24299
rect 56558 -25075 56592 -24299
rect 56492 -25168 56530 -25134
rect 57125 -24223 57159 -24189
rect 57217 -24223 57251 -24189
rect 57309 -24223 57343 -24189
rect 57086 -24310 57376 -24280
rect 57086 -24380 57116 -24310
rect 57116 -24380 57346 -24310
rect 57346 -24380 57376 -24310
rect 57086 -24410 57376 -24380
rect 58926 -24646 58930 -24160
rect 58930 -24646 58964 -24160
rect 58964 -24646 58966 -24160
rect 59044 -24547 59078 -24171
rect 59162 -24547 59196 -24171
rect 59103 -24640 59137 -24606
rect 58926 -24802 58966 -24646
rect 59766 -24134 59772 -23956
rect 59772 -24134 59806 -23956
rect 59958 -24008 60334 -23974
rect 59874 -24062 59908 -24028
rect 60384 -24062 60418 -24028
rect 59958 -24116 60334 -24082
rect 59766 -24140 59806 -24134
rect 59476 -24196 59656 -24190
rect 59476 -24230 59484 -24196
rect 59484 -24230 59642 -24196
rect 59642 -24230 59656 -24196
rect 59386 -24292 59426 -24290
rect 59386 -24648 59388 -24292
rect 59388 -24648 59422 -24292
rect 59422 -24648 59426 -24292
rect 59546 -24332 59580 -24298
rect 59502 -24558 59536 -24382
rect 59590 -24558 59624 -24382
rect 59546 -24642 59580 -24608
rect 59386 -24650 59426 -24648
rect 59862 -24332 59896 -24298
rect 59818 -24558 59852 -24382
rect 59906 -24558 59940 -24382
rect 59862 -24642 59896 -24608
rect 61196 -24420 61366 -24400
rect 61196 -24460 61216 -24420
rect 61216 -24460 61336 -24420
rect 61336 -24460 61366 -24420
rect 61196 -24480 61366 -24460
rect 57056 -24970 57416 -24940
rect 57056 -25050 57096 -24970
rect 57096 -25050 57376 -24970
rect 57376 -25050 57416 -24970
rect 57056 -25080 57416 -25050
rect 57125 -25199 57159 -25165
rect 57217 -25199 57251 -25165
rect 57309 -25199 57343 -25165
rect 58926 -25290 58930 -24802
rect 58930 -25290 58964 -24802
rect 58964 -25290 58966 -24802
rect 60127 -24591 60161 -24557
rect 60366 -24565 60406 -24560
rect 60366 -24599 60393 -24565
rect 60393 -24599 60406 -24565
rect 60366 -24600 60406 -24599
rect 60127 -24683 60161 -24649
rect 59103 -24842 59137 -24808
rect 59044 -25277 59078 -24901
rect 57118 -25397 57168 -25394
rect 57118 -25431 57133 -25397
rect 57133 -25431 57167 -25397
rect 57167 -25431 57168 -25397
rect 57118 -25444 57168 -25431
rect 57326 -25410 57376 -25370
rect 59162 -25277 59196 -24901
rect 59103 -25370 59137 -25336
rect 59386 -24805 59426 -24800
rect 59386 -25161 59387 -24805
rect 59387 -25161 59421 -24805
rect 59421 -25161 59426 -24805
rect 59545 -24845 59579 -24811
rect 59501 -25071 59535 -24895
rect 59589 -25071 59623 -24895
rect 59545 -25155 59579 -25121
rect 59386 -25170 59426 -25161
rect 59476 -25223 59646 -25220
rect 59861 -24845 59895 -24811
rect 59817 -25071 59851 -24895
rect 59905 -25071 59939 -24895
rect 59861 -25155 59895 -25121
rect 60127 -24775 60161 -24741
rect 60127 -24867 60161 -24833
rect 60671 -24591 60705 -24557
rect 60366 -24657 60406 -24650
rect 60366 -24690 60393 -24657
rect 60393 -24690 60406 -24657
rect 60366 -24741 60406 -24740
rect 60366 -24775 60393 -24741
rect 60393 -24775 60406 -24741
rect 60366 -24780 60406 -24775
rect 60366 -24825 60406 -24820
rect 60366 -24859 60393 -24825
rect 60393 -24859 60406 -24825
rect 60366 -24860 60406 -24859
rect 60671 -24683 60705 -24649
rect 60671 -24775 60705 -24741
rect 60671 -24867 60705 -24833
rect 60127 -24959 60161 -24925
rect 60297 -24959 60331 -24925
rect 60369 -24959 60405 -24925
rect 60449 -24959 60484 -24925
rect 60671 -24959 60705 -24925
rect 60747 -24591 60781 -24557
rect 61046 -24565 61086 -24560
rect 61046 -24599 61059 -24565
rect 61059 -24599 61086 -24565
rect 61046 -24600 61086 -24599
rect 60747 -24683 60781 -24649
rect 60747 -24775 60781 -24741
rect 60747 -24867 60781 -24833
rect 61291 -24591 61325 -24557
rect 61046 -24657 61086 -24650
rect 61046 -24690 61059 -24657
rect 61059 -24690 61086 -24657
rect 61046 -24741 61086 -24740
rect 61046 -24775 61059 -24741
rect 61059 -24775 61086 -24741
rect 61046 -24780 61086 -24775
rect 61046 -24825 61086 -24820
rect 61046 -24859 61059 -24825
rect 61059 -24859 61086 -24825
rect 61046 -24860 61086 -24859
rect 61291 -24683 61325 -24649
rect 61291 -24775 61325 -24741
rect 61291 -24867 61325 -24833
rect 60747 -24959 60781 -24925
rect 60980 -24959 61015 -24925
rect 61053 -24959 61088 -24925
rect 61129 -24958 61164 -24924
rect 61291 -24959 61325 -24925
rect 60486 -25100 60526 -25060
rect 60626 -25100 60666 -25060
rect 60766 -25100 60806 -25060
rect 60906 -25100 60946 -25060
rect 59476 -25257 59483 -25223
rect 59483 -25257 59641 -25223
rect 59641 -25257 59646 -25223
rect 59476 -25260 59646 -25257
rect 59766 -25322 59806 -25320
rect 58926 -25536 58966 -25510
rect 59766 -25500 59772 -25322
rect 59772 -25500 59806 -25322
rect 59958 -25374 60334 -25340
rect 59874 -25428 59908 -25394
rect 60384 -25428 60418 -25394
rect 59958 -25482 60334 -25448
rect 57125 -25743 57159 -25709
rect 57217 -25743 57251 -25709
rect 57309 -25743 57343 -25709
rect 54081 -25978 54857 -25944
rect 53988 -26044 54022 -26006
rect 54916 -26044 54950 -26006
rect 54081 -26106 54857 -26072
rect 56020 -26008 56080 -25858
rect 58926 -25822 58930 -25536
rect 58930 -25822 58964 -25536
rect 58964 -25822 58966 -25536
rect 59656 -25536 59706 -25530
rect 59125 -25588 59501 -25554
rect 59560 -25642 59594 -25608
rect 59125 -25696 59501 -25662
rect 59032 -25750 59066 -25716
rect 59125 -25804 59501 -25770
rect 57156 -25890 57316 -25860
rect 57156 -25990 57186 -25890
rect 57186 -25990 57286 -25890
rect 57286 -25990 57316 -25890
rect 58926 -25900 58966 -25822
rect 59656 -25822 59662 -25536
rect 59662 -25822 59696 -25536
rect 59696 -25822 59706 -25536
rect 59866 -25562 60426 -25560
rect 59866 -25596 59868 -25562
rect 59868 -25596 60424 -25562
rect 60424 -25596 60426 -25562
rect 59866 -25600 60426 -25596
rect 59656 -25830 59706 -25822
rect 57156 -26020 57316 -25990
rect 54150 -26220 54840 -26188
rect 54150 -26308 54840 -26220
rect 55300 -26192 55476 -26158
rect 55526 -26236 55560 -26202
rect 55300 -26280 55476 -26246
rect 55320 -26360 55470 -26348
rect 55320 -26394 55470 -26360
rect 55320 -26408 55470 -26394
rect 54150 -28558 54850 -28508
rect 54150 -28592 54850 -28558
rect 54150 -28598 54850 -28592
rect 54091 -28706 54867 -28672
rect 53998 -28772 54032 -28734
rect 54926 -28772 54960 -28734
rect 54091 -28834 54867 -28800
rect 55960 -28898 56040 -28728
rect 53526 -29140 53614 -29106
rect 53330 -30518 53350 -29168
rect 53350 -30518 53384 -29168
rect 53384 -30518 53400 -29168
rect 53464 -29966 53498 -29190
rect 53642 -29966 53676 -29190
rect 57126 -28900 57356 -28870
rect 54091 -29062 54867 -29028
rect 53998 -29128 54032 -29090
rect 54926 -29128 54960 -29090
rect 54091 -29190 54867 -29156
rect 55334 -29202 55368 -29168
rect 55290 -29428 55324 -29252
rect 55378 -29428 55412 -29252
rect 55142 -29708 55494 -29674
rect 53942 -29812 54718 -29778
rect 53858 -29928 53892 -29840
rect 54768 -29928 54802 -29840
rect 53942 -29990 54718 -29956
rect 53526 -30050 53614 -30016
rect 55046 -29794 55080 -29760
rect 55556 -29794 55590 -29760
rect 55142 -29880 55494 -29846
rect 57126 -28970 57156 -28900
rect 57156 -28970 57316 -28900
rect 57316 -28970 57356 -28900
rect 57126 -29000 57356 -28970
rect 58926 -29029 58966 -29020
rect 55882 -29090 55970 -29056
rect 55820 -29916 55854 -29140
rect 55998 -29916 56032 -29140
rect 55882 -30000 55970 -29966
rect 57125 -29079 57159 -29045
rect 57217 -29079 57251 -29045
rect 57309 -29079 57343 -29045
rect 57118 -29357 57178 -29344
rect 57118 -29391 57133 -29357
rect 57133 -29391 57167 -29357
rect 57167 -29391 57178 -29357
rect 57118 -29394 57178 -29391
rect 58926 -29315 58930 -29029
rect 58930 -29315 58964 -29029
rect 58964 -29315 58966 -29029
rect 59125 -29081 59501 -29047
rect 59560 -29135 59594 -29101
rect 59125 -29189 59501 -29155
rect 59032 -29243 59066 -29209
rect 59125 -29297 59501 -29263
rect 58926 -29320 58966 -29315
rect 59656 -29315 59662 -29030
rect 59662 -29315 59696 -29030
rect 59656 -29320 59696 -29315
rect 57326 -29380 57366 -29340
rect 53526 -30158 53614 -30124
rect 55030 -30128 55110 -30048
rect 55740 -30068 55810 -30048
rect 55740 -30102 55802 -30068
rect 55802 -30102 55810 -30068
rect 55740 -30128 55810 -30102
rect 25700 -31094 25780 -31020
rect 25700 -32530 25738 -31094
rect 25738 -32530 25772 -31094
rect 25772 -32530 25780 -31094
rect 25884 -31543 26998 -31146
rect 27126 -31543 28240 -31146
rect 28368 -31543 29482 -31146
rect 29610 -31543 30724 -31146
rect 30852 -31543 31966 -31146
rect 32094 -31543 33208 -31146
rect 33336 -31543 34450 -31146
rect 34578 -31543 35692 -31146
rect 25884 -32478 26998 -32081
rect 27126 -32478 28240 -32081
rect 28368 -32478 29482 -32081
rect 29610 -32478 30724 -32081
rect 30852 -32478 31966 -32081
rect 32094 -32478 33208 -32081
rect 33336 -32478 34450 -32081
rect 34578 -32478 35692 -32081
rect 25700 -32692 25780 -32530
rect 53464 -30984 53498 -30208
rect 53642 -30984 53676 -30208
rect 53942 -30218 54718 -30184
rect 53858 -30334 53892 -30246
rect 54768 -30334 54802 -30246
rect 53942 -30396 54718 -30362
rect 55142 -30330 55494 -30296
rect 55046 -30416 55080 -30382
rect 55556 -30416 55590 -30382
rect 55142 -30502 55494 -30468
rect 53526 -31068 53614 -31034
rect 54081 -31022 54857 -30988
rect 53988 -31088 54022 -31050
rect 54916 -31088 54950 -31050
rect 54081 -31150 54857 -31116
rect 55280 -30924 55314 -30748
rect 55368 -30924 55402 -30748
rect 55324 -31008 55358 -30974
rect 56280 -29600 56350 -29518
rect 56280 -30148 56316 -29600
rect 56316 -30148 56350 -29600
rect 59866 -29294 59868 -29260
rect 59868 -29294 60424 -29260
rect 60424 -29294 60426 -29260
rect 59866 -29300 60426 -29294
rect 59766 -29356 59806 -29350
rect 59103 -29512 59137 -29478
rect 56492 -29640 56530 -29606
rect 55882 -30204 55970 -30170
rect 55820 -31030 55854 -30254
rect 55998 -31030 56032 -30254
rect 55882 -31114 55970 -31080
rect 56430 -30475 56464 -29699
rect 56558 -30475 56592 -29699
rect 56492 -30568 56530 -30534
rect 57125 -29623 57159 -29589
rect 57217 -29623 57251 -29589
rect 57309 -29623 57343 -29589
rect 57086 -29710 57376 -29680
rect 57086 -29780 57116 -29710
rect 57116 -29780 57346 -29710
rect 57346 -29780 57376 -29710
rect 57086 -29810 57376 -29780
rect 58926 -30046 58930 -29560
rect 58930 -30046 58964 -29560
rect 58964 -30046 58966 -29560
rect 59044 -29947 59078 -29571
rect 59162 -29947 59196 -29571
rect 59103 -30040 59137 -30006
rect 58926 -30202 58966 -30046
rect 59766 -29534 59772 -29356
rect 59772 -29534 59806 -29356
rect 59958 -29408 60334 -29374
rect 59874 -29462 59908 -29428
rect 60384 -29462 60418 -29428
rect 59958 -29516 60334 -29482
rect 59766 -29540 59806 -29534
rect 59476 -29596 59656 -29590
rect 59476 -29630 59484 -29596
rect 59484 -29630 59642 -29596
rect 59642 -29630 59656 -29596
rect 59386 -29692 59426 -29690
rect 59386 -30048 59388 -29692
rect 59388 -30048 59422 -29692
rect 59422 -30048 59426 -29692
rect 59546 -29732 59580 -29698
rect 59502 -29958 59536 -29782
rect 59590 -29958 59624 -29782
rect 59546 -30042 59580 -30008
rect 59386 -30050 59426 -30048
rect 59862 -29732 59896 -29698
rect 59818 -29958 59852 -29782
rect 59906 -29958 59940 -29782
rect 59862 -30042 59896 -30008
rect 61196 -29820 61366 -29800
rect 61196 -29860 61216 -29820
rect 61216 -29860 61336 -29820
rect 61336 -29860 61366 -29820
rect 61196 -29880 61366 -29860
rect 57056 -30370 57416 -30340
rect 57056 -30450 57096 -30370
rect 57096 -30450 57376 -30370
rect 57376 -30450 57416 -30370
rect 57056 -30480 57416 -30450
rect 57125 -30599 57159 -30565
rect 57217 -30599 57251 -30565
rect 57309 -30599 57343 -30565
rect 58926 -30690 58930 -30202
rect 58930 -30690 58964 -30202
rect 58964 -30690 58966 -30202
rect 60127 -29991 60161 -29957
rect 60366 -29965 60406 -29960
rect 60366 -29999 60393 -29965
rect 60393 -29999 60406 -29965
rect 60366 -30000 60406 -29999
rect 60127 -30083 60161 -30049
rect 59103 -30242 59137 -30208
rect 59044 -30677 59078 -30301
rect 57118 -30797 57168 -30794
rect 57118 -30831 57133 -30797
rect 57133 -30831 57167 -30797
rect 57167 -30831 57168 -30797
rect 57118 -30844 57168 -30831
rect 57326 -30810 57376 -30770
rect 59162 -30677 59196 -30301
rect 59103 -30770 59137 -30736
rect 59386 -30205 59426 -30200
rect 59386 -30561 59387 -30205
rect 59387 -30561 59421 -30205
rect 59421 -30561 59426 -30205
rect 59545 -30245 59579 -30211
rect 59501 -30471 59535 -30295
rect 59589 -30471 59623 -30295
rect 59545 -30555 59579 -30521
rect 59386 -30570 59426 -30561
rect 59476 -30623 59646 -30620
rect 59861 -30245 59895 -30211
rect 59817 -30471 59851 -30295
rect 59905 -30471 59939 -30295
rect 59861 -30555 59895 -30521
rect 60127 -30175 60161 -30141
rect 60127 -30267 60161 -30233
rect 60671 -29991 60705 -29957
rect 60366 -30057 60406 -30050
rect 60366 -30090 60393 -30057
rect 60393 -30090 60406 -30057
rect 60366 -30141 60406 -30140
rect 60366 -30175 60393 -30141
rect 60393 -30175 60406 -30141
rect 60366 -30180 60406 -30175
rect 60366 -30225 60406 -30220
rect 60366 -30259 60393 -30225
rect 60393 -30259 60406 -30225
rect 60366 -30260 60406 -30259
rect 60671 -30083 60705 -30049
rect 60671 -30175 60705 -30141
rect 60671 -30267 60705 -30233
rect 60127 -30359 60161 -30325
rect 60297 -30359 60331 -30325
rect 60369 -30359 60405 -30325
rect 60449 -30359 60484 -30325
rect 60671 -30359 60705 -30325
rect 60747 -29991 60781 -29957
rect 61046 -29965 61086 -29960
rect 61046 -29999 61059 -29965
rect 61059 -29999 61086 -29965
rect 61046 -30000 61086 -29999
rect 60747 -30083 60781 -30049
rect 60747 -30175 60781 -30141
rect 60747 -30267 60781 -30233
rect 61291 -29991 61325 -29957
rect 61046 -30057 61086 -30050
rect 61046 -30090 61059 -30057
rect 61059 -30090 61086 -30057
rect 61046 -30141 61086 -30140
rect 61046 -30175 61059 -30141
rect 61059 -30175 61086 -30141
rect 61046 -30180 61086 -30175
rect 61046 -30225 61086 -30220
rect 61046 -30259 61059 -30225
rect 61059 -30259 61086 -30225
rect 61046 -30260 61086 -30259
rect 61291 -30083 61325 -30049
rect 61291 -30175 61325 -30141
rect 61291 -30267 61325 -30233
rect 60747 -30359 60781 -30325
rect 60980 -30359 61015 -30325
rect 61053 -30359 61088 -30325
rect 61129 -30358 61164 -30324
rect 61291 -30359 61325 -30325
rect 60486 -30500 60526 -30460
rect 60626 -30500 60666 -30460
rect 60766 -30500 60806 -30460
rect 60906 -30500 60946 -30460
rect 59476 -30657 59483 -30623
rect 59483 -30657 59641 -30623
rect 59641 -30657 59646 -30623
rect 59476 -30660 59646 -30657
rect 59766 -30722 59806 -30720
rect 58926 -30936 58966 -30910
rect 59766 -30900 59772 -30722
rect 59772 -30900 59806 -30722
rect 59958 -30774 60334 -30740
rect 59874 -30828 59908 -30794
rect 60384 -30828 60418 -30794
rect 59958 -30882 60334 -30848
rect 57125 -31143 57159 -31109
rect 57217 -31143 57251 -31109
rect 57309 -31143 57343 -31109
rect 54081 -31378 54857 -31344
rect 53988 -31444 54022 -31406
rect 54916 -31444 54950 -31406
rect 54081 -31506 54857 -31472
rect 56020 -31408 56080 -31258
rect 58926 -31222 58930 -30936
rect 58930 -31222 58964 -30936
rect 58964 -31222 58966 -30936
rect 59656 -30936 59706 -30930
rect 59125 -30988 59501 -30954
rect 59560 -31042 59594 -31008
rect 59125 -31096 59501 -31062
rect 59032 -31150 59066 -31116
rect 59125 -31204 59501 -31170
rect 57156 -31290 57316 -31260
rect 57156 -31390 57186 -31290
rect 57186 -31390 57286 -31290
rect 57286 -31390 57316 -31290
rect 58926 -31300 58966 -31222
rect 59656 -31222 59662 -30936
rect 59662 -31222 59696 -30936
rect 59696 -31222 59706 -30936
rect 59866 -30962 60426 -30960
rect 59866 -30996 59868 -30962
rect 59868 -30996 60424 -30962
rect 60424 -30996 60426 -30962
rect 59866 -31000 60426 -30996
rect 59656 -31230 59706 -31222
rect 57156 -31420 57316 -31390
rect 54150 -31620 54840 -31588
rect 54150 -31708 54840 -31620
rect 55300 -31592 55476 -31558
rect 55526 -31636 55560 -31602
rect 55300 -31680 55476 -31646
rect 55320 -31760 55470 -31748
rect 55320 -31794 55470 -31760
rect 55320 -31808 55470 -31794
rect 25700 -34128 25736 -32692
rect 25736 -34128 25770 -32692
rect 25770 -34128 25780 -32692
rect 25882 -33141 26996 -32744
rect 27124 -33141 28238 -32744
rect 28366 -33141 29480 -32744
rect 29608 -33141 30722 -32744
rect 30850 -33141 31964 -32744
rect 32092 -33141 33206 -32744
rect 33334 -33141 34448 -32744
rect 34576 -33141 35690 -32744
rect 25882 -34076 26996 -33679
rect 27124 -34076 28238 -33679
rect 28366 -34076 29480 -33679
rect 29608 -34076 30722 -33679
rect 30850 -34076 31964 -33679
rect 32092 -34076 33206 -33679
rect 33334 -34076 34448 -33679
rect 34576 -34076 35690 -33679
rect 25700 -34290 25780 -34128
rect 54150 -33958 54850 -33908
rect 25700 -35726 25736 -34290
rect 25736 -35726 25770 -34290
rect 25770 -35726 25780 -34290
rect 25882 -34739 26996 -34342
rect 27124 -34739 28238 -34342
rect 28366 -34739 29480 -34342
rect 29608 -34739 30722 -34342
rect 30850 -34739 31964 -34342
rect 32092 -34739 33206 -34342
rect 33334 -34739 34448 -34342
rect 34576 -34739 35690 -34342
rect 25882 -35674 26996 -35277
rect 27124 -35674 28238 -35277
rect 28366 -35674 29480 -35277
rect 29608 -35674 30722 -35277
rect 30850 -35674 31964 -35277
rect 32092 -35674 33206 -35277
rect 33334 -35674 34448 -35277
rect 34576 -35674 35690 -35277
rect 25700 -35892 25780 -35726
rect 54150 -33992 54850 -33958
rect 54150 -33998 54850 -33992
rect 54091 -34106 54867 -34072
rect 53998 -34172 54032 -34134
rect 54926 -34172 54960 -34134
rect 54091 -34234 54867 -34200
rect 55960 -34298 56040 -34128
rect 53526 -34540 53614 -34506
rect 25700 -37328 25736 -35892
rect 25736 -37328 25770 -35892
rect 25770 -37328 25780 -35892
rect 25882 -36341 26996 -35944
rect 27124 -36341 28238 -35944
rect 28366 -36341 29480 -35944
rect 29608 -36341 30722 -35944
rect 30850 -36341 31964 -35944
rect 32092 -36341 33206 -35944
rect 33334 -36341 34448 -35944
rect 34576 -36341 35690 -35944
rect 25882 -37276 26996 -36879
rect 27124 -37276 28238 -36879
rect 28366 -37276 29480 -36879
rect 29608 -37276 30722 -36879
rect 30850 -37276 31964 -36879
rect 32092 -37276 33206 -36879
rect 33334 -37276 34448 -36879
rect 34576 -37276 35690 -36879
rect 25700 -37492 25780 -37328
rect 53330 -35918 53350 -34568
rect 53350 -35918 53384 -34568
rect 53384 -35918 53400 -34568
rect 53464 -35366 53498 -34590
rect 53642 -35366 53676 -34590
rect 57126 -34300 57356 -34270
rect 54091 -34462 54867 -34428
rect 53998 -34528 54032 -34490
rect 54926 -34528 54960 -34490
rect 54091 -34590 54867 -34556
rect 55334 -34602 55368 -34568
rect 55290 -34828 55324 -34652
rect 55378 -34828 55412 -34652
rect 55142 -35108 55494 -35074
rect 53942 -35212 54718 -35178
rect 53858 -35328 53892 -35240
rect 54768 -35328 54802 -35240
rect 53942 -35390 54718 -35356
rect 53526 -35450 53614 -35416
rect 55046 -35194 55080 -35160
rect 55556 -35194 55590 -35160
rect 55142 -35280 55494 -35246
rect 57126 -34370 57156 -34300
rect 57156 -34370 57316 -34300
rect 57316 -34370 57356 -34300
rect 57126 -34400 57356 -34370
rect 58926 -34429 58966 -34420
rect 55882 -34490 55970 -34456
rect 55820 -35316 55854 -34540
rect 55998 -35316 56032 -34540
rect 55882 -35400 55970 -35366
rect 57125 -34479 57159 -34445
rect 57217 -34479 57251 -34445
rect 57309 -34479 57343 -34445
rect 57118 -34757 57178 -34744
rect 57118 -34791 57133 -34757
rect 57133 -34791 57167 -34757
rect 57167 -34791 57178 -34757
rect 57118 -34794 57178 -34791
rect 58926 -34715 58930 -34429
rect 58930 -34715 58964 -34429
rect 58964 -34715 58966 -34429
rect 59125 -34481 59501 -34447
rect 59560 -34535 59594 -34501
rect 59125 -34589 59501 -34555
rect 59032 -34643 59066 -34609
rect 59125 -34697 59501 -34663
rect 58926 -34720 58966 -34715
rect 59656 -34715 59662 -34430
rect 59662 -34715 59696 -34430
rect 59656 -34720 59696 -34715
rect 57326 -34780 57366 -34740
rect 53526 -35558 53614 -35524
rect 55030 -35528 55110 -35448
rect 55740 -35468 55810 -35448
rect 55740 -35502 55802 -35468
rect 55802 -35502 55810 -35468
rect 55740 -35528 55810 -35502
rect 53464 -36384 53498 -35608
rect 53642 -36384 53676 -35608
rect 53942 -35618 54718 -35584
rect 53858 -35734 53892 -35646
rect 54768 -35734 54802 -35646
rect 53942 -35796 54718 -35762
rect 55142 -35730 55494 -35696
rect 55046 -35816 55080 -35782
rect 55556 -35816 55590 -35782
rect 55142 -35902 55494 -35868
rect 53526 -36468 53614 -36434
rect 54081 -36422 54857 -36388
rect 53988 -36488 54022 -36450
rect 54916 -36488 54950 -36450
rect 54081 -36550 54857 -36516
rect 55280 -36324 55314 -36148
rect 55368 -36324 55402 -36148
rect 55324 -36408 55358 -36374
rect 56280 -35000 56350 -34918
rect 56280 -35548 56316 -35000
rect 56316 -35548 56350 -35000
rect 59866 -34694 59868 -34660
rect 59868 -34694 60424 -34660
rect 60424 -34694 60426 -34660
rect 59866 -34700 60426 -34694
rect 59766 -34756 59806 -34750
rect 59103 -34912 59137 -34878
rect 56492 -35040 56530 -35006
rect 55882 -35604 55970 -35570
rect 55820 -36430 55854 -35654
rect 55998 -36430 56032 -35654
rect 55882 -36514 55970 -36480
rect 56430 -35875 56464 -35099
rect 56558 -35875 56592 -35099
rect 56492 -35968 56530 -35934
rect 57125 -35023 57159 -34989
rect 57217 -35023 57251 -34989
rect 57309 -35023 57343 -34989
rect 57086 -35110 57376 -35080
rect 57086 -35180 57116 -35110
rect 57116 -35180 57346 -35110
rect 57346 -35180 57376 -35110
rect 57086 -35210 57376 -35180
rect 58926 -35446 58930 -34960
rect 58930 -35446 58964 -34960
rect 58964 -35446 58966 -34960
rect 59044 -35347 59078 -34971
rect 59162 -35347 59196 -34971
rect 59103 -35440 59137 -35406
rect 58926 -35602 58966 -35446
rect 59766 -34934 59772 -34756
rect 59772 -34934 59806 -34756
rect 59958 -34808 60334 -34774
rect 59874 -34862 59908 -34828
rect 60384 -34862 60418 -34828
rect 59958 -34916 60334 -34882
rect 59766 -34940 59806 -34934
rect 59476 -34996 59656 -34990
rect 59476 -35030 59484 -34996
rect 59484 -35030 59642 -34996
rect 59642 -35030 59656 -34996
rect 59386 -35092 59426 -35090
rect 59386 -35448 59388 -35092
rect 59388 -35448 59422 -35092
rect 59422 -35448 59426 -35092
rect 59546 -35132 59580 -35098
rect 59502 -35358 59536 -35182
rect 59590 -35358 59624 -35182
rect 59546 -35442 59580 -35408
rect 59386 -35450 59426 -35448
rect 59862 -35132 59896 -35098
rect 59818 -35358 59852 -35182
rect 59906 -35358 59940 -35182
rect 59862 -35442 59896 -35408
rect 61196 -35220 61366 -35200
rect 61196 -35260 61216 -35220
rect 61216 -35260 61336 -35220
rect 61336 -35260 61366 -35220
rect 61196 -35280 61366 -35260
rect 57056 -35770 57416 -35740
rect 57056 -35850 57096 -35770
rect 57096 -35850 57376 -35770
rect 57376 -35850 57416 -35770
rect 57056 -35880 57416 -35850
rect 57125 -35999 57159 -35965
rect 57217 -35999 57251 -35965
rect 57309 -35999 57343 -35965
rect 58926 -36090 58930 -35602
rect 58930 -36090 58964 -35602
rect 58964 -36090 58966 -35602
rect 60127 -35391 60161 -35357
rect 60366 -35365 60406 -35360
rect 60366 -35399 60393 -35365
rect 60393 -35399 60406 -35365
rect 60366 -35400 60406 -35399
rect 60127 -35483 60161 -35449
rect 59103 -35642 59137 -35608
rect 59044 -36077 59078 -35701
rect 57118 -36197 57168 -36194
rect 57118 -36231 57133 -36197
rect 57133 -36231 57167 -36197
rect 57167 -36231 57168 -36197
rect 57118 -36244 57168 -36231
rect 57326 -36210 57376 -36170
rect 59162 -36077 59196 -35701
rect 59103 -36170 59137 -36136
rect 59386 -35605 59426 -35600
rect 59386 -35961 59387 -35605
rect 59387 -35961 59421 -35605
rect 59421 -35961 59426 -35605
rect 59545 -35645 59579 -35611
rect 59501 -35871 59535 -35695
rect 59589 -35871 59623 -35695
rect 59545 -35955 59579 -35921
rect 59386 -35970 59426 -35961
rect 59476 -36023 59646 -36020
rect 59861 -35645 59895 -35611
rect 59817 -35871 59851 -35695
rect 59905 -35871 59939 -35695
rect 59861 -35955 59895 -35921
rect 60127 -35575 60161 -35541
rect 60127 -35667 60161 -35633
rect 60671 -35391 60705 -35357
rect 60366 -35457 60406 -35450
rect 60366 -35490 60393 -35457
rect 60393 -35490 60406 -35457
rect 60366 -35541 60406 -35540
rect 60366 -35575 60393 -35541
rect 60393 -35575 60406 -35541
rect 60366 -35580 60406 -35575
rect 60366 -35625 60406 -35620
rect 60366 -35659 60393 -35625
rect 60393 -35659 60406 -35625
rect 60366 -35660 60406 -35659
rect 60671 -35483 60705 -35449
rect 60671 -35575 60705 -35541
rect 60671 -35667 60705 -35633
rect 60127 -35759 60161 -35725
rect 60297 -35759 60331 -35725
rect 60369 -35759 60405 -35725
rect 60449 -35759 60484 -35725
rect 60671 -35759 60705 -35725
rect 60747 -35391 60781 -35357
rect 61046 -35365 61086 -35360
rect 61046 -35399 61059 -35365
rect 61059 -35399 61086 -35365
rect 61046 -35400 61086 -35399
rect 60747 -35483 60781 -35449
rect 60747 -35575 60781 -35541
rect 60747 -35667 60781 -35633
rect 61291 -35391 61325 -35357
rect 61046 -35457 61086 -35450
rect 61046 -35490 61059 -35457
rect 61059 -35490 61086 -35457
rect 61046 -35541 61086 -35540
rect 61046 -35575 61059 -35541
rect 61059 -35575 61086 -35541
rect 61046 -35580 61086 -35575
rect 61046 -35625 61086 -35620
rect 61046 -35659 61059 -35625
rect 61059 -35659 61086 -35625
rect 61046 -35660 61086 -35659
rect 61291 -35483 61325 -35449
rect 61291 -35575 61325 -35541
rect 61291 -35667 61325 -35633
rect 60747 -35759 60781 -35725
rect 60980 -35759 61015 -35725
rect 61053 -35759 61088 -35725
rect 61129 -35758 61164 -35724
rect 61291 -35759 61325 -35725
rect 60486 -35900 60526 -35860
rect 60626 -35900 60666 -35860
rect 60766 -35900 60806 -35860
rect 60906 -35900 60946 -35860
rect 59476 -36057 59483 -36023
rect 59483 -36057 59641 -36023
rect 59641 -36057 59646 -36023
rect 59476 -36060 59646 -36057
rect 59766 -36122 59806 -36120
rect 58926 -36336 58966 -36310
rect 59766 -36300 59772 -36122
rect 59772 -36300 59806 -36122
rect 59958 -36174 60334 -36140
rect 59874 -36228 59908 -36194
rect 60384 -36228 60418 -36194
rect 59958 -36282 60334 -36248
rect 57125 -36543 57159 -36509
rect 57217 -36543 57251 -36509
rect 57309 -36543 57343 -36509
rect 54081 -36778 54857 -36744
rect 53988 -36844 54022 -36806
rect 54916 -36844 54950 -36806
rect 54081 -36906 54857 -36872
rect 56020 -36808 56080 -36658
rect 58926 -36622 58930 -36336
rect 58930 -36622 58964 -36336
rect 58964 -36622 58966 -36336
rect 59656 -36336 59706 -36330
rect 59125 -36388 59501 -36354
rect 59560 -36442 59594 -36408
rect 59125 -36496 59501 -36462
rect 59032 -36550 59066 -36516
rect 59125 -36604 59501 -36570
rect 57156 -36690 57316 -36660
rect 57156 -36790 57186 -36690
rect 57186 -36790 57286 -36690
rect 57286 -36790 57316 -36690
rect 58926 -36700 58966 -36622
rect 59656 -36622 59662 -36336
rect 59662 -36622 59696 -36336
rect 59696 -36622 59706 -36336
rect 59866 -36362 60426 -36360
rect 59866 -36396 59868 -36362
rect 59868 -36396 60424 -36362
rect 60424 -36396 60426 -36362
rect 59866 -36400 60426 -36396
rect 59656 -36630 59706 -36622
rect 57156 -36820 57316 -36790
rect 54150 -37020 54840 -36988
rect 54150 -37108 54840 -37020
rect 55300 -36992 55476 -36958
rect 55526 -37036 55560 -37002
rect 55300 -37080 55476 -37046
rect 55320 -37160 55470 -37148
rect 55320 -37194 55470 -37160
rect 55320 -37208 55470 -37194
rect 25700 -38928 25736 -37492
rect 25736 -38928 25770 -37492
rect 25770 -38928 25780 -37492
rect 25882 -37941 26996 -37544
rect 27124 -37941 28238 -37544
rect 28366 -37941 29480 -37544
rect 29608 -37941 30722 -37544
rect 30850 -37941 31964 -37544
rect 32092 -37941 33206 -37544
rect 33334 -37941 34448 -37544
rect 34576 -37941 35690 -37544
rect 25882 -38876 26996 -38479
rect 27124 -38876 28238 -38479
rect 28366 -38876 29480 -38479
rect 29608 -38876 30722 -38479
rect 30850 -38876 31964 -38479
rect 32092 -38876 33206 -38479
rect 33334 -38876 34448 -38479
rect 34576 -38876 35690 -38479
rect 25700 -39094 25780 -38928
rect 77110 -38370 77220 -38350
rect 75535 -38405 75569 -38371
rect 75627 -38405 75661 -38371
rect 75719 -38405 75753 -38371
rect 75811 -38405 75845 -38371
rect 75903 -38405 75937 -38371
rect 75995 -38405 76029 -38371
rect 76085 -38405 76119 -38371
rect 76177 -38405 76211 -38371
rect 76269 -38405 76303 -38371
rect 76361 -38405 76395 -38371
rect 76453 -38405 76487 -38371
rect 76545 -38405 76579 -38371
rect 76637 -38405 76671 -38371
rect 76729 -38405 76763 -38371
rect 76821 -38405 76855 -38371
rect 75670 -38519 75704 -38517
rect 75670 -38551 75700 -38519
rect 75700 -38551 75704 -38519
rect 75580 -38637 75586 -38610
rect 75586 -38637 75620 -38610
rect 75580 -38650 75620 -38637
rect 75942 -38553 75976 -38520
rect 75942 -38554 75976 -38553
rect 75670 -38643 75704 -38609
rect 75862 -38637 75896 -38603
rect 76217 -38553 76250 -38519
rect 76250 -38553 76251 -38519
rect 75947 -38643 75981 -38609
rect 76128 -38637 76136 -38610
rect 76136 -38637 76162 -38610
rect 76128 -38644 76162 -38637
rect 76492 -38553 76526 -38519
rect 76224 -38644 76258 -38610
rect 76404 -38637 76412 -38609
rect 76412 -38637 76438 -38609
rect 76404 -38643 76438 -38637
rect 77110 -38420 77140 -38370
rect 77140 -38420 77190 -38370
rect 77190 -38420 77220 -38370
rect 76768 -38553 76802 -38521
rect 76768 -38555 76802 -38553
rect 76497 -38643 76531 -38609
rect 76680 -38637 76688 -38609
rect 76688 -38637 76714 -38609
rect 76680 -38643 76714 -38637
rect 77110 -38490 77220 -38420
rect 77110 -38540 77140 -38490
rect 77140 -38540 77190 -38490
rect 77190 -38540 77220 -38490
rect 77110 -38570 77220 -38540
rect 76772 -38644 76806 -38610
rect 75670 -38703 75704 -38698
rect 75670 -38732 75700 -38703
rect 75700 -38732 75704 -38703
rect 75943 -38737 75976 -38703
rect 75976 -38737 75977 -38703
rect 76215 -38737 76216 -38704
rect 76216 -38737 76249 -38704
rect 76215 -38738 76249 -38737
rect 76218 -38805 76250 -38776
rect 76250 -38805 76252 -38776
rect 76218 -38810 76252 -38805
rect 76492 -38737 76526 -38703
rect 76768 -38737 76802 -38703
rect 76930 -38830 77040 -38800
rect 76930 -38880 76960 -38830
rect 76960 -38880 77010 -38830
rect 77010 -38880 77040 -38830
rect 75535 -38949 75569 -38915
rect 75627 -38949 75661 -38915
rect 75719 -38949 75753 -38915
rect 75811 -38949 75845 -38915
rect 75903 -38949 75937 -38915
rect 75995 -38949 76029 -38915
rect 76085 -38949 76119 -38915
rect 76177 -38949 76211 -38915
rect 76269 -38949 76303 -38915
rect 76361 -38949 76395 -38915
rect 76453 -38949 76487 -38915
rect 76545 -38949 76579 -38915
rect 76637 -38949 76671 -38915
rect 76729 -38949 76763 -38915
rect 76821 -38949 76855 -38915
rect 76930 -38960 77040 -38880
rect 80890 -38820 81070 -38790
rect 80890 -38930 80920 -38820
rect 80920 -38930 81030 -38820
rect 81030 -38930 81070 -38820
rect 80890 -38960 81070 -38930
rect 81500 -38820 81680 -38790
rect 81500 -38930 81540 -38820
rect 81540 -38930 81650 -38820
rect 81650 -38930 81680 -38820
rect 81500 -38960 81680 -38930
rect 82110 -38830 82290 -38800
rect 82110 -38940 82140 -38830
rect 82140 -38940 82250 -38830
rect 82250 -38940 82290 -38830
rect 25700 -40530 25738 -39094
rect 25738 -40530 25772 -39094
rect 25772 -40530 25780 -39094
rect 76930 -39010 76960 -38960
rect 76960 -39010 77010 -38960
rect 77010 -39010 77040 -38960
rect 82110 -38970 82290 -38940
rect 82760 -38840 82940 -38810
rect 82760 -38950 82790 -38840
rect 82790 -38950 82900 -38840
rect 82900 -38950 82940 -38840
rect 82760 -38980 82940 -38950
rect 83470 -38830 83650 -38800
rect 83470 -38940 83510 -38830
rect 83510 -38940 83620 -38830
rect 83620 -38940 83650 -38830
rect 83470 -38970 83650 -38940
rect 84190 -38830 84370 -38800
rect 84190 -38940 84220 -38830
rect 84220 -38940 84330 -38830
rect 84330 -38940 84370 -38830
rect 84190 -38970 84370 -38940
rect 85840 -38850 86020 -38820
rect 85840 -38960 85880 -38850
rect 85880 -38960 85990 -38850
rect 85990 -38960 86020 -38850
rect 85840 -38990 86020 -38960
rect 87280 -38860 87460 -38830
rect 87280 -38970 87320 -38860
rect 87320 -38970 87430 -38860
rect 87430 -38970 87460 -38860
rect 87280 -39000 87460 -38970
rect 76930 -39040 77040 -39010
rect 77607 -39075 77641 -39041
rect 77699 -39075 77733 -39041
rect 77791 -39075 77825 -39041
rect 77883 -39075 77917 -39041
rect 77975 -39075 78009 -39041
rect 78067 -39075 78101 -39041
rect 78159 -39075 78193 -39041
rect 78251 -39075 78285 -39041
rect 78343 -39075 78377 -39041
rect 78435 -39075 78469 -39041
rect 78527 -39075 78561 -39041
rect 78619 -39075 78653 -39041
rect 78711 -39075 78745 -39041
rect 78803 -39075 78837 -39041
rect 78895 -39075 78929 -39041
rect 78987 -39075 79021 -39041
rect 25884 -39543 26998 -39146
rect 27126 -39543 28240 -39146
rect 28368 -39543 29482 -39146
rect 29610 -39543 30724 -39146
rect 30852 -39543 31966 -39146
rect 32094 -39543 33208 -39146
rect 33336 -39543 34450 -39146
rect 34578 -39543 35692 -39146
rect 25884 -40478 26998 -40081
rect 27126 -40478 28240 -40081
rect 28368 -40478 29482 -40081
rect 29610 -40478 30724 -40081
rect 30852 -40478 31966 -40081
rect 32094 -40478 33208 -40081
rect 33336 -40478 34450 -40081
rect 34578 -40478 35692 -40081
rect 25700 -40692 25780 -40530
rect 77430 -39170 77520 -39130
rect 54150 -39358 54850 -39308
rect 77780 -39320 77820 -39280
rect 80767 -39125 80801 -39091
rect 80859 -39125 80893 -39091
rect 80951 -39125 80985 -39091
rect 81043 -39125 81077 -39091
rect 81135 -39125 81169 -39091
rect 81227 -39125 81261 -39091
rect 81319 -39125 81353 -39091
rect 81411 -39125 81445 -39091
rect 81503 -39125 81537 -39091
rect 81595 -39125 81629 -39091
rect 81687 -39125 81721 -39091
rect 81779 -39125 81813 -39091
rect 81871 -39125 81905 -39091
rect 81963 -39125 81997 -39091
rect 82055 -39125 82089 -39091
rect 82147 -39125 82181 -39091
rect 82239 -39125 82273 -39091
rect 82331 -39125 82365 -39091
rect 82423 -39125 82457 -39091
rect 82515 -39125 82549 -39091
rect 82607 -39125 82641 -39091
rect 82699 -39125 82733 -39091
rect 82791 -39125 82825 -39091
rect 82883 -39125 82917 -39091
rect 82975 -39125 83009 -39091
rect 83067 -39125 83101 -39091
rect 83159 -39125 83193 -39091
rect 83251 -39125 83285 -39091
rect 83343 -39125 83377 -39091
rect 83435 -39125 83469 -39091
rect 83527 -39125 83561 -39091
rect 83619 -39125 83653 -39091
rect 83711 -39125 83745 -39091
rect 83803 -39125 83837 -39091
rect 83895 -39125 83929 -39091
rect 83987 -39125 84021 -39091
rect 84079 -39125 84113 -39091
rect 84171 -39125 84205 -39091
rect 84263 -39125 84297 -39091
rect 84355 -39125 84389 -39091
rect 84447 -39125 84481 -39091
rect 84539 -39125 84573 -39091
rect 84631 -39125 84665 -39091
rect 84723 -39125 84757 -39091
rect 84815 -39125 84849 -39091
rect 84907 -39125 84941 -39091
rect 84999 -39125 85033 -39091
rect 85091 -39125 85125 -39091
rect 85183 -39125 85217 -39091
rect 85275 -39125 85309 -39091
rect 85367 -39125 85401 -39091
rect 85459 -39125 85493 -39091
rect 85551 -39125 85585 -39091
rect 85643 -39125 85677 -39091
rect 85735 -39125 85769 -39091
rect 85827 -39125 85861 -39091
rect 85919 -39125 85953 -39091
rect 86011 -39125 86045 -39091
rect 86103 -39125 86137 -39091
rect 86195 -39125 86229 -39091
rect 86287 -39125 86321 -39091
rect 86379 -39125 86413 -39091
rect 86471 -39125 86505 -39091
rect 86563 -39125 86597 -39091
rect 86655 -39125 86689 -39091
rect 86747 -39125 86781 -39091
rect 86839 -39125 86873 -39091
rect 86931 -39125 86965 -39091
rect 87023 -39125 87057 -39091
rect 87115 -39125 87149 -39091
rect 87207 -39125 87241 -39091
rect 87299 -39125 87333 -39091
rect 87391 -39125 87425 -39091
rect 87483 -39125 87517 -39091
rect 87575 -39125 87609 -39091
rect 87667 -39125 87701 -39091
rect 87759 -39125 87793 -39091
rect 87851 -39125 87885 -39091
rect 87943 -39125 87977 -39091
rect 88035 -39125 88069 -39091
rect 88127 -39125 88161 -39091
rect 88219 -39125 88253 -39091
rect 88311 -39125 88345 -39091
rect 88403 -39125 88437 -39091
rect 88495 -39125 88529 -39091
rect 88587 -39125 88621 -39091
rect 88679 -39125 88713 -39091
rect 88771 -39125 88805 -39091
rect 54150 -39392 54850 -39358
rect 54150 -39398 54850 -39392
rect 54091 -39506 54867 -39472
rect 53998 -39572 54032 -39534
rect 54926 -39572 54960 -39534
rect 54091 -39634 54867 -39600
rect 77900 -39353 77940 -39350
rect 77900 -39387 77915 -39353
rect 77915 -39387 77940 -39353
rect 77900 -39390 77940 -39387
rect 77240 -39490 77300 -39450
rect 77420 -39490 77540 -39460
rect 78160 -39353 78200 -39350
rect 78160 -39387 78164 -39353
rect 78164 -39387 78198 -39353
rect 78198 -39387 78200 -39353
rect 78160 -39390 78200 -39387
rect 78290 -39390 78330 -39350
rect 78370 -39353 78410 -39350
rect 78370 -39387 78374 -39353
rect 78374 -39387 78408 -39353
rect 78408 -39387 78410 -39353
rect 78370 -39390 78410 -39387
rect 78590 -39370 78630 -39330
rect 78800 -39353 78850 -39340
rect 78800 -39380 78805 -39353
rect 78805 -39380 78839 -39353
rect 78839 -39380 78850 -39353
rect 55960 -39698 56040 -39528
rect 77420 -39550 77450 -39490
rect 77450 -39550 77510 -39490
rect 77510 -39550 77540 -39490
rect 77420 -39580 77540 -39550
rect 79080 -39400 79140 -39340
rect 79080 -39510 79140 -39450
rect 80480 -39510 80640 -39350
rect 82780 -39269 82782 -39240
rect 82782 -39269 82816 -39240
rect 82816 -39269 82820 -39240
rect 82780 -39280 82820 -39269
rect 82780 -39339 82782 -39320
rect 82782 -39339 82816 -39320
rect 82816 -39339 82820 -39320
rect 82780 -39360 82820 -39339
rect 84250 -39269 84254 -39260
rect 84254 -39269 84288 -39260
rect 84288 -39269 84290 -39260
rect 84250 -39305 84290 -39269
rect 84250 -39339 84254 -39305
rect 84254 -39339 84288 -39305
rect 84288 -39339 84290 -39305
rect 82780 -39440 82820 -39400
rect 83368 -39403 83773 -39394
rect 83368 -39434 83499 -39403
rect 83499 -39434 83533 -39403
rect 83533 -39434 83666 -39403
rect 83666 -39434 83700 -39403
rect 83700 -39434 83773 -39403
rect 77607 -39619 77641 -39585
rect 77699 -39619 77733 -39585
rect 77791 -39619 77825 -39585
rect 77883 -39619 77917 -39585
rect 77975 -39619 78009 -39585
rect 78067 -39619 78101 -39585
rect 78159 -39619 78193 -39585
rect 78251 -39619 78285 -39585
rect 78343 -39619 78377 -39585
rect 78435 -39619 78469 -39585
rect 78527 -39619 78561 -39585
rect 78619 -39619 78653 -39585
rect 78711 -39619 78745 -39585
rect 78803 -39619 78837 -39585
rect 78895 -39619 78929 -39585
rect 78987 -39619 79021 -39585
rect 82780 -39491 82820 -39490
rect 82780 -39525 82782 -39491
rect 82782 -39525 82816 -39491
rect 82816 -39525 82820 -39491
rect 82780 -39530 82820 -39525
rect 84250 -39491 84290 -39339
rect 84250 -39525 84254 -39491
rect 84254 -39525 84288 -39491
rect 84288 -39525 84290 -39491
rect 84250 -39530 84290 -39525
rect 85730 -39305 85770 -39270
rect 85730 -39339 85760 -39305
rect 85760 -39339 85770 -39305
rect 84870 -39403 85240 -39397
rect 84870 -39437 84971 -39403
rect 84971 -39437 85005 -39403
rect 85005 -39437 85138 -39403
rect 85138 -39437 85172 -39403
rect 85172 -39437 85240 -39403
rect 85730 -39491 85770 -39339
rect 85730 -39525 85760 -39491
rect 85760 -39525 85770 -39491
rect 85730 -39540 85770 -39525
rect 87200 -39269 87232 -39240
rect 87232 -39269 87240 -39240
rect 87200 -39305 87240 -39269
rect 87200 -39339 87232 -39305
rect 87232 -39339 87240 -39305
rect 86329 -39403 86699 -39394
rect 86329 -39434 86443 -39403
rect 86443 -39434 86477 -39403
rect 86477 -39434 86610 -39403
rect 86610 -39434 86644 -39403
rect 86644 -39434 86699 -39403
rect 87200 -39491 87240 -39339
rect 87200 -39510 87232 -39491
rect 87232 -39510 87240 -39491
rect 88670 -39269 88704 -39260
rect 88704 -39269 88710 -39260
rect 88670 -39305 88710 -39269
rect 88670 -39339 88704 -39305
rect 88704 -39339 88710 -39305
rect 87469 -39403 87749 -39395
rect 87469 -39435 87578 -39403
rect 87578 -39435 87612 -39403
rect 87612 -39435 87746 -39403
rect 87746 -39435 87749 -39403
rect 88670 -39491 88710 -39339
rect 88670 -39525 88704 -39491
rect 88704 -39525 88710 -39491
rect 88670 -39530 88710 -39525
rect 53526 -39940 53614 -39906
rect 25700 -42128 25736 -40692
rect 25736 -42128 25770 -40692
rect 25770 -42128 25780 -40692
rect 25882 -41141 26996 -40744
rect 27124 -41141 28238 -40744
rect 28366 -41141 29480 -40744
rect 29608 -41141 30722 -40744
rect 30850 -41141 31964 -40744
rect 32092 -41141 33206 -40744
rect 33334 -41141 34448 -40744
rect 34576 -41141 35690 -40744
rect 25882 -42076 26996 -41679
rect 27124 -42076 28238 -41679
rect 28366 -42076 29480 -41679
rect 29608 -42076 30722 -41679
rect 30850 -42076 31964 -41679
rect 32092 -42076 33206 -41679
rect 33334 -42076 34448 -41679
rect 34576 -42076 35690 -41679
rect 25700 -42290 25780 -42128
rect 53330 -41318 53350 -39968
rect 53350 -41318 53384 -39968
rect 53384 -41318 53400 -39968
rect 53464 -40766 53498 -39990
rect 53642 -40766 53676 -39990
rect 57126 -39700 57356 -39670
rect 54091 -39862 54867 -39828
rect 53998 -39928 54032 -39890
rect 54926 -39928 54960 -39890
rect 54091 -39990 54867 -39956
rect 55334 -40002 55368 -39968
rect 55290 -40228 55324 -40052
rect 55378 -40228 55412 -40052
rect 55142 -40508 55494 -40474
rect 53942 -40612 54718 -40578
rect 53858 -40728 53892 -40640
rect 54768 -40728 54802 -40640
rect 53942 -40790 54718 -40756
rect 53526 -40850 53614 -40816
rect 55046 -40594 55080 -40560
rect 55556 -40594 55590 -40560
rect 55142 -40680 55494 -40646
rect 57126 -39770 57156 -39700
rect 57156 -39770 57316 -39700
rect 57316 -39770 57356 -39700
rect 77420 -39690 77540 -39660
rect 80767 -39669 80801 -39635
rect 80859 -39669 80893 -39635
rect 80951 -39669 80985 -39635
rect 81043 -39669 81077 -39635
rect 81135 -39669 81169 -39635
rect 81227 -39669 81261 -39635
rect 81319 -39669 81353 -39635
rect 81411 -39669 81445 -39635
rect 81503 -39669 81537 -39635
rect 81595 -39669 81629 -39635
rect 81687 -39669 81721 -39635
rect 81779 -39669 81813 -39635
rect 81871 -39669 81905 -39635
rect 81963 -39669 81997 -39635
rect 82055 -39669 82089 -39635
rect 82147 -39669 82181 -39635
rect 82239 -39669 82273 -39635
rect 82331 -39669 82365 -39635
rect 82423 -39669 82457 -39635
rect 82515 -39669 82549 -39635
rect 82607 -39669 82641 -39635
rect 82699 -39669 82733 -39635
rect 82791 -39669 82825 -39635
rect 82883 -39669 82917 -39635
rect 82975 -39669 83009 -39635
rect 83067 -39669 83101 -39635
rect 83159 -39669 83193 -39635
rect 83251 -39669 83285 -39635
rect 83343 -39669 83377 -39635
rect 83435 -39669 83469 -39635
rect 83527 -39669 83561 -39635
rect 83619 -39669 83653 -39635
rect 83711 -39669 83745 -39635
rect 83803 -39669 83837 -39635
rect 83895 -39669 83929 -39635
rect 83987 -39669 84021 -39635
rect 84079 -39669 84113 -39635
rect 84171 -39669 84205 -39635
rect 84263 -39669 84297 -39635
rect 84355 -39669 84389 -39635
rect 84447 -39669 84481 -39635
rect 84539 -39669 84573 -39635
rect 84631 -39669 84665 -39635
rect 84723 -39669 84757 -39635
rect 84815 -39669 84849 -39635
rect 84907 -39669 84941 -39635
rect 84999 -39669 85033 -39635
rect 85091 -39669 85125 -39635
rect 85183 -39669 85217 -39635
rect 85275 -39669 85309 -39635
rect 85367 -39669 85401 -39635
rect 85459 -39669 85493 -39635
rect 85551 -39669 85585 -39635
rect 85643 -39669 85677 -39635
rect 85735 -39669 85769 -39635
rect 85827 -39669 85861 -39635
rect 85919 -39669 85953 -39635
rect 86011 -39669 86045 -39635
rect 86103 -39669 86137 -39635
rect 86195 -39669 86229 -39635
rect 86287 -39669 86321 -39635
rect 86379 -39669 86413 -39635
rect 86471 -39669 86505 -39635
rect 86563 -39669 86597 -39635
rect 86655 -39669 86689 -39635
rect 86747 -39669 86781 -39635
rect 86839 -39669 86873 -39635
rect 86931 -39669 86965 -39635
rect 87023 -39669 87057 -39635
rect 87115 -39669 87149 -39635
rect 87207 -39669 87241 -39635
rect 87299 -39669 87333 -39635
rect 87391 -39669 87425 -39635
rect 87483 -39669 87517 -39635
rect 87575 -39669 87609 -39635
rect 87667 -39669 87701 -39635
rect 87759 -39669 87793 -39635
rect 87851 -39669 87885 -39635
rect 87943 -39669 87977 -39635
rect 88035 -39669 88069 -39635
rect 88127 -39669 88161 -39635
rect 88219 -39669 88253 -39635
rect 88311 -39669 88345 -39635
rect 88403 -39669 88437 -39635
rect 88495 -39669 88529 -39635
rect 88587 -39669 88621 -39635
rect 88679 -39669 88713 -39635
rect 88771 -39669 88805 -39635
rect 57126 -39800 57356 -39770
rect 77420 -39750 77450 -39690
rect 77450 -39750 77510 -39690
rect 77510 -39750 77540 -39690
rect 77607 -39705 77641 -39671
rect 77699 -39705 77733 -39671
rect 77791 -39705 77825 -39671
rect 77883 -39705 77917 -39671
rect 77975 -39705 78009 -39671
rect 78067 -39705 78101 -39671
rect 58926 -39829 58966 -39820
rect 55882 -39890 55970 -39856
rect 55820 -40716 55854 -39940
rect 55998 -40716 56032 -39940
rect 55882 -40800 55970 -40766
rect 57125 -39879 57159 -39845
rect 57217 -39879 57251 -39845
rect 57309 -39879 57343 -39845
rect 57118 -40157 57178 -40144
rect 57118 -40191 57133 -40157
rect 57133 -40191 57167 -40157
rect 57167 -40191 57178 -40157
rect 57118 -40194 57178 -40191
rect 58926 -40115 58930 -39829
rect 58930 -40115 58964 -39829
rect 58964 -40115 58966 -39829
rect 59125 -39881 59501 -39847
rect 59560 -39935 59594 -39901
rect 59125 -39989 59501 -39955
rect 59032 -40043 59066 -40009
rect 59125 -40097 59501 -40063
rect 58926 -40120 58966 -40115
rect 59656 -40115 59662 -39830
rect 59662 -40115 59696 -39830
rect 77420 -39780 77540 -39750
rect 77170 -39840 77260 -39790
rect 80817 -39745 80851 -39711
rect 80909 -39745 80943 -39711
rect 81001 -39745 81035 -39711
rect 78160 -39830 78200 -39790
rect 77900 -39903 77940 -39900
rect 77900 -39937 77915 -39903
rect 77915 -39937 77940 -39903
rect 77900 -39940 77940 -39937
rect 78160 -39940 78200 -39900
rect 77770 -40000 77810 -39960
rect 80480 -39960 80640 -39800
rect 82490 -39770 82660 -39740
rect 59656 -40120 59696 -40115
rect 57326 -40180 57366 -40140
rect 53526 -40958 53614 -40924
rect 55030 -40928 55110 -40848
rect 55740 -40868 55810 -40848
rect 55740 -40902 55802 -40868
rect 55802 -40902 55810 -40868
rect 55740 -40928 55810 -40902
rect 53464 -41784 53498 -41008
rect 53642 -41784 53676 -41008
rect 53942 -41018 54718 -40984
rect 53858 -41134 53892 -41046
rect 54768 -41134 54802 -41046
rect 53942 -41196 54718 -41162
rect 55142 -41130 55494 -41096
rect 55046 -41216 55080 -41182
rect 55556 -41216 55590 -41182
rect 55142 -41302 55494 -41268
rect 53526 -41868 53614 -41834
rect 54081 -41822 54857 -41788
rect 53988 -41888 54022 -41850
rect 54916 -41888 54950 -41850
rect 54081 -41950 54857 -41916
rect 25700 -43726 25736 -42290
rect 25736 -43726 25770 -42290
rect 25770 -43726 25780 -42290
rect 25882 -42739 26996 -42342
rect 27124 -42739 28238 -42342
rect 28366 -42739 29480 -42342
rect 29608 -42739 30722 -42342
rect 30850 -42739 31964 -42342
rect 32092 -42739 33206 -42342
rect 33334 -42739 34448 -42342
rect 34576 -42739 35690 -42342
rect 25882 -43674 26996 -43277
rect 27124 -43674 28238 -43277
rect 28366 -43674 29480 -43277
rect 29608 -43674 30722 -43277
rect 30850 -43674 31964 -43277
rect 32092 -43674 33206 -43277
rect 33334 -43674 34448 -43277
rect 34576 -43674 35690 -43277
rect 25700 -43892 25780 -43726
rect 55280 -41724 55314 -41548
rect 55368 -41724 55402 -41548
rect 55324 -41808 55358 -41774
rect 56280 -40400 56350 -40318
rect 56280 -40948 56316 -40400
rect 56316 -40948 56350 -40400
rect 59866 -40094 59868 -40060
rect 59868 -40094 60424 -40060
rect 60424 -40094 60426 -40060
rect 59866 -40100 60426 -40094
rect 59766 -40156 59806 -40150
rect 59103 -40312 59137 -40278
rect 56492 -40440 56530 -40406
rect 55882 -41004 55970 -40970
rect 55820 -41830 55854 -41054
rect 55998 -41830 56032 -41054
rect 55882 -41914 55970 -41880
rect 56430 -41275 56464 -40499
rect 56558 -41275 56592 -40499
rect 56492 -41368 56530 -41334
rect 57125 -40423 57159 -40389
rect 57217 -40423 57251 -40389
rect 57309 -40423 57343 -40389
rect 57086 -40510 57376 -40480
rect 57086 -40580 57116 -40510
rect 57116 -40580 57346 -40510
rect 57346 -40580 57376 -40510
rect 57086 -40610 57376 -40580
rect 58926 -40846 58930 -40360
rect 58930 -40846 58964 -40360
rect 58964 -40846 58966 -40360
rect 59044 -40747 59078 -40371
rect 59162 -40747 59196 -40371
rect 59103 -40840 59137 -40806
rect 58926 -41002 58966 -40846
rect 59766 -40334 59772 -40156
rect 59772 -40334 59806 -40156
rect 59958 -40208 60334 -40174
rect 59874 -40262 59908 -40228
rect 60384 -40262 60418 -40228
rect 59958 -40316 60334 -40282
rect 59766 -40340 59806 -40334
rect 59476 -40396 59656 -40390
rect 77420 -40170 77470 -40120
rect 78160 -40060 78200 -40020
rect 81590 -39800 81760 -39770
rect 81590 -39910 81620 -39800
rect 81620 -39910 81730 -39800
rect 81730 -39910 81760 -39800
rect 82490 -39880 82520 -39770
rect 82520 -39880 82630 -39770
rect 82630 -39880 82660 -39770
rect 82490 -39910 82660 -39880
rect 83750 -39780 83920 -39750
rect 83750 -39890 83780 -39780
rect 83780 -39890 83890 -39780
rect 83890 -39890 83920 -39780
rect 81590 -39940 81760 -39910
rect 83750 -39920 83920 -39890
rect 85160 -39770 85330 -39740
rect 85160 -39880 85190 -39770
rect 85190 -39880 85300 -39770
rect 85300 -39880 85330 -39770
rect 85160 -39910 85330 -39880
rect 86320 -39780 86490 -39750
rect 86320 -39890 86350 -39780
rect 86350 -39890 86460 -39780
rect 86460 -39890 86490 -39780
rect 86320 -39920 86490 -39890
rect 87390 -39770 87560 -39740
rect 87390 -39880 87420 -39770
rect 87420 -39880 87530 -39770
rect 87530 -39880 87560 -39770
rect 87390 -39910 87560 -39880
rect 88500 -39760 88670 -39730
rect 88500 -39870 88530 -39760
rect 88530 -39870 88640 -39760
rect 88640 -39870 88670 -39760
rect 88500 -39900 88670 -39870
rect 77607 -40249 77641 -40215
rect 77699 -40249 77733 -40215
rect 77791 -40249 77825 -40215
rect 77883 -40249 77917 -40215
rect 77975 -40249 78009 -40215
rect 78067 -40249 78101 -40215
rect 78250 -40250 78360 -40220
rect 77607 -40325 77641 -40291
rect 77699 -40325 77733 -40291
rect 77791 -40325 77825 -40291
rect 77883 -40325 77917 -40291
rect 77975 -40325 78009 -40291
rect 78250 -40300 78280 -40250
rect 78280 -40300 78330 -40250
rect 78330 -40300 78360 -40250
rect 59476 -40430 59484 -40396
rect 59484 -40430 59642 -40396
rect 59642 -40430 59656 -40396
rect 78250 -40330 78360 -40300
rect 78560 -40250 78670 -40220
rect 78560 -40300 78590 -40250
rect 78590 -40300 78640 -40250
rect 78640 -40300 78670 -40250
rect 78560 -40330 78670 -40300
rect 78800 -40250 78910 -40220
rect 78800 -40300 78830 -40250
rect 78830 -40300 78880 -40250
rect 78880 -40300 78910 -40250
rect 78800 -40330 78910 -40300
rect 79060 -40250 79170 -40220
rect 79060 -40300 79090 -40250
rect 79090 -40300 79140 -40250
rect 79140 -40300 79170 -40250
rect 80940 -40077 80948 -40050
rect 80948 -40077 80982 -40050
rect 80982 -40077 80990 -40050
rect 80940 -40111 80990 -40077
rect 80940 -40145 80948 -40111
rect 80948 -40145 80982 -40111
rect 80982 -40145 80990 -40111
rect 80940 -40160 80990 -40145
rect 80817 -40289 80851 -40255
rect 80909 -40289 80943 -40255
rect 81001 -40289 81035 -40255
rect 79060 -40330 79170 -40300
rect 59386 -40492 59426 -40490
rect 59386 -40848 59388 -40492
rect 59388 -40848 59422 -40492
rect 59422 -40848 59426 -40492
rect 59546 -40532 59580 -40498
rect 59502 -40758 59536 -40582
rect 59590 -40758 59624 -40582
rect 59546 -40842 59580 -40808
rect 59386 -40850 59426 -40848
rect 59862 -40532 59896 -40498
rect 59818 -40758 59852 -40582
rect 59906 -40758 59940 -40582
rect 59862 -40842 59896 -40808
rect 80850 -40360 81020 -40330
rect 77460 -40600 77510 -40550
rect 80850 -40470 80880 -40360
rect 80880 -40470 80990 -40360
rect 80990 -40470 81020 -40360
rect 80850 -40500 81020 -40470
rect 78000 -40570 78040 -40530
rect 61196 -40620 61366 -40600
rect 61196 -40660 61216 -40620
rect 61216 -40660 61336 -40620
rect 61336 -40660 61366 -40620
rect 77790 -40603 77830 -40590
rect 77790 -40630 77793 -40603
rect 77793 -40630 77827 -40603
rect 77827 -40630 77830 -40603
rect 61196 -40680 61366 -40660
rect 57056 -41170 57416 -41140
rect 57056 -41250 57096 -41170
rect 57096 -41250 57376 -41170
rect 57376 -41250 57416 -41170
rect 57056 -41280 57416 -41250
rect 57125 -41399 57159 -41365
rect 57217 -41399 57251 -41365
rect 57309 -41399 57343 -41365
rect 58926 -41490 58930 -41002
rect 58930 -41490 58964 -41002
rect 58964 -41490 58966 -41002
rect 60127 -40791 60161 -40757
rect 60366 -40765 60406 -40760
rect 60366 -40799 60393 -40765
rect 60393 -40799 60406 -40765
rect 60366 -40800 60406 -40799
rect 60127 -40883 60161 -40849
rect 59103 -41042 59137 -41008
rect 59044 -41477 59078 -41101
rect 57118 -41597 57168 -41594
rect 57118 -41631 57133 -41597
rect 57133 -41631 57167 -41597
rect 57167 -41631 57168 -41597
rect 57118 -41644 57168 -41631
rect 57326 -41610 57376 -41570
rect 59162 -41477 59196 -41101
rect 59103 -41570 59137 -41536
rect 59386 -41005 59426 -41000
rect 59386 -41361 59387 -41005
rect 59387 -41361 59421 -41005
rect 59421 -41361 59426 -41005
rect 59545 -41045 59579 -41011
rect 59501 -41271 59535 -41095
rect 59589 -41271 59623 -41095
rect 59545 -41355 59579 -41321
rect 59386 -41370 59426 -41361
rect 59476 -41423 59646 -41420
rect 59861 -41045 59895 -41011
rect 59817 -41271 59851 -41095
rect 59905 -41271 59939 -41095
rect 59861 -41355 59895 -41321
rect 60127 -40975 60161 -40941
rect 60127 -41067 60161 -41033
rect 60671 -40791 60705 -40757
rect 60366 -40857 60406 -40850
rect 60366 -40890 60393 -40857
rect 60393 -40890 60406 -40857
rect 60366 -40941 60406 -40940
rect 60366 -40975 60393 -40941
rect 60393 -40975 60406 -40941
rect 60366 -40980 60406 -40975
rect 60366 -41025 60406 -41020
rect 60366 -41059 60393 -41025
rect 60393 -41059 60406 -41025
rect 60366 -41060 60406 -41059
rect 60671 -40883 60705 -40849
rect 60671 -40975 60705 -40941
rect 60671 -41067 60705 -41033
rect 60127 -41159 60161 -41125
rect 60297 -41159 60331 -41125
rect 60369 -41159 60405 -41125
rect 60449 -41159 60484 -41125
rect 60671 -41159 60705 -41125
rect 60747 -40791 60781 -40757
rect 61046 -40765 61086 -40760
rect 61046 -40799 61059 -40765
rect 61059 -40799 61086 -40765
rect 61046 -40800 61086 -40799
rect 60747 -40883 60781 -40849
rect 60747 -40975 60781 -40941
rect 60747 -41067 60781 -41033
rect 61291 -40791 61325 -40757
rect 61046 -40857 61086 -40850
rect 61046 -40890 61059 -40857
rect 61059 -40890 61086 -40857
rect 61046 -40941 61086 -40940
rect 61046 -40975 61059 -40941
rect 61059 -40975 61086 -40941
rect 61046 -40980 61086 -40975
rect 61046 -41025 61086 -41020
rect 61046 -41059 61059 -41025
rect 61059 -41059 61086 -41025
rect 61046 -41060 61086 -41059
rect 77400 -40730 77520 -40700
rect 77400 -40790 77430 -40730
rect 77430 -40790 77490 -40730
rect 77490 -40790 77520 -40730
rect 78000 -40660 78040 -40620
rect 78000 -40740 78040 -40700
rect 77400 -40820 77520 -40790
rect 61291 -40883 61325 -40849
rect 77607 -40869 77641 -40835
rect 77699 -40869 77733 -40835
rect 77791 -40869 77825 -40835
rect 77883 -40869 77917 -40835
rect 77975 -40869 78009 -40835
rect 61291 -40975 61325 -40941
rect 77607 -40945 77641 -40911
rect 77699 -40945 77733 -40911
rect 77791 -40945 77825 -40911
rect 77883 -40945 77917 -40911
rect 77975 -40945 78009 -40911
rect 78067 -40945 78101 -40911
rect 78159 -40945 78193 -40911
rect 78251 -40945 78285 -40911
rect 78343 -40945 78377 -40911
rect 78435 -40945 78469 -40911
rect 78527 -40945 78561 -40911
rect 61291 -41067 61325 -41033
rect 77400 -40980 77520 -40950
rect 77400 -41040 77430 -40980
rect 77430 -41040 77490 -40980
rect 77490 -41040 77520 -40980
rect 77400 -41070 77520 -41040
rect 60747 -41159 60781 -41125
rect 60980 -41159 61015 -41125
rect 61053 -41159 61088 -41125
rect 61129 -41158 61164 -41124
rect 61291 -41159 61325 -41125
rect 77470 -41220 77510 -41180
rect 77790 -41177 77793 -41150
rect 77793 -41177 77827 -41150
rect 77827 -41177 77830 -41150
rect 77790 -41190 77830 -41177
rect 60486 -41300 60526 -41260
rect 60626 -41300 60666 -41260
rect 60766 -41300 60806 -41260
rect 60906 -41300 60946 -41260
rect 59476 -41457 59483 -41423
rect 59483 -41457 59641 -41423
rect 59641 -41457 59646 -41423
rect 78070 -41143 78110 -41090
rect 78070 -41177 78073 -41143
rect 78073 -41177 78107 -41143
rect 78107 -41177 78110 -41143
rect 78070 -41180 78110 -41177
rect 78570 -41100 78640 -41030
rect 78190 -41143 78280 -41140
rect 78190 -41177 78199 -41143
rect 78199 -41177 78233 -41143
rect 78233 -41177 78280 -41143
rect 78190 -41230 78280 -41177
rect 78360 -41143 78400 -41140
rect 78360 -41177 78375 -41143
rect 78375 -41177 78400 -41143
rect 78360 -41180 78400 -41177
rect 78570 -41240 78640 -41170
rect 78570 -41380 78640 -41310
rect 59476 -41460 59646 -41457
rect 59766 -41522 59806 -41520
rect 58926 -41736 58966 -41710
rect 59766 -41700 59772 -41522
rect 59772 -41700 59806 -41522
rect 77607 -41489 77641 -41455
rect 77699 -41489 77733 -41455
rect 77791 -41489 77825 -41455
rect 77883 -41489 77917 -41455
rect 77975 -41489 78009 -41455
rect 78067 -41489 78101 -41455
rect 78159 -41489 78193 -41455
rect 78251 -41489 78285 -41455
rect 78343 -41489 78377 -41455
rect 78435 -41489 78469 -41455
rect 78527 -41489 78561 -41455
rect 59958 -41574 60334 -41540
rect 59874 -41628 59908 -41594
rect 60384 -41628 60418 -41594
rect 59958 -41682 60334 -41648
rect 57125 -41943 57159 -41909
rect 57217 -41943 57251 -41909
rect 57309 -41943 57343 -41909
rect 54081 -42178 54857 -42144
rect 53988 -42244 54022 -42206
rect 54916 -42244 54950 -42206
rect 54081 -42306 54857 -42272
rect 56020 -42208 56080 -42058
rect 58926 -42022 58930 -41736
rect 58930 -42022 58964 -41736
rect 58964 -42022 58966 -41736
rect 59656 -41736 59706 -41730
rect 59125 -41788 59501 -41754
rect 59560 -41842 59594 -41808
rect 59125 -41896 59501 -41862
rect 59032 -41950 59066 -41916
rect 59125 -42004 59501 -41970
rect 57156 -42090 57316 -42060
rect 57156 -42190 57186 -42090
rect 57186 -42190 57286 -42090
rect 57286 -42190 57316 -42090
rect 58926 -42100 58966 -42022
rect 59656 -42022 59662 -41736
rect 59662 -42022 59696 -41736
rect 59696 -42022 59706 -41736
rect 78630 -41490 78740 -41460
rect 77607 -41565 77641 -41531
rect 77699 -41565 77733 -41531
rect 77791 -41565 77825 -41531
rect 77883 -41565 77917 -41531
rect 77975 -41565 78009 -41531
rect 78630 -41540 78660 -41490
rect 78660 -41540 78710 -41490
rect 78710 -41540 78740 -41490
rect 78630 -41570 78740 -41540
rect 78850 -41490 78960 -41460
rect 78850 -41540 78880 -41490
rect 78880 -41540 78930 -41490
rect 78930 -41540 78960 -41490
rect 78850 -41570 78960 -41540
rect 79090 -41490 79200 -41460
rect 79090 -41540 79120 -41490
rect 79120 -41540 79170 -41490
rect 79170 -41540 79200 -41490
rect 79090 -41570 79200 -41540
rect 59866 -41762 60426 -41760
rect 59866 -41796 59868 -41762
rect 59868 -41796 60424 -41762
rect 60424 -41796 60426 -41762
rect 59866 -41800 60426 -41796
rect 77510 -41840 77560 -41790
rect 77980 -41780 78020 -41740
rect 77790 -41843 77830 -41830
rect 77790 -41870 77793 -41843
rect 77793 -41870 77827 -41843
rect 77827 -41870 77830 -41843
rect 77980 -41900 78020 -41860
rect 59656 -42030 59706 -42022
rect 77420 -41990 77540 -41960
rect 77420 -42050 77450 -41990
rect 77450 -42050 77510 -41990
rect 77510 -42050 77540 -41990
rect 57156 -42220 57316 -42190
rect 77420 -42160 77540 -42050
rect 77980 -42000 78020 -41960
rect 77607 -42109 77641 -42075
rect 77699 -42109 77733 -42075
rect 77791 -42109 77825 -42075
rect 77883 -42109 77917 -42075
rect 77975 -42109 78009 -42075
rect 77420 -42220 77450 -42160
rect 77450 -42220 77510 -42160
rect 77510 -42220 77540 -42160
rect 77609 -42199 77643 -42165
rect 77701 -42199 77735 -42165
rect 77793 -42199 77827 -42165
rect 77885 -42199 77919 -42165
rect 77977 -42199 78011 -42165
rect 54150 -42420 54840 -42388
rect 77420 -42250 77540 -42220
rect 54150 -42508 54840 -42420
rect 55300 -42392 55476 -42358
rect 55526 -42436 55560 -42402
rect 55300 -42480 55476 -42446
rect 77980 -42380 78020 -42340
rect 55320 -42560 55470 -42548
rect 77490 -42480 77540 -42430
rect 77790 -42431 77795 -42400
rect 77795 -42431 77829 -42400
rect 77829 -42431 77830 -42400
rect 77790 -42440 77830 -42431
rect 55320 -42594 55470 -42560
rect 77980 -42460 78020 -42420
rect 55320 -42608 55470 -42594
rect 77980 -42560 78020 -42520
rect 77980 -42633 78020 -42600
rect 77980 -42640 77981 -42633
rect 77981 -42640 78020 -42633
rect 77609 -42743 77643 -42709
rect 77701 -42743 77735 -42709
rect 77793 -42743 77827 -42709
rect 77885 -42743 77919 -42709
rect 77977 -42743 78011 -42709
rect 78940 -42740 79050 -42710
rect 77607 -42815 77641 -42781
rect 77699 -42815 77733 -42781
rect 77791 -42815 77825 -42781
rect 77883 -42815 77917 -42781
rect 77975 -42815 78009 -42781
rect 78067 -42815 78101 -42781
rect 78159 -42815 78193 -42781
rect 78351 -42815 78385 -42781
rect 78443 -42815 78477 -42781
rect 78535 -42815 78569 -42781
rect 78627 -42815 78661 -42781
rect 78719 -42815 78753 -42781
rect 78811 -42815 78845 -42781
rect 78940 -42790 78970 -42740
rect 78970 -42790 79020 -42740
rect 79020 -42790 79050 -42740
rect 77580 -42990 77630 -42940
rect 78940 -42820 79050 -42790
rect 79130 -42740 79240 -42710
rect 79130 -42790 79160 -42740
rect 79160 -42790 79210 -42740
rect 79210 -42790 79240 -42740
rect 79130 -42820 79240 -42790
rect 78250 -42923 78290 -42889
rect 77410 -43240 77530 -43210
rect 78170 -43027 78187 -43010
rect 78187 -43027 78220 -43010
rect 77410 -43300 77440 -43240
rect 77440 -43300 77500 -43240
rect 77500 -43300 77530 -43240
rect 77770 -43093 77810 -43090
rect 77770 -43127 77789 -43093
rect 77789 -43127 77810 -43093
rect 77770 -43130 77810 -43127
rect 77870 -43127 77895 -43120
rect 77895 -43127 77910 -43120
rect 77870 -43160 77910 -43127
rect 77870 -43240 77910 -43200
rect 77970 -43250 78010 -43210
rect 78170 -43180 78220 -43027
rect 78850 -42970 78900 -42920
rect 78350 -43180 78400 -43140
rect 78470 -43090 78560 -43040
rect 78640 -43093 78690 -43090
rect 78640 -43127 78659 -43093
rect 78659 -43127 78690 -43093
rect 78640 -43130 78690 -43127
rect 78850 -43090 78900 -43040
rect 77410 -43330 77530 -43300
rect 78850 -43210 78900 -43160
rect 77607 -43359 77641 -43325
rect 77699 -43359 77733 -43325
rect 77791 -43359 77825 -43325
rect 77883 -43359 77917 -43325
rect 77975 -43359 78009 -43325
rect 78067 -43359 78101 -43325
rect 78159 -43359 78193 -43325
rect 78351 -43359 78385 -43325
rect 78443 -43359 78477 -43325
rect 78535 -43359 78569 -43325
rect 78627 -43359 78661 -43325
rect 78719 -43359 78753 -43325
rect 78811 -43359 78845 -43325
rect 77410 -43420 77530 -43390
rect 77410 -43480 77440 -43420
rect 77440 -43480 77500 -43420
rect 77500 -43480 77530 -43420
rect 77607 -43431 77641 -43397
rect 77699 -43431 77733 -43397
rect 77791 -43431 77825 -43397
rect 77883 -43431 77917 -43397
rect 77975 -43431 78009 -43397
rect 78067 -43431 78101 -43397
rect 78159 -43431 78193 -43397
rect 83450 -43410 83620 -43380
rect 77410 -43510 77530 -43480
rect 25700 -45328 25736 -43892
rect 25736 -45328 25770 -43892
rect 25770 -45328 25780 -43892
rect 77770 -43560 77810 -43520
rect 77770 -43629 77810 -43610
rect 77770 -43650 77789 -43629
rect 77789 -43650 77810 -43629
rect 77870 -43580 77910 -43540
rect 77870 -43629 77910 -43620
rect 77870 -43660 77895 -43629
rect 77895 -43660 77910 -43629
rect 78200 -43560 78280 -43510
rect 83450 -43520 83480 -43410
rect 83480 -43520 83590 -43410
rect 83590 -43520 83620 -43410
rect 83450 -43550 83620 -43520
rect 85150 -43410 85320 -43380
rect 85150 -43520 85180 -43410
rect 85180 -43520 85290 -43410
rect 85290 -43520 85320 -43410
rect 85150 -43550 85320 -43520
rect 86530 -43410 86700 -43380
rect 86530 -43520 86560 -43410
rect 86560 -43520 86670 -43410
rect 86670 -43520 86700 -43410
rect 86530 -43550 86700 -43520
rect 87820 -43410 87990 -43380
rect 87820 -43520 87850 -43410
rect 87850 -43520 87960 -43410
rect 87960 -43520 87990 -43410
rect 87820 -43550 87990 -43520
rect 89340 -43410 89510 -43380
rect 89340 -43520 89370 -43410
rect 89370 -43520 89480 -43410
rect 89480 -43520 89510 -43410
rect 89340 -43550 89510 -43520
rect 90750 -43410 90920 -43380
rect 90750 -43520 90780 -43410
rect 90780 -43520 90890 -43410
rect 90890 -43520 90920 -43410
rect 90750 -43550 90920 -43520
rect 77970 -43663 77991 -43630
rect 77991 -43663 78010 -43630
rect 77970 -43670 78010 -43663
rect 82867 -43625 82901 -43591
rect 82959 -43625 82993 -43591
rect 83051 -43625 83085 -43591
rect 83143 -43625 83177 -43591
rect 83235 -43625 83269 -43591
rect 83327 -43625 83361 -43591
rect 83419 -43625 83453 -43591
rect 83511 -43625 83545 -43591
rect 83603 -43625 83637 -43591
rect 83695 -43625 83729 -43591
rect 83787 -43625 83821 -43591
rect 83879 -43625 83913 -43591
rect 83971 -43625 84005 -43591
rect 84063 -43625 84097 -43591
rect 84155 -43625 84189 -43591
rect 84247 -43625 84281 -43591
rect 84339 -43625 84373 -43591
rect 84431 -43625 84465 -43591
rect 84523 -43625 84557 -43591
rect 84615 -43625 84649 -43591
rect 84707 -43625 84741 -43591
rect 84799 -43625 84833 -43591
rect 84891 -43625 84925 -43591
rect 84983 -43625 85017 -43591
rect 85075 -43625 85109 -43591
rect 85167 -43625 85201 -43591
rect 85259 -43625 85293 -43591
rect 85351 -43625 85385 -43591
rect 85443 -43625 85477 -43591
rect 85535 -43625 85569 -43591
rect 85627 -43625 85661 -43591
rect 85719 -43625 85753 -43591
rect 85811 -43625 85845 -43591
rect 85903 -43625 85937 -43591
rect 85995 -43625 86029 -43591
rect 86087 -43625 86121 -43591
rect 86179 -43625 86213 -43591
rect 86271 -43625 86305 -43591
rect 86363 -43625 86397 -43591
rect 86455 -43625 86489 -43591
rect 86547 -43625 86581 -43591
rect 86639 -43625 86673 -43591
rect 86731 -43625 86765 -43591
rect 86823 -43625 86857 -43591
rect 86915 -43625 86949 -43591
rect 87007 -43625 87041 -43591
rect 87099 -43625 87133 -43591
rect 87191 -43625 87225 -43591
rect 87283 -43625 87317 -43591
rect 87375 -43625 87409 -43591
rect 87467 -43625 87501 -43591
rect 87559 -43625 87593 -43591
rect 87651 -43625 87685 -43591
rect 87743 -43625 87777 -43591
rect 87835 -43625 87869 -43591
rect 87927 -43625 87961 -43591
rect 88019 -43625 88053 -43591
rect 88111 -43625 88145 -43591
rect 88203 -43625 88237 -43591
rect 88295 -43625 88329 -43591
rect 88387 -43625 88421 -43591
rect 88479 -43625 88513 -43591
rect 88571 -43625 88605 -43591
rect 88663 -43625 88697 -43591
rect 88755 -43625 88789 -43591
rect 88847 -43625 88881 -43591
rect 88939 -43625 88973 -43591
rect 89031 -43625 89065 -43591
rect 89123 -43625 89157 -43591
rect 89215 -43625 89249 -43591
rect 89307 -43625 89341 -43591
rect 89399 -43625 89433 -43591
rect 89491 -43625 89525 -43591
rect 89583 -43625 89617 -43591
rect 89675 -43625 89709 -43591
rect 89767 -43625 89801 -43591
rect 89859 -43625 89893 -43591
rect 89951 -43625 89985 -43591
rect 90043 -43625 90077 -43591
rect 90135 -43625 90169 -43591
rect 90227 -43625 90261 -43591
rect 90319 -43625 90353 -43591
rect 90411 -43625 90445 -43591
rect 90503 -43625 90537 -43591
rect 90595 -43625 90629 -43591
rect 90687 -43625 90721 -43591
rect 90779 -43625 90813 -43591
rect 90871 -43625 90905 -43591
rect 90963 -43625 90997 -43591
rect 91055 -43625 91089 -43591
rect 91147 -43625 91181 -43591
rect 91239 -43625 91273 -43591
rect 91331 -43625 91365 -43591
rect 78200 -43700 78280 -43650
rect 77440 -43820 77490 -43770
rect 25882 -44341 26996 -43944
rect 27124 -44341 28238 -43944
rect 28366 -44341 29480 -43944
rect 29608 -44341 30722 -43944
rect 30850 -44341 31964 -43944
rect 32092 -44341 33206 -43944
rect 33334 -44341 34448 -43944
rect 34576 -44341 35690 -43944
rect 25882 -45276 26996 -44879
rect 27124 -45276 28238 -44879
rect 28366 -45276 29480 -44879
rect 29608 -45276 30722 -44879
rect 30850 -45276 31964 -44879
rect 32092 -45276 33206 -44879
rect 33334 -45276 34448 -44879
rect 34576 -45276 35690 -44879
rect 25700 -45490 25780 -45328
rect 78200 -43840 78280 -43790
rect 77607 -43975 77641 -43941
rect 77699 -43975 77733 -43941
rect 77791 -43975 77825 -43941
rect 77883 -43975 77917 -43941
rect 77975 -43975 78009 -43941
rect 78067 -43975 78101 -43941
rect 78159 -43975 78193 -43941
rect 78280 -43970 78390 -43940
rect 77607 -44047 77641 -44013
rect 77699 -44047 77733 -44013
rect 77791 -44047 77825 -44013
rect 77883 -44047 77917 -44013
rect 77975 -44047 78009 -44013
rect 78067 -44047 78101 -44013
rect 78159 -44047 78193 -44013
rect 78280 -44020 78310 -43970
rect 78310 -44020 78360 -43970
rect 78360 -44020 78390 -43970
rect 77470 -44220 77510 -44170
rect 78280 -44050 78390 -44020
rect 78580 -43970 78690 -43940
rect 78580 -44020 78610 -43970
rect 78610 -44020 78660 -43970
rect 78660 -44020 78690 -43970
rect 78580 -44050 78690 -44020
rect 78880 -43970 78990 -43940
rect 78880 -44020 78910 -43970
rect 78910 -44020 78960 -43970
rect 78960 -44020 78990 -43970
rect 82880 -43903 82930 -43900
rect 82880 -43937 82904 -43903
rect 82904 -43937 82930 -43903
rect 82880 -43990 82930 -43937
rect 78880 -44050 78990 -44020
rect 83050 -43937 83074 -43910
rect 83074 -43937 83090 -43910
rect 83050 -43990 83090 -43937
rect 85330 -43839 85342 -43820
rect 85342 -43839 85376 -43820
rect 85376 -43839 85380 -43820
rect 85330 -43990 85380 -43839
rect 86810 -43805 86860 -43800
rect 86810 -43839 86814 -43805
rect 86814 -43839 86848 -43805
rect 86848 -43839 86860 -43805
rect 85610 -43903 86471 -43897
rect 85610 -43931 85722 -43903
rect 85722 -43931 85756 -43903
rect 85756 -43931 85890 -43903
rect 85890 -43931 85924 -43903
rect 85924 -43931 86059 -43903
rect 86059 -43931 86093 -43903
rect 86093 -43931 86226 -43903
rect 86226 -43931 86260 -43903
rect 86260 -43931 86394 -43903
rect 86394 -43931 86428 -43903
rect 86428 -43931 86471 -43903
rect 86810 -43990 86860 -43839
rect 88280 -43839 88286 -43810
rect 88286 -43839 88320 -43810
rect 88320 -43839 88330 -43810
rect 87044 -43903 87905 -43896
rect 87044 -43930 87054 -43903
rect 87054 -43930 87194 -43903
rect 87194 -43930 87228 -43903
rect 87228 -43930 87362 -43903
rect 87362 -43930 87396 -43903
rect 87396 -43930 87531 -43903
rect 87531 -43930 87565 -43903
rect 87565 -43930 87698 -43903
rect 87698 -43930 87732 -43903
rect 87732 -43930 87866 -43903
rect 87866 -43930 87900 -43903
rect 87900 -43930 87905 -43903
rect 88280 -43990 88330 -43839
rect 89750 -43839 89758 -43810
rect 89758 -43839 89792 -43810
rect 89792 -43839 89800 -43810
rect 88523 -43903 89384 -43896
rect 88523 -43930 88526 -43903
rect 88526 -43930 88666 -43903
rect 88666 -43930 88700 -43903
rect 88700 -43930 88834 -43903
rect 88834 -43930 88868 -43903
rect 88868 -43930 89003 -43903
rect 89003 -43930 89037 -43903
rect 89037 -43930 89170 -43903
rect 89170 -43930 89204 -43903
rect 89204 -43930 89338 -43903
rect 89338 -43930 89372 -43903
rect 89372 -43930 89384 -43903
rect 89750 -43991 89800 -43839
rect 89750 -44000 89758 -43991
rect 89758 -44000 89792 -43991
rect 89792 -44000 89800 -43991
rect 91220 -43839 91230 -43810
rect 91230 -43839 91264 -43810
rect 91264 -43839 91270 -43810
rect 89980 -43899 90747 -43897
rect 89978 -43903 90748 -43899
rect 89978 -43933 89998 -43903
rect 89998 -43933 90138 -43903
rect 90138 -43933 90172 -43903
rect 90172 -43933 90306 -43903
rect 90306 -43933 90340 -43903
rect 90340 -43933 90475 -43903
rect 90475 -43933 90509 -43903
rect 90509 -43933 90642 -43903
rect 90642 -43933 90676 -43903
rect 90676 -43933 90748 -43903
rect 91220 -43991 91270 -43839
rect 91220 -44000 91230 -43991
rect 91230 -44000 91264 -43991
rect 91264 -44000 91270 -43991
rect 78180 -44157 78290 -44140
rect 78180 -44191 78187 -44157
rect 78187 -44191 78290 -44157
rect 78180 -44225 78290 -44191
rect 77400 -44410 77520 -44380
rect 77400 -44470 77430 -44410
rect 77430 -44470 77490 -44410
rect 77490 -44470 77520 -44410
rect 78180 -44259 78187 -44225
rect 78187 -44259 78290 -44225
rect 77400 -44500 77520 -44470
rect 77770 -44480 77810 -44440
rect 77870 -44325 77910 -44320
rect 77870 -44359 77895 -44325
rect 77895 -44359 77910 -44325
rect 77870 -44360 77910 -44359
rect 77870 -44470 77910 -44410
rect 77970 -44460 78010 -44360
rect 78180 -44413 78290 -44259
rect 78180 -44447 78187 -44413
rect 78187 -44447 78290 -44413
rect 78180 -44460 78290 -44447
rect 82867 -44169 82901 -44135
rect 82959 -44169 82993 -44135
rect 83051 -44169 83085 -44135
rect 83143 -44169 83177 -44135
rect 83235 -44169 83269 -44135
rect 83327 -44169 83361 -44135
rect 83419 -44169 83453 -44135
rect 83511 -44169 83545 -44135
rect 83603 -44169 83637 -44135
rect 83695 -44169 83729 -44135
rect 83787 -44169 83821 -44135
rect 83879 -44169 83913 -44135
rect 83971 -44169 84005 -44135
rect 84063 -44169 84097 -44135
rect 84155 -44169 84189 -44135
rect 84247 -44169 84281 -44135
rect 84339 -44169 84373 -44135
rect 84431 -44169 84465 -44135
rect 84523 -44169 84557 -44135
rect 84615 -44169 84649 -44135
rect 84707 -44169 84741 -44135
rect 84799 -44169 84833 -44135
rect 84891 -44169 84925 -44135
rect 84983 -44169 85017 -44135
rect 85075 -44169 85109 -44135
rect 85167 -44169 85201 -44135
rect 85259 -44169 85293 -44135
rect 85351 -44169 85385 -44135
rect 85443 -44169 85477 -44135
rect 85535 -44169 85569 -44135
rect 85627 -44169 85661 -44135
rect 85719 -44169 85753 -44135
rect 85811 -44169 85845 -44135
rect 85903 -44169 85937 -44135
rect 85995 -44169 86029 -44135
rect 86087 -44169 86121 -44135
rect 86179 -44169 86213 -44135
rect 86271 -44169 86305 -44135
rect 86363 -44169 86397 -44135
rect 86455 -44169 86489 -44135
rect 86547 -44169 86581 -44135
rect 86639 -44169 86673 -44135
rect 86731 -44169 86765 -44135
rect 86823 -44169 86857 -44135
rect 86915 -44169 86949 -44135
rect 87007 -44169 87041 -44135
rect 87099 -44169 87133 -44135
rect 87191 -44169 87225 -44135
rect 87283 -44169 87317 -44135
rect 87375 -44169 87409 -44135
rect 87467 -44169 87501 -44135
rect 87559 -44169 87593 -44135
rect 87651 -44169 87685 -44135
rect 87743 -44169 87777 -44135
rect 87835 -44169 87869 -44135
rect 87927 -44169 87961 -44135
rect 88019 -44169 88053 -44135
rect 88111 -44169 88145 -44135
rect 88203 -44169 88237 -44135
rect 88295 -44169 88329 -44135
rect 88387 -44169 88421 -44135
rect 88479 -44169 88513 -44135
rect 88571 -44169 88605 -44135
rect 88663 -44169 88697 -44135
rect 88755 -44169 88789 -44135
rect 88847 -44169 88881 -44135
rect 88939 -44169 88973 -44135
rect 89031 -44169 89065 -44135
rect 89123 -44169 89157 -44135
rect 89215 -44169 89249 -44135
rect 89307 -44169 89341 -44135
rect 89399 -44169 89433 -44135
rect 89491 -44169 89525 -44135
rect 89583 -44169 89617 -44135
rect 89675 -44169 89709 -44135
rect 89767 -44169 89801 -44135
rect 89859 -44169 89893 -44135
rect 89951 -44169 89985 -44135
rect 90043 -44169 90077 -44135
rect 90135 -44169 90169 -44135
rect 90227 -44169 90261 -44135
rect 90319 -44169 90353 -44135
rect 90411 -44169 90445 -44135
rect 90503 -44169 90537 -44135
rect 90595 -44169 90629 -44135
rect 90687 -44169 90721 -44135
rect 90779 -44169 90813 -44135
rect 90871 -44169 90905 -44135
rect 90963 -44169 90997 -44135
rect 91055 -44169 91089 -44135
rect 91147 -44169 91181 -44135
rect 91239 -44169 91273 -44135
rect 91331 -44169 91365 -44135
rect 83480 -44240 83650 -44210
rect 83480 -44350 83510 -44240
rect 83510 -44350 83620 -44240
rect 83620 -44350 83650 -44240
rect 83480 -44380 83650 -44350
rect 85120 -44250 85290 -44220
rect 85120 -44360 85150 -44250
rect 85150 -44360 85260 -44250
rect 85260 -44360 85290 -44250
rect 85120 -44390 85290 -44360
rect 86530 -44240 86700 -44210
rect 86530 -44350 86560 -44240
rect 86560 -44350 86670 -44240
rect 86670 -44350 86700 -44240
rect 86530 -44380 86700 -44350
rect 87910 -44240 88080 -44210
rect 87910 -44350 87940 -44240
rect 87940 -44350 88050 -44240
rect 88050 -44350 88080 -44240
rect 87910 -44380 88080 -44350
rect 89450 -44250 89620 -44220
rect 89450 -44360 89480 -44250
rect 89480 -44360 89590 -44250
rect 89590 -44360 89620 -44250
rect 89450 -44390 89620 -44360
rect 90730 -44250 90900 -44220
rect 90730 -44360 90760 -44250
rect 90760 -44360 90870 -44250
rect 90870 -44360 90900 -44250
rect 90730 -44390 90900 -44360
rect 77607 -44591 77641 -44557
rect 77699 -44591 77733 -44557
rect 77791 -44591 77825 -44557
rect 77883 -44591 77917 -44557
rect 77975 -44591 78009 -44557
rect 78067 -44591 78101 -44557
rect 78159 -44591 78193 -44557
rect 77400 -44660 77520 -44630
rect 54150 -44758 54850 -44708
rect 77400 -44720 77430 -44660
rect 77430 -44720 77490 -44660
rect 77490 -44720 77520 -44660
rect 77607 -44665 77641 -44631
rect 77699 -44665 77733 -44631
rect 77791 -44665 77825 -44631
rect 77883 -44665 77917 -44631
rect 77975 -44665 78009 -44631
rect 78067 -44665 78101 -44631
rect 78159 -44665 78193 -44631
rect 77400 -44750 77520 -44720
rect 54150 -44792 54850 -44758
rect 54150 -44798 54850 -44792
rect 54091 -44906 54867 -44872
rect 53998 -44972 54032 -44934
rect 54926 -44972 54960 -44934
rect 54091 -45034 54867 -45000
rect 55960 -45098 56040 -44928
rect 77580 -45040 77630 -44950
rect 77770 -44780 77810 -44740
rect 77870 -44863 77910 -44850
rect 77870 -44890 77895 -44863
rect 77895 -44890 77910 -44863
rect 77960 -44863 78010 -44860
rect 77960 -44897 77991 -44863
rect 77991 -44897 78010 -44863
rect 77960 -44910 78010 -44897
rect 53526 -45340 53614 -45306
rect 25700 -46926 25736 -45490
rect 25736 -46926 25770 -45490
rect 25770 -46926 25780 -45490
rect 25882 -45939 26996 -45542
rect 27124 -45939 28238 -45542
rect 28366 -45939 29480 -45542
rect 29608 -45939 30722 -45542
rect 30850 -45939 31964 -45542
rect 32092 -45939 33206 -45542
rect 33334 -45939 34448 -45542
rect 34576 -45939 35690 -45542
rect 25882 -46874 26996 -46477
rect 27124 -46874 28238 -46477
rect 28366 -46874 29480 -46477
rect 29608 -46874 30722 -46477
rect 30850 -46874 31964 -46477
rect 32092 -46874 33206 -46477
rect 33334 -46874 34448 -46477
rect 34576 -46874 35690 -46477
rect 25700 -47084 25780 -46926
rect 53330 -46718 53350 -45368
rect 53350 -46718 53384 -45368
rect 53384 -46718 53400 -45368
rect 53464 -46166 53498 -45390
rect 53642 -46166 53676 -45390
rect 57126 -45100 57356 -45070
rect 54091 -45262 54867 -45228
rect 53998 -45328 54032 -45290
rect 54926 -45328 54960 -45290
rect 54091 -45390 54867 -45356
rect 55334 -45402 55368 -45368
rect 55290 -45628 55324 -45452
rect 55378 -45628 55412 -45452
rect 55142 -45908 55494 -45874
rect 53942 -46012 54718 -45978
rect 53858 -46128 53892 -46040
rect 54768 -46128 54802 -46040
rect 53942 -46190 54718 -46156
rect 53526 -46250 53614 -46216
rect 55046 -45994 55080 -45960
rect 55556 -45994 55590 -45960
rect 55142 -46080 55494 -46046
rect 57126 -45170 57156 -45100
rect 57156 -45170 57316 -45100
rect 57316 -45170 57356 -45100
rect 57126 -45200 57356 -45170
rect 58926 -45229 58966 -45220
rect 55882 -45290 55970 -45256
rect 55820 -46116 55854 -45340
rect 55998 -46116 56032 -45340
rect 55882 -46200 55970 -46166
rect 57125 -45279 57159 -45245
rect 57217 -45279 57251 -45245
rect 57309 -45279 57343 -45245
rect 57118 -45557 57178 -45544
rect 57118 -45591 57133 -45557
rect 57133 -45591 57167 -45557
rect 57167 -45591 57178 -45557
rect 57118 -45594 57178 -45591
rect 58926 -45515 58930 -45229
rect 58930 -45515 58964 -45229
rect 58964 -45515 58966 -45229
rect 78190 -45080 78260 -44950
rect 77607 -45209 77641 -45175
rect 77699 -45209 77733 -45175
rect 77791 -45209 77825 -45175
rect 77883 -45209 77917 -45175
rect 77975 -45209 78009 -45175
rect 78067 -45209 78101 -45175
rect 78159 -45209 78193 -45175
rect 59125 -45281 59501 -45247
rect 59560 -45335 59594 -45301
rect 59125 -45389 59501 -45355
rect 59032 -45443 59066 -45409
rect 59125 -45497 59501 -45463
rect 58926 -45520 58966 -45515
rect 59656 -45515 59662 -45230
rect 59662 -45515 59696 -45230
rect 79120 -45210 79230 -45180
rect 77607 -45285 77641 -45251
rect 77699 -45285 77733 -45251
rect 77791 -45285 77825 -45251
rect 77883 -45285 77917 -45251
rect 77975 -45285 78009 -45251
rect 78067 -45285 78101 -45251
rect 78159 -45285 78193 -45251
rect 78251 -45285 78285 -45251
rect 78343 -45285 78377 -45251
rect 78435 -45285 78469 -45251
rect 78527 -45285 78561 -45251
rect 78619 -45285 78653 -45251
rect 78711 -45285 78745 -45251
rect 78803 -45285 78837 -45251
rect 78895 -45285 78929 -45251
rect 78987 -45285 79021 -45251
rect 79120 -45260 79150 -45210
rect 79150 -45260 79200 -45210
rect 79200 -45260 79230 -45210
rect 77770 -45370 77785 -45352
rect 77785 -45370 77830 -45352
rect 77770 -45392 77830 -45370
rect 59656 -45520 59696 -45515
rect 57326 -45580 57366 -45540
rect 53526 -46358 53614 -46324
rect 55030 -46328 55110 -46248
rect 55740 -46268 55810 -46248
rect 55740 -46302 55802 -46268
rect 55802 -46302 55810 -46268
rect 55740 -46328 55810 -46302
rect 25700 -48520 25736 -47084
rect 25736 -48520 25770 -47084
rect 25770 -48520 25780 -47084
rect 25882 -47533 26996 -47136
rect 27124 -47533 28238 -47136
rect 28366 -47533 29480 -47136
rect 29608 -47533 30722 -47136
rect 30850 -47533 31964 -47136
rect 32092 -47533 33206 -47136
rect 33334 -47533 34448 -47136
rect 34576 -47533 35690 -47136
rect 25882 -48468 26996 -48071
rect 27124 -48468 28238 -48071
rect 28366 -48468 29480 -48071
rect 29608 -48468 30722 -48071
rect 30850 -48468 31964 -48071
rect 32092 -48468 33206 -48071
rect 33334 -48468 34448 -48071
rect 34576 -48468 35690 -48071
rect 25700 -48682 25780 -48520
rect 53464 -47184 53498 -46408
rect 53642 -47184 53676 -46408
rect 53942 -46418 54718 -46384
rect 53858 -46534 53892 -46446
rect 54768 -46534 54802 -46446
rect 53942 -46596 54718 -46562
rect 55142 -46530 55494 -46496
rect 55046 -46616 55080 -46582
rect 55556 -46616 55590 -46582
rect 55142 -46702 55494 -46668
rect 53526 -47268 53614 -47234
rect 54081 -47222 54857 -47188
rect 53988 -47288 54022 -47250
rect 54916 -47288 54950 -47250
rect 54081 -47350 54857 -47316
rect 55280 -47124 55314 -46948
rect 55368 -47124 55402 -46948
rect 55324 -47208 55358 -47174
rect 56280 -45800 56350 -45718
rect 56280 -46348 56316 -45800
rect 56316 -46348 56350 -45800
rect 59866 -45494 59868 -45460
rect 59868 -45494 60424 -45460
rect 60424 -45494 60426 -45460
rect 59866 -45500 60426 -45494
rect 59766 -45556 59806 -45550
rect 59103 -45712 59137 -45678
rect 56492 -45840 56530 -45806
rect 55882 -46404 55970 -46370
rect 55820 -47230 55854 -46454
rect 55998 -47230 56032 -46454
rect 55882 -47314 55970 -47280
rect 56430 -46675 56464 -45899
rect 56558 -46675 56592 -45899
rect 56492 -46768 56530 -46734
rect 57125 -45823 57159 -45789
rect 57217 -45823 57251 -45789
rect 57309 -45823 57343 -45789
rect 57086 -45910 57376 -45880
rect 57086 -45980 57116 -45910
rect 57116 -45980 57346 -45910
rect 57346 -45980 57376 -45910
rect 57086 -46010 57376 -45980
rect 58926 -46246 58930 -45760
rect 58930 -46246 58964 -45760
rect 58964 -46246 58966 -45760
rect 59044 -46147 59078 -45771
rect 59162 -46147 59196 -45771
rect 59103 -46240 59137 -46206
rect 58926 -46402 58966 -46246
rect 59766 -45734 59772 -45556
rect 59772 -45734 59806 -45556
rect 59958 -45608 60334 -45574
rect 59874 -45662 59908 -45628
rect 60384 -45662 60418 -45628
rect 59958 -45716 60334 -45682
rect 59766 -45740 59806 -45734
rect 59476 -45796 59656 -45790
rect 77390 -45660 77510 -45630
rect 77390 -45720 77420 -45660
rect 77420 -45720 77480 -45660
rect 77480 -45720 77510 -45660
rect 77620 -45643 77647 -45620
rect 77647 -45643 77690 -45620
rect 77620 -45670 77690 -45643
rect 77390 -45750 77510 -45720
rect 77820 -45603 77823 -45590
rect 77823 -45603 77857 -45590
rect 77857 -45603 77860 -45590
rect 77820 -45640 77860 -45603
rect 79120 -45290 79230 -45260
rect 78080 -45563 78130 -45490
rect 78080 -45580 78112 -45563
rect 78112 -45580 78130 -45563
rect 78250 -45563 78290 -45550
rect 78250 -45590 78253 -45563
rect 78253 -45590 78287 -45563
rect 78287 -45590 78290 -45563
rect 77990 -45693 78030 -45680
rect 77990 -45720 78003 -45693
rect 78003 -45720 78030 -45693
rect 78530 -45563 78570 -45560
rect 78530 -45597 78533 -45563
rect 78533 -45597 78567 -45563
rect 78567 -45597 78570 -45563
rect 78530 -45640 78570 -45597
rect 78650 -45563 78730 -45520
rect 78650 -45590 78659 -45563
rect 78659 -45590 78693 -45563
rect 78693 -45590 78730 -45563
rect 78820 -45563 78860 -45560
rect 78820 -45597 78835 -45563
rect 78835 -45597 78860 -45563
rect 78820 -45600 78860 -45597
rect 79020 -45680 79070 -45370
rect 59476 -45830 59484 -45796
rect 59484 -45830 59642 -45796
rect 59642 -45830 59656 -45796
rect 77607 -45829 77641 -45795
rect 77699 -45829 77733 -45795
rect 77791 -45829 77825 -45795
rect 77883 -45829 77917 -45795
rect 77975 -45829 78009 -45795
rect 78067 -45829 78101 -45795
rect 78159 -45829 78193 -45795
rect 78251 -45829 78285 -45795
rect 78343 -45829 78377 -45795
rect 78435 -45829 78469 -45795
rect 78527 -45829 78561 -45795
rect 78619 -45829 78653 -45795
rect 78711 -45829 78745 -45795
rect 78803 -45829 78837 -45795
rect 78895 -45829 78929 -45795
rect 78987 -45829 79021 -45795
rect 59386 -45892 59426 -45890
rect 59386 -46248 59388 -45892
rect 59388 -46248 59422 -45892
rect 59422 -46248 59426 -45892
rect 59546 -45932 59580 -45898
rect 59502 -46158 59536 -45982
rect 59590 -46158 59624 -45982
rect 59546 -46242 59580 -46208
rect 59386 -46250 59426 -46248
rect 59862 -45932 59896 -45898
rect 59818 -46158 59852 -45982
rect 59906 -46158 59940 -45982
rect 59862 -46242 59896 -46208
rect 61196 -46020 61366 -46000
rect 61196 -46060 61216 -46020
rect 61216 -46060 61336 -46020
rect 61336 -46060 61366 -46020
rect 61196 -46080 61366 -46060
rect 57056 -46570 57416 -46540
rect 57056 -46650 57096 -46570
rect 57096 -46650 57376 -46570
rect 57376 -46650 57416 -46570
rect 57056 -46680 57416 -46650
rect 57125 -46799 57159 -46765
rect 57217 -46799 57251 -46765
rect 57309 -46799 57343 -46765
rect 58926 -46890 58930 -46402
rect 58930 -46890 58964 -46402
rect 58964 -46890 58966 -46402
rect 60127 -46191 60161 -46157
rect 60366 -46165 60406 -46160
rect 60366 -46199 60393 -46165
rect 60393 -46199 60406 -46165
rect 60366 -46200 60406 -46199
rect 60127 -46283 60161 -46249
rect 59103 -46442 59137 -46408
rect 59044 -46877 59078 -46501
rect 57118 -46997 57168 -46994
rect 57118 -47031 57133 -46997
rect 57133 -47031 57167 -46997
rect 57167 -47031 57168 -46997
rect 57118 -47044 57168 -47031
rect 57326 -47010 57376 -46970
rect 59162 -46877 59196 -46501
rect 59103 -46970 59137 -46936
rect 59386 -46405 59426 -46400
rect 59386 -46761 59387 -46405
rect 59387 -46761 59421 -46405
rect 59421 -46761 59426 -46405
rect 59545 -46445 59579 -46411
rect 59501 -46671 59535 -46495
rect 59589 -46671 59623 -46495
rect 59545 -46755 59579 -46721
rect 59386 -46770 59426 -46761
rect 59476 -46823 59646 -46820
rect 59861 -46445 59895 -46411
rect 59817 -46671 59851 -46495
rect 59905 -46671 59939 -46495
rect 59861 -46755 59895 -46721
rect 60127 -46375 60161 -46341
rect 60127 -46467 60161 -46433
rect 60671 -46191 60705 -46157
rect 60366 -46257 60406 -46250
rect 60366 -46290 60393 -46257
rect 60393 -46290 60406 -46257
rect 60366 -46341 60406 -46340
rect 60366 -46375 60393 -46341
rect 60393 -46375 60406 -46341
rect 60366 -46380 60406 -46375
rect 60366 -46425 60406 -46420
rect 60366 -46459 60393 -46425
rect 60393 -46459 60406 -46425
rect 60366 -46460 60406 -46459
rect 60671 -46283 60705 -46249
rect 60671 -46375 60705 -46341
rect 60671 -46467 60705 -46433
rect 60127 -46559 60161 -46525
rect 60297 -46559 60331 -46525
rect 60369 -46559 60405 -46525
rect 60449 -46559 60484 -46525
rect 60671 -46559 60705 -46525
rect 60747 -46191 60781 -46157
rect 61046 -46165 61086 -46160
rect 61046 -46199 61059 -46165
rect 61059 -46199 61086 -46165
rect 61046 -46200 61086 -46199
rect 60747 -46283 60781 -46249
rect 60747 -46375 60781 -46341
rect 60747 -46467 60781 -46433
rect 61291 -46191 61325 -46157
rect 61046 -46257 61086 -46250
rect 61046 -46290 61059 -46257
rect 61059 -46290 61086 -46257
rect 61046 -46341 61086 -46340
rect 61046 -46375 61059 -46341
rect 61059 -46375 61086 -46341
rect 61046 -46380 61086 -46375
rect 61046 -46425 61086 -46420
rect 61046 -46459 61059 -46425
rect 61059 -46459 61086 -46425
rect 61046 -46460 61086 -46459
rect 61291 -46283 61325 -46249
rect 61291 -46375 61325 -46341
rect 77110 -46410 77220 -46390
rect 61291 -46467 61325 -46433
rect 75535 -46445 75569 -46411
rect 75627 -46445 75661 -46411
rect 75719 -46445 75753 -46411
rect 75811 -46445 75845 -46411
rect 75903 -46445 75937 -46411
rect 75995 -46445 76029 -46411
rect 76085 -46445 76119 -46411
rect 76177 -46445 76211 -46411
rect 76269 -46445 76303 -46411
rect 76361 -46445 76395 -46411
rect 76453 -46445 76487 -46411
rect 76545 -46445 76579 -46411
rect 76637 -46445 76671 -46411
rect 76729 -46445 76763 -46411
rect 76821 -46445 76855 -46411
rect 60747 -46559 60781 -46525
rect 60980 -46559 61015 -46525
rect 61053 -46559 61088 -46525
rect 61129 -46558 61164 -46524
rect 61291 -46559 61325 -46525
rect 75670 -46559 75704 -46557
rect 75670 -46591 75700 -46559
rect 75700 -46591 75704 -46559
rect 60486 -46700 60526 -46660
rect 60626 -46700 60666 -46660
rect 60766 -46700 60806 -46660
rect 60906 -46700 60946 -46660
rect 75580 -46677 75586 -46650
rect 75586 -46677 75620 -46650
rect 75580 -46690 75620 -46677
rect 75942 -46593 75976 -46560
rect 75942 -46594 75976 -46593
rect 75670 -46683 75704 -46649
rect 75862 -46677 75896 -46643
rect 76217 -46593 76250 -46559
rect 76250 -46593 76251 -46559
rect 75947 -46683 75981 -46649
rect 76128 -46677 76136 -46650
rect 76136 -46677 76162 -46650
rect 76128 -46684 76162 -46677
rect 76492 -46593 76526 -46559
rect 76224 -46684 76258 -46650
rect 76404 -46677 76412 -46649
rect 76412 -46677 76438 -46649
rect 76404 -46683 76438 -46677
rect 77110 -46460 77140 -46410
rect 77140 -46460 77190 -46410
rect 77190 -46460 77220 -46410
rect 76768 -46593 76802 -46561
rect 76768 -46595 76802 -46593
rect 76497 -46683 76531 -46649
rect 76680 -46677 76688 -46649
rect 76688 -46677 76714 -46649
rect 76680 -46683 76714 -46677
rect 77110 -46530 77220 -46460
rect 77110 -46580 77140 -46530
rect 77140 -46580 77190 -46530
rect 77190 -46580 77220 -46530
rect 77110 -46610 77220 -46580
rect 76772 -46684 76806 -46650
rect 59476 -46857 59483 -46823
rect 59483 -46857 59641 -46823
rect 59641 -46857 59646 -46823
rect 59476 -46860 59646 -46857
rect 59766 -46922 59806 -46920
rect 58926 -47136 58966 -47110
rect 59766 -47100 59772 -46922
rect 59772 -47100 59806 -46922
rect 59958 -46974 60334 -46940
rect 59874 -47028 59908 -46994
rect 60384 -47028 60418 -46994
rect 59958 -47082 60334 -47048
rect 57125 -47343 57159 -47309
rect 57217 -47343 57251 -47309
rect 57309 -47343 57343 -47309
rect 54081 -47578 54857 -47544
rect 53988 -47644 54022 -47606
rect 54916 -47644 54950 -47606
rect 54081 -47706 54857 -47672
rect 56020 -47608 56080 -47458
rect 58926 -47422 58930 -47136
rect 58930 -47422 58964 -47136
rect 58964 -47422 58966 -47136
rect 59656 -47136 59706 -47130
rect 59125 -47188 59501 -47154
rect 59560 -47242 59594 -47208
rect 59125 -47296 59501 -47262
rect 59032 -47350 59066 -47316
rect 59125 -47404 59501 -47370
rect 57156 -47490 57316 -47460
rect 57156 -47590 57186 -47490
rect 57186 -47590 57286 -47490
rect 57286 -47590 57316 -47490
rect 58926 -47500 58966 -47422
rect 59656 -47422 59662 -47136
rect 59662 -47422 59696 -47136
rect 59696 -47422 59706 -47136
rect 75670 -46743 75704 -46738
rect 75670 -46772 75700 -46743
rect 75700 -46772 75704 -46743
rect 75943 -46777 75976 -46743
rect 75976 -46777 75977 -46743
rect 76215 -46777 76216 -46744
rect 76216 -46777 76249 -46744
rect 76215 -46778 76249 -46777
rect 76218 -46845 76250 -46816
rect 76250 -46845 76252 -46816
rect 76218 -46850 76252 -46845
rect 76492 -46777 76526 -46743
rect 76768 -46777 76802 -46743
rect 76930 -46870 77040 -46840
rect 76930 -46920 76960 -46870
rect 76960 -46920 77010 -46870
rect 77010 -46920 77040 -46870
rect 75535 -46989 75569 -46955
rect 75627 -46989 75661 -46955
rect 75719 -46989 75753 -46955
rect 75811 -46989 75845 -46955
rect 75903 -46989 75937 -46955
rect 75995 -46989 76029 -46955
rect 76085 -46989 76119 -46955
rect 76177 -46989 76211 -46955
rect 76269 -46989 76303 -46955
rect 76361 -46989 76395 -46955
rect 76453 -46989 76487 -46955
rect 76545 -46989 76579 -46955
rect 76637 -46989 76671 -46955
rect 76729 -46989 76763 -46955
rect 76821 -46989 76855 -46955
rect 76930 -47000 77040 -46920
rect 76930 -47050 76960 -47000
rect 76960 -47050 77010 -47000
rect 77010 -47050 77040 -47000
rect 76930 -47080 77040 -47050
rect 59866 -47162 60426 -47160
rect 77607 -47115 77641 -47081
rect 77699 -47115 77733 -47081
rect 77791 -47115 77825 -47081
rect 77883 -47115 77917 -47081
rect 77975 -47115 78009 -47081
rect 78067 -47115 78101 -47081
rect 78159 -47115 78193 -47081
rect 78251 -47115 78285 -47081
rect 78343 -47115 78377 -47081
rect 78435 -47115 78469 -47081
rect 78527 -47115 78561 -47081
rect 78619 -47115 78653 -47081
rect 78711 -47115 78745 -47081
rect 78803 -47115 78837 -47081
rect 78895 -47115 78929 -47081
rect 78987 -47115 79021 -47081
rect 59866 -47196 59868 -47162
rect 59868 -47196 60424 -47162
rect 60424 -47196 60426 -47162
rect 59866 -47200 60426 -47196
rect 77430 -47210 77520 -47170
rect 77780 -47360 77820 -47320
rect 59656 -47430 59706 -47422
rect 77900 -47393 77940 -47390
rect 77900 -47427 77915 -47393
rect 77915 -47427 77940 -47393
rect 77900 -47430 77940 -47427
rect 77240 -47530 77300 -47490
rect 77420 -47530 77540 -47500
rect 78160 -47393 78200 -47390
rect 78160 -47427 78164 -47393
rect 78164 -47427 78198 -47393
rect 78198 -47427 78200 -47393
rect 78160 -47430 78200 -47427
rect 78290 -47430 78330 -47390
rect 78370 -47393 78410 -47390
rect 78370 -47427 78374 -47393
rect 78374 -47427 78408 -47393
rect 78408 -47427 78410 -47393
rect 78370 -47430 78410 -47427
rect 78590 -47410 78630 -47370
rect 78800 -47393 78850 -47380
rect 78800 -47420 78805 -47393
rect 78805 -47420 78839 -47393
rect 78839 -47420 78850 -47393
rect 57156 -47620 57316 -47590
rect 77420 -47590 77450 -47530
rect 77450 -47590 77510 -47530
rect 77510 -47590 77540 -47530
rect 77420 -47620 77540 -47590
rect 79080 -47440 79140 -47380
rect 79080 -47550 79140 -47490
rect 83454 -47548 83624 -47518
rect 54150 -47820 54840 -47788
rect 77607 -47659 77641 -47625
rect 77699 -47659 77733 -47625
rect 77791 -47659 77825 -47625
rect 77883 -47659 77917 -47625
rect 77975 -47659 78009 -47625
rect 78067 -47659 78101 -47625
rect 78159 -47659 78193 -47625
rect 78251 -47659 78285 -47625
rect 78343 -47659 78377 -47625
rect 78435 -47659 78469 -47625
rect 78527 -47659 78561 -47625
rect 78619 -47659 78653 -47625
rect 78711 -47659 78745 -47625
rect 78803 -47659 78837 -47625
rect 78895 -47659 78929 -47625
rect 78987 -47659 79021 -47625
rect 83454 -47658 83484 -47548
rect 83484 -47658 83594 -47548
rect 83594 -47658 83624 -47548
rect 54150 -47908 54840 -47820
rect 83454 -47688 83624 -47658
rect 85154 -47548 85324 -47518
rect 85154 -47658 85184 -47548
rect 85184 -47658 85294 -47548
rect 85294 -47658 85324 -47548
rect 85154 -47688 85324 -47658
rect 86534 -47548 86704 -47518
rect 86534 -47658 86564 -47548
rect 86564 -47658 86674 -47548
rect 86674 -47658 86704 -47548
rect 86534 -47688 86704 -47658
rect 87824 -47548 87994 -47518
rect 87824 -47658 87854 -47548
rect 87854 -47658 87964 -47548
rect 87964 -47658 87994 -47548
rect 87824 -47688 87994 -47658
rect 89344 -47548 89514 -47518
rect 89344 -47658 89374 -47548
rect 89374 -47658 89484 -47548
rect 89484 -47658 89514 -47548
rect 89344 -47688 89514 -47658
rect 90754 -47548 90924 -47518
rect 90754 -47658 90784 -47548
rect 90784 -47658 90894 -47548
rect 90894 -47658 90924 -47548
rect 90754 -47688 90924 -47658
rect 55300 -47792 55476 -47758
rect 55526 -47836 55560 -47802
rect 55300 -47880 55476 -47846
rect 77420 -47730 77540 -47700
rect 77420 -47790 77450 -47730
rect 77450 -47790 77510 -47730
rect 77510 -47790 77540 -47730
rect 77607 -47745 77641 -47711
rect 77699 -47745 77733 -47711
rect 77791 -47745 77825 -47711
rect 77883 -47745 77917 -47711
rect 77975 -47745 78009 -47711
rect 78067 -47745 78101 -47711
rect 55320 -47960 55470 -47948
rect 55320 -47994 55470 -47960
rect 77420 -47820 77540 -47790
rect 77170 -47880 77260 -47830
rect 82867 -47765 82901 -47731
rect 82959 -47765 82993 -47731
rect 83051 -47765 83085 -47731
rect 83143 -47765 83177 -47731
rect 83235 -47765 83269 -47731
rect 83327 -47765 83361 -47731
rect 83419 -47765 83453 -47731
rect 83511 -47765 83545 -47731
rect 83603 -47765 83637 -47731
rect 83695 -47765 83729 -47731
rect 83787 -47765 83821 -47731
rect 83879 -47765 83913 -47731
rect 83971 -47765 84005 -47731
rect 84063 -47765 84097 -47731
rect 84155 -47765 84189 -47731
rect 84247 -47765 84281 -47731
rect 84339 -47765 84373 -47731
rect 84431 -47765 84465 -47731
rect 84523 -47765 84557 -47731
rect 84615 -47765 84649 -47731
rect 84707 -47765 84741 -47731
rect 84799 -47765 84833 -47731
rect 84891 -47765 84925 -47731
rect 84983 -47765 85017 -47731
rect 85075 -47765 85109 -47731
rect 85167 -47765 85201 -47731
rect 85259 -47765 85293 -47731
rect 85351 -47765 85385 -47731
rect 85443 -47765 85477 -47731
rect 85535 -47765 85569 -47731
rect 85627 -47765 85661 -47731
rect 85719 -47765 85753 -47731
rect 85811 -47765 85845 -47731
rect 85903 -47765 85937 -47731
rect 85995 -47765 86029 -47731
rect 86087 -47765 86121 -47731
rect 86179 -47765 86213 -47731
rect 86271 -47765 86305 -47731
rect 86363 -47765 86397 -47731
rect 86455 -47765 86489 -47731
rect 86547 -47765 86581 -47731
rect 86639 -47765 86673 -47731
rect 86731 -47765 86765 -47731
rect 86823 -47765 86857 -47731
rect 86915 -47765 86949 -47731
rect 87007 -47765 87041 -47731
rect 87099 -47765 87133 -47731
rect 87191 -47765 87225 -47731
rect 87283 -47765 87317 -47731
rect 87375 -47765 87409 -47731
rect 87467 -47765 87501 -47731
rect 87559 -47765 87593 -47731
rect 87651 -47765 87685 -47731
rect 87743 -47765 87777 -47731
rect 87835 -47765 87869 -47731
rect 87927 -47765 87961 -47731
rect 88019 -47765 88053 -47731
rect 88111 -47765 88145 -47731
rect 88203 -47765 88237 -47731
rect 88295 -47765 88329 -47731
rect 88387 -47765 88421 -47731
rect 88479 -47765 88513 -47731
rect 88571 -47765 88605 -47731
rect 88663 -47765 88697 -47731
rect 88755 -47765 88789 -47731
rect 88847 -47765 88881 -47731
rect 88939 -47765 88973 -47731
rect 89031 -47765 89065 -47731
rect 89123 -47765 89157 -47731
rect 89215 -47765 89249 -47731
rect 89307 -47765 89341 -47731
rect 89399 -47765 89433 -47731
rect 89491 -47765 89525 -47731
rect 89583 -47765 89617 -47731
rect 89675 -47765 89709 -47731
rect 89767 -47765 89801 -47731
rect 89859 -47765 89893 -47731
rect 89951 -47765 89985 -47731
rect 90043 -47765 90077 -47731
rect 90135 -47765 90169 -47731
rect 90227 -47765 90261 -47731
rect 90319 -47765 90353 -47731
rect 90411 -47765 90445 -47731
rect 90503 -47765 90537 -47731
rect 90595 -47765 90629 -47731
rect 90687 -47765 90721 -47731
rect 90779 -47765 90813 -47731
rect 90871 -47765 90905 -47731
rect 90963 -47765 90997 -47731
rect 91055 -47765 91089 -47731
rect 91147 -47765 91181 -47731
rect 91239 -47765 91273 -47731
rect 91331 -47765 91365 -47731
rect 78160 -47870 78200 -47830
rect 55320 -48008 55470 -47994
rect 77900 -47943 77940 -47940
rect 77900 -47977 77915 -47943
rect 77915 -47977 77940 -47943
rect 77900 -47980 77940 -47977
rect 78160 -47980 78200 -47940
rect 77770 -48040 77810 -48000
rect 77420 -48210 77470 -48160
rect 78160 -48100 78200 -48060
rect 82870 -48043 82930 -48040
rect 82870 -48077 82904 -48043
rect 82904 -48077 82930 -48043
rect 82870 -48130 82930 -48077
rect 83050 -48043 83090 -48040
rect 83050 -48077 83074 -48043
rect 83074 -48077 83090 -48043
rect 83050 -48130 83090 -48077
rect 85334 -47979 85342 -47958
rect 85342 -47979 85376 -47958
rect 85376 -47979 85384 -47958
rect 77607 -48289 77641 -48255
rect 77699 -48289 77733 -48255
rect 77791 -48289 77825 -48255
rect 77883 -48289 77917 -48255
rect 77975 -48289 78009 -48255
rect 78067 -48289 78101 -48255
rect 78250 -48290 78360 -48260
rect 77607 -48365 77641 -48331
rect 77699 -48365 77733 -48331
rect 77791 -48365 77825 -48331
rect 77883 -48365 77917 -48331
rect 77975 -48365 78009 -48331
rect 78250 -48340 78280 -48290
rect 78280 -48340 78330 -48290
rect 78330 -48340 78360 -48290
rect 78250 -48370 78360 -48340
rect 78560 -48290 78670 -48260
rect 78560 -48340 78590 -48290
rect 78590 -48340 78640 -48290
rect 78640 -48340 78670 -48290
rect 78560 -48370 78670 -48340
rect 78800 -48290 78910 -48260
rect 78800 -48340 78830 -48290
rect 78830 -48340 78880 -48290
rect 78880 -48340 78910 -48290
rect 78800 -48370 78910 -48340
rect 79060 -48290 79170 -48260
rect 85334 -48128 85384 -47979
rect 86814 -47945 86864 -47938
rect 86814 -47979 86848 -47945
rect 86848 -47979 86864 -47945
rect 85614 -48043 86475 -48035
rect 85614 -48069 85722 -48043
rect 85722 -48069 85756 -48043
rect 85756 -48069 85890 -48043
rect 85890 -48069 85924 -48043
rect 85924 -48069 86059 -48043
rect 86059 -48069 86093 -48043
rect 86093 -48069 86226 -48043
rect 86226 -48069 86260 -48043
rect 86260 -48069 86394 -48043
rect 86394 -48069 86428 -48043
rect 86428 -48069 86475 -48043
rect 86814 -48128 86864 -47979
rect 88284 -47979 88286 -47948
rect 88286 -47979 88320 -47948
rect 88320 -47979 88334 -47948
rect 87048 -48043 87909 -48034
rect 87048 -48068 87054 -48043
rect 87054 -48068 87194 -48043
rect 87194 -48068 87228 -48043
rect 87228 -48068 87362 -48043
rect 87362 -48068 87396 -48043
rect 87396 -48068 87531 -48043
rect 87531 -48068 87565 -48043
rect 87565 -48068 87698 -48043
rect 87698 -48068 87732 -48043
rect 87732 -48068 87866 -48043
rect 87866 -48068 87900 -48043
rect 87900 -48068 87909 -48043
rect 88284 -48128 88334 -47979
rect 89754 -47979 89758 -47948
rect 89758 -47979 89792 -47948
rect 89792 -47979 89804 -47948
rect 88527 -48043 89388 -48034
rect 88527 -48068 88666 -48043
rect 88666 -48068 88700 -48043
rect 88700 -48068 88834 -48043
rect 88834 -48068 88868 -48043
rect 88868 -48068 89003 -48043
rect 89003 -48068 89037 -48043
rect 89037 -48068 89170 -48043
rect 89170 -48068 89204 -48043
rect 89204 -48068 89338 -48043
rect 89338 -48068 89372 -48043
rect 89372 -48068 89388 -48043
rect 89754 -48131 89804 -47979
rect 89754 -48138 89758 -48131
rect 89758 -48138 89792 -48131
rect 89792 -48138 89804 -48131
rect 91224 -47979 91230 -47948
rect 91230 -47979 91264 -47948
rect 91264 -47979 91274 -47948
rect 89984 -48037 90751 -48035
rect 89982 -48043 90752 -48037
rect 89982 -48071 89998 -48043
rect 89998 -48071 90138 -48043
rect 90138 -48071 90172 -48043
rect 90172 -48071 90306 -48043
rect 90306 -48071 90340 -48043
rect 90340 -48071 90475 -48043
rect 90475 -48071 90509 -48043
rect 90509 -48071 90642 -48043
rect 90642 -48071 90676 -48043
rect 90676 -48071 90752 -48043
rect 91224 -48131 91274 -47979
rect 91224 -48138 91230 -48131
rect 91230 -48138 91264 -48131
rect 91264 -48138 91274 -48131
rect 79060 -48340 79090 -48290
rect 79090 -48340 79140 -48290
rect 79140 -48340 79170 -48290
rect 82867 -48309 82901 -48275
rect 82959 -48309 82993 -48275
rect 83051 -48309 83085 -48275
rect 83143 -48309 83177 -48275
rect 83235 -48309 83269 -48275
rect 83327 -48309 83361 -48275
rect 83419 -48309 83453 -48275
rect 83511 -48309 83545 -48275
rect 83603 -48309 83637 -48275
rect 83695 -48309 83729 -48275
rect 83787 -48309 83821 -48275
rect 83879 -48309 83913 -48275
rect 83971 -48309 84005 -48275
rect 84063 -48309 84097 -48275
rect 84155 -48309 84189 -48275
rect 84247 -48309 84281 -48275
rect 84339 -48309 84373 -48275
rect 84431 -48309 84465 -48275
rect 84523 -48309 84557 -48275
rect 84615 -48309 84649 -48275
rect 84707 -48309 84741 -48275
rect 84799 -48309 84833 -48275
rect 84891 -48309 84925 -48275
rect 84983 -48309 85017 -48275
rect 85075 -48309 85109 -48275
rect 85167 -48309 85201 -48275
rect 85259 -48309 85293 -48275
rect 85351 -48309 85385 -48275
rect 85443 -48309 85477 -48275
rect 85535 -48309 85569 -48275
rect 85627 -48309 85661 -48275
rect 85719 -48309 85753 -48275
rect 85811 -48309 85845 -48275
rect 85903 -48309 85937 -48275
rect 85995 -48309 86029 -48275
rect 86087 -48309 86121 -48275
rect 86179 -48309 86213 -48275
rect 86271 -48309 86305 -48275
rect 86363 -48309 86397 -48275
rect 86455 -48309 86489 -48275
rect 86547 -48309 86581 -48275
rect 86639 -48309 86673 -48275
rect 86731 -48309 86765 -48275
rect 86823 -48309 86857 -48275
rect 86915 -48309 86949 -48275
rect 87007 -48309 87041 -48275
rect 87099 -48309 87133 -48275
rect 87191 -48309 87225 -48275
rect 87283 -48309 87317 -48275
rect 87375 -48309 87409 -48275
rect 87467 -48309 87501 -48275
rect 87559 -48309 87593 -48275
rect 87651 -48309 87685 -48275
rect 87743 -48309 87777 -48275
rect 87835 -48309 87869 -48275
rect 87927 -48309 87961 -48275
rect 88019 -48309 88053 -48275
rect 88111 -48309 88145 -48275
rect 88203 -48309 88237 -48275
rect 88295 -48309 88329 -48275
rect 88387 -48309 88421 -48275
rect 88479 -48309 88513 -48275
rect 88571 -48309 88605 -48275
rect 88663 -48309 88697 -48275
rect 88755 -48309 88789 -48275
rect 88847 -48309 88881 -48275
rect 88939 -48309 88973 -48275
rect 89031 -48309 89065 -48275
rect 89123 -48309 89157 -48275
rect 89215 -48309 89249 -48275
rect 89307 -48309 89341 -48275
rect 89399 -48309 89433 -48275
rect 89491 -48309 89525 -48275
rect 89583 -48309 89617 -48275
rect 89675 -48309 89709 -48275
rect 89767 -48309 89801 -48275
rect 89859 -48309 89893 -48275
rect 89951 -48309 89985 -48275
rect 90043 -48309 90077 -48275
rect 90135 -48309 90169 -48275
rect 90227 -48309 90261 -48275
rect 90319 -48309 90353 -48275
rect 90411 -48309 90445 -48275
rect 90503 -48309 90537 -48275
rect 90595 -48309 90629 -48275
rect 90687 -48309 90721 -48275
rect 90779 -48309 90813 -48275
rect 90871 -48309 90905 -48275
rect 90963 -48309 90997 -48275
rect 91055 -48309 91089 -48275
rect 91147 -48309 91181 -48275
rect 91239 -48309 91273 -48275
rect 91331 -48309 91365 -48275
rect 79060 -48370 79170 -48340
rect 83484 -48378 83654 -48348
rect 25700 -50118 25736 -48682
rect 25736 -50118 25770 -48682
rect 25770 -50118 25780 -48682
rect 77460 -48640 77510 -48590
rect 83484 -48488 83514 -48378
rect 83514 -48488 83624 -48378
rect 83624 -48488 83654 -48378
rect 83484 -48518 83654 -48488
rect 85124 -48388 85294 -48358
rect 85124 -48498 85154 -48388
rect 85154 -48498 85264 -48388
rect 85264 -48498 85294 -48388
rect 85124 -48528 85294 -48498
rect 86534 -48378 86704 -48348
rect 86534 -48488 86564 -48378
rect 86564 -48488 86674 -48378
rect 86674 -48488 86704 -48378
rect 86534 -48518 86704 -48488
rect 87914 -48378 88084 -48348
rect 87914 -48488 87944 -48378
rect 87944 -48488 88054 -48378
rect 88054 -48488 88084 -48378
rect 87914 -48518 88084 -48488
rect 89454 -48388 89624 -48358
rect 89454 -48498 89484 -48388
rect 89484 -48498 89594 -48388
rect 89594 -48498 89624 -48388
rect 89454 -48528 89624 -48498
rect 90734 -48388 90904 -48358
rect 90734 -48498 90764 -48388
rect 90764 -48498 90874 -48388
rect 90874 -48498 90904 -48388
rect 90734 -48528 90904 -48498
rect 78000 -48610 78040 -48570
rect 77790 -48643 77830 -48630
rect 77790 -48670 77793 -48643
rect 77793 -48670 77827 -48643
rect 77827 -48670 77830 -48643
rect 25882 -49131 26996 -48734
rect 27124 -49131 28238 -48734
rect 28366 -49131 29480 -48734
rect 29608 -49131 30722 -48734
rect 30850 -49131 31964 -48734
rect 32092 -49131 33206 -48734
rect 33334 -49131 34448 -48734
rect 34576 -49131 35690 -48734
rect 25882 -50066 26996 -49669
rect 27124 -50066 28238 -49669
rect 28366 -50066 29480 -49669
rect 29608 -50066 30722 -49669
rect 30850 -50066 31964 -49669
rect 32092 -50066 33206 -49669
rect 33334 -50066 34448 -49669
rect 34576 -50066 35690 -49669
rect 25700 -50284 25780 -50118
rect 77400 -48770 77520 -48740
rect 77400 -48830 77430 -48770
rect 77430 -48830 77490 -48770
rect 77490 -48830 77520 -48770
rect 78000 -48700 78040 -48660
rect 78000 -48780 78040 -48740
rect 77400 -48860 77520 -48830
rect 77607 -48909 77641 -48875
rect 77699 -48909 77733 -48875
rect 77791 -48909 77825 -48875
rect 77883 -48909 77917 -48875
rect 77975 -48909 78009 -48875
rect 77607 -48985 77641 -48951
rect 77699 -48985 77733 -48951
rect 77791 -48985 77825 -48951
rect 77883 -48985 77917 -48951
rect 77975 -48985 78009 -48951
rect 78067 -48985 78101 -48951
rect 78159 -48985 78193 -48951
rect 78251 -48985 78285 -48951
rect 78343 -48985 78377 -48951
rect 78435 -48985 78469 -48951
rect 78527 -48985 78561 -48951
rect 77400 -49020 77520 -48990
rect 77400 -49080 77430 -49020
rect 77430 -49080 77490 -49020
rect 77490 -49080 77520 -49020
rect 77400 -49110 77520 -49080
rect 77470 -49260 77510 -49220
rect 77790 -49217 77793 -49190
rect 77793 -49217 77827 -49190
rect 77827 -49217 77830 -49190
rect 77790 -49230 77830 -49217
rect 78070 -49183 78110 -49130
rect 78070 -49217 78073 -49183
rect 78073 -49217 78107 -49183
rect 78107 -49217 78110 -49183
rect 78070 -49220 78110 -49217
rect 78570 -49140 78640 -49070
rect 78190 -49183 78280 -49180
rect 78190 -49217 78199 -49183
rect 78199 -49217 78233 -49183
rect 78233 -49217 78280 -49183
rect 78190 -49270 78280 -49217
rect 78360 -49183 78400 -49180
rect 78360 -49217 78375 -49183
rect 78375 -49217 78400 -49183
rect 78360 -49220 78400 -49217
rect 78570 -49280 78640 -49210
rect 78570 -49420 78640 -49350
rect 77607 -49529 77641 -49495
rect 77699 -49529 77733 -49495
rect 77791 -49529 77825 -49495
rect 77883 -49529 77917 -49495
rect 77975 -49529 78009 -49495
rect 78067 -49529 78101 -49495
rect 78159 -49529 78193 -49495
rect 78251 -49529 78285 -49495
rect 78343 -49529 78377 -49495
rect 78435 -49529 78469 -49495
rect 78527 -49529 78561 -49495
rect 78630 -49530 78740 -49500
rect 77607 -49605 77641 -49571
rect 77699 -49605 77733 -49571
rect 77791 -49605 77825 -49571
rect 77883 -49605 77917 -49571
rect 77975 -49605 78009 -49571
rect 78630 -49580 78660 -49530
rect 78660 -49580 78710 -49530
rect 78710 -49580 78740 -49530
rect 78630 -49610 78740 -49580
rect 78850 -49530 78960 -49500
rect 78850 -49580 78880 -49530
rect 78880 -49580 78930 -49530
rect 78930 -49580 78960 -49530
rect 78850 -49610 78960 -49580
rect 79090 -49530 79200 -49500
rect 79090 -49580 79120 -49530
rect 79120 -49580 79170 -49530
rect 79170 -49580 79200 -49530
rect 79090 -49610 79200 -49580
rect 77510 -49880 77560 -49830
rect 77980 -49820 78020 -49780
rect 77790 -49883 77830 -49870
rect 77790 -49910 77793 -49883
rect 77793 -49910 77827 -49883
rect 77827 -49910 77830 -49883
rect 77980 -49940 78020 -49900
rect 77420 -50030 77540 -50000
rect 77420 -50090 77450 -50030
rect 77450 -50090 77510 -50030
rect 77510 -50090 77540 -50030
rect 54150 -50158 54850 -50108
rect 25700 -51720 25736 -50284
rect 25736 -51720 25770 -50284
rect 25770 -51720 25780 -50284
rect 25882 -50733 26996 -50336
rect 27124 -50733 28238 -50336
rect 28366 -50733 29480 -50336
rect 29608 -50733 30722 -50336
rect 30850 -50733 31964 -50336
rect 32092 -50733 33206 -50336
rect 33334 -50733 34448 -50336
rect 34576 -50733 35690 -50336
rect 25882 -51668 26996 -51271
rect 27124 -51668 28238 -51271
rect 28366 -51668 29480 -51271
rect 29608 -51668 30722 -51271
rect 30850 -51668 31964 -51271
rect 32092 -51668 33206 -51271
rect 33334 -51668 34448 -51271
rect 34576 -51668 35690 -51271
rect 25700 -51882 25780 -51720
rect 54150 -50192 54850 -50158
rect 54150 -50198 54850 -50192
rect 54091 -50306 54867 -50272
rect 53998 -50372 54032 -50334
rect 54926 -50372 54960 -50334
rect 54091 -50434 54867 -50400
rect 77420 -50200 77540 -50090
rect 77980 -50040 78020 -50000
rect 77607 -50149 77641 -50115
rect 77699 -50149 77733 -50115
rect 77791 -50149 77825 -50115
rect 77883 -50149 77917 -50115
rect 77975 -50149 78009 -50115
rect 77420 -50260 77450 -50200
rect 77450 -50260 77510 -50200
rect 77510 -50260 77540 -50200
rect 77609 -50239 77643 -50205
rect 77701 -50239 77735 -50205
rect 77793 -50239 77827 -50205
rect 77885 -50239 77919 -50205
rect 77977 -50239 78011 -50205
rect 77420 -50290 77540 -50260
rect 55960 -50498 56040 -50328
rect 77980 -50420 78020 -50380
rect 53526 -50740 53614 -50706
rect 25700 -53318 25736 -51882
rect 25736 -53318 25770 -51882
rect 25770 -53318 25780 -51882
rect 25882 -52331 26996 -51934
rect 27124 -52331 28238 -51934
rect 28366 -52331 29480 -51934
rect 29608 -52331 30722 -51934
rect 30850 -52331 31964 -51934
rect 32092 -52331 33206 -51934
rect 33334 -52331 34448 -51934
rect 34576 -52331 35690 -51934
rect 25882 -53266 26996 -52869
rect 27124 -53266 28238 -52869
rect 28366 -53266 29480 -52869
rect 29608 -53266 30722 -52869
rect 30850 -53266 31964 -52869
rect 32092 -53266 33206 -52869
rect 33334 -53266 34448 -52869
rect 34576 -53266 35690 -52869
rect 25700 -53484 25780 -53318
rect 53330 -52118 53350 -50768
rect 53350 -52118 53384 -50768
rect 53384 -52118 53400 -50768
rect 53464 -51566 53498 -50790
rect 53642 -51566 53676 -50790
rect 57126 -50500 57356 -50470
rect 54091 -50662 54867 -50628
rect 53998 -50728 54032 -50690
rect 54926 -50728 54960 -50690
rect 54091 -50790 54867 -50756
rect 55334 -50802 55368 -50768
rect 55290 -51028 55324 -50852
rect 55378 -51028 55412 -50852
rect 55142 -51308 55494 -51274
rect 53942 -51412 54718 -51378
rect 53858 -51528 53892 -51440
rect 54768 -51528 54802 -51440
rect 53942 -51590 54718 -51556
rect 53526 -51650 53614 -51616
rect 55046 -51394 55080 -51360
rect 55556 -51394 55590 -51360
rect 55142 -51480 55494 -51446
rect 57126 -50570 57156 -50500
rect 57156 -50570 57316 -50500
rect 57316 -50570 57356 -50500
rect 77490 -50520 77540 -50470
rect 77790 -50471 77795 -50440
rect 77795 -50471 77829 -50440
rect 77829 -50471 77830 -50440
rect 77790 -50480 77830 -50471
rect 57126 -50600 57356 -50570
rect 58926 -50629 58966 -50620
rect 55882 -50690 55970 -50656
rect 55820 -51516 55854 -50740
rect 55998 -51516 56032 -50740
rect 55882 -51600 55970 -51566
rect 57125 -50679 57159 -50645
rect 57217 -50679 57251 -50645
rect 57309 -50679 57343 -50645
rect 57118 -50957 57178 -50944
rect 57118 -50991 57133 -50957
rect 57133 -50991 57167 -50957
rect 57167 -50991 57178 -50957
rect 57118 -50994 57178 -50991
rect 58926 -50915 58930 -50629
rect 58930 -50915 58964 -50629
rect 58964 -50915 58966 -50629
rect 77980 -50500 78020 -50460
rect 59125 -50681 59501 -50647
rect 59560 -50735 59594 -50701
rect 59125 -50789 59501 -50755
rect 59032 -50843 59066 -50809
rect 59125 -50897 59501 -50863
rect 58926 -50920 58966 -50915
rect 59656 -50915 59662 -50630
rect 59662 -50915 59696 -50630
rect 77980 -50600 78020 -50560
rect 77980 -50673 78020 -50640
rect 77980 -50680 77981 -50673
rect 77981 -50680 78020 -50673
rect 77609 -50783 77643 -50749
rect 77701 -50783 77735 -50749
rect 77793 -50783 77827 -50749
rect 77885 -50783 77919 -50749
rect 77977 -50783 78011 -50749
rect 78940 -50780 79050 -50750
rect 77607 -50855 77641 -50821
rect 77699 -50855 77733 -50821
rect 77791 -50855 77825 -50821
rect 77883 -50855 77917 -50821
rect 77975 -50855 78009 -50821
rect 78067 -50855 78101 -50821
rect 78159 -50855 78193 -50821
rect 78351 -50855 78385 -50821
rect 78443 -50855 78477 -50821
rect 78535 -50855 78569 -50821
rect 78627 -50855 78661 -50821
rect 78719 -50855 78753 -50821
rect 78811 -50855 78845 -50821
rect 78940 -50830 78970 -50780
rect 78970 -50830 79020 -50780
rect 79020 -50830 79050 -50780
rect 59656 -50920 59696 -50915
rect 57326 -50980 57366 -50940
rect 53526 -51758 53614 -51724
rect 55030 -51728 55110 -51648
rect 55740 -51668 55810 -51648
rect 55740 -51702 55802 -51668
rect 55802 -51702 55810 -51668
rect 55740 -51728 55810 -51702
rect 53464 -52584 53498 -51808
rect 53642 -52584 53676 -51808
rect 53942 -51818 54718 -51784
rect 53858 -51934 53892 -51846
rect 54768 -51934 54802 -51846
rect 53942 -51996 54718 -51962
rect 55142 -51930 55494 -51896
rect 55046 -52016 55080 -51982
rect 55556 -52016 55590 -51982
rect 55142 -52102 55494 -52068
rect 53526 -52668 53614 -52634
rect 54081 -52622 54857 -52588
rect 53988 -52688 54022 -52650
rect 54916 -52688 54950 -52650
rect 54081 -52750 54857 -52716
rect 55280 -52524 55314 -52348
rect 55368 -52524 55402 -52348
rect 55324 -52608 55358 -52574
rect 56280 -51200 56350 -51118
rect 56280 -51748 56316 -51200
rect 56316 -51748 56350 -51200
rect 59866 -50894 59868 -50860
rect 59868 -50894 60424 -50860
rect 60424 -50894 60426 -50860
rect 59866 -50900 60426 -50894
rect 59766 -50956 59806 -50950
rect 59103 -51112 59137 -51078
rect 56492 -51240 56530 -51206
rect 55882 -51804 55970 -51770
rect 55820 -52630 55854 -51854
rect 55998 -52630 56032 -51854
rect 55882 -52714 55970 -52680
rect 56430 -52075 56464 -51299
rect 56558 -52075 56592 -51299
rect 56492 -52168 56530 -52134
rect 57125 -51223 57159 -51189
rect 57217 -51223 57251 -51189
rect 57309 -51223 57343 -51189
rect 57086 -51310 57376 -51280
rect 57086 -51380 57116 -51310
rect 57116 -51380 57346 -51310
rect 57346 -51380 57376 -51310
rect 57086 -51410 57376 -51380
rect 58926 -51646 58930 -51160
rect 58930 -51646 58964 -51160
rect 58964 -51646 58966 -51160
rect 59044 -51547 59078 -51171
rect 59162 -51547 59196 -51171
rect 59103 -51640 59137 -51606
rect 58926 -51802 58966 -51646
rect 59766 -51134 59772 -50956
rect 59772 -51134 59806 -50956
rect 59958 -51008 60334 -50974
rect 59874 -51062 59908 -51028
rect 60384 -51062 60418 -51028
rect 59958 -51116 60334 -51082
rect 59766 -51140 59806 -51134
rect 59476 -51196 59656 -51190
rect 59476 -51230 59484 -51196
rect 59484 -51230 59642 -51196
rect 59642 -51230 59656 -51196
rect 77580 -51030 77630 -50980
rect 78940 -50860 79050 -50830
rect 79130 -50780 79240 -50750
rect 79130 -50830 79160 -50780
rect 79160 -50830 79210 -50780
rect 79210 -50830 79240 -50780
rect 79130 -50860 79240 -50830
rect 78250 -50963 78290 -50929
rect 59386 -51292 59426 -51290
rect 59386 -51648 59388 -51292
rect 59388 -51648 59422 -51292
rect 59422 -51648 59426 -51292
rect 59546 -51332 59580 -51298
rect 59502 -51558 59536 -51382
rect 59590 -51558 59624 -51382
rect 59546 -51642 59580 -51608
rect 59386 -51650 59426 -51648
rect 59862 -51332 59896 -51298
rect 59818 -51558 59852 -51382
rect 59906 -51558 59940 -51382
rect 59862 -51642 59896 -51608
rect 77410 -51280 77530 -51250
rect 78170 -51067 78187 -51050
rect 78187 -51067 78220 -51050
rect 77410 -51340 77440 -51280
rect 77440 -51340 77500 -51280
rect 77500 -51340 77530 -51280
rect 77770 -51133 77810 -51130
rect 77770 -51167 77789 -51133
rect 77789 -51167 77810 -51133
rect 77770 -51170 77810 -51167
rect 77870 -51167 77895 -51160
rect 77895 -51167 77910 -51160
rect 77870 -51200 77910 -51167
rect 77870 -51280 77910 -51240
rect 77970 -51290 78010 -51250
rect 78170 -51220 78220 -51067
rect 78850 -51010 78900 -50960
rect 78350 -51220 78400 -51180
rect 78470 -51130 78560 -51080
rect 78640 -51133 78690 -51130
rect 78640 -51167 78659 -51133
rect 78659 -51167 78690 -51133
rect 78640 -51170 78690 -51167
rect 78850 -51130 78900 -51080
rect 77410 -51370 77530 -51340
rect 78850 -51250 78900 -51200
rect 83450 -51200 83620 -51170
rect 83450 -51310 83480 -51200
rect 83480 -51310 83590 -51200
rect 83590 -51310 83620 -51200
rect 83450 -51340 83620 -51310
rect 85150 -51200 85320 -51170
rect 85150 -51310 85180 -51200
rect 85180 -51310 85290 -51200
rect 85290 -51310 85320 -51200
rect 85150 -51340 85320 -51310
rect 86530 -51200 86700 -51170
rect 86530 -51310 86560 -51200
rect 86560 -51310 86670 -51200
rect 86670 -51310 86700 -51200
rect 86530 -51340 86700 -51310
rect 87820 -51200 87990 -51170
rect 87820 -51310 87850 -51200
rect 87850 -51310 87960 -51200
rect 87960 -51310 87990 -51200
rect 87820 -51340 87990 -51310
rect 89340 -51200 89510 -51170
rect 89340 -51310 89370 -51200
rect 89370 -51310 89480 -51200
rect 89480 -51310 89510 -51200
rect 89340 -51340 89510 -51310
rect 90750 -51200 90920 -51170
rect 90750 -51310 90780 -51200
rect 90780 -51310 90890 -51200
rect 90890 -51310 90920 -51200
rect 90750 -51340 90920 -51310
rect 77607 -51399 77641 -51365
rect 77699 -51399 77733 -51365
rect 77791 -51399 77825 -51365
rect 77883 -51399 77917 -51365
rect 77975 -51399 78009 -51365
rect 78067 -51399 78101 -51365
rect 78159 -51399 78193 -51365
rect 78351 -51399 78385 -51365
rect 78443 -51399 78477 -51365
rect 78535 -51399 78569 -51365
rect 78627 -51399 78661 -51365
rect 78719 -51399 78753 -51365
rect 78811 -51399 78845 -51365
rect 61196 -51420 61366 -51400
rect 82867 -51415 82901 -51381
rect 82959 -51415 82993 -51381
rect 83051 -51415 83085 -51381
rect 83143 -51415 83177 -51381
rect 83235 -51415 83269 -51381
rect 83327 -51415 83361 -51381
rect 83419 -51415 83453 -51381
rect 83511 -51415 83545 -51381
rect 83603 -51415 83637 -51381
rect 83695 -51415 83729 -51381
rect 83787 -51415 83821 -51381
rect 83879 -51415 83913 -51381
rect 83971 -51415 84005 -51381
rect 84063 -51415 84097 -51381
rect 84155 -51415 84189 -51381
rect 84247 -51415 84281 -51381
rect 84339 -51415 84373 -51381
rect 84431 -51415 84465 -51381
rect 84523 -51415 84557 -51381
rect 84615 -51415 84649 -51381
rect 84707 -51415 84741 -51381
rect 84799 -51415 84833 -51381
rect 84891 -51415 84925 -51381
rect 84983 -51415 85017 -51381
rect 85075 -51415 85109 -51381
rect 85167 -51415 85201 -51381
rect 85259 -51415 85293 -51381
rect 85351 -51415 85385 -51381
rect 85443 -51415 85477 -51381
rect 85535 -51415 85569 -51381
rect 85627 -51415 85661 -51381
rect 85719 -51415 85753 -51381
rect 85811 -51415 85845 -51381
rect 85903 -51415 85937 -51381
rect 85995 -51415 86029 -51381
rect 86087 -51415 86121 -51381
rect 86179 -51415 86213 -51381
rect 86271 -51415 86305 -51381
rect 86363 -51415 86397 -51381
rect 86455 -51415 86489 -51381
rect 86547 -51415 86581 -51381
rect 86639 -51415 86673 -51381
rect 86731 -51415 86765 -51381
rect 86823 -51415 86857 -51381
rect 86915 -51415 86949 -51381
rect 87007 -51415 87041 -51381
rect 87099 -51415 87133 -51381
rect 87191 -51415 87225 -51381
rect 87283 -51415 87317 -51381
rect 87375 -51415 87409 -51381
rect 87467 -51415 87501 -51381
rect 87559 -51415 87593 -51381
rect 87651 -51415 87685 -51381
rect 87743 -51415 87777 -51381
rect 87835 -51415 87869 -51381
rect 87927 -51415 87961 -51381
rect 88019 -51415 88053 -51381
rect 88111 -51415 88145 -51381
rect 88203 -51415 88237 -51381
rect 88295 -51415 88329 -51381
rect 88387 -51415 88421 -51381
rect 88479 -51415 88513 -51381
rect 88571 -51415 88605 -51381
rect 88663 -51415 88697 -51381
rect 88755 -51415 88789 -51381
rect 88847 -51415 88881 -51381
rect 88939 -51415 88973 -51381
rect 89031 -51415 89065 -51381
rect 89123 -51415 89157 -51381
rect 89215 -51415 89249 -51381
rect 89307 -51415 89341 -51381
rect 89399 -51415 89433 -51381
rect 89491 -51415 89525 -51381
rect 89583 -51415 89617 -51381
rect 89675 -51415 89709 -51381
rect 89767 -51415 89801 -51381
rect 89859 -51415 89893 -51381
rect 89951 -51415 89985 -51381
rect 90043 -51415 90077 -51381
rect 90135 -51415 90169 -51381
rect 90227 -51415 90261 -51381
rect 90319 -51415 90353 -51381
rect 90411 -51415 90445 -51381
rect 90503 -51415 90537 -51381
rect 90595 -51415 90629 -51381
rect 90687 -51415 90721 -51381
rect 90779 -51415 90813 -51381
rect 90871 -51415 90905 -51381
rect 90963 -51415 90997 -51381
rect 91055 -51415 91089 -51381
rect 91147 -51415 91181 -51381
rect 91239 -51415 91273 -51381
rect 91331 -51415 91365 -51381
rect 61196 -51460 61216 -51420
rect 61216 -51460 61336 -51420
rect 61336 -51460 61366 -51420
rect 61196 -51480 61366 -51460
rect 77410 -51460 77530 -51430
rect 77410 -51520 77440 -51460
rect 77440 -51520 77500 -51460
rect 77500 -51520 77530 -51460
rect 77607 -51471 77641 -51437
rect 77699 -51471 77733 -51437
rect 77791 -51471 77825 -51437
rect 77883 -51471 77917 -51437
rect 77975 -51471 78009 -51437
rect 78067 -51471 78101 -51437
rect 78159 -51471 78193 -51437
rect 57056 -51970 57416 -51940
rect 57056 -52050 57096 -51970
rect 57096 -52050 57376 -51970
rect 57376 -52050 57416 -51970
rect 57056 -52080 57416 -52050
rect 57125 -52199 57159 -52165
rect 57217 -52199 57251 -52165
rect 57309 -52199 57343 -52165
rect 58926 -52290 58930 -51802
rect 58930 -52290 58964 -51802
rect 58964 -52290 58966 -51802
rect 60127 -51591 60161 -51557
rect 60366 -51565 60406 -51560
rect 60366 -51599 60393 -51565
rect 60393 -51599 60406 -51565
rect 60366 -51600 60406 -51599
rect 60127 -51683 60161 -51649
rect 59103 -51842 59137 -51808
rect 59044 -52277 59078 -51901
rect 57118 -52397 57168 -52394
rect 57118 -52431 57133 -52397
rect 57133 -52431 57167 -52397
rect 57167 -52431 57168 -52397
rect 57118 -52444 57168 -52431
rect 57326 -52410 57376 -52370
rect 59162 -52277 59196 -51901
rect 59103 -52370 59137 -52336
rect 59386 -51805 59426 -51800
rect 59386 -52161 59387 -51805
rect 59387 -52161 59421 -51805
rect 59421 -52161 59426 -51805
rect 59545 -51845 59579 -51811
rect 59501 -52071 59535 -51895
rect 59589 -52071 59623 -51895
rect 59545 -52155 59579 -52121
rect 59386 -52170 59426 -52161
rect 59476 -52223 59646 -52220
rect 59861 -51845 59895 -51811
rect 59817 -52071 59851 -51895
rect 59905 -52071 59939 -51895
rect 59861 -52155 59895 -52121
rect 60127 -51775 60161 -51741
rect 60127 -51867 60161 -51833
rect 60671 -51591 60705 -51557
rect 60366 -51657 60406 -51650
rect 60366 -51690 60393 -51657
rect 60393 -51690 60406 -51657
rect 60366 -51741 60406 -51740
rect 60366 -51775 60393 -51741
rect 60393 -51775 60406 -51741
rect 60366 -51780 60406 -51775
rect 60366 -51825 60406 -51820
rect 60366 -51859 60393 -51825
rect 60393 -51859 60406 -51825
rect 60366 -51860 60406 -51859
rect 60671 -51683 60705 -51649
rect 60671 -51775 60705 -51741
rect 60671 -51867 60705 -51833
rect 60127 -51959 60161 -51925
rect 60297 -51959 60331 -51925
rect 60369 -51959 60405 -51925
rect 60449 -51959 60484 -51925
rect 60671 -51959 60705 -51925
rect 60747 -51591 60781 -51557
rect 77410 -51550 77530 -51520
rect 61046 -51565 61086 -51560
rect 61046 -51599 61059 -51565
rect 61059 -51599 61086 -51565
rect 61046 -51600 61086 -51599
rect 60747 -51683 60781 -51649
rect 60747 -51775 60781 -51741
rect 60747 -51867 60781 -51833
rect 61291 -51591 61325 -51557
rect 61046 -51657 61086 -51650
rect 61046 -51690 61059 -51657
rect 61059 -51690 61086 -51657
rect 61046 -51741 61086 -51740
rect 61046 -51775 61059 -51741
rect 61059 -51775 61086 -51741
rect 61046 -51780 61086 -51775
rect 61046 -51825 61086 -51820
rect 61046 -51859 61059 -51825
rect 61059 -51859 61086 -51825
rect 61046 -51860 61086 -51859
rect 61291 -51683 61325 -51649
rect 61291 -51775 61325 -51741
rect 61291 -51867 61325 -51833
rect 77770 -51600 77810 -51560
rect 77770 -51669 77810 -51650
rect 77770 -51690 77789 -51669
rect 77789 -51690 77810 -51669
rect 77870 -51620 77910 -51580
rect 77870 -51669 77910 -51660
rect 77870 -51700 77895 -51669
rect 77895 -51700 77910 -51669
rect 78200 -51600 78280 -51550
rect 77970 -51703 77991 -51670
rect 77991 -51703 78010 -51670
rect 77970 -51710 78010 -51703
rect 78200 -51740 78280 -51690
rect 77440 -51860 77490 -51810
rect 60747 -51959 60781 -51925
rect 60980 -51959 61015 -51925
rect 61053 -51959 61088 -51925
rect 61129 -51958 61164 -51924
rect 61291 -51959 61325 -51925
rect 82870 -51693 82930 -51690
rect 82870 -51727 82904 -51693
rect 82904 -51727 82930 -51693
rect 82870 -51780 82930 -51727
rect 83040 -51693 83090 -51690
rect 83040 -51727 83074 -51693
rect 83074 -51727 83090 -51693
rect 83040 -51780 83090 -51727
rect 85330 -51629 85342 -51610
rect 85342 -51629 85376 -51610
rect 85376 -51629 85380 -51610
rect 78200 -51880 78280 -51830
rect 85330 -51780 85380 -51629
rect 86810 -51595 86860 -51590
rect 86810 -51629 86814 -51595
rect 86814 -51629 86848 -51595
rect 86848 -51629 86860 -51595
rect 85610 -51693 86471 -51687
rect 85610 -51721 85722 -51693
rect 85722 -51721 85756 -51693
rect 85756 -51721 85890 -51693
rect 85890 -51721 85924 -51693
rect 85924 -51721 86059 -51693
rect 86059 -51721 86093 -51693
rect 86093 -51721 86226 -51693
rect 86226 -51721 86260 -51693
rect 86260 -51721 86394 -51693
rect 86394 -51721 86428 -51693
rect 86428 -51721 86471 -51693
rect 86810 -51780 86860 -51629
rect 88280 -51629 88286 -51600
rect 88286 -51629 88320 -51600
rect 88320 -51629 88330 -51600
rect 87044 -51693 87905 -51686
rect 87044 -51720 87054 -51693
rect 87054 -51720 87194 -51693
rect 87194 -51720 87228 -51693
rect 87228 -51720 87362 -51693
rect 87362 -51720 87396 -51693
rect 87396 -51720 87531 -51693
rect 87531 -51720 87565 -51693
rect 87565 -51720 87698 -51693
rect 87698 -51720 87732 -51693
rect 87732 -51720 87866 -51693
rect 87866 -51720 87900 -51693
rect 87900 -51720 87905 -51693
rect 88280 -51780 88330 -51629
rect 89750 -51629 89758 -51600
rect 89758 -51629 89792 -51600
rect 89792 -51629 89800 -51600
rect 88523 -51693 89384 -51686
rect 88523 -51720 88526 -51693
rect 88526 -51720 88666 -51693
rect 88666 -51720 88700 -51693
rect 88700 -51720 88834 -51693
rect 88834 -51720 88868 -51693
rect 88868 -51720 89003 -51693
rect 89003 -51720 89037 -51693
rect 89037 -51720 89170 -51693
rect 89170 -51720 89204 -51693
rect 89204 -51720 89338 -51693
rect 89338 -51720 89372 -51693
rect 89372 -51720 89384 -51693
rect 89750 -51781 89800 -51629
rect 89750 -51790 89758 -51781
rect 89758 -51790 89792 -51781
rect 89792 -51790 89800 -51781
rect 91220 -51629 91230 -51600
rect 91230 -51629 91264 -51600
rect 91264 -51629 91270 -51600
rect 89980 -51689 90747 -51687
rect 89978 -51693 90748 -51689
rect 89978 -51723 89998 -51693
rect 89998 -51723 90138 -51693
rect 90138 -51723 90172 -51693
rect 90172 -51723 90306 -51693
rect 90306 -51723 90340 -51693
rect 90340 -51723 90475 -51693
rect 90475 -51723 90509 -51693
rect 90509 -51723 90642 -51693
rect 90642 -51723 90676 -51693
rect 90676 -51723 90748 -51693
rect 91220 -51781 91270 -51629
rect 91220 -51790 91230 -51781
rect 91230 -51790 91264 -51781
rect 91264 -51790 91270 -51781
rect 82867 -51959 82901 -51925
rect 82959 -51959 82993 -51925
rect 83051 -51959 83085 -51925
rect 83143 -51959 83177 -51925
rect 83235 -51959 83269 -51925
rect 83327 -51959 83361 -51925
rect 83419 -51959 83453 -51925
rect 83511 -51959 83545 -51925
rect 83603 -51959 83637 -51925
rect 83695 -51959 83729 -51925
rect 83787 -51959 83821 -51925
rect 83879 -51959 83913 -51925
rect 83971 -51959 84005 -51925
rect 84063 -51959 84097 -51925
rect 84155 -51959 84189 -51925
rect 84247 -51959 84281 -51925
rect 84339 -51959 84373 -51925
rect 84431 -51959 84465 -51925
rect 84523 -51959 84557 -51925
rect 84615 -51959 84649 -51925
rect 84707 -51959 84741 -51925
rect 84799 -51959 84833 -51925
rect 84891 -51959 84925 -51925
rect 84983 -51959 85017 -51925
rect 85075 -51959 85109 -51925
rect 85167 -51959 85201 -51925
rect 85259 -51959 85293 -51925
rect 85351 -51959 85385 -51925
rect 85443 -51959 85477 -51925
rect 85535 -51959 85569 -51925
rect 85627 -51959 85661 -51925
rect 85719 -51959 85753 -51925
rect 85811 -51959 85845 -51925
rect 85903 -51959 85937 -51925
rect 85995 -51959 86029 -51925
rect 86087 -51959 86121 -51925
rect 86179 -51959 86213 -51925
rect 86271 -51959 86305 -51925
rect 86363 -51959 86397 -51925
rect 86455 -51959 86489 -51925
rect 86547 -51959 86581 -51925
rect 86639 -51959 86673 -51925
rect 86731 -51959 86765 -51925
rect 86823 -51959 86857 -51925
rect 86915 -51959 86949 -51925
rect 87007 -51959 87041 -51925
rect 87099 -51959 87133 -51925
rect 87191 -51959 87225 -51925
rect 87283 -51959 87317 -51925
rect 87375 -51959 87409 -51925
rect 87467 -51959 87501 -51925
rect 87559 -51959 87593 -51925
rect 87651 -51959 87685 -51925
rect 87743 -51959 87777 -51925
rect 87835 -51959 87869 -51925
rect 87927 -51959 87961 -51925
rect 88019 -51959 88053 -51925
rect 88111 -51959 88145 -51925
rect 88203 -51959 88237 -51925
rect 88295 -51959 88329 -51925
rect 88387 -51959 88421 -51925
rect 88479 -51959 88513 -51925
rect 88571 -51959 88605 -51925
rect 88663 -51959 88697 -51925
rect 88755 -51959 88789 -51925
rect 88847 -51959 88881 -51925
rect 88939 -51959 88973 -51925
rect 89031 -51959 89065 -51925
rect 89123 -51959 89157 -51925
rect 89215 -51959 89249 -51925
rect 89307 -51959 89341 -51925
rect 89399 -51959 89433 -51925
rect 89491 -51959 89525 -51925
rect 89583 -51959 89617 -51925
rect 89675 -51959 89709 -51925
rect 89767 -51959 89801 -51925
rect 89859 -51959 89893 -51925
rect 89951 -51959 89985 -51925
rect 90043 -51959 90077 -51925
rect 90135 -51959 90169 -51925
rect 90227 -51959 90261 -51925
rect 90319 -51959 90353 -51925
rect 90411 -51959 90445 -51925
rect 90503 -51959 90537 -51925
rect 90595 -51959 90629 -51925
rect 90687 -51959 90721 -51925
rect 90779 -51959 90813 -51925
rect 90871 -51959 90905 -51925
rect 90963 -51959 90997 -51925
rect 91055 -51959 91089 -51925
rect 91147 -51959 91181 -51925
rect 91239 -51959 91273 -51925
rect 91331 -51959 91365 -51925
rect 77607 -52015 77641 -51981
rect 77699 -52015 77733 -51981
rect 77791 -52015 77825 -51981
rect 77883 -52015 77917 -51981
rect 77975 -52015 78009 -51981
rect 78067 -52015 78101 -51981
rect 78159 -52015 78193 -51981
rect 78280 -52010 78390 -51980
rect 60486 -52100 60526 -52060
rect 60626 -52100 60666 -52060
rect 60766 -52100 60806 -52060
rect 60906 -52100 60946 -52060
rect 77607 -52087 77641 -52053
rect 77699 -52087 77733 -52053
rect 77791 -52087 77825 -52053
rect 77883 -52087 77917 -52053
rect 77975 -52087 78009 -52053
rect 78067 -52087 78101 -52053
rect 78159 -52087 78193 -52053
rect 78280 -52060 78310 -52010
rect 78310 -52060 78360 -52010
rect 78360 -52060 78390 -52010
rect 59476 -52257 59483 -52223
rect 59483 -52257 59641 -52223
rect 59641 -52257 59646 -52223
rect 59476 -52260 59646 -52257
rect 59766 -52322 59806 -52320
rect 58926 -52536 58966 -52510
rect 59766 -52500 59772 -52322
rect 59772 -52500 59806 -52322
rect 77470 -52260 77510 -52210
rect 59958 -52374 60334 -52340
rect 59874 -52428 59908 -52394
rect 60384 -52428 60418 -52394
rect 59958 -52482 60334 -52448
rect 57125 -52743 57159 -52709
rect 57217 -52743 57251 -52709
rect 57309 -52743 57343 -52709
rect 54081 -52978 54857 -52944
rect 53988 -53044 54022 -53006
rect 54916 -53044 54950 -53006
rect 54081 -53106 54857 -53072
rect 56020 -53008 56080 -52858
rect 58926 -52822 58930 -52536
rect 58930 -52822 58964 -52536
rect 58964 -52822 58966 -52536
rect 59656 -52536 59706 -52530
rect 59125 -52588 59501 -52554
rect 59560 -52642 59594 -52608
rect 59125 -52696 59501 -52662
rect 59032 -52750 59066 -52716
rect 59125 -52804 59501 -52770
rect 57156 -52890 57316 -52860
rect 57156 -52990 57186 -52890
rect 57186 -52990 57286 -52890
rect 57286 -52990 57316 -52890
rect 58926 -52900 58966 -52822
rect 59656 -52822 59662 -52536
rect 59662 -52822 59696 -52536
rect 59696 -52822 59706 -52536
rect 78280 -52090 78390 -52060
rect 78580 -52010 78690 -51980
rect 78580 -52060 78610 -52010
rect 78610 -52060 78660 -52010
rect 78660 -52060 78690 -52010
rect 78580 -52090 78690 -52060
rect 78880 -52010 78990 -51980
rect 78880 -52060 78910 -52010
rect 78910 -52060 78960 -52010
rect 78960 -52060 78990 -52010
rect 78880 -52090 78990 -52060
rect 83480 -52030 83650 -52000
rect 83480 -52140 83510 -52030
rect 83510 -52140 83620 -52030
rect 83620 -52140 83650 -52030
rect 83480 -52170 83650 -52140
rect 85120 -52040 85290 -52010
rect 85120 -52150 85150 -52040
rect 85150 -52150 85260 -52040
rect 85260 -52150 85290 -52040
rect 85120 -52180 85290 -52150
rect 86530 -52030 86700 -52000
rect 86530 -52140 86560 -52030
rect 86560 -52140 86670 -52030
rect 86670 -52140 86700 -52030
rect 86530 -52170 86700 -52140
rect 87910 -52030 88080 -52000
rect 87910 -52140 87940 -52030
rect 87940 -52140 88050 -52030
rect 88050 -52140 88080 -52030
rect 87910 -52170 88080 -52140
rect 89450 -52040 89620 -52010
rect 89450 -52150 89480 -52040
rect 89480 -52150 89590 -52040
rect 89590 -52150 89620 -52040
rect 89450 -52180 89620 -52150
rect 90730 -52040 90900 -52010
rect 90730 -52150 90760 -52040
rect 90760 -52150 90870 -52040
rect 90870 -52150 90900 -52040
rect 90730 -52180 90900 -52150
rect 78180 -52197 78290 -52180
rect 78180 -52231 78187 -52197
rect 78187 -52231 78290 -52197
rect 78180 -52265 78290 -52231
rect 59866 -52562 60426 -52560
rect 77400 -52450 77520 -52420
rect 77400 -52510 77430 -52450
rect 77430 -52510 77490 -52450
rect 77490 -52510 77520 -52450
rect 78180 -52299 78187 -52265
rect 78187 -52299 78290 -52265
rect 77400 -52540 77520 -52510
rect 59866 -52596 59868 -52562
rect 59868 -52596 60424 -52562
rect 60424 -52596 60426 -52562
rect 77770 -52520 77810 -52480
rect 77870 -52365 77910 -52360
rect 77870 -52399 77895 -52365
rect 77895 -52399 77910 -52365
rect 77870 -52400 77910 -52399
rect 77870 -52510 77910 -52450
rect 77970 -52500 78010 -52400
rect 78180 -52453 78290 -52299
rect 78180 -52487 78187 -52453
rect 78187 -52487 78290 -52453
rect 78180 -52500 78290 -52487
rect 59866 -52600 60426 -52596
rect 77607 -52631 77641 -52597
rect 77699 -52631 77733 -52597
rect 77791 -52631 77825 -52597
rect 77883 -52631 77917 -52597
rect 77975 -52631 78009 -52597
rect 78067 -52631 78101 -52597
rect 78159 -52631 78193 -52597
rect 77400 -52700 77520 -52670
rect 77400 -52760 77430 -52700
rect 77430 -52760 77490 -52700
rect 77490 -52760 77520 -52700
rect 77607 -52705 77641 -52671
rect 77699 -52705 77733 -52671
rect 77791 -52705 77825 -52671
rect 77883 -52705 77917 -52671
rect 77975 -52705 78009 -52671
rect 78067 -52705 78101 -52671
rect 78159 -52705 78193 -52671
rect 77400 -52790 77520 -52760
rect 59656 -52830 59706 -52822
rect 57156 -53020 57316 -52990
rect 54150 -53220 54840 -53188
rect 54150 -53308 54840 -53220
rect 77580 -53080 77630 -52990
rect 77770 -52820 77810 -52780
rect 77870 -52903 77910 -52890
rect 77870 -52930 77895 -52903
rect 77895 -52930 77910 -52903
rect 77960 -52903 78010 -52900
rect 77960 -52937 77991 -52903
rect 77991 -52937 78010 -52903
rect 77960 -52950 78010 -52937
rect 55300 -53192 55476 -53158
rect 55526 -53236 55560 -53202
rect 55300 -53280 55476 -53246
rect 78190 -53120 78260 -52990
rect 77607 -53249 77641 -53215
rect 77699 -53249 77733 -53215
rect 77791 -53249 77825 -53215
rect 77883 -53249 77917 -53215
rect 77975 -53249 78009 -53215
rect 78067 -53249 78101 -53215
rect 78159 -53249 78193 -53215
rect 79120 -53250 79230 -53220
rect 55320 -53360 55470 -53348
rect 77607 -53325 77641 -53291
rect 77699 -53325 77733 -53291
rect 77791 -53325 77825 -53291
rect 77883 -53325 77917 -53291
rect 77975 -53325 78009 -53291
rect 78067 -53325 78101 -53291
rect 78159 -53325 78193 -53291
rect 78251 -53325 78285 -53291
rect 78343 -53325 78377 -53291
rect 78435 -53325 78469 -53291
rect 78527 -53325 78561 -53291
rect 78619 -53325 78653 -53291
rect 78711 -53325 78745 -53291
rect 78803 -53325 78837 -53291
rect 78895 -53325 78929 -53291
rect 78987 -53325 79021 -53291
rect 79120 -53300 79150 -53250
rect 79150 -53300 79200 -53250
rect 79200 -53300 79230 -53250
rect 55320 -53394 55470 -53360
rect 55320 -53408 55470 -53394
rect 25700 -54920 25738 -53484
rect 25738 -54920 25772 -53484
rect 25772 -54920 25780 -53484
rect 77770 -53410 77785 -53392
rect 77785 -53410 77830 -53392
rect 77770 -53432 77830 -53410
rect 25884 -53933 26998 -53536
rect 27126 -53933 28240 -53536
rect 28368 -53933 29482 -53536
rect 29610 -53933 30724 -53536
rect 30852 -53933 31966 -53536
rect 32094 -53933 33208 -53536
rect 33336 -53933 34450 -53536
rect 34578 -53933 35692 -53536
rect 25884 -54868 26998 -54471
rect 27126 -54868 28240 -54471
rect 28368 -54868 29482 -54471
rect 29610 -54868 30724 -54471
rect 30852 -54868 31966 -54471
rect 32094 -54868 33208 -54471
rect 33336 -54868 34450 -54471
rect 34578 -54868 35692 -54471
rect 25700 -55082 25780 -54920
rect 77390 -53700 77510 -53670
rect 77390 -53760 77420 -53700
rect 77420 -53760 77480 -53700
rect 77480 -53760 77510 -53700
rect 77620 -53683 77647 -53660
rect 77647 -53683 77690 -53660
rect 77620 -53710 77690 -53683
rect 77390 -53790 77510 -53760
rect 77820 -53643 77823 -53630
rect 77823 -53643 77857 -53630
rect 77857 -53643 77860 -53630
rect 77820 -53680 77860 -53643
rect 79120 -53330 79230 -53300
rect 78080 -53603 78130 -53530
rect 78080 -53620 78112 -53603
rect 78112 -53620 78130 -53603
rect 78250 -53603 78290 -53590
rect 78250 -53630 78253 -53603
rect 78253 -53630 78287 -53603
rect 78287 -53630 78290 -53603
rect 77990 -53733 78030 -53720
rect 77990 -53760 78003 -53733
rect 78003 -53760 78030 -53733
rect 78530 -53603 78570 -53600
rect 78530 -53637 78533 -53603
rect 78533 -53637 78567 -53603
rect 78567 -53637 78570 -53603
rect 78530 -53680 78570 -53637
rect 78650 -53603 78730 -53560
rect 78650 -53630 78659 -53603
rect 78659 -53630 78693 -53603
rect 78693 -53630 78730 -53603
rect 78820 -53603 78860 -53600
rect 78820 -53637 78835 -53603
rect 78835 -53637 78860 -53603
rect 78820 -53640 78860 -53637
rect 79020 -53720 79070 -53410
rect 77607 -53869 77641 -53835
rect 77699 -53869 77733 -53835
rect 77791 -53869 77825 -53835
rect 77883 -53869 77917 -53835
rect 77975 -53869 78009 -53835
rect 78067 -53869 78101 -53835
rect 78159 -53869 78193 -53835
rect 78251 -53869 78285 -53835
rect 78343 -53869 78377 -53835
rect 78435 -53869 78469 -53835
rect 78527 -53869 78561 -53835
rect 78619 -53869 78653 -53835
rect 78711 -53869 78745 -53835
rect 78803 -53869 78837 -53835
rect 78895 -53869 78929 -53835
rect 78987 -53869 79021 -53835
rect 25700 -56518 25736 -55082
rect 25736 -56518 25770 -55082
rect 25770 -56518 25780 -55082
rect 25882 -55531 26996 -55134
rect 27124 -55531 28238 -55134
rect 28366 -55531 29480 -55134
rect 29608 -55531 30722 -55134
rect 30850 -55531 31964 -55134
rect 32092 -55531 33206 -55134
rect 33334 -55531 34448 -55134
rect 34576 -55531 35690 -55134
rect 25882 -56466 26996 -56069
rect 27124 -56466 28238 -56069
rect 28366 -56466 29480 -56069
rect 29608 -56466 30722 -56069
rect 30850 -56466 31964 -56069
rect 32092 -56466 33206 -56069
rect 33334 -56466 34448 -56069
rect 34576 -56466 35690 -56069
rect 25700 -56682 25780 -56518
rect 54150 -55558 54850 -55508
rect 54150 -55592 54850 -55558
rect 54150 -55598 54850 -55592
rect 54091 -55706 54867 -55672
rect 53998 -55772 54032 -55734
rect 54926 -55772 54960 -55734
rect 54091 -55834 54867 -55800
rect 55960 -55898 56040 -55728
rect 53526 -56140 53614 -56106
rect 25700 -57980 25736 -56682
rect 25736 -57980 25770 -56682
rect 25770 -57980 25780 -56682
rect 25882 -57131 26996 -56734
rect 27124 -57131 28238 -56734
rect 28366 -57131 29480 -56734
rect 29608 -57131 30722 -56734
rect 30850 -57131 31964 -56734
rect 32092 -57131 33206 -56734
rect 33334 -57131 34448 -56734
rect 34576 -57131 35690 -56734
rect 25882 -58066 26996 -57669
rect 27124 -58066 28238 -57669
rect 28366 -58066 29480 -57669
rect 29608 -58066 30722 -57669
rect 30850 -58066 31964 -57669
rect 32092 -58066 33206 -57669
rect 33334 -58066 34448 -57669
rect 34576 -58066 35690 -57669
rect 53330 -57518 53350 -56168
rect 53350 -57518 53384 -56168
rect 53384 -57518 53400 -56168
rect 53464 -56966 53498 -56190
rect 53642 -56966 53676 -56190
rect 57126 -55900 57356 -55870
rect 54091 -56062 54867 -56028
rect 53998 -56128 54032 -56090
rect 54926 -56128 54960 -56090
rect 54091 -56190 54867 -56156
rect 55334 -56202 55368 -56168
rect 55290 -56428 55324 -56252
rect 55378 -56428 55412 -56252
rect 55142 -56708 55494 -56674
rect 53942 -56812 54718 -56778
rect 53858 -56928 53892 -56840
rect 54768 -56928 54802 -56840
rect 53942 -56990 54718 -56956
rect 53526 -57050 53614 -57016
rect 55046 -56794 55080 -56760
rect 55556 -56794 55590 -56760
rect 55142 -56880 55494 -56846
rect 57126 -55970 57156 -55900
rect 57156 -55970 57316 -55900
rect 57316 -55970 57356 -55900
rect 57126 -56000 57356 -55970
rect 58926 -56029 58966 -56020
rect 55882 -56090 55970 -56056
rect 55820 -56916 55854 -56140
rect 55998 -56916 56032 -56140
rect 55882 -57000 55970 -56966
rect 57125 -56079 57159 -56045
rect 57217 -56079 57251 -56045
rect 57309 -56079 57343 -56045
rect 57118 -56357 57178 -56344
rect 57118 -56391 57133 -56357
rect 57133 -56391 57167 -56357
rect 57167 -56391 57178 -56357
rect 57118 -56394 57178 -56391
rect 58926 -56315 58930 -56029
rect 58930 -56315 58964 -56029
rect 58964 -56315 58966 -56029
rect 59125 -56081 59501 -56047
rect 59560 -56135 59594 -56101
rect 59125 -56189 59501 -56155
rect 59032 -56243 59066 -56209
rect 59125 -56297 59501 -56263
rect 58926 -56320 58966 -56315
rect 59656 -56315 59662 -56030
rect 59662 -56315 59696 -56030
rect 59656 -56320 59696 -56315
rect 57326 -56380 57366 -56340
rect 53526 -57158 53614 -57124
rect 55030 -57128 55110 -57048
rect 55740 -57068 55810 -57048
rect 55740 -57102 55802 -57068
rect 55802 -57102 55810 -57068
rect 55740 -57128 55810 -57102
rect 53464 -57984 53498 -57208
rect 53642 -57984 53676 -57208
rect 53942 -57218 54718 -57184
rect 53858 -57334 53892 -57246
rect 54768 -57334 54802 -57246
rect 53942 -57396 54718 -57362
rect 55142 -57330 55494 -57296
rect 55046 -57416 55080 -57382
rect 55556 -57416 55590 -57382
rect 55142 -57502 55494 -57468
rect 53526 -58068 53614 -58034
rect 54081 -58022 54857 -57988
rect 53988 -58088 54022 -58050
rect 54916 -58088 54950 -58050
rect 54081 -58150 54857 -58116
rect 55280 -57924 55314 -57748
rect 55368 -57924 55402 -57748
rect 55324 -58008 55358 -57974
rect 56280 -56600 56350 -56518
rect 56280 -57148 56316 -56600
rect 56316 -57148 56350 -56600
rect 59866 -56294 59868 -56260
rect 59868 -56294 60424 -56260
rect 60424 -56294 60426 -56260
rect 59866 -56300 60426 -56294
rect 59766 -56356 59806 -56350
rect 59103 -56512 59137 -56478
rect 56492 -56640 56530 -56606
rect 55882 -57204 55970 -57170
rect 55820 -58030 55854 -57254
rect 55998 -58030 56032 -57254
rect 55882 -58114 55970 -58080
rect 56430 -57475 56464 -56699
rect 56558 -57475 56592 -56699
rect 56492 -57568 56530 -57534
rect 57125 -56623 57159 -56589
rect 57217 -56623 57251 -56589
rect 57309 -56623 57343 -56589
rect 57086 -56710 57376 -56680
rect 57086 -56780 57116 -56710
rect 57116 -56780 57346 -56710
rect 57346 -56780 57376 -56710
rect 57086 -56810 57376 -56780
rect 58926 -57046 58930 -56560
rect 58930 -57046 58964 -56560
rect 58964 -57046 58966 -56560
rect 59044 -56947 59078 -56571
rect 59162 -56947 59196 -56571
rect 59103 -57040 59137 -57006
rect 58926 -57202 58966 -57046
rect 59766 -56534 59772 -56356
rect 59772 -56534 59806 -56356
rect 59958 -56408 60334 -56374
rect 59874 -56462 59908 -56428
rect 60384 -56462 60418 -56428
rect 59958 -56516 60334 -56482
rect 59766 -56540 59806 -56534
rect 59476 -56596 59656 -56590
rect 59476 -56630 59484 -56596
rect 59484 -56630 59642 -56596
rect 59642 -56630 59656 -56596
rect 59386 -56692 59426 -56690
rect 59386 -57048 59388 -56692
rect 59388 -57048 59422 -56692
rect 59422 -57048 59426 -56692
rect 59546 -56732 59580 -56698
rect 59502 -56958 59536 -56782
rect 59590 -56958 59624 -56782
rect 59546 -57042 59580 -57008
rect 59386 -57050 59426 -57048
rect 59862 -56732 59896 -56698
rect 59818 -56958 59852 -56782
rect 59906 -56958 59940 -56782
rect 59862 -57042 59896 -57008
rect 61196 -56820 61366 -56800
rect 61196 -56860 61216 -56820
rect 61216 -56860 61336 -56820
rect 61336 -56860 61366 -56820
rect 61196 -56880 61366 -56860
rect 57056 -57370 57416 -57340
rect 57056 -57450 57096 -57370
rect 57096 -57450 57376 -57370
rect 57376 -57450 57416 -57370
rect 57056 -57480 57416 -57450
rect 57125 -57599 57159 -57565
rect 57217 -57599 57251 -57565
rect 57309 -57599 57343 -57565
rect 58926 -57690 58930 -57202
rect 58930 -57690 58964 -57202
rect 58964 -57690 58966 -57202
rect 60127 -56991 60161 -56957
rect 60366 -56965 60406 -56960
rect 60366 -56999 60393 -56965
rect 60393 -56999 60406 -56965
rect 60366 -57000 60406 -56999
rect 60127 -57083 60161 -57049
rect 59103 -57242 59137 -57208
rect 59044 -57677 59078 -57301
rect 57118 -57797 57168 -57794
rect 57118 -57831 57133 -57797
rect 57133 -57831 57167 -57797
rect 57167 -57831 57168 -57797
rect 57118 -57844 57168 -57831
rect 57326 -57810 57376 -57770
rect 59162 -57677 59196 -57301
rect 59103 -57770 59137 -57736
rect 59386 -57205 59426 -57200
rect 59386 -57561 59387 -57205
rect 59387 -57561 59421 -57205
rect 59421 -57561 59426 -57205
rect 59545 -57245 59579 -57211
rect 59501 -57471 59535 -57295
rect 59589 -57471 59623 -57295
rect 59545 -57555 59579 -57521
rect 59386 -57570 59426 -57561
rect 59476 -57623 59646 -57620
rect 59861 -57245 59895 -57211
rect 59817 -57471 59851 -57295
rect 59905 -57471 59939 -57295
rect 59861 -57555 59895 -57521
rect 60127 -57175 60161 -57141
rect 60127 -57267 60161 -57233
rect 60671 -56991 60705 -56957
rect 60366 -57057 60406 -57050
rect 60366 -57090 60393 -57057
rect 60393 -57090 60406 -57057
rect 60366 -57141 60406 -57140
rect 60366 -57175 60393 -57141
rect 60393 -57175 60406 -57141
rect 60366 -57180 60406 -57175
rect 60366 -57225 60406 -57220
rect 60366 -57259 60393 -57225
rect 60393 -57259 60406 -57225
rect 60366 -57260 60406 -57259
rect 60671 -57083 60705 -57049
rect 60671 -57175 60705 -57141
rect 60671 -57267 60705 -57233
rect 60127 -57359 60161 -57325
rect 60297 -57359 60331 -57325
rect 60369 -57359 60405 -57325
rect 60449 -57359 60484 -57325
rect 60671 -57359 60705 -57325
rect 60747 -56991 60781 -56957
rect 61046 -56965 61086 -56960
rect 61046 -56999 61059 -56965
rect 61059 -56999 61086 -56965
rect 61046 -57000 61086 -56999
rect 60747 -57083 60781 -57049
rect 60747 -57175 60781 -57141
rect 60747 -57267 60781 -57233
rect 61291 -56991 61325 -56957
rect 61046 -57057 61086 -57050
rect 61046 -57090 61059 -57057
rect 61059 -57090 61086 -57057
rect 61046 -57141 61086 -57140
rect 61046 -57175 61059 -57141
rect 61059 -57175 61086 -57141
rect 61046 -57180 61086 -57175
rect 61046 -57225 61086 -57220
rect 61046 -57259 61059 -57225
rect 61059 -57259 61086 -57225
rect 61046 -57260 61086 -57259
rect 61291 -57083 61325 -57049
rect 61291 -57175 61325 -57141
rect 61291 -57267 61325 -57233
rect 60747 -57359 60781 -57325
rect 60980 -57359 61015 -57325
rect 61053 -57359 61088 -57325
rect 61129 -57358 61164 -57324
rect 61291 -57359 61325 -57325
rect 60486 -57500 60526 -57460
rect 60626 -57500 60666 -57460
rect 60766 -57500 60806 -57460
rect 60906 -57500 60946 -57460
rect 59476 -57657 59483 -57623
rect 59483 -57657 59641 -57623
rect 59641 -57657 59646 -57623
rect 59476 -57660 59646 -57657
rect 59766 -57722 59806 -57720
rect 58926 -57936 58966 -57910
rect 59766 -57900 59772 -57722
rect 59772 -57900 59806 -57722
rect 59958 -57774 60334 -57740
rect 59874 -57828 59908 -57794
rect 60384 -57828 60418 -57794
rect 59958 -57882 60334 -57848
rect 57125 -58143 57159 -58109
rect 57217 -58143 57251 -58109
rect 57309 -58143 57343 -58109
rect 54081 -58378 54857 -58344
rect 53988 -58444 54022 -58406
rect 54916 -58444 54950 -58406
rect 54081 -58506 54857 -58472
rect 56020 -58408 56080 -58258
rect 58926 -58222 58930 -57936
rect 58930 -58222 58964 -57936
rect 58964 -58222 58966 -57936
rect 59656 -57936 59706 -57930
rect 59125 -57988 59501 -57954
rect 59560 -58042 59594 -58008
rect 59125 -58096 59501 -58062
rect 59032 -58150 59066 -58116
rect 59125 -58204 59501 -58170
rect 57156 -58290 57316 -58260
rect 57156 -58390 57186 -58290
rect 57186 -58390 57286 -58290
rect 57286 -58390 57316 -58290
rect 58926 -58300 58966 -58222
rect 59656 -58222 59662 -57936
rect 59662 -58222 59696 -57936
rect 59696 -58222 59706 -57936
rect 59866 -57962 60426 -57960
rect 59866 -57996 59868 -57962
rect 59868 -57996 60424 -57962
rect 60424 -57996 60426 -57962
rect 59866 -58000 60426 -57996
rect 59656 -58230 59706 -58222
rect 57156 -58420 57316 -58390
rect 54150 -58620 54840 -58588
rect 54150 -58708 54840 -58620
rect 55300 -58592 55476 -58558
rect 55526 -58636 55560 -58602
rect 55300 -58680 55476 -58646
rect 55320 -58760 55470 -58748
rect 55320 -58794 55470 -58760
rect 55320 -58808 55470 -58794
rect 54150 -60958 54850 -60908
rect 54150 -60992 54850 -60958
rect 54150 -60998 54850 -60992
rect 54091 -61106 54867 -61072
rect 53998 -61172 54032 -61134
rect 54926 -61172 54960 -61134
rect 54091 -61234 54867 -61200
rect 55960 -61298 56040 -61128
rect 53526 -61540 53614 -61506
rect 53330 -62918 53350 -61568
rect 53350 -62918 53384 -61568
rect 53384 -62918 53400 -61568
rect 53464 -62366 53498 -61590
rect 53642 -62366 53676 -61590
rect 57126 -61300 57356 -61270
rect 54091 -61462 54867 -61428
rect 53998 -61528 54032 -61490
rect 54926 -61528 54960 -61490
rect 54091 -61590 54867 -61556
rect 55334 -61602 55368 -61568
rect 55290 -61828 55324 -61652
rect 55378 -61828 55412 -61652
rect 55142 -62108 55494 -62074
rect 53942 -62212 54718 -62178
rect 53858 -62328 53892 -62240
rect 54768 -62328 54802 -62240
rect 53942 -62390 54718 -62356
rect 53526 -62450 53614 -62416
rect 55046 -62194 55080 -62160
rect 55556 -62194 55590 -62160
rect 55142 -62280 55494 -62246
rect 57126 -61370 57156 -61300
rect 57156 -61370 57316 -61300
rect 57316 -61370 57356 -61300
rect 57126 -61400 57356 -61370
rect 58926 -61429 58966 -61420
rect 55882 -61490 55970 -61456
rect 55820 -62316 55854 -61540
rect 55998 -62316 56032 -61540
rect 55882 -62400 55970 -62366
rect 57125 -61479 57159 -61445
rect 57217 -61479 57251 -61445
rect 57309 -61479 57343 -61445
rect 57118 -61757 57178 -61744
rect 57118 -61791 57133 -61757
rect 57133 -61791 57167 -61757
rect 57167 -61791 57178 -61757
rect 57118 -61794 57178 -61791
rect 58926 -61715 58930 -61429
rect 58930 -61715 58964 -61429
rect 58964 -61715 58966 -61429
rect 59125 -61481 59501 -61447
rect 59560 -61535 59594 -61501
rect 59125 -61589 59501 -61555
rect 59032 -61643 59066 -61609
rect 59125 -61697 59501 -61663
rect 58926 -61720 58966 -61715
rect 59656 -61715 59662 -61430
rect 59662 -61715 59696 -61430
rect 59656 -61720 59696 -61715
rect 57326 -61780 57366 -61740
rect 53526 -62558 53614 -62524
rect 55030 -62528 55110 -62448
rect 55740 -62468 55810 -62448
rect 55740 -62502 55802 -62468
rect 55802 -62502 55810 -62468
rect 55740 -62528 55810 -62502
rect 53464 -63384 53498 -62608
rect 53642 -63384 53676 -62608
rect 53942 -62618 54718 -62584
rect 53858 -62734 53892 -62646
rect 54768 -62734 54802 -62646
rect 53942 -62796 54718 -62762
rect 55142 -62730 55494 -62696
rect 55046 -62816 55080 -62782
rect 55556 -62816 55590 -62782
rect 55142 -62902 55494 -62868
rect 53526 -63468 53614 -63434
rect 54081 -63422 54857 -63388
rect 53988 -63488 54022 -63450
rect 54916 -63488 54950 -63450
rect 54081 -63550 54857 -63516
rect 55280 -63324 55314 -63148
rect 55368 -63324 55402 -63148
rect 55324 -63408 55358 -63374
rect 56280 -62000 56350 -61918
rect 56280 -62548 56316 -62000
rect 56316 -62548 56350 -62000
rect 59866 -61694 59868 -61660
rect 59868 -61694 60424 -61660
rect 60424 -61694 60426 -61660
rect 59866 -61700 60426 -61694
rect 59766 -61756 59806 -61750
rect 59103 -61912 59137 -61878
rect 56492 -62040 56530 -62006
rect 55882 -62604 55970 -62570
rect 55820 -63430 55854 -62654
rect 55998 -63430 56032 -62654
rect 55882 -63514 55970 -63480
rect 56430 -62875 56464 -62099
rect 56558 -62875 56592 -62099
rect 56492 -62968 56530 -62934
rect 57125 -62023 57159 -61989
rect 57217 -62023 57251 -61989
rect 57309 -62023 57343 -61989
rect 57086 -62110 57376 -62080
rect 57086 -62180 57116 -62110
rect 57116 -62180 57346 -62110
rect 57346 -62180 57376 -62110
rect 57086 -62210 57376 -62180
rect 58926 -62446 58930 -61960
rect 58930 -62446 58964 -61960
rect 58964 -62446 58966 -61960
rect 59044 -62347 59078 -61971
rect 59162 -62347 59196 -61971
rect 59103 -62440 59137 -62406
rect 58926 -62602 58966 -62446
rect 59766 -61934 59772 -61756
rect 59772 -61934 59806 -61756
rect 59958 -61808 60334 -61774
rect 59874 -61862 59908 -61828
rect 60384 -61862 60418 -61828
rect 59958 -61916 60334 -61882
rect 59766 -61940 59806 -61934
rect 59476 -61996 59656 -61990
rect 59476 -62030 59484 -61996
rect 59484 -62030 59642 -61996
rect 59642 -62030 59656 -61996
rect 59386 -62092 59426 -62090
rect 59386 -62448 59388 -62092
rect 59388 -62448 59422 -62092
rect 59422 -62448 59426 -62092
rect 59546 -62132 59580 -62098
rect 59502 -62358 59536 -62182
rect 59590 -62358 59624 -62182
rect 59546 -62442 59580 -62408
rect 59386 -62450 59426 -62448
rect 59862 -62132 59896 -62098
rect 59818 -62358 59852 -62182
rect 59906 -62358 59940 -62182
rect 59862 -62442 59896 -62408
rect 61196 -62220 61366 -62200
rect 61196 -62260 61216 -62220
rect 61216 -62260 61336 -62220
rect 61336 -62260 61366 -62220
rect 61196 -62280 61366 -62260
rect 57056 -62770 57416 -62740
rect 57056 -62850 57096 -62770
rect 57096 -62850 57376 -62770
rect 57376 -62850 57416 -62770
rect 57056 -62880 57416 -62850
rect 57125 -62999 57159 -62965
rect 57217 -62999 57251 -62965
rect 57309 -62999 57343 -62965
rect 58926 -63090 58930 -62602
rect 58930 -63090 58964 -62602
rect 58964 -63090 58966 -62602
rect 60127 -62391 60161 -62357
rect 60366 -62365 60406 -62360
rect 60366 -62399 60393 -62365
rect 60393 -62399 60406 -62365
rect 60366 -62400 60406 -62399
rect 60127 -62483 60161 -62449
rect 59103 -62642 59137 -62608
rect 59044 -63077 59078 -62701
rect 57118 -63197 57168 -63194
rect 57118 -63231 57133 -63197
rect 57133 -63231 57167 -63197
rect 57167 -63231 57168 -63197
rect 57118 -63244 57168 -63231
rect 57326 -63210 57376 -63170
rect 59162 -63077 59196 -62701
rect 59103 -63170 59137 -63136
rect 59386 -62605 59426 -62600
rect 59386 -62961 59387 -62605
rect 59387 -62961 59421 -62605
rect 59421 -62961 59426 -62605
rect 59545 -62645 59579 -62611
rect 59501 -62871 59535 -62695
rect 59589 -62871 59623 -62695
rect 59545 -62955 59579 -62921
rect 59386 -62970 59426 -62961
rect 59476 -63023 59646 -63020
rect 59861 -62645 59895 -62611
rect 59817 -62871 59851 -62695
rect 59905 -62871 59939 -62695
rect 59861 -62955 59895 -62921
rect 60127 -62575 60161 -62541
rect 60127 -62667 60161 -62633
rect 60671 -62391 60705 -62357
rect 60366 -62457 60406 -62450
rect 60366 -62490 60393 -62457
rect 60393 -62490 60406 -62457
rect 60366 -62541 60406 -62540
rect 60366 -62575 60393 -62541
rect 60393 -62575 60406 -62541
rect 60366 -62580 60406 -62575
rect 60366 -62625 60406 -62620
rect 60366 -62659 60393 -62625
rect 60393 -62659 60406 -62625
rect 60366 -62660 60406 -62659
rect 60671 -62483 60705 -62449
rect 60671 -62575 60705 -62541
rect 60671 -62667 60705 -62633
rect 60127 -62759 60161 -62725
rect 60297 -62759 60331 -62725
rect 60369 -62759 60405 -62725
rect 60449 -62759 60484 -62725
rect 60671 -62759 60705 -62725
rect 60747 -62391 60781 -62357
rect 61046 -62365 61086 -62360
rect 61046 -62399 61059 -62365
rect 61059 -62399 61086 -62365
rect 61046 -62400 61086 -62399
rect 60747 -62483 60781 -62449
rect 60747 -62575 60781 -62541
rect 60747 -62667 60781 -62633
rect 61291 -62391 61325 -62357
rect 61046 -62457 61086 -62450
rect 61046 -62490 61059 -62457
rect 61059 -62490 61086 -62457
rect 61046 -62541 61086 -62540
rect 61046 -62575 61059 -62541
rect 61059 -62575 61086 -62541
rect 61046 -62580 61086 -62575
rect 61046 -62625 61086 -62620
rect 61046 -62659 61059 -62625
rect 61059 -62659 61086 -62625
rect 61046 -62660 61086 -62659
rect 61291 -62483 61325 -62449
rect 61291 -62575 61325 -62541
rect 61291 -62667 61325 -62633
rect 60747 -62759 60781 -62725
rect 60980 -62759 61015 -62725
rect 61053 -62759 61088 -62725
rect 61129 -62758 61164 -62724
rect 61291 -62759 61325 -62725
rect 60486 -62900 60526 -62860
rect 60626 -62900 60666 -62860
rect 60766 -62900 60806 -62860
rect 60906 -62900 60946 -62860
rect 59476 -63057 59483 -63023
rect 59483 -63057 59641 -63023
rect 59641 -63057 59646 -63023
rect 59476 -63060 59646 -63057
rect 59766 -63122 59806 -63120
rect 58926 -63336 58966 -63310
rect 59766 -63300 59772 -63122
rect 59772 -63300 59806 -63122
rect 59958 -63174 60334 -63140
rect 59874 -63228 59908 -63194
rect 60384 -63228 60418 -63194
rect 59958 -63282 60334 -63248
rect 57125 -63543 57159 -63509
rect 57217 -63543 57251 -63509
rect 57309 -63543 57343 -63509
rect 54081 -63778 54857 -63744
rect 53988 -63844 54022 -63806
rect 54916 -63844 54950 -63806
rect 54081 -63906 54857 -63872
rect 56020 -63808 56080 -63658
rect 58926 -63622 58930 -63336
rect 58930 -63622 58964 -63336
rect 58964 -63622 58966 -63336
rect 59656 -63336 59706 -63330
rect 59125 -63388 59501 -63354
rect 59560 -63442 59594 -63408
rect 59125 -63496 59501 -63462
rect 59032 -63550 59066 -63516
rect 59125 -63604 59501 -63570
rect 57156 -63690 57316 -63660
rect 57156 -63790 57186 -63690
rect 57186 -63790 57286 -63690
rect 57286 -63790 57316 -63690
rect 58926 -63700 58966 -63622
rect 59656 -63622 59662 -63336
rect 59662 -63622 59696 -63336
rect 59696 -63622 59706 -63336
rect 59866 -63362 60426 -63360
rect 59866 -63396 59868 -63362
rect 59868 -63396 60424 -63362
rect 60424 -63396 60426 -63362
rect 59866 -63400 60426 -63396
rect 59656 -63630 59706 -63622
rect 57156 -63820 57316 -63790
rect 54150 -64020 54840 -63988
rect 54150 -64108 54840 -64020
rect 55300 -63992 55476 -63958
rect 55526 -64036 55560 -64002
rect 55300 -64080 55476 -64046
rect 55320 -64160 55470 -64148
rect 55320 -64194 55470 -64160
rect 55320 -64208 55470 -64194
rect 54150 -66358 54850 -66308
rect 54150 -66392 54850 -66358
rect 54150 -66398 54850 -66392
rect 54091 -66506 54867 -66472
rect 53998 -66572 54032 -66534
rect 54926 -66572 54960 -66534
rect 54091 -66634 54867 -66600
rect 55960 -66698 56040 -66528
rect 53526 -66940 53614 -66906
rect 53330 -68318 53350 -66968
rect 53350 -68318 53384 -66968
rect 53384 -68318 53400 -66968
rect 53464 -67766 53498 -66990
rect 53642 -67766 53676 -66990
rect 57126 -66700 57356 -66670
rect 54091 -66862 54867 -66828
rect 53998 -66928 54032 -66890
rect 54926 -66928 54960 -66890
rect 54091 -66990 54867 -66956
rect 55334 -67002 55368 -66968
rect 55290 -67228 55324 -67052
rect 55378 -67228 55412 -67052
rect 55142 -67508 55494 -67474
rect 53942 -67612 54718 -67578
rect 53858 -67728 53892 -67640
rect 54768 -67728 54802 -67640
rect 53942 -67790 54718 -67756
rect 53526 -67850 53614 -67816
rect 55046 -67594 55080 -67560
rect 55556 -67594 55590 -67560
rect 55142 -67680 55494 -67646
rect 57126 -66770 57156 -66700
rect 57156 -66770 57316 -66700
rect 57316 -66770 57356 -66700
rect 57126 -66800 57356 -66770
rect 58926 -66829 58966 -66820
rect 55882 -66890 55970 -66856
rect 55820 -67716 55854 -66940
rect 55998 -67716 56032 -66940
rect 55882 -67800 55970 -67766
rect 57125 -66879 57159 -66845
rect 57217 -66879 57251 -66845
rect 57309 -66879 57343 -66845
rect 57118 -67157 57178 -67144
rect 57118 -67191 57133 -67157
rect 57133 -67191 57167 -67157
rect 57167 -67191 57178 -67157
rect 57118 -67194 57178 -67191
rect 58926 -67115 58930 -66829
rect 58930 -67115 58964 -66829
rect 58964 -67115 58966 -66829
rect 59125 -66881 59501 -66847
rect 59560 -66935 59594 -66901
rect 59125 -66989 59501 -66955
rect 59032 -67043 59066 -67009
rect 59125 -67097 59501 -67063
rect 58926 -67120 58966 -67115
rect 59656 -67115 59662 -66830
rect 59662 -67115 59696 -66830
rect 59656 -67120 59696 -67115
rect 57326 -67180 57366 -67140
rect 53526 -67958 53614 -67924
rect 55030 -67928 55110 -67848
rect 55740 -67868 55810 -67848
rect 55740 -67902 55802 -67868
rect 55802 -67902 55810 -67868
rect 55740 -67928 55810 -67902
rect 53464 -68784 53498 -68008
rect 53642 -68784 53676 -68008
rect 53942 -68018 54718 -67984
rect 53858 -68134 53892 -68046
rect 54768 -68134 54802 -68046
rect 53942 -68196 54718 -68162
rect 55142 -68130 55494 -68096
rect 55046 -68216 55080 -68182
rect 55556 -68216 55590 -68182
rect 55142 -68302 55494 -68268
rect 53526 -68868 53614 -68834
rect 54081 -68822 54857 -68788
rect 53988 -68888 54022 -68850
rect 54916 -68888 54950 -68850
rect 54081 -68950 54857 -68916
rect 55280 -68724 55314 -68548
rect 55368 -68724 55402 -68548
rect 55324 -68808 55358 -68774
rect 56280 -67400 56350 -67318
rect 56280 -67948 56316 -67400
rect 56316 -67948 56350 -67400
rect 59866 -67094 59868 -67060
rect 59868 -67094 60424 -67060
rect 60424 -67094 60426 -67060
rect 59866 -67100 60426 -67094
rect 59766 -67156 59806 -67150
rect 59103 -67312 59137 -67278
rect 56492 -67440 56530 -67406
rect 55882 -68004 55970 -67970
rect 55820 -68830 55854 -68054
rect 55998 -68830 56032 -68054
rect 55882 -68914 55970 -68880
rect 56430 -68275 56464 -67499
rect 56558 -68275 56592 -67499
rect 56492 -68368 56530 -68334
rect 57125 -67423 57159 -67389
rect 57217 -67423 57251 -67389
rect 57309 -67423 57343 -67389
rect 57086 -67510 57376 -67480
rect 57086 -67580 57116 -67510
rect 57116 -67580 57346 -67510
rect 57346 -67580 57376 -67510
rect 57086 -67610 57376 -67580
rect 58926 -67846 58930 -67360
rect 58930 -67846 58964 -67360
rect 58964 -67846 58966 -67360
rect 59044 -67747 59078 -67371
rect 59162 -67747 59196 -67371
rect 59103 -67840 59137 -67806
rect 58926 -68002 58966 -67846
rect 59766 -67334 59772 -67156
rect 59772 -67334 59806 -67156
rect 59958 -67208 60334 -67174
rect 59874 -67262 59908 -67228
rect 60384 -67262 60418 -67228
rect 59958 -67316 60334 -67282
rect 59766 -67340 59806 -67334
rect 59476 -67396 59656 -67390
rect 59476 -67430 59484 -67396
rect 59484 -67430 59642 -67396
rect 59642 -67430 59656 -67396
rect 59386 -67492 59426 -67490
rect 59386 -67848 59388 -67492
rect 59388 -67848 59422 -67492
rect 59422 -67848 59426 -67492
rect 59546 -67532 59580 -67498
rect 59502 -67758 59536 -67582
rect 59590 -67758 59624 -67582
rect 59546 -67842 59580 -67808
rect 59386 -67850 59426 -67848
rect 59862 -67532 59896 -67498
rect 59818 -67758 59852 -67582
rect 59906 -67758 59940 -67582
rect 59862 -67842 59896 -67808
rect 61196 -67620 61366 -67600
rect 61196 -67660 61216 -67620
rect 61216 -67660 61336 -67620
rect 61336 -67660 61366 -67620
rect 61196 -67680 61366 -67660
rect 57056 -68170 57416 -68140
rect 57056 -68250 57096 -68170
rect 57096 -68250 57376 -68170
rect 57376 -68250 57416 -68170
rect 57056 -68280 57416 -68250
rect 57125 -68399 57159 -68365
rect 57217 -68399 57251 -68365
rect 57309 -68399 57343 -68365
rect 58926 -68490 58930 -68002
rect 58930 -68490 58964 -68002
rect 58964 -68490 58966 -68002
rect 60127 -67791 60161 -67757
rect 60366 -67765 60406 -67760
rect 60366 -67799 60393 -67765
rect 60393 -67799 60406 -67765
rect 60366 -67800 60406 -67799
rect 60127 -67883 60161 -67849
rect 59103 -68042 59137 -68008
rect 59044 -68477 59078 -68101
rect 57118 -68597 57168 -68594
rect 57118 -68631 57133 -68597
rect 57133 -68631 57167 -68597
rect 57167 -68631 57168 -68597
rect 57118 -68644 57168 -68631
rect 57326 -68610 57376 -68570
rect 59162 -68477 59196 -68101
rect 59103 -68570 59137 -68536
rect 59386 -68005 59426 -68000
rect 59386 -68361 59387 -68005
rect 59387 -68361 59421 -68005
rect 59421 -68361 59426 -68005
rect 59545 -68045 59579 -68011
rect 59501 -68271 59535 -68095
rect 59589 -68271 59623 -68095
rect 59545 -68355 59579 -68321
rect 59386 -68370 59426 -68361
rect 59476 -68423 59646 -68420
rect 59861 -68045 59895 -68011
rect 59817 -68271 59851 -68095
rect 59905 -68271 59939 -68095
rect 59861 -68355 59895 -68321
rect 60127 -67975 60161 -67941
rect 60127 -68067 60161 -68033
rect 60671 -67791 60705 -67757
rect 60366 -67857 60406 -67850
rect 60366 -67890 60393 -67857
rect 60393 -67890 60406 -67857
rect 60366 -67941 60406 -67940
rect 60366 -67975 60393 -67941
rect 60393 -67975 60406 -67941
rect 60366 -67980 60406 -67975
rect 60366 -68025 60406 -68020
rect 60366 -68059 60393 -68025
rect 60393 -68059 60406 -68025
rect 60366 -68060 60406 -68059
rect 60671 -67883 60705 -67849
rect 60671 -67975 60705 -67941
rect 60671 -68067 60705 -68033
rect 60127 -68159 60161 -68125
rect 60297 -68159 60331 -68125
rect 60369 -68159 60405 -68125
rect 60449 -68159 60484 -68125
rect 60671 -68159 60705 -68125
rect 60747 -67791 60781 -67757
rect 61046 -67765 61086 -67760
rect 61046 -67799 61059 -67765
rect 61059 -67799 61086 -67765
rect 61046 -67800 61086 -67799
rect 60747 -67883 60781 -67849
rect 60747 -67975 60781 -67941
rect 60747 -68067 60781 -68033
rect 61291 -67791 61325 -67757
rect 61046 -67857 61086 -67850
rect 61046 -67890 61059 -67857
rect 61059 -67890 61086 -67857
rect 61046 -67941 61086 -67940
rect 61046 -67975 61059 -67941
rect 61059 -67975 61086 -67941
rect 61046 -67980 61086 -67975
rect 61046 -68025 61086 -68020
rect 61046 -68059 61059 -68025
rect 61059 -68059 61086 -68025
rect 61046 -68060 61086 -68059
rect 61291 -67883 61325 -67849
rect 61291 -67975 61325 -67941
rect 61291 -68067 61325 -68033
rect 60747 -68159 60781 -68125
rect 60980 -68159 61015 -68125
rect 61053 -68159 61088 -68125
rect 61129 -68158 61164 -68124
rect 61291 -68159 61325 -68125
rect 60486 -68300 60526 -68260
rect 60626 -68300 60666 -68260
rect 60766 -68300 60806 -68260
rect 60906 -68300 60946 -68260
rect 59476 -68457 59483 -68423
rect 59483 -68457 59641 -68423
rect 59641 -68457 59646 -68423
rect 59476 -68460 59646 -68457
rect 59766 -68522 59806 -68520
rect 58926 -68736 58966 -68710
rect 59766 -68700 59772 -68522
rect 59772 -68700 59806 -68522
rect 59958 -68574 60334 -68540
rect 59874 -68628 59908 -68594
rect 60384 -68628 60418 -68594
rect 59958 -68682 60334 -68648
rect 57125 -68943 57159 -68909
rect 57217 -68943 57251 -68909
rect 57309 -68943 57343 -68909
rect 54081 -69178 54857 -69144
rect 53988 -69244 54022 -69206
rect 54916 -69244 54950 -69206
rect 54081 -69306 54857 -69272
rect 56020 -69208 56080 -69058
rect 58926 -69022 58930 -68736
rect 58930 -69022 58964 -68736
rect 58964 -69022 58966 -68736
rect 59656 -68736 59706 -68730
rect 59125 -68788 59501 -68754
rect 59560 -68842 59594 -68808
rect 59125 -68896 59501 -68862
rect 59032 -68950 59066 -68916
rect 59125 -69004 59501 -68970
rect 57156 -69090 57316 -69060
rect 57156 -69190 57186 -69090
rect 57186 -69190 57286 -69090
rect 57286 -69190 57316 -69090
rect 58926 -69100 58966 -69022
rect 59656 -69022 59662 -68736
rect 59662 -69022 59696 -68736
rect 59696 -69022 59706 -68736
rect 59866 -68762 60426 -68760
rect 59866 -68796 59868 -68762
rect 59868 -68796 60424 -68762
rect 60424 -68796 60426 -68762
rect 59866 -68800 60426 -68796
rect 59656 -69030 59706 -69022
rect 57156 -69220 57316 -69190
rect 54150 -69420 54840 -69388
rect 54150 -69508 54840 -69420
rect 55300 -69392 55476 -69358
rect 55526 -69436 55560 -69402
rect 55300 -69480 55476 -69446
rect 55320 -69560 55470 -69548
rect 55320 -69594 55470 -69560
rect 55320 -69608 55470 -69594
rect 54150 -71758 54850 -71708
rect 54150 -71792 54850 -71758
rect 54150 -71798 54850 -71792
rect 54091 -71906 54867 -71872
rect 53998 -71972 54032 -71934
rect 54926 -71972 54960 -71934
rect 54091 -72034 54867 -72000
rect 55960 -72098 56040 -71928
rect 53526 -72340 53614 -72306
rect 53330 -73718 53350 -72368
rect 53350 -73718 53384 -72368
rect 53384 -73718 53400 -72368
rect 53464 -73166 53498 -72390
rect 53642 -73166 53676 -72390
rect 57126 -72100 57356 -72070
rect 54091 -72262 54867 -72228
rect 53998 -72328 54032 -72290
rect 54926 -72328 54960 -72290
rect 54091 -72390 54867 -72356
rect 55334 -72402 55368 -72368
rect 55290 -72628 55324 -72452
rect 55378 -72628 55412 -72452
rect 55142 -72908 55494 -72874
rect 53942 -73012 54718 -72978
rect 53858 -73128 53892 -73040
rect 54768 -73128 54802 -73040
rect 53942 -73190 54718 -73156
rect 53526 -73250 53614 -73216
rect 55046 -72994 55080 -72960
rect 55556 -72994 55590 -72960
rect 55142 -73080 55494 -73046
rect 57126 -72170 57156 -72100
rect 57156 -72170 57316 -72100
rect 57316 -72170 57356 -72100
rect 57126 -72200 57356 -72170
rect 58926 -72229 58966 -72220
rect 55882 -72290 55970 -72256
rect 55820 -73116 55854 -72340
rect 55998 -73116 56032 -72340
rect 55882 -73200 55970 -73166
rect 57125 -72279 57159 -72245
rect 57217 -72279 57251 -72245
rect 57309 -72279 57343 -72245
rect 57118 -72557 57178 -72544
rect 57118 -72591 57133 -72557
rect 57133 -72591 57167 -72557
rect 57167 -72591 57178 -72557
rect 57118 -72594 57178 -72591
rect 58926 -72515 58930 -72229
rect 58930 -72515 58964 -72229
rect 58964 -72515 58966 -72229
rect 59125 -72281 59501 -72247
rect 59560 -72335 59594 -72301
rect 59125 -72389 59501 -72355
rect 59032 -72443 59066 -72409
rect 59125 -72497 59501 -72463
rect 58926 -72520 58966 -72515
rect 59656 -72515 59662 -72230
rect 59662 -72515 59696 -72230
rect 59656 -72520 59696 -72515
rect 57326 -72580 57366 -72540
rect 53526 -73358 53614 -73324
rect 55030 -73328 55110 -73248
rect 55740 -73268 55810 -73248
rect 55740 -73302 55802 -73268
rect 55802 -73302 55810 -73268
rect 55740 -73328 55810 -73302
rect 53464 -74184 53498 -73408
rect 53642 -74184 53676 -73408
rect 53942 -73418 54718 -73384
rect 53858 -73534 53892 -73446
rect 54768 -73534 54802 -73446
rect 53942 -73596 54718 -73562
rect 55142 -73530 55494 -73496
rect 55046 -73616 55080 -73582
rect 55556 -73616 55590 -73582
rect 55142 -73702 55494 -73668
rect 53526 -74268 53614 -74234
rect 54081 -74222 54857 -74188
rect 53988 -74288 54022 -74250
rect 54916 -74288 54950 -74250
rect 54081 -74350 54857 -74316
rect 55280 -74124 55314 -73948
rect 55368 -74124 55402 -73948
rect 55324 -74208 55358 -74174
rect 56280 -72800 56350 -72718
rect 56280 -73348 56316 -72800
rect 56316 -73348 56350 -72800
rect 59866 -72494 59868 -72460
rect 59868 -72494 60424 -72460
rect 60424 -72494 60426 -72460
rect 59866 -72500 60426 -72494
rect 59766 -72556 59806 -72550
rect 59103 -72712 59137 -72678
rect 56492 -72840 56530 -72806
rect 55882 -73404 55970 -73370
rect 55820 -74230 55854 -73454
rect 55998 -74230 56032 -73454
rect 55882 -74314 55970 -74280
rect 56430 -73675 56464 -72899
rect 56558 -73675 56592 -72899
rect 56492 -73768 56530 -73734
rect 57125 -72823 57159 -72789
rect 57217 -72823 57251 -72789
rect 57309 -72823 57343 -72789
rect 57086 -72910 57376 -72880
rect 57086 -72980 57116 -72910
rect 57116 -72980 57346 -72910
rect 57346 -72980 57376 -72910
rect 57086 -73010 57376 -72980
rect 58926 -73246 58930 -72760
rect 58930 -73246 58964 -72760
rect 58964 -73246 58966 -72760
rect 59044 -73147 59078 -72771
rect 59162 -73147 59196 -72771
rect 59103 -73240 59137 -73206
rect 58926 -73402 58966 -73246
rect 59766 -72734 59772 -72556
rect 59772 -72734 59806 -72556
rect 59958 -72608 60334 -72574
rect 59874 -72662 59908 -72628
rect 60384 -72662 60418 -72628
rect 59958 -72716 60334 -72682
rect 59766 -72740 59806 -72734
rect 59476 -72796 59656 -72790
rect 59476 -72830 59484 -72796
rect 59484 -72830 59642 -72796
rect 59642 -72830 59656 -72796
rect 59386 -72892 59426 -72890
rect 59386 -73248 59388 -72892
rect 59388 -73248 59422 -72892
rect 59422 -73248 59426 -72892
rect 59546 -72932 59580 -72898
rect 59502 -73158 59536 -72982
rect 59590 -73158 59624 -72982
rect 59546 -73242 59580 -73208
rect 59386 -73250 59426 -73248
rect 59862 -72932 59896 -72898
rect 59818 -73158 59852 -72982
rect 59906 -73158 59940 -72982
rect 59862 -73242 59896 -73208
rect 61196 -73020 61366 -73000
rect 61196 -73060 61216 -73020
rect 61216 -73060 61336 -73020
rect 61336 -73060 61366 -73020
rect 61196 -73080 61366 -73060
rect 57056 -73570 57416 -73540
rect 57056 -73650 57096 -73570
rect 57096 -73650 57376 -73570
rect 57376 -73650 57416 -73570
rect 57056 -73680 57416 -73650
rect 57125 -73799 57159 -73765
rect 57217 -73799 57251 -73765
rect 57309 -73799 57343 -73765
rect 58926 -73890 58930 -73402
rect 58930 -73890 58964 -73402
rect 58964 -73890 58966 -73402
rect 60127 -73191 60161 -73157
rect 60366 -73165 60406 -73160
rect 60366 -73199 60393 -73165
rect 60393 -73199 60406 -73165
rect 60366 -73200 60406 -73199
rect 60127 -73283 60161 -73249
rect 59103 -73442 59137 -73408
rect 59044 -73877 59078 -73501
rect 57118 -73997 57168 -73994
rect 57118 -74031 57133 -73997
rect 57133 -74031 57167 -73997
rect 57167 -74031 57168 -73997
rect 57118 -74044 57168 -74031
rect 57326 -74010 57376 -73970
rect 59162 -73877 59196 -73501
rect 59103 -73970 59137 -73936
rect 59386 -73405 59426 -73400
rect 59386 -73761 59387 -73405
rect 59387 -73761 59421 -73405
rect 59421 -73761 59426 -73405
rect 59545 -73445 59579 -73411
rect 59501 -73671 59535 -73495
rect 59589 -73671 59623 -73495
rect 59545 -73755 59579 -73721
rect 59386 -73770 59426 -73761
rect 59476 -73823 59646 -73820
rect 59861 -73445 59895 -73411
rect 59817 -73671 59851 -73495
rect 59905 -73671 59939 -73495
rect 59861 -73755 59895 -73721
rect 60127 -73375 60161 -73341
rect 60127 -73467 60161 -73433
rect 60671 -73191 60705 -73157
rect 60366 -73257 60406 -73250
rect 60366 -73290 60393 -73257
rect 60393 -73290 60406 -73257
rect 60366 -73341 60406 -73340
rect 60366 -73375 60393 -73341
rect 60393 -73375 60406 -73341
rect 60366 -73380 60406 -73375
rect 60366 -73425 60406 -73420
rect 60366 -73459 60393 -73425
rect 60393 -73459 60406 -73425
rect 60366 -73460 60406 -73459
rect 60671 -73283 60705 -73249
rect 60671 -73375 60705 -73341
rect 60671 -73467 60705 -73433
rect 60127 -73559 60161 -73525
rect 60297 -73559 60331 -73525
rect 60369 -73559 60405 -73525
rect 60449 -73559 60484 -73525
rect 60671 -73559 60705 -73525
rect 60747 -73191 60781 -73157
rect 61046 -73165 61086 -73160
rect 61046 -73199 61059 -73165
rect 61059 -73199 61086 -73165
rect 61046 -73200 61086 -73199
rect 60747 -73283 60781 -73249
rect 60747 -73375 60781 -73341
rect 60747 -73467 60781 -73433
rect 61291 -73191 61325 -73157
rect 61046 -73257 61086 -73250
rect 61046 -73290 61059 -73257
rect 61059 -73290 61086 -73257
rect 61046 -73341 61086 -73340
rect 61046 -73375 61059 -73341
rect 61059 -73375 61086 -73341
rect 61046 -73380 61086 -73375
rect 61046 -73425 61086 -73420
rect 61046 -73459 61059 -73425
rect 61059 -73459 61086 -73425
rect 61046 -73460 61086 -73459
rect 61291 -73283 61325 -73249
rect 61291 -73375 61325 -73341
rect 61291 -73467 61325 -73433
rect 60747 -73559 60781 -73525
rect 60980 -73559 61015 -73525
rect 61053 -73559 61088 -73525
rect 61129 -73558 61164 -73524
rect 61291 -73559 61325 -73525
rect 60486 -73700 60526 -73660
rect 60626 -73700 60666 -73660
rect 60766 -73700 60806 -73660
rect 60906 -73700 60946 -73660
rect 59476 -73857 59483 -73823
rect 59483 -73857 59641 -73823
rect 59641 -73857 59646 -73823
rect 59476 -73860 59646 -73857
rect 59766 -73922 59806 -73920
rect 58926 -74136 58966 -74110
rect 59766 -74100 59772 -73922
rect 59772 -74100 59806 -73922
rect 59958 -73974 60334 -73940
rect 59874 -74028 59908 -73994
rect 60384 -74028 60418 -73994
rect 59958 -74082 60334 -74048
rect 57125 -74343 57159 -74309
rect 57217 -74343 57251 -74309
rect 57309 -74343 57343 -74309
rect 54081 -74578 54857 -74544
rect 53988 -74644 54022 -74606
rect 54916 -74644 54950 -74606
rect 54081 -74706 54857 -74672
rect 56020 -74608 56080 -74458
rect 58926 -74422 58930 -74136
rect 58930 -74422 58964 -74136
rect 58964 -74422 58966 -74136
rect 59656 -74136 59706 -74130
rect 59125 -74188 59501 -74154
rect 59560 -74242 59594 -74208
rect 59125 -74296 59501 -74262
rect 59032 -74350 59066 -74316
rect 59125 -74404 59501 -74370
rect 57156 -74490 57316 -74460
rect 57156 -74590 57186 -74490
rect 57186 -74590 57286 -74490
rect 57286 -74590 57316 -74490
rect 58926 -74500 58966 -74422
rect 59656 -74422 59662 -74136
rect 59662 -74422 59696 -74136
rect 59696 -74422 59706 -74136
rect 59866 -74162 60426 -74160
rect 59866 -74196 59868 -74162
rect 59868 -74196 60424 -74162
rect 60424 -74196 60426 -74162
rect 59866 -74200 60426 -74196
rect 59656 -74430 59706 -74422
rect 57156 -74620 57316 -74590
rect 54150 -74820 54840 -74788
rect 54150 -74908 54840 -74820
rect 55300 -74792 55476 -74758
rect 55526 -74836 55560 -74802
rect 55300 -74880 55476 -74846
rect 55320 -74960 55470 -74948
rect 55320 -74994 55470 -74960
rect 55320 -75008 55470 -74994
rect 54150 -77158 54850 -77108
rect 54150 -77192 54850 -77158
rect 54150 -77198 54850 -77192
rect 54091 -77306 54867 -77272
rect 53998 -77372 54032 -77334
rect 54926 -77372 54960 -77334
rect 54091 -77434 54867 -77400
rect 55960 -77498 56040 -77328
rect 53526 -77740 53614 -77706
rect 53330 -79118 53350 -77768
rect 53350 -79118 53384 -77768
rect 53384 -79118 53400 -77768
rect 53464 -78566 53498 -77790
rect 53642 -78566 53676 -77790
rect 57126 -77500 57356 -77470
rect 54091 -77662 54867 -77628
rect 53998 -77728 54032 -77690
rect 54926 -77728 54960 -77690
rect 54091 -77790 54867 -77756
rect 55334 -77802 55368 -77768
rect 55290 -78028 55324 -77852
rect 55378 -78028 55412 -77852
rect 55142 -78308 55494 -78274
rect 53942 -78412 54718 -78378
rect 53858 -78528 53892 -78440
rect 54768 -78528 54802 -78440
rect 53942 -78590 54718 -78556
rect 53526 -78650 53614 -78616
rect 55046 -78394 55080 -78360
rect 55556 -78394 55590 -78360
rect 55142 -78480 55494 -78446
rect 57126 -77570 57156 -77500
rect 57156 -77570 57316 -77500
rect 57316 -77570 57356 -77500
rect 57126 -77600 57356 -77570
rect 58926 -77629 58966 -77620
rect 55882 -77690 55970 -77656
rect 55820 -78516 55854 -77740
rect 55998 -78516 56032 -77740
rect 55882 -78600 55970 -78566
rect 57125 -77679 57159 -77645
rect 57217 -77679 57251 -77645
rect 57309 -77679 57343 -77645
rect 57118 -77957 57178 -77944
rect 57118 -77991 57133 -77957
rect 57133 -77991 57167 -77957
rect 57167 -77991 57178 -77957
rect 57118 -77994 57178 -77991
rect 58926 -77915 58930 -77629
rect 58930 -77915 58964 -77629
rect 58964 -77915 58966 -77629
rect 59125 -77681 59501 -77647
rect 59560 -77735 59594 -77701
rect 59125 -77789 59501 -77755
rect 59032 -77843 59066 -77809
rect 59125 -77897 59501 -77863
rect 58926 -77920 58966 -77915
rect 59656 -77915 59662 -77630
rect 59662 -77915 59696 -77630
rect 59656 -77920 59696 -77915
rect 57326 -77980 57366 -77940
rect 53526 -78758 53614 -78724
rect 55030 -78728 55110 -78648
rect 55740 -78668 55810 -78648
rect 55740 -78702 55802 -78668
rect 55802 -78702 55810 -78668
rect 55740 -78728 55810 -78702
rect 53464 -79584 53498 -78808
rect 53642 -79584 53676 -78808
rect 53942 -78818 54718 -78784
rect 53858 -78934 53892 -78846
rect 54768 -78934 54802 -78846
rect 53942 -78996 54718 -78962
rect 55142 -78930 55494 -78896
rect 55046 -79016 55080 -78982
rect 55556 -79016 55590 -78982
rect 55142 -79102 55494 -79068
rect 53526 -79668 53614 -79634
rect 54081 -79622 54857 -79588
rect 53988 -79688 54022 -79650
rect 54916 -79688 54950 -79650
rect 54081 -79750 54857 -79716
rect 55280 -79524 55314 -79348
rect 55368 -79524 55402 -79348
rect 55324 -79608 55358 -79574
rect 56280 -78200 56350 -78118
rect 56280 -78748 56316 -78200
rect 56316 -78748 56350 -78200
rect 59866 -77894 59868 -77860
rect 59868 -77894 60424 -77860
rect 60424 -77894 60426 -77860
rect 59866 -77900 60426 -77894
rect 59766 -77956 59806 -77950
rect 59103 -78112 59137 -78078
rect 56492 -78240 56530 -78206
rect 55882 -78804 55970 -78770
rect 55820 -79630 55854 -78854
rect 55998 -79630 56032 -78854
rect 55882 -79714 55970 -79680
rect 56430 -79075 56464 -78299
rect 56558 -79075 56592 -78299
rect 56492 -79168 56530 -79134
rect 57125 -78223 57159 -78189
rect 57217 -78223 57251 -78189
rect 57309 -78223 57343 -78189
rect 57086 -78310 57376 -78280
rect 57086 -78380 57116 -78310
rect 57116 -78380 57346 -78310
rect 57346 -78380 57376 -78310
rect 57086 -78410 57376 -78380
rect 58926 -78646 58930 -78160
rect 58930 -78646 58964 -78160
rect 58964 -78646 58966 -78160
rect 59044 -78547 59078 -78171
rect 59162 -78547 59196 -78171
rect 59103 -78640 59137 -78606
rect 58926 -78802 58966 -78646
rect 59766 -78134 59772 -77956
rect 59772 -78134 59806 -77956
rect 59958 -78008 60334 -77974
rect 59874 -78062 59908 -78028
rect 60384 -78062 60418 -78028
rect 59958 -78116 60334 -78082
rect 59766 -78140 59806 -78134
rect 59476 -78196 59656 -78190
rect 59476 -78230 59484 -78196
rect 59484 -78230 59642 -78196
rect 59642 -78230 59656 -78196
rect 59386 -78292 59426 -78290
rect 59386 -78648 59388 -78292
rect 59388 -78648 59422 -78292
rect 59422 -78648 59426 -78292
rect 59546 -78332 59580 -78298
rect 59502 -78558 59536 -78382
rect 59590 -78558 59624 -78382
rect 59546 -78642 59580 -78608
rect 59386 -78650 59426 -78648
rect 59862 -78332 59896 -78298
rect 59818 -78558 59852 -78382
rect 59906 -78558 59940 -78382
rect 59862 -78642 59896 -78608
rect 61196 -78420 61366 -78400
rect 61196 -78460 61216 -78420
rect 61216 -78460 61336 -78420
rect 61336 -78460 61366 -78420
rect 61196 -78480 61366 -78460
rect 57056 -78970 57416 -78940
rect 57056 -79050 57096 -78970
rect 57096 -79050 57376 -78970
rect 57376 -79050 57416 -78970
rect 57056 -79080 57416 -79050
rect 57125 -79199 57159 -79165
rect 57217 -79199 57251 -79165
rect 57309 -79199 57343 -79165
rect 58926 -79290 58930 -78802
rect 58930 -79290 58964 -78802
rect 58964 -79290 58966 -78802
rect 60127 -78591 60161 -78557
rect 60366 -78565 60406 -78560
rect 60366 -78599 60393 -78565
rect 60393 -78599 60406 -78565
rect 60366 -78600 60406 -78599
rect 60127 -78683 60161 -78649
rect 59103 -78842 59137 -78808
rect 59044 -79277 59078 -78901
rect 57118 -79397 57168 -79394
rect 57118 -79431 57133 -79397
rect 57133 -79431 57167 -79397
rect 57167 -79431 57168 -79397
rect 57118 -79444 57168 -79431
rect 57326 -79410 57376 -79370
rect 59162 -79277 59196 -78901
rect 59103 -79370 59137 -79336
rect 59386 -78805 59426 -78800
rect 59386 -79161 59387 -78805
rect 59387 -79161 59421 -78805
rect 59421 -79161 59426 -78805
rect 59545 -78845 59579 -78811
rect 59501 -79071 59535 -78895
rect 59589 -79071 59623 -78895
rect 59545 -79155 59579 -79121
rect 59386 -79170 59426 -79161
rect 59476 -79223 59646 -79220
rect 59861 -78845 59895 -78811
rect 59817 -79071 59851 -78895
rect 59905 -79071 59939 -78895
rect 59861 -79155 59895 -79121
rect 60127 -78775 60161 -78741
rect 60127 -78867 60161 -78833
rect 60671 -78591 60705 -78557
rect 60366 -78657 60406 -78650
rect 60366 -78690 60393 -78657
rect 60393 -78690 60406 -78657
rect 60366 -78741 60406 -78740
rect 60366 -78775 60393 -78741
rect 60393 -78775 60406 -78741
rect 60366 -78780 60406 -78775
rect 60366 -78825 60406 -78820
rect 60366 -78859 60393 -78825
rect 60393 -78859 60406 -78825
rect 60366 -78860 60406 -78859
rect 60671 -78683 60705 -78649
rect 60671 -78775 60705 -78741
rect 60671 -78867 60705 -78833
rect 60127 -78959 60161 -78925
rect 60297 -78959 60331 -78925
rect 60369 -78959 60405 -78925
rect 60449 -78959 60484 -78925
rect 60671 -78959 60705 -78925
rect 60747 -78591 60781 -78557
rect 61046 -78565 61086 -78560
rect 61046 -78599 61059 -78565
rect 61059 -78599 61086 -78565
rect 61046 -78600 61086 -78599
rect 60747 -78683 60781 -78649
rect 60747 -78775 60781 -78741
rect 60747 -78867 60781 -78833
rect 61291 -78591 61325 -78557
rect 61046 -78657 61086 -78650
rect 61046 -78690 61059 -78657
rect 61059 -78690 61086 -78657
rect 61046 -78741 61086 -78740
rect 61046 -78775 61059 -78741
rect 61059 -78775 61086 -78741
rect 61046 -78780 61086 -78775
rect 61046 -78825 61086 -78820
rect 61046 -78859 61059 -78825
rect 61059 -78859 61086 -78825
rect 61046 -78860 61086 -78859
rect 61291 -78683 61325 -78649
rect 61291 -78775 61325 -78741
rect 61291 -78867 61325 -78833
rect 60747 -78959 60781 -78925
rect 60980 -78959 61015 -78925
rect 61053 -78959 61088 -78925
rect 61129 -78958 61164 -78924
rect 61291 -78959 61325 -78925
rect 60486 -79100 60526 -79060
rect 60626 -79100 60666 -79060
rect 60766 -79100 60806 -79060
rect 60906 -79100 60946 -79060
rect 59476 -79257 59483 -79223
rect 59483 -79257 59641 -79223
rect 59641 -79257 59646 -79223
rect 59476 -79260 59646 -79257
rect 59766 -79322 59806 -79320
rect 58926 -79536 58966 -79510
rect 59766 -79500 59772 -79322
rect 59772 -79500 59806 -79322
rect 59958 -79374 60334 -79340
rect 59874 -79428 59908 -79394
rect 60384 -79428 60418 -79394
rect 59958 -79482 60334 -79448
rect 57125 -79743 57159 -79709
rect 57217 -79743 57251 -79709
rect 57309 -79743 57343 -79709
rect 54081 -79978 54857 -79944
rect 53988 -80044 54022 -80006
rect 54916 -80044 54950 -80006
rect 54081 -80106 54857 -80072
rect 56020 -80008 56080 -79858
rect 58926 -79822 58930 -79536
rect 58930 -79822 58964 -79536
rect 58964 -79822 58966 -79536
rect 59656 -79536 59706 -79530
rect 59125 -79588 59501 -79554
rect 59560 -79642 59594 -79608
rect 59125 -79696 59501 -79662
rect 59032 -79750 59066 -79716
rect 59125 -79804 59501 -79770
rect 57156 -79890 57316 -79860
rect 57156 -79990 57186 -79890
rect 57186 -79990 57286 -79890
rect 57286 -79990 57316 -79890
rect 58926 -79900 58966 -79822
rect 59656 -79822 59662 -79536
rect 59662 -79822 59696 -79536
rect 59696 -79822 59706 -79536
rect 59866 -79562 60426 -79560
rect 59866 -79596 59868 -79562
rect 59868 -79596 60424 -79562
rect 60424 -79596 60426 -79562
rect 59866 -79600 60426 -79596
rect 59656 -79830 59706 -79822
rect 57156 -80020 57316 -79990
rect 54150 -80220 54840 -80188
rect 54150 -80308 54840 -80220
rect 55300 -80192 55476 -80158
rect 55526 -80236 55560 -80202
rect 55300 -80280 55476 -80246
rect 55320 -80360 55470 -80348
rect 55320 -80394 55470 -80360
rect 55320 -80408 55470 -80394
rect 54150 -82558 54850 -82508
rect 54150 -82592 54850 -82558
rect 54150 -82598 54850 -82592
rect 54091 -82706 54867 -82672
rect 53998 -82772 54032 -82734
rect 54926 -82772 54960 -82734
rect 54091 -82834 54867 -82800
rect 55960 -82898 56040 -82728
rect 53526 -83140 53614 -83106
rect 53330 -84518 53350 -83168
rect 53350 -84518 53384 -83168
rect 53384 -84518 53400 -83168
rect 53464 -83966 53498 -83190
rect 53642 -83966 53676 -83190
rect 57126 -82900 57356 -82870
rect 54091 -83062 54867 -83028
rect 53998 -83128 54032 -83090
rect 54926 -83128 54960 -83090
rect 54091 -83190 54867 -83156
rect 55334 -83202 55368 -83168
rect 55290 -83428 55324 -83252
rect 55378 -83428 55412 -83252
rect 55142 -83708 55494 -83674
rect 53942 -83812 54718 -83778
rect 53858 -83928 53892 -83840
rect 54768 -83928 54802 -83840
rect 53942 -83990 54718 -83956
rect 53526 -84050 53614 -84016
rect 55046 -83794 55080 -83760
rect 55556 -83794 55590 -83760
rect 55142 -83880 55494 -83846
rect 57126 -82970 57156 -82900
rect 57156 -82970 57316 -82900
rect 57316 -82970 57356 -82900
rect 57126 -83000 57356 -82970
rect 58926 -83029 58966 -83020
rect 55882 -83090 55970 -83056
rect 55820 -83916 55854 -83140
rect 55998 -83916 56032 -83140
rect 55882 -84000 55970 -83966
rect 57125 -83079 57159 -83045
rect 57217 -83079 57251 -83045
rect 57309 -83079 57343 -83045
rect 57118 -83357 57178 -83344
rect 57118 -83391 57133 -83357
rect 57133 -83391 57167 -83357
rect 57167 -83391 57178 -83357
rect 57118 -83394 57178 -83391
rect 58926 -83315 58930 -83029
rect 58930 -83315 58964 -83029
rect 58964 -83315 58966 -83029
rect 59125 -83081 59501 -83047
rect 59560 -83135 59594 -83101
rect 59125 -83189 59501 -83155
rect 59032 -83243 59066 -83209
rect 59125 -83297 59501 -83263
rect 58926 -83320 58966 -83315
rect 59656 -83315 59662 -83030
rect 59662 -83315 59696 -83030
rect 59656 -83320 59696 -83315
rect 57326 -83380 57366 -83340
rect 53526 -84158 53614 -84124
rect 55030 -84128 55110 -84048
rect 55740 -84068 55810 -84048
rect 55740 -84102 55802 -84068
rect 55802 -84102 55810 -84068
rect 55740 -84128 55810 -84102
rect 53464 -84984 53498 -84208
rect 53642 -84984 53676 -84208
rect 53942 -84218 54718 -84184
rect 53858 -84334 53892 -84246
rect 54768 -84334 54802 -84246
rect 53942 -84396 54718 -84362
rect 55142 -84330 55494 -84296
rect 55046 -84416 55080 -84382
rect 55556 -84416 55590 -84382
rect 55142 -84502 55494 -84468
rect 53526 -85068 53614 -85034
rect 54081 -85022 54857 -84988
rect 53988 -85088 54022 -85050
rect 54916 -85088 54950 -85050
rect 54081 -85150 54857 -85116
rect 55280 -84924 55314 -84748
rect 55368 -84924 55402 -84748
rect 55324 -85008 55358 -84974
rect 56280 -83600 56350 -83518
rect 56280 -84148 56316 -83600
rect 56316 -84148 56350 -83600
rect 59866 -83294 59868 -83260
rect 59868 -83294 60424 -83260
rect 60424 -83294 60426 -83260
rect 59866 -83300 60426 -83294
rect 59766 -83356 59806 -83350
rect 59103 -83512 59137 -83478
rect 56492 -83640 56530 -83606
rect 55882 -84204 55970 -84170
rect 55820 -85030 55854 -84254
rect 55998 -85030 56032 -84254
rect 55882 -85114 55970 -85080
rect 56430 -84475 56464 -83699
rect 56558 -84475 56592 -83699
rect 56492 -84568 56530 -84534
rect 57125 -83623 57159 -83589
rect 57217 -83623 57251 -83589
rect 57309 -83623 57343 -83589
rect 57086 -83710 57376 -83680
rect 57086 -83780 57116 -83710
rect 57116 -83780 57346 -83710
rect 57346 -83780 57376 -83710
rect 57086 -83810 57376 -83780
rect 58926 -84046 58930 -83560
rect 58930 -84046 58964 -83560
rect 58964 -84046 58966 -83560
rect 59044 -83947 59078 -83571
rect 59162 -83947 59196 -83571
rect 59103 -84040 59137 -84006
rect 58926 -84202 58966 -84046
rect 59766 -83534 59772 -83356
rect 59772 -83534 59806 -83356
rect 59958 -83408 60334 -83374
rect 59874 -83462 59908 -83428
rect 60384 -83462 60418 -83428
rect 59958 -83516 60334 -83482
rect 59766 -83540 59806 -83534
rect 59476 -83596 59656 -83590
rect 59476 -83630 59484 -83596
rect 59484 -83630 59642 -83596
rect 59642 -83630 59656 -83596
rect 59386 -83692 59426 -83690
rect 59386 -84048 59388 -83692
rect 59388 -84048 59422 -83692
rect 59422 -84048 59426 -83692
rect 59546 -83732 59580 -83698
rect 59502 -83958 59536 -83782
rect 59590 -83958 59624 -83782
rect 59546 -84042 59580 -84008
rect 59386 -84050 59426 -84048
rect 59862 -83732 59896 -83698
rect 59818 -83958 59852 -83782
rect 59906 -83958 59940 -83782
rect 59862 -84042 59896 -84008
rect 61196 -83820 61366 -83800
rect 61196 -83860 61216 -83820
rect 61216 -83860 61336 -83820
rect 61336 -83860 61366 -83820
rect 61196 -83880 61366 -83860
rect 57056 -84370 57416 -84340
rect 57056 -84450 57096 -84370
rect 57096 -84450 57376 -84370
rect 57376 -84450 57416 -84370
rect 57056 -84480 57416 -84450
rect 57125 -84599 57159 -84565
rect 57217 -84599 57251 -84565
rect 57309 -84599 57343 -84565
rect 58926 -84690 58930 -84202
rect 58930 -84690 58964 -84202
rect 58964 -84690 58966 -84202
rect 60127 -83991 60161 -83957
rect 60366 -83965 60406 -83960
rect 60366 -83999 60393 -83965
rect 60393 -83999 60406 -83965
rect 60366 -84000 60406 -83999
rect 60127 -84083 60161 -84049
rect 59103 -84242 59137 -84208
rect 59044 -84677 59078 -84301
rect 57118 -84797 57168 -84794
rect 57118 -84831 57133 -84797
rect 57133 -84831 57167 -84797
rect 57167 -84831 57168 -84797
rect 57118 -84844 57168 -84831
rect 57326 -84810 57376 -84770
rect 59162 -84677 59196 -84301
rect 59103 -84770 59137 -84736
rect 59386 -84205 59426 -84200
rect 59386 -84561 59387 -84205
rect 59387 -84561 59421 -84205
rect 59421 -84561 59426 -84205
rect 59545 -84245 59579 -84211
rect 59501 -84471 59535 -84295
rect 59589 -84471 59623 -84295
rect 59545 -84555 59579 -84521
rect 59386 -84570 59426 -84561
rect 59476 -84623 59646 -84620
rect 59861 -84245 59895 -84211
rect 59817 -84471 59851 -84295
rect 59905 -84471 59939 -84295
rect 59861 -84555 59895 -84521
rect 60127 -84175 60161 -84141
rect 60127 -84267 60161 -84233
rect 60671 -83991 60705 -83957
rect 60366 -84057 60406 -84050
rect 60366 -84090 60393 -84057
rect 60393 -84090 60406 -84057
rect 60366 -84141 60406 -84140
rect 60366 -84175 60393 -84141
rect 60393 -84175 60406 -84141
rect 60366 -84180 60406 -84175
rect 60366 -84225 60406 -84220
rect 60366 -84259 60393 -84225
rect 60393 -84259 60406 -84225
rect 60366 -84260 60406 -84259
rect 60671 -84083 60705 -84049
rect 60671 -84175 60705 -84141
rect 60671 -84267 60705 -84233
rect 60127 -84359 60161 -84325
rect 60297 -84359 60331 -84325
rect 60369 -84359 60405 -84325
rect 60449 -84359 60484 -84325
rect 60671 -84359 60705 -84325
rect 60747 -83991 60781 -83957
rect 61046 -83965 61086 -83960
rect 61046 -83999 61059 -83965
rect 61059 -83999 61086 -83965
rect 61046 -84000 61086 -83999
rect 60747 -84083 60781 -84049
rect 60747 -84175 60781 -84141
rect 60747 -84267 60781 -84233
rect 61291 -83991 61325 -83957
rect 61046 -84057 61086 -84050
rect 61046 -84090 61059 -84057
rect 61059 -84090 61086 -84057
rect 61046 -84141 61086 -84140
rect 61046 -84175 61059 -84141
rect 61059 -84175 61086 -84141
rect 61046 -84180 61086 -84175
rect 61046 -84225 61086 -84220
rect 61046 -84259 61059 -84225
rect 61059 -84259 61086 -84225
rect 61046 -84260 61086 -84259
rect 61291 -84083 61325 -84049
rect 61291 -84175 61325 -84141
rect 61291 -84267 61325 -84233
rect 60747 -84359 60781 -84325
rect 60980 -84359 61015 -84325
rect 61053 -84359 61088 -84325
rect 61129 -84358 61164 -84324
rect 61291 -84359 61325 -84325
rect 60486 -84500 60526 -84460
rect 60626 -84500 60666 -84460
rect 60766 -84500 60806 -84460
rect 60906 -84500 60946 -84460
rect 59476 -84657 59483 -84623
rect 59483 -84657 59641 -84623
rect 59641 -84657 59646 -84623
rect 59476 -84660 59646 -84657
rect 59766 -84722 59806 -84720
rect 58926 -84936 58966 -84910
rect 59766 -84900 59772 -84722
rect 59772 -84900 59806 -84722
rect 59958 -84774 60334 -84740
rect 59874 -84828 59908 -84794
rect 60384 -84828 60418 -84794
rect 59958 -84882 60334 -84848
rect 57125 -85143 57159 -85109
rect 57217 -85143 57251 -85109
rect 57309 -85143 57343 -85109
rect 54081 -85378 54857 -85344
rect 53988 -85444 54022 -85406
rect 54916 -85444 54950 -85406
rect 54081 -85506 54857 -85472
rect 56020 -85408 56080 -85258
rect 58926 -85222 58930 -84936
rect 58930 -85222 58964 -84936
rect 58964 -85222 58966 -84936
rect 59656 -84936 59706 -84930
rect 59125 -84988 59501 -84954
rect 59560 -85042 59594 -85008
rect 59125 -85096 59501 -85062
rect 59032 -85150 59066 -85116
rect 59125 -85204 59501 -85170
rect 57156 -85290 57316 -85260
rect 57156 -85390 57186 -85290
rect 57186 -85390 57286 -85290
rect 57286 -85390 57316 -85290
rect 58926 -85300 58966 -85222
rect 59656 -85222 59662 -84936
rect 59662 -85222 59696 -84936
rect 59696 -85222 59706 -84936
rect 59866 -84962 60426 -84960
rect 59866 -84996 59868 -84962
rect 59868 -84996 60424 -84962
rect 60424 -84996 60426 -84962
rect 59866 -85000 60426 -84996
rect 59656 -85230 59706 -85222
rect 57156 -85420 57316 -85390
rect 54150 -85620 54840 -85588
rect 54150 -85708 54840 -85620
rect 55300 -85592 55476 -85558
rect 55526 -85636 55560 -85602
rect 55300 -85680 55476 -85646
rect 55320 -85760 55470 -85748
rect 55320 -85794 55470 -85760
rect 55320 -85808 55470 -85794
<< metal1 >>
rect 37800 2800 41600 3000
rect 37800 1400 38000 2800
rect 41400 1400 41600 2800
rect 37800 -400 41600 1400
rect 37800 -3600 37900 -400
rect 41500 -3600 41600 -400
rect 42800 2400 46600 2600
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 0 46600 1000
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 50700 820 53300 2600
rect 50700 -20 50900 820
rect 53100 -20 53300 820
rect 50700 -100 53300 -20
rect 56720 1020 59220 2600
rect 56720 -40 56880 1020
rect 59080 -40 59220 1020
rect 56720 -100 59220 -40
rect 55300 -600 55800 -500
rect 55300 -1000 55400 -600
rect 55700 -1000 55800 -600
rect 42800 -1600 46600 -1400
rect 53300 -1400 53800 -1300
rect 53300 -1600 53400 -1400
rect 53700 -1600 53800 -1400
rect 54090 -1338 54890 -1298
rect 55300 -1300 55800 -1000
rect 54090 -1468 54150 -1338
rect 53300 -1700 53800 -1600
rect 54080 -1598 54150 -1468
rect 54860 -1578 54890 -1338
rect 54850 -1598 54890 -1578
rect 54080 -1666 54880 -1598
rect 53500 -1858 53800 -1700
rect 54079 -1672 54880 -1666
rect 54079 -1706 54091 -1672
rect 54867 -1698 54880 -1672
rect 54867 -1706 54879 -1698
rect 54079 -1712 54879 -1706
rect 53500 -1860 53520 -1858
rect 53002 -2020 53480 -1958
rect 37800 -3700 41600 -3600
rect 53000 -2158 53480 -2020
rect 53510 -1968 53520 -1860
rect 53640 -1968 53800 -1858
rect 53510 -2088 53800 -1968
rect 53970 -1734 54040 -1718
rect 53970 -1772 53998 -1734
rect 54032 -1772 54040 -1734
rect 53970 -1968 54040 -1772
rect 54920 -1734 54990 -1718
rect 54920 -1772 54926 -1734
rect 54960 -1772 54990 -1734
rect 54079 -1800 54879 -1794
rect 54079 -1834 54091 -1800
rect 54867 -1834 54879 -1800
rect 54079 -1838 54879 -1834
rect 54079 -1840 54750 -1838
rect 54090 -1888 54750 -1840
rect 54740 -1918 54750 -1888
rect 54850 -1840 54879 -1838
rect 54850 -1908 54860 -1840
rect 54840 -1918 54860 -1908
rect 54750 -1928 54860 -1918
rect 54920 -1968 54990 -1772
rect 55430 -1818 55520 -1808
rect 55290 -1928 55390 -1918
rect 53970 -1998 55290 -1968
rect 55430 -1958 55520 -1888
rect 53970 -2008 55390 -1998
rect 54050 -2018 55380 -2008
rect 54050 -2028 54880 -2018
rect 54050 -2038 54091 -2028
rect 54079 -2062 54091 -2038
rect 54867 -2038 54880 -2028
rect 54867 -2062 54879 -2038
rect 54079 -2068 54879 -2062
rect 54920 -2078 54990 -2068
rect 53510 -2106 53630 -2088
rect 53510 -2138 53526 -2106
rect 53514 -2140 53526 -2138
rect 53614 -2138 53630 -2106
rect 53940 -2090 54038 -2078
rect 53940 -2098 53998 -2090
rect 53614 -2140 53626 -2138
rect 53514 -2146 53626 -2140
rect 53000 -3908 53050 -2158
rect 53250 -2168 53480 -2158
rect 53250 -3518 53330 -2168
rect 53400 -2178 53480 -2168
rect 53400 -2190 53504 -2178
rect 53400 -2966 53464 -2190
rect 53498 -2966 53504 -2190
rect 53400 -2978 53504 -2966
rect 53636 -2188 53682 -2178
rect 53636 -2190 53760 -2188
rect 53636 -2966 53642 -2190
rect 53676 -2966 53760 -2190
rect 53940 -2198 53950 -2098
rect 54032 -2128 54038 -2090
rect 54020 -2140 54038 -2128
rect 54020 -2198 54030 -2140
rect 54079 -2156 54879 -2150
rect 54079 -2190 54091 -2156
rect 54867 -2190 54879 -2156
rect 54920 -2178 54990 -2168
rect 55320 -2168 55380 -2018
rect 54079 -2196 54879 -2190
rect 53940 -2218 54030 -2198
rect 54090 -2228 54870 -2196
rect 55320 -2202 55334 -2168
rect 55368 -2202 55380 -2168
rect 55320 -2208 55380 -2202
rect 53840 -2528 53920 -2518
rect 53840 -2638 53860 -2528
rect 53840 -2648 53920 -2638
rect 53840 -2840 53900 -2648
rect 54320 -2728 54510 -2228
rect 55440 -2238 55520 -1958
rect 55410 -2240 55520 -2238
rect 55284 -2248 55330 -2240
rect 55230 -2252 55330 -2248
rect 55230 -2258 55290 -2252
rect 55324 -2428 55330 -2252
rect 55230 -2438 55330 -2428
rect 55284 -2440 55330 -2438
rect 55372 -2248 55520 -2240
rect 55372 -2252 55430 -2248
rect 55372 -2428 55378 -2252
rect 55412 -2418 55430 -2252
rect 55510 -2418 55520 -2248
rect 55412 -2428 55520 -2418
rect 55372 -2440 55418 -2428
rect 55580 -2528 55720 -1300
rect 58776 -1470 59306 -1350
rect 58776 -1480 58966 -1470
rect 56146 -1580 57366 -1530
rect 55954 -1728 56046 -1716
rect 56146 -1728 56506 -1580
rect 55954 -1898 55960 -1728
rect 56040 -1898 56046 -1728
rect 55954 -1910 56046 -1898
rect 56120 -1758 56506 -1728
rect 56120 -1968 56190 -1758
rect 56390 -1830 56506 -1758
rect 57016 -1734 57366 -1580
rect 57586 -1630 58966 -1480
rect 59126 -1630 59306 -1470
rect 57586 -1650 59306 -1630
rect 59946 -1500 60386 -1400
rect 57586 -1680 58986 -1650
rect 59946 -1660 59956 -1500
rect 60166 -1660 60386 -1500
rect 57016 -1830 57368 -1734
rect 56390 -1870 57368 -1830
rect 56390 -1968 57126 -1870
rect 56120 -1974 57126 -1968
rect 56120 -1978 56750 -1974
rect 55880 -2018 55970 -2008
rect 55870 -2096 55880 -2050
rect 55970 -2096 55982 -2050
rect 55880 -2108 55970 -2098
rect 55000 -2538 55090 -2528
rect 55000 -2648 55090 -2638
rect 54710 -2728 54960 -2708
rect 53940 -2768 54960 -2728
rect 53940 -2772 54730 -2768
rect 53930 -2778 54730 -2772
rect 53930 -2812 53942 -2778
rect 54718 -2812 54730 -2778
rect 53930 -2818 54730 -2812
rect 53840 -2928 53858 -2840
rect 53892 -2928 53900 -2840
rect 53840 -2948 53900 -2928
rect 54762 -2838 54850 -2828
rect 54762 -2840 54770 -2838
rect 54762 -2928 54768 -2840
rect 54840 -2928 54850 -2838
rect 54762 -2940 54850 -2928
rect 54770 -2948 54850 -2940
rect 53636 -2978 53760 -2966
rect 53400 -3196 53480 -2978
rect 53514 -3016 53626 -3010
rect 53514 -3018 53526 -3016
rect 53510 -3050 53526 -3018
rect 53614 -3018 53626 -3016
rect 53614 -3050 53630 -3018
rect 53510 -3124 53630 -3050
rect 53510 -3158 53526 -3124
rect 53614 -3158 53630 -3124
rect 53680 -3038 53760 -2978
rect 53930 -2956 54730 -2950
rect 53930 -2990 53942 -2956
rect 54718 -2990 54730 -2956
rect 53930 -2996 54730 -2990
rect 53940 -3028 54720 -2996
rect 53920 -3038 54720 -3028
rect 53680 -3128 54720 -3038
rect 53514 -3164 53626 -3158
rect 53680 -3196 53760 -3128
rect 53920 -3138 54720 -3128
rect 53940 -3178 54720 -3138
rect 54900 -3168 54960 -2768
rect 55010 -2760 55090 -2648
rect 55540 -2538 55720 -2528
rect 55630 -2638 55720 -2538
rect 55130 -2674 55506 -2668
rect 55130 -2708 55142 -2674
rect 55494 -2708 55506 -2674
rect 55130 -2714 55506 -2708
rect 55010 -2794 55046 -2760
rect 55080 -2794 55090 -2760
rect 55010 -2808 55090 -2794
rect 55142 -2840 55494 -2714
rect 55540 -2760 55720 -2638
rect 55540 -2794 55556 -2760
rect 55590 -2794 55720 -2760
rect 55540 -2808 55720 -2794
rect 55780 -2140 55860 -2128
rect 55130 -2846 55506 -2840
rect 55130 -2880 55142 -2846
rect 55494 -2878 55506 -2846
rect 55494 -2880 55510 -2878
rect 55130 -2886 55510 -2880
rect 55140 -2898 55510 -2886
rect 55780 -2898 55820 -2140
rect 55140 -2916 55820 -2898
rect 55854 -2916 55860 -2140
rect 55140 -2928 55860 -2916
rect 55992 -2140 56038 -2128
rect 55992 -2916 55998 -2140
rect 56032 -2148 56038 -2140
rect 56120 -2148 56300 -1978
rect 57098 -2000 57126 -1974
rect 57356 -2000 57368 -1870
rect 57098 -2014 57368 -2000
rect 57096 -2045 57372 -2014
rect 57096 -2079 57125 -2045
rect 57159 -2079 57217 -2045
rect 57251 -2079 57309 -2045
rect 57343 -2079 57372 -2045
rect 57096 -2110 57372 -2079
rect 56032 -2506 56300 -2148
rect 56590 -2268 56660 -2258
rect 56660 -2334 57000 -2268
rect 57586 -2330 57706 -1680
rect 59946 -1690 60386 -1660
rect 57366 -2334 57706 -2330
rect 56660 -2338 57188 -2334
rect 56660 -2344 57190 -2338
rect 56660 -2394 57118 -2344
rect 57178 -2394 57190 -2344
rect 57314 -2340 57706 -2334
rect 57314 -2380 57326 -2340
rect 57366 -2380 57706 -2340
rect 57314 -2386 57706 -2380
rect 57366 -2390 57706 -2386
rect 58896 -1970 58986 -1950
rect 58896 -2030 58906 -1970
rect 58896 -2320 58926 -2030
rect 58966 -2320 58986 -1970
rect 59106 -1970 59516 -1960
rect 59106 -2030 59216 -1970
rect 59276 -2030 59326 -1970
rect 59386 -2030 59436 -1970
rect 59496 -2030 59516 -1970
rect 59106 -2047 59516 -2030
rect 59626 -1970 59706 -1930
rect 59626 -2030 59636 -1970
rect 59626 -2040 59656 -2030
rect 59106 -2080 59125 -2047
rect 59113 -2081 59125 -2080
rect 59501 -2080 59516 -2047
rect 59501 -2081 59513 -2080
rect 59113 -2087 59513 -2081
rect 59546 -2090 59616 -2080
rect 59276 -2130 59356 -2120
rect 59276 -2149 59286 -2130
rect 59113 -2155 59286 -2149
rect 59346 -2149 59356 -2130
rect 59346 -2155 59513 -2149
rect 59113 -2189 59125 -2155
rect 59501 -2189 59513 -2155
rect 59606 -2150 59616 -2090
rect 59546 -2160 59616 -2150
rect 59113 -2190 59286 -2189
rect 59346 -2190 59513 -2189
rect 59016 -2200 59076 -2190
rect 59113 -2195 59513 -2190
rect 59276 -2200 59356 -2195
rect 59546 -2210 59616 -2200
rect 59016 -2270 59076 -2260
rect 59113 -2263 59513 -2257
rect 59113 -2297 59125 -2263
rect 59501 -2297 59513 -2263
rect 59606 -2270 59616 -2210
rect 59546 -2280 59616 -2270
rect 59113 -2300 59513 -2297
rect 59113 -2303 59516 -2300
rect 58896 -2330 58986 -2320
rect 58896 -2390 58906 -2330
rect 58966 -2390 58986 -2330
rect 58896 -2392 58986 -2390
rect 59116 -2320 59516 -2303
rect 59646 -2310 59656 -2040
rect 59116 -2380 59216 -2320
rect 59276 -2380 59336 -2320
rect 59396 -2380 59436 -2320
rect 59496 -2380 59516 -2320
rect 56660 -2398 57190 -2394
rect 56590 -2400 57190 -2398
rect 56590 -2404 57188 -2400
rect 56590 -2468 57000 -2404
rect 56032 -2518 56356 -2506
rect 56032 -2916 56280 -2518
rect 55992 -2928 56280 -2916
rect 55140 -2938 55200 -2928
rect 55450 -2958 55810 -2928
rect 55870 -2966 55982 -2960
rect 55870 -3000 55882 -2966
rect 55970 -3000 55982 -2966
rect 55870 -3006 55982 -3000
rect 55140 -3018 55200 -3008
rect 55024 -3048 55116 -3036
rect 55024 -3128 55030 -3048
rect 55110 -3128 55116 -3048
rect 55024 -3140 55116 -3128
rect 55734 -3048 55816 -3036
rect 55734 -3128 55740 -3048
rect 55810 -3128 55816 -3048
rect 55734 -3140 55816 -3128
rect 55880 -3038 55970 -3006
rect 55880 -3164 55970 -3128
rect 56060 -3148 56280 -2928
rect 56350 -3148 56356 -2518
rect 56480 -2588 56550 -2578
rect 56480 -2658 56550 -2648
rect 56590 -2687 56750 -2468
rect 58894 -2486 58988 -2392
rect 59116 -2400 59516 -2380
rect 59636 -2320 59656 -2310
rect 59696 -2320 59706 -1970
rect 59856 -2140 59976 -2130
rect 59856 -2230 59866 -2140
rect 59966 -2230 59976 -2140
rect 59856 -2240 59976 -2230
rect 60436 -2220 60446 -2120
rect 60526 -2220 60536 -2120
rect 60436 -2240 60536 -2220
rect 59636 -2330 59706 -2320
rect 59696 -2390 59706 -2330
rect 59636 -2410 59706 -2390
rect 59756 -2260 60536 -2240
rect 59756 -2300 59866 -2260
rect 60426 -2300 60536 -2260
rect 59756 -2310 60536 -2300
rect 59756 -2350 59826 -2310
rect 59066 -2440 59176 -2430
rect 58896 -2550 58986 -2486
rect 59066 -2510 59076 -2440
rect 59166 -2510 59176 -2440
rect 59066 -2512 59103 -2510
rect 59137 -2512 59176 -2510
rect 59066 -2520 59176 -2512
rect 59756 -2540 59766 -2350
rect 59806 -2540 59826 -2350
rect 59956 -2368 60046 -2340
rect 59946 -2374 60046 -2368
rect 60126 -2368 60336 -2340
rect 60126 -2374 60346 -2368
rect 59856 -2410 59916 -2400
rect 59946 -2408 59958 -2374
rect 60334 -2408 60346 -2374
rect 59946 -2414 60346 -2408
rect 60376 -2420 60446 -2410
rect 59856 -2490 59916 -2480
rect 59946 -2482 60346 -2476
rect 59946 -2516 59958 -2482
rect 60334 -2516 60346 -2482
rect 60376 -2490 60446 -2480
rect 59946 -2522 59976 -2516
rect 57098 -2558 57368 -2554
rect 57096 -2564 57372 -2558
rect 57096 -2650 57098 -2564
rect 56424 -2688 56470 -2687
rect 56060 -3160 56356 -3148
rect 56410 -2699 56470 -2688
rect 53400 -3208 53504 -3196
rect 53400 -3518 53464 -3208
rect 53250 -3908 53464 -3518
rect 53000 -3984 53464 -3908
rect 53498 -3984 53504 -3208
rect 53000 -3988 53504 -3984
rect 53458 -3996 53504 -3988
rect 53636 -3208 53760 -3196
rect 53636 -3984 53642 -3208
rect 53676 -3984 53760 -3208
rect 53930 -3184 54730 -3178
rect 53930 -3218 53942 -3184
rect 54718 -3218 54730 -3184
rect 53930 -3224 54730 -3218
rect 53830 -3246 53900 -3228
rect 53830 -3334 53858 -3246
rect 53892 -3334 53900 -3246
rect 53830 -3528 53900 -3334
rect 54760 -3246 54850 -3228
rect 54760 -3334 54768 -3246
rect 54802 -3248 54850 -3246
rect 54900 -3238 55200 -3168
rect 55870 -3170 55982 -3164
rect 55870 -3204 55882 -3170
rect 55970 -3204 55982 -3170
rect 55450 -3238 55810 -3208
rect 55870 -3210 55982 -3204
rect 56060 -3238 56300 -3160
rect 54900 -3242 55820 -3238
rect 56000 -3242 56300 -3238
rect 54900 -3248 55860 -3242
rect 54840 -3328 54850 -3248
rect 54802 -3334 54850 -3328
rect 54760 -3348 54850 -3334
rect 55130 -3254 55860 -3248
rect 55130 -3278 55820 -3254
rect 55130 -3296 55510 -3278
rect 55130 -3330 55142 -3296
rect 55494 -3298 55510 -3296
rect 55494 -3330 55506 -3298
rect 55130 -3336 55506 -3330
rect 53930 -3362 54730 -3356
rect 53930 -3396 53942 -3362
rect 54718 -3396 54730 -3362
rect 55020 -3382 55090 -3368
rect 53930 -3402 54730 -3396
rect 53940 -3408 54730 -3402
rect 54920 -3398 54980 -3388
rect 53940 -3448 54920 -3408
rect 53830 -3538 53920 -3528
rect 53830 -3648 53850 -3538
rect 53830 -3658 53920 -3648
rect 54320 -3948 54510 -3448
rect 54710 -3468 54920 -3448
rect 54910 -3478 54980 -3468
rect 55020 -3416 55046 -3382
rect 55080 -3416 55090 -3382
rect 55020 -3528 55090 -3416
rect 55142 -3462 55494 -3336
rect 55540 -3382 55620 -3368
rect 55540 -3416 55556 -3382
rect 55590 -3416 55620 -3382
rect 55130 -3468 55506 -3462
rect 55130 -3502 55142 -3468
rect 55494 -3502 55506 -3468
rect 55130 -3508 55506 -3502
rect 55000 -3538 55090 -3528
rect 55000 -3648 55090 -3638
rect 55540 -3528 55620 -3416
rect 55540 -3538 55630 -3528
rect 55630 -3638 55680 -3548
rect 55540 -3648 55680 -3638
rect 55274 -3738 55320 -3736
rect 55220 -3748 55320 -3738
rect 55220 -3924 55280 -3918
rect 55314 -3924 55320 -3748
rect 55220 -3928 55320 -3924
rect 55274 -3936 55320 -3928
rect 55362 -3748 55408 -3736
rect 55362 -3924 55368 -3748
rect 55402 -3758 55510 -3748
rect 55402 -3924 55410 -3758
rect 55362 -3928 55410 -3924
rect 55500 -3928 55510 -3758
rect 55362 -3936 55510 -3928
rect 55390 -3938 55510 -3936
rect 53636 -3988 53760 -3984
rect 53636 -3996 53682 -3988
rect 53940 -4008 54020 -3968
rect 54080 -3982 54860 -3948
rect 55311 -3974 55371 -3968
rect 53514 -4034 53626 -4028
rect 53514 -4038 53526 -4034
rect 53510 -4068 53526 -4038
rect 53614 -4038 53626 -4034
rect 53614 -4068 53630 -4038
rect 53510 -4128 53630 -4068
rect 53940 -4088 53950 -4008
rect 54010 -4038 54020 -4008
rect 54069 -3988 54869 -3982
rect 54069 -4022 54081 -3988
rect 54857 -4022 54869 -3988
rect 54069 -4028 54869 -4022
rect 54910 -3998 54980 -3988
rect 54010 -4050 54028 -4038
rect 54022 -4088 54028 -4050
rect 53940 -4100 54028 -4088
rect 53940 -4108 54020 -4100
rect 54910 -4108 54980 -4098
rect 55311 -4008 55324 -3974
rect 55358 -4008 55371 -3974
rect 54070 -4110 54870 -4108
rect 54069 -4116 54870 -4110
rect 54069 -4138 54081 -4116
rect 54041 -4150 54081 -4138
rect 54857 -4118 54870 -4116
rect 54857 -4150 54880 -4118
rect 55311 -4148 55371 -4008
rect 54041 -4158 54880 -4150
rect 55240 -4158 55371 -4148
rect 54041 -4168 55240 -4158
rect 53510 -4258 53630 -4248
rect 53961 -4208 55240 -4168
rect 53961 -4406 54031 -4208
rect 54730 -4268 54860 -4258
rect 54730 -4288 54740 -4268
rect 54080 -4338 54740 -4288
rect 54069 -4344 54740 -4338
rect 54850 -4338 54860 -4268
rect 54850 -4344 54869 -4338
rect 54069 -4378 54081 -4344
rect 54857 -4378 54869 -4344
rect 54069 -4384 54869 -4378
rect 54911 -4394 54981 -4208
rect 55370 -4208 55371 -4158
rect 55240 -4228 55370 -4218
rect 55410 -4248 55510 -3938
rect 55410 -4358 55510 -4338
rect 55570 -4268 55680 -3648
rect 55780 -4030 55820 -3278
rect 55854 -4030 55860 -3254
rect 55780 -4038 55860 -4030
rect 55814 -4042 55860 -4038
rect 55992 -3254 56300 -3242
rect 55992 -4030 55998 -3254
rect 56032 -4028 56300 -3254
rect 56410 -3298 56430 -2699
rect 56380 -3475 56430 -3298
rect 56464 -3475 56470 -2699
rect 56380 -3487 56470 -3475
rect 56552 -2699 56750 -2687
rect 56552 -3475 56558 -2699
rect 56592 -2838 56750 -2699
rect 57066 -2680 57098 -2650
rect 57368 -2650 57372 -2564
rect 58896 -2559 59076 -2550
rect 58896 -2560 59084 -2559
rect 59156 -2560 59202 -2559
rect 57368 -2680 57396 -2650
rect 57066 -2810 57086 -2680
rect 57376 -2810 57396 -2680
rect 56592 -3475 56610 -2838
rect 57066 -2840 57396 -2810
rect 56860 -2990 57060 -2978
rect 56860 -3018 57236 -2990
rect 56860 -3148 56900 -3018
rect 57020 -3148 57236 -3018
rect 56860 -3188 57236 -3148
rect 57036 -3190 57236 -3188
rect 58556 -3080 58756 -3060
rect 58556 -3240 58576 -3080
rect 58736 -3240 58756 -3080
rect 58556 -3260 58756 -3240
rect 56552 -3478 56610 -3475
rect 57036 -3340 57446 -3330
rect 56552 -3487 56598 -3478
rect 57036 -3480 57056 -3340
rect 57416 -3480 57446 -3340
rect 56380 -3758 56440 -3487
rect 57036 -3500 57098 -3480
rect 56480 -3528 56550 -3518
rect 56480 -3598 56550 -3588
rect 57096 -3614 57098 -3534
rect 57368 -3500 57446 -3480
rect 57368 -3614 57372 -3534
rect 57096 -3630 57372 -3614
rect 58896 -3690 58926 -2560
rect 58966 -2571 59086 -2560
rect 58966 -2947 59044 -2571
rect 59078 -2947 59086 -2571
rect 58966 -2970 59086 -2947
rect 59156 -2571 59256 -2560
rect 59756 -2570 59826 -2540
rect 59966 -2552 59976 -2522
rect 60316 -2522 60346 -2516
rect 61036 -2520 61466 -2510
rect 60316 -2552 60326 -2522
rect 59966 -2560 60326 -2552
rect 59156 -2947 59162 -2571
rect 59196 -2640 59256 -2571
rect 59236 -2720 59256 -2640
rect 59196 -2840 59256 -2720
rect 59236 -2920 59256 -2840
rect 59196 -2947 59256 -2920
rect 59156 -2960 59256 -2947
rect 58966 -3280 59036 -2970
rect 59066 -3006 59176 -3000
rect 59066 -3010 59103 -3006
rect 59137 -3010 59176 -3006
rect 59066 -3080 59076 -3010
rect 59166 -3080 59176 -3010
rect 59066 -3090 59176 -3080
rect 59206 -3160 59256 -2960
rect 59376 -2590 59826 -2570
rect 59376 -2630 59476 -2590
rect 59656 -2630 59826 -2590
rect 59376 -2640 59826 -2630
rect 59376 -2690 59436 -2640
rect 59376 -3050 59386 -2690
rect 59426 -3050 59436 -2690
rect 59526 -2698 59576 -2670
rect 59526 -2732 59546 -2698
rect 59636 -2730 59706 -2670
rect 59580 -2732 59706 -2730
rect 59526 -2740 59706 -2732
rect 59476 -2782 59546 -2770
rect 59476 -2850 59502 -2782
rect 59476 -2958 59502 -2920
rect 59536 -2958 59546 -2782
rect 59476 -2970 59546 -2958
rect 59576 -2782 59636 -2770
rect 59576 -2790 59590 -2782
rect 59624 -2790 59636 -2782
rect 59576 -2970 59636 -2960
rect 59534 -3008 59592 -3002
rect 59534 -3010 59546 -3008
rect 59066 -3170 59176 -3160
rect 59066 -3240 59076 -3170
rect 59166 -3240 59176 -3170
rect 59066 -3242 59103 -3240
rect 59137 -3242 59176 -3240
rect 59066 -3250 59176 -3242
rect 59206 -3170 59266 -3160
rect 59206 -3250 59266 -3240
rect 59376 -3200 59436 -3050
rect 59516 -3042 59546 -3010
rect 59580 -3010 59592 -3008
rect 59666 -3010 59706 -2740
rect 59580 -3042 59706 -3010
rect 59516 -3080 59706 -3042
rect 59746 -2698 59936 -2670
rect 59746 -2732 59862 -2698
rect 59896 -2732 59936 -2698
rect 59746 -2740 59936 -2732
rect 61036 -2700 61206 -2520
rect 61346 -2700 61466 -2520
rect 61036 -2740 61466 -2700
rect 59746 -3000 59776 -2740
rect 60286 -2750 60476 -2740
rect 59806 -2782 59866 -2770
rect 59806 -2800 59818 -2782
rect 59852 -2800 59866 -2782
rect 59806 -2958 59818 -2940
rect 59852 -2958 59866 -2940
rect 59806 -2970 59866 -2958
rect 59900 -2780 60016 -2770
rect 59900 -2782 59916 -2780
rect 59900 -2958 59906 -2782
rect 59900 -2960 59916 -2958
rect 60006 -2960 60016 -2780
rect 60286 -2890 60306 -2750
rect 60456 -2890 60476 -2750
rect 61176 -2800 61386 -2780
rect 60286 -2900 60476 -2890
rect 61026 -2820 61136 -2810
rect 59900 -2970 60016 -2960
rect 60076 -2957 60196 -2920
rect 60076 -2991 60127 -2957
rect 60161 -2991 60196 -2957
rect 59746 -3008 59926 -3000
rect 59746 -3010 59862 -3008
rect 59896 -3010 59926 -3008
rect 59746 -3080 59826 -3010
rect 59916 -3080 59926 -3010
rect 59746 -3090 59926 -3080
rect 60076 -3049 60196 -2991
rect 60336 -2960 60446 -2900
rect 60336 -3000 60366 -2960
rect 60406 -3000 60446 -2960
rect 60636 -2957 60816 -2920
rect 60636 -2991 60671 -2957
rect 60705 -2991 60747 -2957
rect 60781 -2991 60816 -2957
rect 60076 -3080 60127 -3049
rect 60161 -3080 60196 -3049
rect 59736 -3170 59936 -3160
rect 58966 -3301 59086 -3280
rect 58966 -3677 59044 -3301
rect 59078 -3677 59086 -3301
rect 58966 -3690 59086 -3677
rect 59156 -3290 59202 -3289
rect 59156 -3301 59236 -3290
rect 59156 -3677 59162 -3301
rect 59196 -3330 59236 -3301
rect 59226 -3410 59236 -3330
rect 59196 -3560 59236 -3410
rect 59226 -3640 59236 -3560
rect 59196 -3677 59236 -3640
rect 59376 -3570 59386 -3200
rect 59426 -3570 59436 -3200
rect 59516 -3211 59706 -3170
rect 59516 -3245 59545 -3211
rect 59579 -3245 59706 -3211
rect 59516 -3250 59706 -3245
rect 59533 -3251 59591 -3250
rect 59466 -3295 59546 -3280
rect 59586 -3283 59646 -3280
rect 59466 -3330 59501 -3295
rect 59466 -3471 59501 -3410
rect 59535 -3471 59546 -3295
rect 59466 -3480 59546 -3471
rect 59583 -3295 59646 -3283
rect 59583 -3310 59589 -3295
rect 59623 -3310 59646 -3295
rect 59583 -3450 59586 -3310
rect 59583 -3471 59589 -3450
rect 59623 -3471 59646 -3450
rect 59583 -3480 59646 -3471
rect 59495 -3483 59541 -3480
rect 59583 -3483 59629 -3480
rect 59533 -3520 59591 -3515
rect 59676 -3520 59706 -3250
rect 59376 -3610 59436 -3570
rect 59506 -3580 59516 -3520
rect 59596 -3580 59706 -3520
rect 59736 -3240 59826 -3170
rect 59926 -3240 59936 -3170
rect 59736 -3245 59861 -3240
rect 59895 -3245 59936 -3240
rect 59736 -3250 59936 -3245
rect 60076 -3240 60096 -3080
rect 60176 -3240 60196 -3080
rect 59736 -3520 59766 -3250
rect 59849 -3251 59907 -3250
rect 60076 -3267 60127 -3240
rect 60161 -3267 60196 -3240
rect 59796 -3283 59856 -3280
rect 59796 -3290 59857 -3283
rect 59856 -3470 59857 -3290
rect 59796 -3471 59817 -3470
rect 59851 -3471 59857 -3470
rect 59796 -3480 59857 -3471
rect 59811 -3483 59857 -3480
rect 59899 -3290 59945 -3283
rect 59899 -3295 59916 -3290
rect 59899 -3471 59905 -3295
rect 59899 -3480 59916 -3471
rect 60006 -3480 60016 -3290
rect 60076 -3325 60196 -3267
rect 60346 -3050 60426 -3000
rect 60346 -3090 60366 -3050
rect 60406 -3090 60426 -3050
rect 60346 -3140 60426 -3090
rect 60346 -3180 60366 -3140
rect 60406 -3180 60426 -3140
rect 60346 -3220 60426 -3180
rect 60346 -3260 60366 -3220
rect 60406 -3260 60426 -3220
rect 60346 -3270 60426 -3260
rect 60636 -3049 60816 -2991
rect 60636 -3083 60671 -3049
rect 60705 -3083 60747 -3049
rect 60781 -3083 60816 -3049
rect 60636 -3141 60816 -3083
rect 60636 -3175 60671 -3141
rect 60705 -3175 60747 -3141
rect 60781 -3175 60816 -3141
rect 60636 -3233 60816 -3175
rect 60636 -3267 60671 -3233
rect 60705 -3267 60747 -3233
rect 60781 -3267 60816 -3233
rect 60076 -3359 60127 -3325
rect 60161 -3359 60196 -3325
rect 60076 -3390 60196 -3359
rect 60276 -3310 60546 -3300
rect 60276 -3325 60476 -3310
rect 60276 -3359 60297 -3325
rect 60331 -3359 60369 -3325
rect 60405 -3359 60449 -3325
rect 60276 -3370 60476 -3359
rect 60536 -3370 60546 -3310
rect 60276 -3380 60546 -3370
rect 60636 -3325 60816 -3267
rect 61026 -2930 61036 -2820
rect 61126 -2930 61136 -2820
rect 61176 -2880 61196 -2800
rect 61366 -2880 61386 -2800
rect 61176 -2900 61386 -2880
rect 61026 -2960 61136 -2930
rect 61026 -3000 61046 -2960
rect 61086 -3000 61136 -2960
rect 61026 -3050 61136 -3000
rect 61026 -3090 61046 -3050
rect 61086 -3090 61136 -3050
rect 61026 -3140 61136 -3090
rect 61026 -3180 61046 -3140
rect 61086 -3180 61136 -3140
rect 61026 -3220 61136 -3180
rect 61026 -3260 61046 -3220
rect 61086 -3260 61136 -3220
rect 61026 -3280 61136 -3260
rect 61256 -2957 61366 -2900
rect 61256 -2991 61291 -2957
rect 61325 -2991 61366 -2957
rect 61256 -3049 61366 -2991
rect 61256 -3050 61291 -3049
rect 61325 -3050 61366 -3049
rect 61256 -3260 61276 -3050
rect 61356 -3260 61366 -3050
rect 61256 -3267 61291 -3260
rect 61325 -3267 61366 -3260
rect 60636 -3359 60671 -3325
rect 60705 -3359 60747 -3325
rect 60781 -3359 60816 -3325
rect 60636 -3440 60816 -3359
rect 60966 -3324 61177 -3310
rect 60966 -3325 61129 -3324
rect 60966 -3359 60980 -3325
rect 61015 -3359 61053 -3325
rect 61088 -3358 61129 -3325
rect 61164 -3358 61177 -3324
rect 61088 -3359 61177 -3358
rect 60966 -3390 61177 -3359
rect 61256 -3325 61366 -3267
rect 61256 -3359 61291 -3325
rect 61325 -3359 61366 -3325
rect 61256 -3390 61366 -3359
rect 60466 -3450 60546 -3440
rect 59899 -3483 59945 -3480
rect 60466 -3510 60476 -3450
rect 60536 -3510 60546 -3450
rect 59849 -3520 59907 -3515
rect 60466 -3520 60546 -3510
rect 60606 -3450 60826 -3440
rect 60606 -3510 60616 -3450
rect 60736 -3510 60756 -3450
rect 60816 -3510 60826 -3450
rect 60606 -3520 60826 -3510
rect 60886 -3450 60966 -3440
rect 60886 -3510 60896 -3450
rect 60956 -3510 60966 -3450
rect 60886 -3520 60966 -3510
rect 59736 -3521 59926 -3520
rect 59736 -3555 59861 -3521
rect 59895 -3555 59926 -3521
rect 59736 -3580 59926 -3555
rect 60636 -3570 60816 -3520
rect 59376 -3620 59826 -3610
rect 59376 -3660 59476 -3620
rect 59646 -3660 59826 -3620
rect 59376 -3670 59826 -3660
rect 59156 -3690 59236 -3677
rect 58896 -3700 59086 -3690
rect 56380 -3768 57000 -3758
rect 57356 -3764 57676 -3750
rect 56440 -3774 57000 -3768
rect 57314 -3770 57676 -3764
rect 56440 -3794 57178 -3774
rect 56440 -3844 57118 -3794
rect 57168 -3844 57178 -3794
rect 57314 -3810 57326 -3770
rect 57376 -3810 57676 -3770
rect 57314 -3816 57676 -3810
rect 57356 -3830 57676 -3816
rect 56440 -3854 57178 -3844
rect 56440 -3888 57000 -3854
rect 57112 -3856 57174 -3854
rect 56380 -3958 57000 -3888
rect 56032 -4030 56038 -4028
rect 55992 -4042 56038 -4030
rect 55880 -4074 55970 -4068
rect 55870 -4078 55982 -4074
rect 55870 -4120 55880 -4078
rect 55970 -4120 55982 -4078
rect 55880 -4168 55970 -4158
rect 56120 -4198 56300 -4028
rect 57096 -4109 57372 -4078
rect 57096 -4143 57125 -4109
rect 57159 -4143 57217 -4109
rect 57251 -4143 57309 -4109
rect 57343 -4120 57372 -4109
rect 57343 -4143 57376 -4120
rect 57096 -4180 57376 -4143
rect 57066 -4190 57376 -4180
rect 56426 -4198 57376 -4190
rect 56120 -4208 57376 -4198
rect 56014 -4258 56086 -4246
rect 55570 -4378 55830 -4268
rect 53961 -4444 53988 -4406
rect 54022 -4444 54031 -4406
rect 53961 -4458 54031 -4444
rect 54910 -4406 54981 -4394
rect 54910 -4444 54916 -4406
rect 54950 -4444 54981 -4406
rect 54910 -4456 54981 -4444
rect 54911 -4458 54981 -4456
rect 55220 -4418 55330 -4408
rect 54069 -4472 54869 -4466
rect 54069 -4506 54081 -4472
rect 54857 -4478 54869 -4472
rect 54857 -4506 54880 -4478
rect 54069 -4512 54880 -4506
rect 54090 -4588 54880 -4512
rect 55330 -4518 55380 -4418
rect 55330 -4528 55480 -4518
rect 55220 -4538 55480 -4528
rect 55280 -4552 55480 -4538
rect 55280 -4558 55488 -4552
rect 55280 -4578 55300 -4558
rect 54090 -4688 54150 -4588
rect 54840 -4688 54880 -4588
rect 55288 -4592 55300 -4578
rect 55476 -4592 55488 -4558
rect 55530 -4578 55610 -4568
rect 55288 -4598 55488 -4592
rect 55520 -4602 55530 -4590
rect 55520 -4636 55526 -4602
rect 55288 -4646 55488 -4640
rect 55288 -4680 55300 -4646
rect 55476 -4680 55488 -4646
rect 55520 -4648 55530 -4636
rect 55530 -4678 55610 -4668
rect 55288 -4686 55488 -4680
rect 54090 -4708 54140 -4688
rect 54100 -4948 54140 -4708
rect 54850 -4948 54880 -4688
rect 55300 -4728 55470 -4686
rect 55300 -4868 55320 -4728
rect 55470 -4814 55482 -4742
rect 55300 -4878 55470 -4868
rect 54100 -4988 54880 -4948
rect 55710 -5198 55830 -4378
rect 56014 -4408 56020 -4258
rect 56080 -4408 56086 -4258
rect 56014 -4420 56086 -4408
rect 56120 -4408 56170 -4208
rect 56390 -4260 57376 -4208
rect 56390 -4268 57156 -4260
rect 56390 -4408 56654 -4268
rect 56120 -4458 56654 -4408
rect 56306 -4486 56654 -4458
rect 56998 -4420 57156 -4268
rect 57316 -4420 57376 -4260
rect 56998 -4486 57376 -4420
rect 56306 -4900 57376 -4486
rect 57556 -4610 57676 -3830
rect 58896 -3860 58986 -3700
rect 59756 -3720 59826 -3670
rect 59066 -3736 59176 -3730
rect 59066 -3740 59103 -3736
rect 59137 -3740 59176 -3736
rect 59066 -3800 59076 -3740
rect 59166 -3800 59176 -3740
rect 59066 -3810 59176 -3800
rect 58896 -4230 58926 -3860
rect 58966 -4230 58986 -3930
rect 59116 -3860 59506 -3840
rect 59116 -3930 59146 -3860
rect 59226 -3930 59276 -3860
rect 59356 -3930 59396 -3860
rect 59476 -3930 59506 -3860
rect 59116 -3948 59506 -3930
rect 59646 -3860 59716 -3840
rect 59706 -3920 59716 -3860
rect 59646 -3930 59716 -3920
rect 59113 -3954 59513 -3948
rect 59113 -3988 59125 -3954
rect 59501 -3988 59513 -3954
rect 59113 -3994 59513 -3988
rect 59546 -4000 59616 -3990
rect 59246 -4056 59256 -4030
rect 59113 -4062 59256 -4056
rect 59366 -4056 59376 -4030
rect 59366 -4062 59513 -4056
rect 59016 -4100 59076 -4080
rect 59113 -4096 59125 -4062
rect 59501 -4096 59513 -4062
rect 59606 -4060 59616 -4000
rect 59546 -4070 59616 -4060
rect 59113 -4102 59513 -4096
rect 59016 -4190 59076 -4160
rect 59113 -4170 59513 -4164
rect 59113 -4204 59125 -4170
rect 59501 -4204 59513 -4170
rect 59113 -4210 59513 -4204
rect 58896 -4300 58906 -4230
rect 58896 -4320 58986 -4300
rect 59116 -4230 59516 -4210
rect 59116 -4300 59146 -4230
rect 59226 -4300 59276 -4230
rect 59356 -4300 59396 -4230
rect 59476 -4300 59516 -4230
rect 59116 -4320 59516 -4300
rect 59646 -4230 59656 -3930
rect 59706 -4230 59716 -3930
rect 59756 -3900 59766 -3720
rect 59806 -3900 59826 -3720
rect 59956 -3720 60336 -3710
rect 59956 -3734 59966 -3720
rect 59946 -3740 59966 -3734
rect 60326 -3734 60336 -3720
rect 60326 -3740 60346 -3734
rect 59856 -3780 59916 -3770
rect 59946 -3774 59958 -3740
rect 60334 -3774 60346 -3740
rect 61056 -3740 61176 -3390
rect 59946 -3780 59966 -3774
rect 60326 -3780 60346 -3774
rect 60376 -3780 60436 -3760
rect 59956 -3790 60336 -3780
rect 59856 -3860 59916 -3840
rect 59946 -3848 60346 -3842
rect 59756 -3940 59826 -3900
rect 59946 -3882 59958 -3848
rect 60334 -3882 60346 -3848
rect 60376 -3860 60436 -3840
rect 61126 -3840 61176 -3740
rect 61056 -3870 61176 -3840
rect 59946 -3888 60346 -3882
rect 59946 -3940 60336 -3888
rect 59756 -3960 60536 -3940
rect 59756 -4000 59866 -3960
rect 60426 -4000 60536 -3960
rect 59756 -4010 60536 -4000
rect 59796 -4120 59806 -4010
rect 59916 -4120 59926 -4010
rect 59796 -4130 59926 -4120
rect 60436 -4030 60536 -4010
rect 60436 -4150 60446 -4030
rect 60526 -4150 60536 -4030
rect 60436 -4160 60536 -4150
rect 59646 -4240 59716 -4230
rect 59706 -4300 59716 -4240
rect 59646 -4320 59716 -4300
rect 58806 -4610 59356 -4580
rect 57556 -4620 59356 -4610
rect 57556 -4760 58986 -4620
rect 59126 -4760 59356 -4620
rect 59846 -4590 60256 -4580
rect 59846 -4700 59996 -4590
rect 60106 -4700 60256 -4590
rect 57556 -4810 59356 -4760
rect 58806 -4890 59356 -4810
rect 59600 -4900 60500 -4700
rect 55710 -5200 55910 -5198
rect 59600 -5200 59700 -4900
rect 60400 -5200 60500 -4900
rect 55500 -5300 56000 -5200
rect 59600 -5300 60500 -5200
rect 55500 -5600 55600 -5300
rect 55900 -5600 56000 -5300
rect 55500 -5700 56000 -5600
rect 55300 -6200 55800 -6100
rect 20800 -6600 22200 -6400
rect 55300 -6500 55400 -6200
rect 55700 -6500 55800 -6200
rect 55300 -6600 55800 -6500
rect 20800 -7400 21000 -6600
rect 22000 -7400 22200 -6600
rect 55576 -6638 55780 -6600
rect 55576 -6640 55776 -6638
rect 54090 -6738 54890 -6698
rect 53500 -6860 53800 -6840
rect 53500 -7120 53520 -6860
rect 53780 -7120 53800 -6860
rect 54090 -6868 54150 -6738
rect 54080 -6998 54150 -6868
rect 54860 -6978 54890 -6738
rect 54850 -6998 54890 -6978
rect 54080 -7066 54880 -6998
rect 54079 -7072 54880 -7066
rect 54079 -7106 54091 -7072
rect 54867 -7098 54880 -7072
rect 54867 -7106 54879 -7098
rect 54079 -7112 54879 -7106
rect 53500 -7140 53800 -7120
rect 53510 -7258 53800 -7140
rect 20800 -7482 22200 -7400
rect 53002 -7420 53480 -7358
rect 20800 -7600 21390 -7482
rect 21346 -7609 21390 -7600
rect 21380 -7612 21390 -7609
rect 21620 -7600 22200 -7482
rect 53000 -7558 53480 -7420
rect 53510 -7368 53520 -7258
rect 53640 -7368 53800 -7258
rect 53510 -7488 53800 -7368
rect 53970 -7134 54040 -7118
rect 53970 -7172 53998 -7134
rect 54032 -7172 54040 -7134
rect 53970 -7368 54040 -7172
rect 54920 -7134 54990 -7118
rect 54920 -7172 54926 -7134
rect 54960 -7172 54990 -7134
rect 54079 -7200 54879 -7194
rect 54079 -7234 54091 -7200
rect 54867 -7234 54879 -7200
rect 54079 -7238 54879 -7234
rect 54079 -7240 54750 -7238
rect 54090 -7288 54750 -7240
rect 54740 -7318 54750 -7288
rect 54850 -7240 54879 -7238
rect 54850 -7308 54860 -7240
rect 54840 -7318 54860 -7308
rect 54750 -7328 54860 -7318
rect 54920 -7368 54990 -7172
rect 55430 -7218 55520 -7208
rect 55290 -7328 55390 -7318
rect 53970 -7398 55290 -7368
rect 55430 -7358 55520 -7288
rect 53970 -7408 55390 -7398
rect 54050 -7418 55380 -7408
rect 54050 -7428 54880 -7418
rect 54050 -7438 54091 -7428
rect 54079 -7462 54091 -7438
rect 54867 -7438 54880 -7428
rect 54867 -7462 54879 -7438
rect 54079 -7468 54879 -7462
rect 54920 -7478 54990 -7468
rect 53510 -7506 53630 -7488
rect 53510 -7538 53526 -7506
rect 53514 -7540 53526 -7538
rect 53614 -7538 53630 -7506
rect 53940 -7490 54038 -7478
rect 53940 -7498 53998 -7490
rect 53614 -7540 53626 -7538
rect 53514 -7546 53626 -7540
rect 21620 -7609 21666 -7600
rect 21620 -7612 21630 -7609
rect 20886 -7775 22076 -7729
rect 20886 -7809 20908 -7775
rect 21076 -7809 21394 -7775
rect 21562 -7809 21880 -7775
rect 22048 -7809 22076 -7775
rect 20896 -7815 21088 -7809
rect 21382 -7815 21646 -7809
rect 21868 -7815 22060 -7809
rect 20840 -7859 20886 -7856
rect 21098 -7859 21144 -7856
rect 21326 -7859 21372 -7856
rect 20796 -7868 20886 -7859
rect 20796 -7875 20846 -7868
rect 20880 -7875 20886 -7868
rect 21096 -7868 21376 -7859
rect 20794 -11629 20804 -7875
rect 20880 -11629 20888 -7875
rect 20796 -11644 20846 -11629
rect 20880 -11644 20886 -11629
rect 20796 -11659 20886 -11644
rect 21096 -11644 21104 -7868
rect 21138 -7889 21332 -7868
rect 21138 -7969 21206 -7889
rect 21256 -7969 21332 -7889
rect 21138 -11479 21186 -7969
rect 21276 -11479 21332 -7969
rect 21138 -11619 21206 -11479
rect 21256 -11619 21332 -11479
rect 21138 -11644 21332 -11619
rect 21366 -11644 21376 -7868
rect 21096 -11649 21376 -11644
rect 21556 -7868 21646 -7815
rect 21812 -7859 21858 -7856
rect 21556 -11644 21590 -7868
rect 21624 -11644 21646 -7868
rect 21706 -7868 21858 -7859
rect 21706 -7877 21818 -7868
rect 21700 -7889 21818 -7877
rect 21700 -11629 21706 -7889
rect 21756 -7969 21818 -7889
rect 21816 -11479 21818 -7969
rect 21756 -11629 21818 -11479
rect 21700 -11641 21818 -11629
rect 21098 -11656 21144 -11649
rect 21326 -11656 21372 -11649
rect 21556 -11697 21646 -11644
rect 21706 -11644 21818 -11641
rect 21852 -11644 21858 -7868
rect 22070 -7868 22116 -7856
rect 22070 -7872 22076 -7868
rect 22110 -7872 22116 -7868
rect 22060 -11632 22070 -7872
rect 22140 -11632 22150 -7872
rect 53000 -9308 53050 -7558
rect 53250 -7568 53480 -7558
rect 53250 -8918 53330 -7568
rect 53400 -7578 53480 -7568
rect 53400 -7590 53504 -7578
rect 53400 -8366 53464 -7590
rect 53498 -8366 53504 -7590
rect 53400 -8378 53504 -8366
rect 53636 -7588 53682 -7578
rect 53636 -7590 53760 -7588
rect 53636 -8366 53642 -7590
rect 53676 -8366 53760 -7590
rect 53940 -7598 53950 -7498
rect 54032 -7528 54038 -7490
rect 54020 -7540 54038 -7528
rect 54020 -7598 54030 -7540
rect 54079 -7556 54879 -7550
rect 54079 -7590 54091 -7556
rect 54867 -7590 54879 -7556
rect 54920 -7578 54990 -7568
rect 55320 -7568 55380 -7418
rect 54079 -7596 54879 -7590
rect 53940 -7618 54030 -7598
rect 54090 -7628 54870 -7596
rect 55320 -7602 55334 -7568
rect 55368 -7602 55380 -7568
rect 55320 -7608 55380 -7602
rect 53840 -7928 53920 -7918
rect 53840 -8038 53860 -7928
rect 53840 -8048 53920 -8038
rect 53840 -8240 53900 -8048
rect 54320 -8128 54510 -7628
rect 55440 -7638 55520 -7358
rect 55410 -7640 55520 -7638
rect 55284 -7648 55330 -7640
rect 55230 -7652 55330 -7648
rect 55230 -7658 55290 -7652
rect 55324 -7828 55330 -7652
rect 55230 -7838 55330 -7828
rect 55284 -7840 55330 -7838
rect 55372 -7648 55520 -7640
rect 55372 -7652 55430 -7648
rect 55372 -7828 55378 -7652
rect 55412 -7818 55430 -7652
rect 55510 -7818 55520 -7648
rect 55412 -7828 55520 -7818
rect 55372 -7840 55418 -7828
rect 55580 -7928 55720 -6640
rect 58776 -6870 59306 -6750
rect 58776 -6880 58966 -6870
rect 56146 -6980 57366 -6930
rect 55954 -7128 56046 -7116
rect 56146 -7128 56506 -6980
rect 55954 -7298 55960 -7128
rect 56040 -7298 56046 -7128
rect 55954 -7310 56046 -7298
rect 56120 -7158 56506 -7128
rect 56120 -7368 56190 -7158
rect 56390 -7230 56506 -7158
rect 57016 -7134 57366 -6980
rect 57586 -7030 58966 -6880
rect 59126 -7030 59306 -6870
rect 57586 -7050 59306 -7030
rect 59946 -6900 60386 -6800
rect 57586 -7080 58986 -7050
rect 59946 -7060 59956 -6900
rect 60166 -7060 60386 -6900
rect 57016 -7230 57368 -7134
rect 56390 -7270 57368 -7230
rect 56390 -7368 57126 -7270
rect 56120 -7374 57126 -7368
rect 56120 -7378 56750 -7374
rect 55880 -7418 55970 -7408
rect 55870 -7496 55880 -7450
rect 55970 -7496 55982 -7450
rect 55880 -7508 55970 -7498
rect 55000 -7938 55090 -7928
rect 55000 -8048 55090 -8038
rect 54710 -8128 54960 -8108
rect 53940 -8168 54960 -8128
rect 53940 -8172 54730 -8168
rect 53930 -8178 54730 -8172
rect 53930 -8212 53942 -8178
rect 54718 -8212 54730 -8178
rect 53930 -8218 54730 -8212
rect 53840 -8328 53858 -8240
rect 53892 -8328 53900 -8240
rect 53840 -8348 53900 -8328
rect 54762 -8238 54850 -8228
rect 54762 -8240 54770 -8238
rect 54762 -8328 54768 -8240
rect 54840 -8328 54850 -8238
rect 54762 -8340 54850 -8328
rect 54770 -8348 54850 -8340
rect 53636 -8378 53760 -8366
rect 53400 -8596 53480 -8378
rect 53514 -8416 53626 -8410
rect 53514 -8418 53526 -8416
rect 53510 -8450 53526 -8418
rect 53614 -8418 53626 -8416
rect 53614 -8450 53630 -8418
rect 53510 -8524 53630 -8450
rect 53510 -8558 53526 -8524
rect 53614 -8558 53630 -8524
rect 53680 -8438 53760 -8378
rect 53930 -8356 54730 -8350
rect 53930 -8390 53942 -8356
rect 54718 -8390 54730 -8356
rect 53930 -8396 54730 -8390
rect 53940 -8428 54720 -8396
rect 53920 -8438 54720 -8428
rect 53680 -8528 54720 -8438
rect 53514 -8564 53626 -8558
rect 53680 -8596 53760 -8528
rect 53920 -8538 54720 -8528
rect 53940 -8578 54720 -8538
rect 54900 -8568 54960 -8168
rect 55010 -8160 55090 -8048
rect 55540 -7938 55720 -7928
rect 55630 -8038 55720 -7938
rect 55130 -8074 55506 -8068
rect 55130 -8108 55142 -8074
rect 55494 -8108 55506 -8074
rect 55130 -8114 55506 -8108
rect 55010 -8194 55046 -8160
rect 55080 -8194 55090 -8160
rect 55010 -8208 55090 -8194
rect 55142 -8240 55494 -8114
rect 55540 -8160 55720 -8038
rect 55540 -8194 55556 -8160
rect 55590 -8194 55720 -8160
rect 55540 -8208 55720 -8194
rect 55780 -7540 55860 -7528
rect 55130 -8246 55506 -8240
rect 55130 -8280 55142 -8246
rect 55494 -8278 55506 -8246
rect 55494 -8280 55510 -8278
rect 55130 -8286 55510 -8280
rect 55140 -8298 55510 -8286
rect 55780 -8298 55820 -7540
rect 55140 -8316 55820 -8298
rect 55854 -8316 55860 -7540
rect 55140 -8328 55860 -8316
rect 55992 -7540 56038 -7528
rect 55992 -8316 55998 -7540
rect 56032 -7548 56038 -7540
rect 56120 -7548 56300 -7378
rect 57098 -7400 57126 -7374
rect 57356 -7400 57368 -7270
rect 57098 -7414 57368 -7400
rect 57096 -7445 57372 -7414
rect 57096 -7479 57125 -7445
rect 57159 -7479 57217 -7445
rect 57251 -7479 57309 -7445
rect 57343 -7479 57372 -7445
rect 57096 -7510 57372 -7479
rect 56032 -7906 56300 -7548
rect 56590 -7668 56660 -7658
rect 56660 -7734 57000 -7668
rect 57586 -7730 57706 -7080
rect 59946 -7090 60386 -7060
rect 57366 -7734 57706 -7730
rect 56660 -7738 57188 -7734
rect 56660 -7744 57190 -7738
rect 56660 -7794 57118 -7744
rect 57178 -7794 57190 -7744
rect 57314 -7740 57706 -7734
rect 57314 -7780 57326 -7740
rect 57366 -7780 57706 -7740
rect 57314 -7786 57706 -7780
rect 57366 -7790 57706 -7786
rect 58896 -7370 58986 -7350
rect 58896 -7430 58906 -7370
rect 58896 -7720 58926 -7430
rect 58966 -7720 58986 -7370
rect 59106 -7370 59516 -7360
rect 59106 -7430 59216 -7370
rect 59276 -7430 59326 -7370
rect 59386 -7430 59436 -7370
rect 59496 -7430 59516 -7370
rect 59106 -7447 59516 -7430
rect 59626 -7370 59706 -7330
rect 59626 -7430 59636 -7370
rect 59626 -7440 59656 -7430
rect 59106 -7480 59125 -7447
rect 59113 -7481 59125 -7480
rect 59501 -7480 59516 -7447
rect 59501 -7481 59513 -7480
rect 59113 -7487 59513 -7481
rect 59546 -7490 59616 -7480
rect 59276 -7530 59356 -7520
rect 59276 -7549 59286 -7530
rect 59113 -7555 59286 -7549
rect 59346 -7549 59356 -7530
rect 59346 -7555 59513 -7549
rect 59113 -7589 59125 -7555
rect 59501 -7589 59513 -7555
rect 59606 -7550 59616 -7490
rect 59546 -7560 59616 -7550
rect 59113 -7590 59286 -7589
rect 59346 -7590 59513 -7589
rect 59016 -7600 59076 -7590
rect 59113 -7595 59513 -7590
rect 59276 -7600 59356 -7595
rect 59546 -7610 59616 -7600
rect 59016 -7670 59076 -7660
rect 59113 -7663 59513 -7657
rect 59113 -7697 59125 -7663
rect 59501 -7697 59513 -7663
rect 59606 -7670 59616 -7610
rect 59546 -7680 59616 -7670
rect 59113 -7700 59513 -7697
rect 59113 -7703 59516 -7700
rect 58896 -7730 58986 -7720
rect 58896 -7790 58906 -7730
rect 58966 -7790 58986 -7730
rect 58896 -7792 58986 -7790
rect 59116 -7720 59516 -7703
rect 59646 -7710 59656 -7440
rect 59116 -7780 59216 -7720
rect 59276 -7780 59336 -7720
rect 59396 -7780 59436 -7720
rect 59496 -7780 59516 -7720
rect 56660 -7798 57190 -7794
rect 56590 -7800 57190 -7798
rect 56590 -7804 57188 -7800
rect 56590 -7868 57000 -7804
rect 56032 -7918 56356 -7906
rect 56032 -8316 56280 -7918
rect 55992 -8328 56280 -8316
rect 55140 -8338 55200 -8328
rect 55450 -8358 55810 -8328
rect 55870 -8366 55982 -8360
rect 55870 -8400 55882 -8366
rect 55970 -8400 55982 -8366
rect 55870 -8406 55982 -8400
rect 55140 -8418 55200 -8408
rect 55024 -8448 55116 -8436
rect 55024 -8528 55030 -8448
rect 55110 -8528 55116 -8448
rect 55024 -8540 55116 -8528
rect 55734 -8448 55816 -8436
rect 55734 -8528 55740 -8448
rect 55810 -8528 55816 -8448
rect 55734 -8540 55816 -8528
rect 55880 -8438 55970 -8406
rect 55880 -8564 55970 -8528
rect 56060 -8548 56280 -8328
rect 56350 -8548 56356 -7918
rect 56480 -7988 56550 -7978
rect 56480 -8058 56550 -8048
rect 56590 -8087 56750 -7868
rect 58894 -7886 58988 -7792
rect 59116 -7800 59516 -7780
rect 59636 -7720 59656 -7710
rect 59696 -7720 59706 -7370
rect 59856 -7540 59976 -7530
rect 59856 -7630 59866 -7540
rect 59966 -7630 59976 -7540
rect 59856 -7640 59976 -7630
rect 60436 -7620 60446 -7520
rect 60526 -7620 60536 -7520
rect 60436 -7640 60536 -7620
rect 59636 -7730 59706 -7720
rect 59696 -7790 59706 -7730
rect 59636 -7810 59706 -7790
rect 59756 -7660 60536 -7640
rect 59756 -7700 59866 -7660
rect 60426 -7700 60536 -7660
rect 59756 -7710 60536 -7700
rect 59756 -7750 59826 -7710
rect 59066 -7840 59176 -7830
rect 58896 -7950 58986 -7886
rect 59066 -7910 59076 -7840
rect 59166 -7910 59176 -7840
rect 59066 -7912 59103 -7910
rect 59137 -7912 59176 -7910
rect 59066 -7920 59176 -7912
rect 59756 -7940 59766 -7750
rect 59806 -7940 59826 -7750
rect 59956 -7768 60046 -7740
rect 59946 -7774 60046 -7768
rect 60126 -7768 60336 -7740
rect 60126 -7774 60346 -7768
rect 59856 -7810 59916 -7800
rect 59946 -7808 59958 -7774
rect 60334 -7808 60346 -7774
rect 59946 -7814 60346 -7808
rect 60376 -7820 60446 -7810
rect 59856 -7890 59916 -7880
rect 59946 -7882 60346 -7876
rect 59946 -7916 59958 -7882
rect 60334 -7916 60346 -7882
rect 60376 -7890 60446 -7880
rect 59946 -7922 59976 -7916
rect 57098 -7958 57368 -7954
rect 57096 -7964 57372 -7958
rect 57096 -8050 57098 -7964
rect 56424 -8088 56470 -8087
rect 56060 -8560 56356 -8548
rect 56410 -8099 56470 -8088
rect 53400 -8608 53504 -8596
rect 53400 -8918 53464 -8608
rect 53250 -9308 53464 -8918
rect 53000 -9384 53464 -9308
rect 53498 -9384 53504 -8608
rect 53000 -9388 53504 -9384
rect 53458 -9396 53504 -9388
rect 53636 -8608 53760 -8596
rect 53636 -9384 53642 -8608
rect 53676 -9384 53760 -8608
rect 53930 -8584 54730 -8578
rect 53930 -8618 53942 -8584
rect 54718 -8618 54730 -8584
rect 53930 -8624 54730 -8618
rect 53830 -8646 53900 -8628
rect 53830 -8734 53858 -8646
rect 53892 -8734 53900 -8646
rect 53830 -8928 53900 -8734
rect 54760 -8646 54850 -8628
rect 54760 -8734 54768 -8646
rect 54802 -8648 54850 -8646
rect 54900 -8638 55200 -8568
rect 55870 -8570 55982 -8564
rect 55870 -8604 55882 -8570
rect 55970 -8604 55982 -8570
rect 55450 -8638 55810 -8608
rect 55870 -8610 55982 -8604
rect 56060 -8638 56300 -8560
rect 54900 -8642 55820 -8638
rect 56000 -8642 56300 -8638
rect 54900 -8648 55860 -8642
rect 54840 -8728 54850 -8648
rect 54802 -8734 54850 -8728
rect 54760 -8748 54850 -8734
rect 55130 -8654 55860 -8648
rect 55130 -8678 55820 -8654
rect 55130 -8696 55510 -8678
rect 55130 -8730 55142 -8696
rect 55494 -8698 55510 -8696
rect 55494 -8730 55506 -8698
rect 55130 -8736 55506 -8730
rect 53930 -8762 54730 -8756
rect 53930 -8796 53942 -8762
rect 54718 -8796 54730 -8762
rect 55020 -8782 55090 -8768
rect 53930 -8802 54730 -8796
rect 53940 -8808 54730 -8802
rect 54920 -8798 54980 -8788
rect 53940 -8848 54920 -8808
rect 53830 -8938 53920 -8928
rect 53830 -9048 53850 -8938
rect 53830 -9058 53920 -9048
rect 54320 -9348 54510 -8848
rect 54710 -8868 54920 -8848
rect 54910 -8878 54980 -8868
rect 55020 -8816 55046 -8782
rect 55080 -8816 55090 -8782
rect 55020 -8928 55090 -8816
rect 55142 -8862 55494 -8736
rect 55540 -8782 55620 -8768
rect 55540 -8816 55556 -8782
rect 55590 -8816 55620 -8782
rect 55130 -8868 55506 -8862
rect 55130 -8902 55142 -8868
rect 55494 -8902 55506 -8868
rect 55130 -8908 55506 -8902
rect 55000 -8938 55090 -8928
rect 55000 -9048 55090 -9038
rect 55540 -8928 55620 -8816
rect 55540 -8938 55630 -8928
rect 55630 -9038 55680 -8948
rect 55540 -9048 55680 -9038
rect 55274 -9138 55320 -9136
rect 55220 -9148 55320 -9138
rect 55220 -9324 55280 -9318
rect 55314 -9324 55320 -9148
rect 55220 -9328 55320 -9324
rect 55274 -9336 55320 -9328
rect 55362 -9148 55408 -9136
rect 55362 -9324 55368 -9148
rect 55402 -9158 55510 -9148
rect 55402 -9324 55410 -9158
rect 55362 -9328 55410 -9324
rect 55500 -9328 55510 -9158
rect 55362 -9336 55510 -9328
rect 55390 -9338 55510 -9336
rect 53636 -9388 53760 -9384
rect 53636 -9396 53682 -9388
rect 53940 -9408 54020 -9368
rect 54080 -9382 54860 -9348
rect 55311 -9374 55371 -9368
rect 53514 -9434 53626 -9428
rect 53514 -9438 53526 -9434
rect 53510 -9468 53526 -9438
rect 53614 -9438 53626 -9434
rect 53614 -9468 53630 -9438
rect 53510 -9528 53630 -9468
rect 53940 -9488 53950 -9408
rect 54010 -9438 54020 -9408
rect 54069 -9388 54869 -9382
rect 54069 -9422 54081 -9388
rect 54857 -9422 54869 -9388
rect 54069 -9428 54869 -9422
rect 54910 -9398 54980 -9388
rect 54010 -9450 54028 -9438
rect 54022 -9488 54028 -9450
rect 53940 -9500 54028 -9488
rect 53940 -9508 54020 -9500
rect 54910 -9508 54980 -9498
rect 55311 -9408 55324 -9374
rect 55358 -9408 55371 -9374
rect 54070 -9510 54870 -9508
rect 54069 -9516 54870 -9510
rect 54069 -9538 54081 -9516
rect 54041 -9550 54081 -9538
rect 54857 -9518 54870 -9516
rect 54857 -9550 54880 -9518
rect 55311 -9548 55371 -9408
rect 54041 -9558 54880 -9550
rect 55240 -9558 55371 -9548
rect 54041 -9568 55240 -9558
rect 53510 -9658 53630 -9648
rect 53961 -9608 55240 -9568
rect 53961 -9806 54031 -9608
rect 54730 -9668 54860 -9658
rect 54730 -9688 54740 -9668
rect 54080 -9738 54740 -9688
rect 54069 -9744 54740 -9738
rect 54850 -9738 54860 -9668
rect 54850 -9744 54869 -9738
rect 54069 -9778 54081 -9744
rect 54857 -9778 54869 -9744
rect 54069 -9784 54869 -9778
rect 54911 -9794 54981 -9608
rect 55370 -9608 55371 -9558
rect 55240 -9628 55370 -9618
rect 55410 -9648 55510 -9338
rect 55410 -9758 55510 -9738
rect 55570 -9668 55680 -9048
rect 55780 -9430 55820 -8678
rect 55854 -9430 55860 -8654
rect 55780 -9438 55860 -9430
rect 55814 -9442 55860 -9438
rect 55992 -8654 56300 -8642
rect 55992 -9430 55998 -8654
rect 56032 -9428 56300 -8654
rect 56410 -8698 56430 -8099
rect 56380 -8875 56430 -8698
rect 56464 -8875 56470 -8099
rect 56380 -8887 56470 -8875
rect 56552 -8099 56750 -8087
rect 56552 -8875 56558 -8099
rect 56592 -8238 56750 -8099
rect 57066 -8080 57098 -8050
rect 57368 -8050 57372 -7964
rect 58896 -7959 59076 -7950
rect 58896 -7960 59084 -7959
rect 59156 -7960 59202 -7959
rect 57368 -8080 57396 -8050
rect 57066 -8210 57086 -8080
rect 57376 -8210 57396 -8080
rect 56592 -8875 56610 -8238
rect 57066 -8240 57396 -8210
rect 56860 -8390 57060 -8378
rect 56860 -8418 57236 -8390
rect 56860 -8548 56900 -8418
rect 57020 -8548 57236 -8418
rect 56860 -8588 57236 -8548
rect 57036 -8590 57236 -8588
rect 58556 -8480 58756 -8460
rect 58556 -8640 58576 -8480
rect 58736 -8640 58756 -8480
rect 58556 -8660 58756 -8640
rect 56552 -8878 56610 -8875
rect 57036 -8740 57446 -8730
rect 56552 -8887 56598 -8878
rect 57036 -8880 57056 -8740
rect 57416 -8880 57446 -8740
rect 56380 -9158 56440 -8887
rect 57036 -8900 57098 -8880
rect 56480 -8928 56550 -8918
rect 56480 -8998 56550 -8988
rect 57096 -9014 57098 -8934
rect 57368 -8900 57446 -8880
rect 57368 -9014 57372 -8934
rect 57096 -9030 57372 -9014
rect 58896 -9090 58926 -7960
rect 58966 -7971 59086 -7960
rect 58966 -8347 59044 -7971
rect 59078 -8347 59086 -7971
rect 58966 -8370 59086 -8347
rect 59156 -7971 59256 -7960
rect 59756 -7970 59826 -7940
rect 59966 -7952 59976 -7922
rect 60316 -7922 60346 -7916
rect 61036 -7920 61466 -7910
rect 60316 -7952 60326 -7922
rect 59966 -7960 60326 -7952
rect 59156 -8347 59162 -7971
rect 59196 -8040 59256 -7971
rect 59236 -8120 59256 -8040
rect 59196 -8240 59256 -8120
rect 59236 -8320 59256 -8240
rect 59196 -8347 59256 -8320
rect 59156 -8360 59256 -8347
rect 58966 -8680 59036 -8370
rect 59066 -8406 59176 -8400
rect 59066 -8410 59103 -8406
rect 59137 -8410 59176 -8406
rect 59066 -8480 59076 -8410
rect 59166 -8480 59176 -8410
rect 59066 -8490 59176 -8480
rect 59206 -8560 59256 -8360
rect 59376 -7990 59826 -7970
rect 59376 -8030 59476 -7990
rect 59656 -8030 59826 -7990
rect 59376 -8040 59826 -8030
rect 59376 -8090 59436 -8040
rect 59376 -8450 59386 -8090
rect 59426 -8450 59436 -8090
rect 59526 -8098 59576 -8070
rect 59526 -8132 59546 -8098
rect 59636 -8130 59706 -8070
rect 59580 -8132 59706 -8130
rect 59526 -8140 59706 -8132
rect 59476 -8182 59546 -8170
rect 59476 -8250 59502 -8182
rect 59476 -8358 59502 -8320
rect 59536 -8358 59546 -8182
rect 59476 -8370 59546 -8358
rect 59576 -8182 59636 -8170
rect 59576 -8190 59590 -8182
rect 59624 -8190 59636 -8182
rect 59576 -8370 59636 -8360
rect 59534 -8408 59592 -8402
rect 59534 -8410 59546 -8408
rect 59066 -8570 59176 -8560
rect 59066 -8640 59076 -8570
rect 59166 -8640 59176 -8570
rect 59066 -8642 59103 -8640
rect 59137 -8642 59176 -8640
rect 59066 -8650 59176 -8642
rect 59206 -8570 59266 -8560
rect 59206 -8650 59266 -8640
rect 59376 -8600 59436 -8450
rect 59516 -8442 59546 -8410
rect 59580 -8410 59592 -8408
rect 59666 -8410 59706 -8140
rect 59580 -8442 59706 -8410
rect 59516 -8480 59706 -8442
rect 59746 -8098 59936 -8070
rect 59746 -8132 59862 -8098
rect 59896 -8132 59936 -8098
rect 59746 -8140 59936 -8132
rect 61036 -8100 61206 -7920
rect 61346 -8100 61466 -7920
rect 61036 -8140 61466 -8100
rect 59746 -8400 59776 -8140
rect 60286 -8150 60476 -8140
rect 59806 -8182 59866 -8170
rect 59806 -8200 59818 -8182
rect 59852 -8200 59866 -8182
rect 59806 -8358 59818 -8340
rect 59852 -8358 59866 -8340
rect 59806 -8370 59866 -8358
rect 59900 -8180 60016 -8170
rect 59900 -8182 59916 -8180
rect 59900 -8358 59906 -8182
rect 59900 -8360 59916 -8358
rect 60006 -8360 60016 -8180
rect 60286 -8290 60306 -8150
rect 60456 -8290 60476 -8150
rect 61176 -8200 61386 -8180
rect 60286 -8300 60476 -8290
rect 61026 -8220 61136 -8210
rect 59900 -8370 60016 -8360
rect 60076 -8357 60196 -8320
rect 60076 -8391 60127 -8357
rect 60161 -8391 60196 -8357
rect 59746 -8408 59926 -8400
rect 59746 -8410 59862 -8408
rect 59896 -8410 59926 -8408
rect 59746 -8480 59826 -8410
rect 59916 -8480 59926 -8410
rect 59746 -8490 59926 -8480
rect 60076 -8449 60196 -8391
rect 60336 -8360 60446 -8300
rect 60336 -8400 60366 -8360
rect 60406 -8400 60446 -8360
rect 60636 -8357 60816 -8320
rect 60636 -8391 60671 -8357
rect 60705 -8391 60747 -8357
rect 60781 -8391 60816 -8357
rect 60076 -8480 60127 -8449
rect 60161 -8480 60196 -8449
rect 59736 -8570 59936 -8560
rect 58966 -8701 59086 -8680
rect 58966 -9077 59044 -8701
rect 59078 -9077 59086 -8701
rect 58966 -9090 59086 -9077
rect 59156 -8690 59202 -8689
rect 59156 -8701 59236 -8690
rect 59156 -9077 59162 -8701
rect 59196 -8730 59236 -8701
rect 59226 -8810 59236 -8730
rect 59196 -8960 59236 -8810
rect 59226 -9040 59236 -8960
rect 59196 -9077 59236 -9040
rect 59376 -8970 59386 -8600
rect 59426 -8970 59436 -8600
rect 59516 -8611 59706 -8570
rect 59516 -8645 59545 -8611
rect 59579 -8645 59706 -8611
rect 59516 -8650 59706 -8645
rect 59533 -8651 59591 -8650
rect 59466 -8695 59546 -8680
rect 59586 -8683 59646 -8680
rect 59466 -8730 59501 -8695
rect 59466 -8871 59501 -8810
rect 59535 -8871 59546 -8695
rect 59466 -8880 59546 -8871
rect 59583 -8695 59646 -8683
rect 59583 -8710 59589 -8695
rect 59623 -8710 59646 -8695
rect 59583 -8850 59586 -8710
rect 59583 -8871 59589 -8850
rect 59623 -8871 59646 -8850
rect 59583 -8880 59646 -8871
rect 59495 -8883 59541 -8880
rect 59583 -8883 59629 -8880
rect 59533 -8920 59591 -8915
rect 59676 -8920 59706 -8650
rect 59376 -9010 59436 -8970
rect 59506 -8980 59516 -8920
rect 59596 -8980 59706 -8920
rect 59736 -8640 59826 -8570
rect 59926 -8640 59936 -8570
rect 59736 -8645 59861 -8640
rect 59895 -8645 59936 -8640
rect 59736 -8650 59936 -8645
rect 60076 -8640 60096 -8480
rect 60176 -8640 60196 -8480
rect 59736 -8920 59766 -8650
rect 59849 -8651 59907 -8650
rect 60076 -8667 60127 -8640
rect 60161 -8667 60196 -8640
rect 59796 -8683 59856 -8680
rect 59796 -8690 59857 -8683
rect 59856 -8870 59857 -8690
rect 59796 -8871 59817 -8870
rect 59851 -8871 59857 -8870
rect 59796 -8880 59857 -8871
rect 59811 -8883 59857 -8880
rect 59899 -8690 59945 -8683
rect 59899 -8695 59916 -8690
rect 59899 -8871 59905 -8695
rect 59899 -8880 59916 -8871
rect 60006 -8880 60016 -8690
rect 60076 -8725 60196 -8667
rect 60346 -8450 60426 -8400
rect 60346 -8490 60366 -8450
rect 60406 -8490 60426 -8450
rect 60346 -8540 60426 -8490
rect 60346 -8580 60366 -8540
rect 60406 -8580 60426 -8540
rect 60346 -8620 60426 -8580
rect 60346 -8660 60366 -8620
rect 60406 -8660 60426 -8620
rect 60346 -8670 60426 -8660
rect 60636 -8449 60816 -8391
rect 60636 -8483 60671 -8449
rect 60705 -8483 60747 -8449
rect 60781 -8483 60816 -8449
rect 60636 -8541 60816 -8483
rect 60636 -8575 60671 -8541
rect 60705 -8575 60747 -8541
rect 60781 -8575 60816 -8541
rect 60636 -8633 60816 -8575
rect 60636 -8667 60671 -8633
rect 60705 -8667 60747 -8633
rect 60781 -8667 60816 -8633
rect 60076 -8759 60127 -8725
rect 60161 -8759 60196 -8725
rect 60076 -8790 60196 -8759
rect 60276 -8710 60546 -8700
rect 60276 -8725 60476 -8710
rect 60276 -8759 60297 -8725
rect 60331 -8759 60369 -8725
rect 60405 -8759 60449 -8725
rect 60276 -8770 60476 -8759
rect 60536 -8770 60546 -8710
rect 60276 -8780 60546 -8770
rect 60636 -8725 60816 -8667
rect 61026 -8330 61036 -8220
rect 61126 -8330 61136 -8220
rect 61176 -8280 61196 -8200
rect 61366 -8280 61386 -8200
rect 61176 -8300 61386 -8280
rect 61026 -8360 61136 -8330
rect 61026 -8400 61046 -8360
rect 61086 -8400 61136 -8360
rect 61026 -8450 61136 -8400
rect 61026 -8490 61046 -8450
rect 61086 -8490 61136 -8450
rect 61026 -8540 61136 -8490
rect 61026 -8580 61046 -8540
rect 61086 -8580 61136 -8540
rect 61026 -8620 61136 -8580
rect 61026 -8660 61046 -8620
rect 61086 -8660 61136 -8620
rect 61026 -8680 61136 -8660
rect 61256 -8357 61366 -8300
rect 61256 -8391 61291 -8357
rect 61325 -8391 61366 -8357
rect 61256 -8449 61366 -8391
rect 61256 -8450 61291 -8449
rect 61325 -8450 61366 -8449
rect 61256 -8660 61276 -8450
rect 61356 -8660 61366 -8450
rect 61256 -8667 61291 -8660
rect 61325 -8667 61366 -8660
rect 60636 -8759 60671 -8725
rect 60705 -8759 60747 -8725
rect 60781 -8759 60816 -8725
rect 60636 -8840 60816 -8759
rect 60966 -8724 61177 -8710
rect 60966 -8725 61129 -8724
rect 60966 -8759 60980 -8725
rect 61015 -8759 61053 -8725
rect 61088 -8758 61129 -8725
rect 61164 -8758 61177 -8724
rect 61088 -8759 61177 -8758
rect 60966 -8790 61177 -8759
rect 61256 -8725 61366 -8667
rect 61256 -8759 61291 -8725
rect 61325 -8759 61366 -8725
rect 61256 -8790 61366 -8759
rect 60466 -8850 60546 -8840
rect 59899 -8883 59945 -8880
rect 60466 -8910 60476 -8850
rect 60536 -8910 60546 -8850
rect 59849 -8920 59907 -8915
rect 60466 -8920 60546 -8910
rect 60606 -8850 60826 -8840
rect 60606 -8910 60616 -8850
rect 60736 -8910 60756 -8850
rect 60816 -8910 60826 -8850
rect 60606 -8920 60826 -8910
rect 60886 -8850 60966 -8840
rect 60886 -8910 60896 -8850
rect 60956 -8910 60966 -8850
rect 60886 -8920 60966 -8910
rect 59736 -8921 59926 -8920
rect 59736 -8955 59861 -8921
rect 59895 -8955 59926 -8921
rect 59736 -8980 59926 -8955
rect 60636 -8970 60816 -8920
rect 59376 -9020 59826 -9010
rect 59376 -9060 59476 -9020
rect 59646 -9060 59826 -9020
rect 59376 -9070 59826 -9060
rect 59156 -9090 59236 -9077
rect 58896 -9100 59086 -9090
rect 56380 -9168 57000 -9158
rect 57356 -9164 57676 -9150
rect 56440 -9174 57000 -9168
rect 57314 -9170 57676 -9164
rect 56440 -9194 57178 -9174
rect 56440 -9244 57118 -9194
rect 57168 -9244 57178 -9194
rect 57314 -9210 57326 -9170
rect 57376 -9210 57676 -9170
rect 57314 -9216 57676 -9210
rect 57356 -9230 57676 -9216
rect 56440 -9254 57178 -9244
rect 56440 -9288 57000 -9254
rect 57112 -9256 57174 -9254
rect 56380 -9358 57000 -9288
rect 56032 -9430 56038 -9428
rect 55992 -9442 56038 -9430
rect 55880 -9474 55970 -9468
rect 55870 -9478 55982 -9474
rect 55870 -9520 55880 -9478
rect 55970 -9520 55982 -9478
rect 55880 -9568 55970 -9558
rect 56120 -9598 56300 -9428
rect 57096 -9509 57372 -9478
rect 57096 -9543 57125 -9509
rect 57159 -9543 57217 -9509
rect 57251 -9543 57309 -9509
rect 57343 -9520 57372 -9509
rect 57343 -9543 57376 -9520
rect 57096 -9580 57376 -9543
rect 57066 -9590 57376 -9580
rect 56426 -9598 57376 -9590
rect 56120 -9608 57376 -9598
rect 56014 -9658 56086 -9646
rect 55570 -9778 55830 -9668
rect 53961 -9844 53988 -9806
rect 54022 -9844 54031 -9806
rect 53961 -9858 54031 -9844
rect 54910 -9806 54981 -9794
rect 54910 -9844 54916 -9806
rect 54950 -9844 54981 -9806
rect 54910 -9856 54981 -9844
rect 54911 -9858 54981 -9856
rect 55220 -9818 55330 -9808
rect 54069 -9872 54869 -9866
rect 54069 -9906 54081 -9872
rect 54857 -9878 54869 -9872
rect 54857 -9906 54880 -9878
rect 54069 -9912 54880 -9906
rect 54090 -9988 54880 -9912
rect 55330 -9918 55380 -9818
rect 55330 -9928 55480 -9918
rect 55220 -9938 55480 -9928
rect 55280 -9952 55480 -9938
rect 55280 -9958 55488 -9952
rect 55280 -9978 55300 -9958
rect 54090 -10088 54150 -9988
rect 54840 -10088 54880 -9988
rect 55288 -9992 55300 -9978
rect 55476 -9992 55488 -9958
rect 55530 -9978 55610 -9968
rect 55288 -9998 55488 -9992
rect 55520 -10002 55530 -9990
rect 55520 -10036 55526 -10002
rect 55288 -10046 55488 -10040
rect 55288 -10080 55300 -10046
rect 55476 -10080 55488 -10046
rect 55520 -10048 55530 -10036
rect 55530 -10078 55610 -10068
rect 55288 -10086 55488 -10080
rect 54090 -10108 54140 -10088
rect 54100 -10348 54140 -10108
rect 54850 -10348 54880 -10088
rect 55300 -10128 55470 -10086
rect 55300 -10268 55320 -10128
rect 55470 -10214 55482 -10142
rect 55300 -10278 55470 -10268
rect 54100 -10388 54880 -10348
rect 27000 -10600 34600 -10400
rect 55710 -10598 55830 -9778
rect 56014 -9808 56020 -9658
rect 56080 -9808 56086 -9658
rect 56014 -9820 56086 -9808
rect 56120 -9808 56170 -9608
rect 56390 -9660 57376 -9608
rect 56390 -9668 57156 -9660
rect 56390 -9808 56654 -9668
rect 56120 -9858 56654 -9808
rect 56306 -9886 56654 -9858
rect 56998 -9820 57156 -9668
rect 57316 -9820 57376 -9660
rect 56998 -9886 57376 -9820
rect 56306 -10300 57376 -9886
rect 57556 -10010 57676 -9230
rect 58896 -9260 58986 -9100
rect 59756 -9120 59826 -9070
rect 59066 -9136 59176 -9130
rect 59066 -9140 59103 -9136
rect 59137 -9140 59176 -9136
rect 59066 -9200 59076 -9140
rect 59166 -9200 59176 -9140
rect 59066 -9210 59176 -9200
rect 58896 -9630 58926 -9260
rect 58966 -9630 58986 -9330
rect 59116 -9260 59506 -9240
rect 59116 -9330 59146 -9260
rect 59226 -9330 59276 -9260
rect 59356 -9330 59396 -9260
rect 59476 -9330 59506 -9260
rect 59116 -9348 59506 -9330
rect 59646 -9260 59716 -9240
rect 59706 -9320 59716 -9260
rect 59646 -9330 59716 -9320
rect 59113 -9354 59513 -9348
rect 59113 -9388 59125 -9354
rect 59501 -9388 59513 -9354
rect 59113 -9394 59513 -9388
rect 59546 -9400 59616 -9390
rect 59246 -9456 59256 -9430
rect 59113 -9462 59256 -9456
rect 59366 -9456 59376 -9430
rect 59366 -9462 59513 -9456
rect 59016 -9500 59076 -9480
rect 59113 -9496 59125 -9462
rect 59501 -9496 59513 -9462
rect 59606 -9460 59616 -9400
rect 59546 -9470 59616 -9460
rect 59113 -9502 59513 -9496
rect 59016 -9590 59076 -9560
rect 59113 -9570 59513 -9564
rect 59113 -9604 59125 -9570
rect 59501 -9604 59513 -9570
rect 59113 -9610 59513 -9604
rect 58896 -9700 58906 -9630
rect 58896 -9720 58986 -9700
rect 59116 -9630 59516 -9610
rect 59116 -9700 59146 -9630
rect 59226 -9700 59276 -9630
rect 59356 -9700 59396 -9630
rect 59476 -9700 59516 -9630
rect 59116 -9720 59516 -9700
rect 59646 -9630 59656 -9330
rect 59706 -9630 59716 -9330
rect 59756 -9300 59766 -9120
rect 59806 -9300 59826 -9120
rect 59956 -9120 60336 -9110
rect 59956 -9134 59966 -9120
rect 59946 -9140 59966 -9134
rect 60326 -9134 60336 -9120
rect 60326 -9140 60346 -9134
rect 59856 -9180 59916 -9170
rect 59946 -9174 59958 -9140
rect 60334 -9174 60346 -9140
rect 61056 -9140 61176 -8790
rect 59946 -9180 59966 -9174
rect 60326 -9180 60346 -9174
rect 60376 -9180 60436 -9160
rect 59956 -9190 60336 -9180
rect 59856 -9260 59916 -9240
rect 59946 -9248 60346 -9242
rect 59756 -9340 59826 -9300
rect 59946 -9282 59958 -9248
rect 60334 -9282 60346 -9248
rect 60376 -9260 60436 -9240
rect 61126 -9240 61176 -9140
rect 61056 -9270 61176 -9240
rect 59946 -9288 60346 -9282
rect 59946 -9340 60336 -9288
rect 59756 -9360 60536 -9340
rect 59756 -9400 59866 -9360
rect 60426 -9400 60536 -9360
rect 59756 -9410 60536 -9400
rect 59796 -9520 59806 -9410
rect 59916 -9520 59926 -9410
rect 59796 -9530 59926 -9520
rect 60436 -9430 60536 -9410
rect 60436 -9550 60446 -9430
rect 60526 -9550 60536 -9430
rect 60436 -9560 60536 -9550
rect 59646 -9640 59716 -9630
rect 59706 -9700 59716 -9640
rect 59646 -9720 59716 -9700
rect 58806 -10010 59356 -9980
rect 57556 -10020 59356 -10010
rect 57556 -10160 58986 -10020
rect 59126 -10160 59356 -10020
rect 59846 -9990 60256 -9980
rect 59846 -10100 59996 -9990
rect 60106 -10100 60256 -9990
rect 57556 -10210 59356 -10160
rect 58806 -10290 59356 -10210
rect 59600 -10300 60500 -10100
rect 55710 -10600 55910 -10598
rect 24730 -11432 25540 -11382
rect 24720 -11632 24730 -11432
rect 25190 -11632 25540 -11432
rect 21706 -11656 21858 -11644
rect 22070 -11644 22076 -11632
rect 22110 -11644 22116 -11632
rect 24730 -11642 25540 -11632
rect 22070 -11656 22116 -11644
rect 21706 -11659 21856 -11656
rect 20896 -11699 21088 -11697
rect 21382 -11699 21646 -11697
rect 21868 -11699 22060 -11697
rect 20886 -11702 22076 -11699
rect 20380 -11703 21070 -11702
rect 21910 -11703 22076 -11702
rect 20380 -11737 20908 -11703
rect 22048 -11737 22076 -11703
rect 20380 -11772 21070 -11737
rect 21910 -11772 22076 -11737
rect 20380 -11779 22076 -11772
rect 20380 -11782 20980 -11779
rect 20380 -11922 20440 -11782
rect 20280 -11924 20440 -11922
rect 20268 -11930 20440 -11924
rect 20268 -11964 20280 -11930
rect 20340 -11962 20440 -11930
rect 20340 -11964 20352 -11962
rect 20268 -11970 20352 -11964
rect 20380 -11974 20440 -11962
rect 20380 -12008 20390 -11974
rect 20424 -12008 20440 -11974
rect 20268 -12018 20352 -12012
rect 20268 -12022 20280 -12018
rect 20250 -12082 20260 -12022
rect 20340 -12058 20352 -12018
rect 20380 -12022 20440 -12008
rect 20340 -12082 20350 -12058
rect 25354 -12116 25416 -12110
rect 16428 -12122 25422 -12116
rect 16428 -12182 16440 -12122
rect 16428 -12188 25360 -12182
rect 16480 -12232 25030 -12222
rect 16410 -12245 25030 -12232
rect 16410 -12279 16615 -12245
rect 16703 -12279 17021 -12245
rect 17109 -12279 17427 -12245
rect 17515 -12279 17833 -12245
rect 17921 -12279 18239 -12245
rect 18327 -12279 18645 -12245
rect 18733 -12279 19051 -12245
rect 19139 -12279 19457 -12245
rect 19545 -12279 19863 -12245
rect 19951 -12279 20269 -12245
rect 20357 -12279 20675 -12245
rect 20763 -12279 21081 -12245
rect 21169 -12279 21487 -12245
rect 21575 -12279 21893 -12245
rect 21981 -12279 22299 -12245
rect 22387 -12279 22705 -12245
rect 22793 -12279 23111 -12245
rect 23199 -12279 23517 -12245
rect 23605 -12279 23923 -12245
rect 24011 -12279 24329 -12245
rect 24417 -12279 24735 -12245
rect 24823 -12279 25030 -12245
rect 16410 -12282 25030 -12279
rect 16410 -13152 16480 -12282
rect 16603 -12285 16715 -12282
rect 17009 -12285 17121 -12282
rect 17415 -12285 17527 -12282
rect 17821 -12285 17933 -12282
rect 18227 -12285 18339 -12282
rect 18633 -12285 18745 -12282
rect 19039 -12285 19151 -12282
rect 19445 -12285 19557 -12282
rect 19851 -12285 19963 -12282
rect 20257 -12285 20369 -12282
rect 20663 -12285 20775 -12282
rect 20810 -12312 20880 -12282
rect 21069 -12285 21181 -12282
rect 21475 -12285 21587 -12282
rect 21881 -12285 21993 -12282
rect 22287 -12285 22399 -12282
rect 22693 -12285 22805 -12282
rect 23099 -12285 23211 -12282
rect 23505 -12285 23617 -12282
rect 23911 -12285 24023 -12282
rect 24317 -12285 24429 -12282
rect 24723 -12285 24835 -12282
rect 20790 -12317 20880 -12312
rect 16547 -12329 16593 -12317
rect 16725 -12329 16771 -12317
rect 16953 -12329 16999 -12317
rect 17131 -12329 17177 -12317
rect 17359 -12329 17405 -12317
rect 17537 -12329 17583 -12317
rect 17765 -12329 17811 -12317
rect 17943 -12329 17989 -12317
rect 18171 -12329 18217 -12317
rect 18349 -12329 18395 -12317
rect 18577 -12329 18623 -12317
rect 18755 -12329 18801 -12317
rect 18983 -12329 19029 -12317
rect 19161 -12329 19207 -12317
rect 19389 -12329 19435 -12317
rect 19567 -12329 19613 -12317
rect 19795 -12329 19841 -12317
rect 19973 -12329 20019 -12317
rect 20201 -12329 20247 -12317
rect 20379 -12329 20425 -12317
rect 20607 -12329 20653 -12317
rect 20785 -12329 20880 -12317
rect 21013 -12329 21059 -12317
rect 21191 -12329 21237 -12317
rect 21419 -12329 21465 -12317
rect 21597 -12329 21643 -12317
rect 21825 -12329 21871 -12317
rect 22003 -12329 22049 -12317
rect 22231 -12329 22277 -12317
rect 22409 -12329 22455 -12317
rect 22637 -12329 22683 -12317
rect 22815 -12329 22861 -12317
rect 23043 -12329 23089 -12317
rect 23221 -12329 23267 -12317
rect 23449 -12329 23495 -12317
rect 23627 -12329 23673 -12317
rect 23855 -12329 23901 -12317
rect 24033 -12329 24079 -12317
rect 24261 -12329 24307 -12317
rect 24439 -12329 24485 -12317
rect 24667 -12329 24713 -12317
rect 24845 -12329 24891 -12317
rect 16517 -13106 16527 -12329
rect 16587 -13105 16596 -12329
rect 16725 -12330 16731 -12329
rect 16765 -12330 16771 -12329
rect 16586 -13106 16596 -13105
rect 16547 -13117 16593 -13106
rect 16720 -13107 16730 -12330
rect 16789 -13107 16799 -12330
rect 16923 -13106 16933 -12329
rect 16993 -13105 17002 -12329
rect 17131 -12330 17137 -12329
rect 17171 -12330 17177 -12329
rect 16992 -13106 17002 -13105
rect 16725 -13117 16771 -13107
rect 16953 -13117 16999 -13106
rect 17126 -13107 17136 -12330
rect 17195 -13107 17205 -12330
rect 17329 -13106 17339 -12329
rect 17399 -13105 17408 -12329
rect 17537 -12330 17543 -12329
rect 17577 -12330 17583 -12329
rect 17398 -13106 17408 -13105
rect 17131 -13117 17177 -13107
rect 17359 -13117 17405 -13106
rect 17532 -13107 17542 -12330
rect 17601 -13107 17611 -12330
rect 17735 -13106 17745 -12329
rect 17805 -13105 17814 -12329
rect 17943 -12330 17949 -12329
rect 17983 -12330 17989 -12329
rect 17804 -13106 17814 -13105
rect 17537 -13117 17583 -13107
rect 17765 -13117 17811 -13106
rect 17938 -13107 17948 -12330
rect 18007 -13107 18017 -12330
rect 18141 -13106 18151 -12329
rect 18211 -13105 18220 -12329
rect 18349 -12330 18355 -12329
rect 18389 -12330 18395 -12329
rect 18210 -13106 18220 -13105
rect 17943 -13117 17989 -13107
rect 18171 -13117 18217 -13106
rect 18344 -13107 18354 -12330
rect 18413 -13107 18423 -12330
rect 18547 -13106 18557 -12329
rect 18617 -13105 18626 -12329
rect 18755 -12330 18761 -12329
rect 18795 -12330 18801 -12329
rect 18616 -13106 18626 -13105
rect 18349 -13117 18395 -13107
rect 18577 -13117 18623 -13106
rect 18750 -13107 18760 -12330
rect 18819 -13107 18829 -12330
rect 18953 -13106 18963 -12329
rect 19023 -13105 19032 -12329
rect 19161 -12330 19167 -12329
rect 19201 -12330 19207 -12329
rect 19022 -13106 19032 -13105
rect 18755 -13117 18801 -13107
rect 18983 -13117 19029 -13106
rect 19156 -13107 19166 -12330
rect 19225 -13107 19235 -12330
rect 19359 -13106 19369 -12329
rect 19429 -13105 19438 -12329
rect 19567 -12330 19573 -12329
rect 19607 -12330 19613 -12329
rect 19428 -13106 19438 -13105
rect 19161 -13117 19207 -13107
rect 19389 -13117 19435 -13106
rect 19562 -13107 19572 -12330
rect 19631 -13107 19641 -12330
rect 19765 -13106 19775 -12329
rect 19835 -13105 19844 -12329
rect 19973 -12330 19979 -12329
rect 20013 -12330 20019 -12329
rect 19834 -13106 19844 -13105
rect 19567 -13117 19613 -13107
rect 19795 -13117 19841 -13106
rect 19968 -13107 19978 -12330
rect 20037 -13107 20047 -12330
rect 20171 -13106 20181 -12329
rect 20241 -13105 20250 -12329
rect 20379 -12330 20385 -12329
rect 20419 -12330 20425 -12329
rect 20240 -13106 20250 -13105
rect 19973 -13117 20019 -13107
rect 20201 -13117 20247 -13106
rect 20374 -13107 20384 -12330
rect 20443 -13107 20453 -12330
rect 20577 -12352 20613 -12329
rect 20570 -13042 20580 -12352
rect 20577 -13105 20613 -13042
rect 20647 -13105 20656 -12329
rect 20785 -12330 20791 -12329
rect 20577 -13106 20656 -13105
rect 20780 -13105 20791 -12330
rect 20825 -12351 20880 -12329
rect 20861 -13041 20880 -12351
rect 20825 -13105 20880 -13041
rect 20379 -13117 20425 -13107
rect 20607 -13117 20653 -13106
rect 20780 -13107 20880 -13105
rect 20983 -13106 20993 -12329
rect 21053 -13105 21062 -12329
rect 21191 -12330 21197 -12329
rect 21231 -12330 21237 -12329
rect 21052 -13106 21062 -13105
rect 20785 -13117 20880 -13107
rect 21013 -13117 21059 -13106
rect 21186 -13107 21196 -12330
rect 21255 -13107 21265 -12330
rect 21389 -13106 21399 -12329
rect 21459 -13105 21468 -12329
rect 21597 -12330 21603 -12329
rect 21637 -12330 21643 -12329
rect 21458 -13106 21468 -13105
rect 21191 -13117 21237 -13107
rect 21419 -13117 21465 -13106
rect 21592 -13107 21602 -12330
rect 21661 -13107 21671 -12330
rect 21795 -13106 21805 -12329
rect 21865 -13105 21874 -12329
rect 22003 -12330 22009 -12329
rect 22043 -12330 22049 -12329
rect 21864 -13106 21874 -13105
rect 21597 -13117 21643 -13107
rect 21825 -13117 21871 -13106
rect 21998 -13107 22008 -12330
rect 22067 -13107 22077 -12330
rect 22201 -13106 22211 -12329
rect 22271 -13105 22280 -12329
rect 22409 -12330 22415 -12329
rect 22449 -12330 22455 -12329
rect 22270 -13106 22280 -13105
rect 22003 -13117 22049 -13107
rect 22231 -13117 22277 -13106
rect 22404 -13107 22414 -12330
rect 22473 -13107 22483 -12330
rect 22607 -13106 22617 -12329
rect 22677 -13105 22686 -12329
rect 22815 -12330 22821 -12329
rect 22855 -12330 22861 -12329
rect 22676 -13106 22686 -13105
rect 22409 -13117 22455 -13107
rect 22637 -13117 22683 -13106
rect 22810 -13107 22820 -12330
rect 22879 -13107 22889 -12330
rect 23013 -13106 23023 -12329
rect 23083 -13105 23092 -12329
rect 23221 -12330 23227 -12329
rect 23261 -12330 23267 -12329
rect 23082 -13106 23092 -13105
rect 22815 -13117 22861 -13107
rect 23043 -13117 23089 -13106
rect 23216 -13107 23226 -12330
rect 23285 -13107 23295 -12330
rect 23419 -13106 23429 -12329
rect 23489 -13105 23498 -12329
rect 23627 -12330 23633 -12329
rect 23667 -12330 23673 -12329
rect 23488 -13106 23498 -13105
rect 23221 -13117 23267 -13107
rect 23449 -13117 23495 -13106
rect 23622 -13107 23632 -12330
rect 23691 -13107 23701 -12330
rect 23825 -13106 23835 -12329
rect 23895 -13105 23904 -12329
rect 24033 -12330 24039 -12329
rect 24073 -12330 24079 -12329
rect 23894 -13106 23904 -13105
rect 23627 -13117 23673 -13107
rect 23855 -13117 23901 -13106
rect 24028 -13107 24038 -12330
rect 24097 -13107 24107 -12330
rect 24231 -13106 24241 -12329
rect 24301 -13105 24310 -12329
rect 24439 -12330 24445 -12329
rect 24479 -12330 24485 -12329
rect 24300 -13106 24310 -13105
rect 24033 -13117 24079 -13107
rect 24261 -13117 24307 -13106
rect 24434 -13107 24444 -12330
rect 24503 -13107 24513 -12330
rect 24637 -13106 24647 -12329
rect 24707 -13105 24716 -12329
rect 24845 -12330 24851 -12329
rect 24885 -12330 24891 -12329
rect 24706 -13106 24716 -13105
rect 24439 -13117 24485 -13107
rect 24667 -13117 24713 -13106
rect 24840 -13107 24850 -12330
rect 24909 -13107 24919 -12330
rect 24845 -13117 24891 -13107
rect 20790 -13122 20880 -13117
rect 16603 -13152 16715 -13149
rect 17009 -13152 17121 -13149
rect 17415 -13152 17527 -13149
rect 17821 -13152 17933 -13149
rect 18227 -13152 18339 -13149
rect 18633 -13152 18745 -13149
rect 19039 -13152 19151 -13149
rect 19445 -13152 19557 -13149
rect 19851 -13152 19963 -13149
rect 20257 -13152 20369 -13149
rect 20663 -13152 20775 -13149
rect 20810 -13152 20880 -13122
rect 21069 -13152 21181 -13149
rect 21475 -13152 21587 -13149
rect 21881 -13152 21993 -13149
rect 22287 -13152 22399 -13149
rect 22693 -13152 22805 -13149
rect 23099 -13152 23211 -13149
rect 23505 -13152 23617 -13149
rect 23911 -13152 24023 -13149
rect 24317 -13152 24429 -13149
rect 24723 -13152 24835 -13149
rect 16410 -13153 24840 -13152
rect 24960 -13153 25030 -12282
rect 25080 -12292 25090 -12222
rect 25210 -12245 25250 -12222
rect 25229 -12276 25250 -12245
rect 25354 -12276 25360 -12188
rect 25410 -12188 25422 -12122
rect 25410 -12262 25416 -12188
rect 27000 -12262 27200 -10600
rect 25229 -12279 25246 -12276
rect 25210 -12282 25246 -12279
rect 25210 -12285 25241 -12282
rect 25210 -12292 25220 -12285
rect 25080 -12317 25140 -12292
rect 25073 -12329 25140 -12317
rect 25073 -13105 25079 -12329
rect 25113 -13105 25140 -12329
rect 25073 -13117 25140 -13105
rect 25251 -12329 25297 -12317
rect 25251 -13105 25257 -12329
rect 25291 -12368 25297 -12329
rect 25354 -12336 25362 -12276
rect 25353 -12368 25362 -12336
rect 25291 -13036 25362 -12368
rect 25291 -13105 25297 -13036
rect 25251 -13117 25297 -13105
rect 16410 -13155 25030 -13153
rect 16410 -13189 16615 -13155
rect 16703 -13189 17021 -13155
rect 17109 -13189 17427 -13155
rect 17515 -13189 17833 -13155
rect 17921 -13189 18239 -13155
rect 18327 -13189 18645 -13155
rect 18733 -13189 19051 -13155
rect 19139 -13189 19457 -13155
rect 19545 -13189 19863 -13155
rect 19951 -13189 20269 -13155
rect 20357 -13189 20675 -13155
rect 20763 -13189 21081 -13155
rect 21169 -13189 21487 -13155
rect 21575 -13189 21893 -13155
rect 21981 -13189 22299 -13155
rect 22387 -13189 22705 -13155
rect 22793 -13189 23111 -13155
rect 23199 -13189 23517 -13155
rect 23605 -13189 23923 -13155
rect 24011 -13189 24329 -13155
rect 24417 -13189 24735 -13155
rect 24823 -13189 25030 -13155
rect 25080 -13149 25140 -13117
rect 25353 -13149 25362 -13036
rect 25410 -13000 27200 -12262
rect 34400 -12262 34600 -10600
rect 55400 -10700 56100 -10600
rect 55400 -11100 55500 -10700
rect 56000 -11100 56100 -10700
rect 59600 -10700 59700 -10300
rect 60400 -10700 60500 -10300
rect 59600 -10800 60500 -10700
rect 55400 -11200 56100 -11100
rect 55320 -11660 55800 -11600
rect 55320 -11980 55380 -11660
rect 55740 -11980 55800 -11660
rect 55320 -12040 55800 -11980
rect 54090 -12138 54890 -12098
rect 34400 -13000 34730 -12262
rect 54090 -12268 54150 -12138
rect 53510 -12320 53800 -12318
rect 53460 -12340 53800 -12320
rect 53460 -12540 53480 -12340
rect 53780 -12540 53800 -12340
rect 54080 -12398 54150 -12268
rect 54860 -12378 54890 -12138
rect 54850 -12398 54890 -12378
rect 54080 -12466 54880 -12398
rect 54079 -12472 54880 -12466
rect 54079 -12506 54091 -12472
rect 54867 -12498 54880 -12472
rect 54867 -12506 54879 -12498
rect 54079 -12512 54879 -12506
rect 53460 -12560 53800 -12540
rect 53510 -12658 53800 -12560
rect 53002 -12820 53480 -12758
rect 25080 -13155 25241 -13149
rect 25080 -13182 25141 -13155
rect 16410 -13212 25030 -13189
rect 25129 -13189 25141 -13182
rect 25229 -13189 25241 -13155
rect 25129 -13195 25241 -13189
rect 25353 -13219 25361 -13149
rect 25353 -13248 25360 -13219
rect 16436 -13254 25360 -13248
rect 16436 -13314 16448 -13254
rect 25410 -13302 34730 -13000
rect 25400 -13314 34730 -13302
rect 16436 -13320 20570 -13314
rect 16440 -13350 20570 -13320
rect 16414 -13362 20570 -13350
rect 20670 -13362 34730 -13314
rect 16414 -16086 16420 -13362
rect 16490 -13428 34630 -13422
rect 16490 -14736 16496 -13428
rect 16578 -13532 16987 -13520
rect 34160 -13532 34630 -13428
rect 16570 -14642 16580 -13532
rect 16990 -14642 17000 -13532
rect 16578 -14646 16584 -14642
rect 16981 -14646 16987 -14642
rect 16578 -14658 16987 -14646
rect 34160 -14646 34171 -13532
rect 34568 -14646 34630 -13532
rect 34160 -14736 34630 -14646
rect 16490 -14742 34630 -14736
rect 34720 -13428 34730 -13362
rect 53000 -12958 53480 -12820
rect 53510 -12768 53520 -12658
rect 53640 -12768 53800 -12658
rect 53510 -12888 53800 -12768
rect 53970 -12534 54040 -12518
rect 53970 -12572 53998 -12534
rect 54032 -12572 54040 -12534
rect 53970 -12768 54040 -12572
rect 54920 -12534 54990 -12518
rect 54920 -12572 54926 -12534
rect 54960 -12572 54990 -12534
rect 54079 -12600 54879 -12594
rect 54079 -12634 54091 -12600
rect 54867 -12634 54879 -12600
rect 54079 -12638 54879 -12634
rect 54079 -12640 54750 -12638
rect 54090 -12688 54750 -12640
rect 54740 -12718 54750 -12688
rect 54850 -12640 54879 -12638
rect 54850 -12708 54860 -12640
rect 54840 -12718 54860 -12708
rect 54750 -12728 54860 -12718
rect 54920 -12768 54990 -12572
rect 55430 -12618 55520 -12608
rect 55290 -12728 55390 -12718
rect 53970 -12798 55290 -12768
rect 55430 -12758 55520 -12688
rect 53970 -12808 55390 -12798
rect 54050 -12818 55380 -12808
rect 54050 -12828 54880 -12818
rect 54050 -12838 54091 -12828
rect 54079 -12862 54091 -12838
rect 54867 -12838 54880 -12828
rect 54867 -12862 54879 -12838
rect 54079 -12868 54879 -12862
rect 54920 -12878 54990 -12868
rect 53510 -12906 53630 -12888
rect 53510 -12938 53526 -12906
rect 53514 -12940 53526 -12938
rect 53614 -12938 53630 -12906
rect 53940 -12890 54038 -12878
rect 53940 -12898 53998 -12890
rect 53614 -12940 53626 -12938
rect 53514 -12946 53626 -12940
rect 34720 -14736 34726 -13428
rect 53000 -14708 53050 -12958
rect 53250 -12968 53480 -12958
rect 53250 -14318 53330 -12968
rect 53400 -12978 53480 -12968
rect 53400 -12990 53504 -12978
rect 53400 -13766 53464 -12990
rect 53498 -13766 53504 -12990
rect 53400 -13778 53504 -13766
rect 53636 -12988 53682 -12978
rect 53636 -12990 53760 -12988
rect 53636 -13766 53642 -12990
rect 53676 -13766 53760 -12990
rect 53940 -12998 53950 -12898
rect 54032 -12928 54038 -12890
rect 54020 -12940 54038 -12928
rect 54020 -12998 54030 -12940
rect 54079 -12956 54879 -12950
rect 54079 -12990 54091 -12956
rect 54867 -12990 54879 -12956
rect 54920 -12978 54990 -12968
rect 55320 -12968 55380 -12818
rect 54079 -12996 54879 -12990
rect 53940 -13018 54030 -12998
rect 54090 -13028 54870 -12996
rect 55320 -13002 55334 -12968
rect 55368 -13002 55380 -12968
rect 55320 -13008 55380 -13002
rect 53840 -13328 53920 -13318
rect 53840 -13438 53860 -13328
rect 53840 -13448 53920 -13438
rect 53840 -13640 53900 -13448
rect 54320 -13528 54510 -13028
rect 55440 -13038 55520 -12758
rect 55410 -13040 55520 -13038
rect 55284 -13048 55330 -13040
rect 55230 -13052 55330 -13048
rect 55230 -13058 55290 -13052
rect 55324 -13228 55330 -13052
rect 55230 -13238 55330 -13228
rect 55284 -13240 55330 -13238
rect 55372 -13048 55520 -13040
rect 55372 -13052 55430 -13048
rect 55372 -13228 55378 -13052
rect 55412 -13218 55430 -13052
rect 55510 -13218 55520 -13048
rect 55412 -13228 55520 -13218
rect 55372 -13240 55418 -13228
rect 55580 -13328 55720 -12040
rect 58776 -12270 59306 -12150
rect 58776 -12280 58966 -12270
rect 56146 -12380 57366 -12330
rect 55954 -12528 56046 -12516
rect 56146 -12528 56506 -12380
rect 55954 -12698 55960 -12528
rect 56040 -12698 56046 -12528
rect 55954 -12710 56046 -12698
rect 56120 -12558 56506 -12528
rect 56120 -12768 56190 -12558
rect 56390 -12630 56506 -12558
rect 57016 -12534 57366 -12380
rect 57586 -12430 58966 -12280
rect 59126 -12430 59306 -12270
rect 57586 -12450 59306 -12430
rect 59946 -12300 60386 -12200
rect 57586 -12480 58986 -12450
rect 59946 -12460 59956 -12300
rect 60166 -12460 60386 -12300
rect 57016 -12630 57368 -12534
rect 56390 -12670 57368 -12630
rect 56390 -12768 57126 -12670
rect 56120 -12774 57126 -12768
rect 56120 -12778 56750 -12774
rect 55880 -12818 55970 -12808
rect 55870 -12896 55880 -12850
rect 55970 -12896 55982 -12850
rect 55880 -12908 55970 -12898
rect 55000 -13338 55090 -13328
rect 55000 -13448 55090 -13438
rect 54710 -13528 54960 -13508
rect 53940 -13568 54960 -13528
rect 53940 -13572 54730 -13568
rect 53930 -13578 54730 -13572
rect 53930 -13612 53942 -13578
rect 54718 -13612 54730 -13578
rect 53930 -13618 54730 -13612
rect 53840 -13728 53858 -13640
rect 53892 -13728 53900 -13640
rect 53840 -13748 53900 -13728
rect 54762 -13638 54850 -13628
rect 54762 -13640 54770 -13638
rect 54762 -13728 54768 -13640
rect 54840 -13728 54850 -13638
rect 54762 -13740 54850 -13728
rect 54770 -13748 54850 -13740
rect 53636 -13778 53760 -13766
rect 53400 -13996 53480 -13778
rect 53514 -13816 53626 -13810
rect 53514 -13818 53526 -13816
rect 53510 -13850 53526 -13818
rect 53614 -13818 53626 -13816
rect 53614 -13850 53630 -13818
rect 53510 -13924 53630 -13850
rect 53510 -13958 53526 -13924
rect 53614 -13958 53630 -13924
rect 53680 -13838 53760 -13778
rect 53930 -13756 54730 -13750
rect 53930 -13790 53942 -13756
rect 54718 -13790 54730 -13756
rect 53930 -13796 54730 -13790
rect 53940 -13828 54720 -13796
rect 53920 -13838 54720 -13828
rect 53680 -13928 54720 -13838
rect 53514 -13964 53626 -13958
rect 53680 -13996 53760 -13928
rect 53920 -13938 54720 -13928
rect 53940 -13978 54720 -13938
rect 54900 -13968 54960 -13568
rect 55010 -13560 55090 -13448
rect 55540 -13338 55720 -13328
rect 55630 -13438 55720 -13338
rect 55130 -13474 55506 -13468
rect 55130 -13508 55142 -13474
rect 55494 -13508 55506 -13474
rect 55130 -13514 55506 -13508
rect 55010 -13594 55046 -13560
rect 55080 -13594 55090 -13560
rect 55010 -13608 55090 -13594
rect 55142 -13640 55494 -13514
rect 55540 -13560 55720 -13438
rect 55540 -13594 55556 -13560
rect 55590 -13594 55720 -13560
rect 55540 -13608 55720 -13594
rect 55780 -12940 55860 -12928
rect 55130 -13646 55506 -13640
rect 55130 -13680 55142 -13646
rect 55494 -13678 55506 -13646
rect 55494 -13680 55510 -13678
rect 55130 -13686 55510 -13680
rect 55140 -13698 55510 -13686
rect 55780 -13698 55820 -12940
rect 55140 -13716 55820 -13698
rect 55854 -13716 55860 -12940
rect 55140 -13728 55860 -13716
rect 55992 -12940 56038 -12928
rect 55992 -13716 55998 -12940
rect 56032 -12948 56038 -12940
rect 56120 -12948 56300 -12778
rect 57098 -12800 57126 -12774
rect 57356 -12800 57368 -12670
rect 57098 -12814 57368 -12800
rect 57096 -12845 57372 -12814
rect 57096 -12879 57125 -12845
rect 57159 -12879 57217 -12845
rect 57251 -12879 57309 -12845
rect 57343 -12879 57372 -12845
rect 57096 -12910 57372 -12879
rect 56032 -13306 56300 -12948
rect 56590 -13068 56660 -13058
rect 56660 -13134 57000 -13068
rect 57586 -13130 57706 -12480
rect 59946 -12490 60386 -12460
rect 57366 -13134 57706 -13130
rect 56660 -13138 57188 -13134
rect 56660 -13144 57190 -13138
rect 56660 -13194 57118 -13144
rect 57178 -13194 57190 -13144
rect 57314 -13140 57706 -13134
rect 57314 -13180 57326 -13140
rect 57366 -13180 57706 -13140
rect 57314 -13186 57706 -13180
rect 57366 -13190 57706 -13186
rect 58896 -12770 58986 -12750
rect 58896 -12830 58906 -12770
rect 58896 -13120 58926 -12830
rect 58966 -13120 58986 -12770
rect 59106 -12770 59516 -12760
rect 59106 -12830 59216 -12770
rect 59276 -12830 59326 -12770
rect 59386 -12830 59436 -12770
rect 59496 -12830 59516 -12770
rect 59106 -12847 59516 -12830
rect 59626 -12770 59706 -12730
rect 59626 -12830 59636 -12770
rect 59626 -12840 59656 -12830
rect 59106 -12880 59125 -12847
rect 59113 -12881 59125 -12880
rect 59501 -12880 59516 -12847
rect 59501 -12881 59513 -12880
rect 59113 -12887 59513 -12881
rect 59546 -12890 59616 -12880
rect 59276 -12930 59356 -12920
rect 59276 -12949 59286 -12930
rect 59113 -12955 59286 -12949
rect 59346 -12949 59356 -12930
rect 59346 -12955 59513 -12949
rect 59113 -12989 59125 -12955
rect 59501 -12989 59513 -12955
rect 59606 -12950 59616 -12890
rect 59546 -12960 59616 -12950
rect 59113 -12990 59286 -12989
rect 59346 -12990 59513 -12989
rect 59016 -13000 59076 -12990
rect 59113 -12995 59513 -12990
rect 59276 -13000 59356 -12995
rect 59546 -13010 59616 -13000
rect 59016 -13070 59076 -13060
rect 59113 -13063 59513 -13057
rect 59113 -13097 59125 -13063
rect 59501 -13097 59513 -13063
rect 59606 -13070 59616 -13010
rect 59546 -13080 59616 -13070
rect 59113 -13100 59513 -13097
rect 59113 -13103 59516 -13100
rect 58896 -13130 58986 -13120
rect 58896 -13190 58906 -13130
rect 58966 -13190 58986 -13130
rect 58896 -13192 58986 -13190
rect 59116 -13120 59516 -13103
rect 59646 -13110 59656 -12840
rect 59116 -13180 59216 -13120
rect 59276 -13180 59336 -13120
rect 59396 -13180 59436 -13120
rect 59496 -13180 59516 -13120
rect 56660 -13198 57190 -13194
rect 56590 -13200 57190 -13198
rect 56590 -13204 57188 -13200
rect 56590 -13268 57000 -13204
rect 56032 -13318 56356 -13306
rect 56032 -13716 56280 -13318
rect 55992 -13728 56280 -13716
rect 55140 -13738 55200 -13728
rect 55450 -13758 55810 -13728
rect 55870 -13766 55982 -13760
rect 55870 -13800 55882 -13766
rect 55970 -13800 55982 -13766
rect 55870 -13806 55982 -13800
rect 55140 -13818 55200 -13808
rect 55024 -13848 55116 -13836
rect 55024 -13928 55030 -13848
rect 55110 -13928 55116 -13848
rect 55024 -13940 55116 -13928
rect 55734 -13848 55816 -13836
rect 55734 -13928 55740 -13848
rect 55810 -13928 55816 -13848
rect 55734 -13940 55816 -13928
rect 55880 -13838 55970 -13806
rect 55880 -13964 55970 -13928
rect 56060 -13948 56280 -13728
rect 56350 -13948 56356 -13318
rect 56480 -13388 56550 -13378
rect 56480 -13458 56550 -13448
rect 56590 -13487 56750 -13268
rect 58894 -13286 58988 -13192
rect 59116 -13200 59516 -13180
rect 59636 -13120 59656 -13110
rect 59696 -13120 59706 -12770
rect 59856 -12940 59976 -12930
rect 59856 -13030 59866 -12940
rect 59966 -13030 59976 -12940
rect 59856 -13040 59976 -13030
rect 60436 -13020 60446 -12920
rect 60526 -13020 60536 -12920
rect 60436 -13040 60536 -13020
rect 59636 -13130 59706 -13120
rect 59696 -13190 59706 -13130
rect 59636 -13210 59706 -13190
rect 59756 -13060 60536 -13040
rect 59756 -13100 59866 -13060
rect 60426 -13100 60536 -13060
rect 59756 -13110 60536 -13100
rect 59756 -13150 59826 -13110
rect 59066 -13240 59176 -13230
rect 58896 -13350 58986 -13286
rect 59066 -13310 59076 -13240
rect 59166 -13310 59176 -13240
rect 59066 -13312 59103 -13310
rect 59137 -13312 59176 -13310
rect 59066 -13320 59176 -13312
rect 59756 -13340 59766 -13150
rect 59806 -13340 59826 -13150
rect 59956 -13168 60046 -13140
rect 59946 -13174 60046 -13168
rect 60126 -13168 60336 -13140
rect 60126 -13174 60346 -13168
rect 59856 -13210 59916 -13200
rect 59946 -13208 59958 -13174
rect 60334 -13208 60346 -13174
rect 59946 -13214 60346 -13208
rect 60376 -13220 60446 -13210
rect 59856 -13290 59916 -13280
rect 59946 -13282 60346 -13276
rect 59946 -13316 59958 -13282
rect 60334 -13316 60346 -13282
rect 60376 -13290 60446 -13280
rect 59946 -13322 59976 -13316
rect 57098 -13358 57368 -13354
rect 57096 -13364 57372 -13358
rect 57096 -13450 57098 -13364
rect 56424 -13488 56470 -13487
rect 56060 -13960 56356 -13948
rect 56410 -13499 56470 -13488
rect 53400 -14008 53504 -13996
rect 53400 -14318 53464 -14008
rect 53250 -14708 53464 -14318
rect 34720 -14742 34736 -14736
rect 34724 -14802 34736 -14742
rect 53000 -14784 53464 -14708
rect 53498 -14784 53504 -14008
rect 53000 -14788 53504 -14784
rect 53458 -14796 53504 -14788
rect 53636 -14008 53760 -13996
rect 53636 -14784 53642 -14008
rect 53676 -14784 53760 -14008
rect 53930 -13984 54730 -13978
rect 53930 -14018 53942 -13984
rect 54718 -14018 54730 -13984
rect 53930 -14024 54730 -14018
rect 53830 -14046 53900 -14028
rect 53830 -14134 53858 -14046
rect 53892 -14134 53900 -14046
rect 53830 -14328 53900 -14134
rect 54760 -14046 54850 -14028
rect 54760 -14134 54768 -14046
rect 54802 -14048 54850 -14046
rect 54900 -14038 55200 -13968
rect 55870 -13970 55982 -13964
rect 55870 -14004 55882 -13970
rect 55970 -14004 55982 -13970
rect 55450 -14038 55810 -14008
rect 55870 -14010 55982 -14004
rect 56060 -14038 56300 -13960
rect 54900 -14042 55820 -14038
rect 56000 -14042 56300 -14038
rect 54900 -14048 55860 -14042
rect 54840 -14128 54850 -14048
rect 54802 -14134 54850 -14128
rect 54760 -14148 54850 -14134
rect 55130 -14054 55860 -14048
rect 55130 -14078 55820 -14054
rect 55130 -14096 55510 -14078
rect 55130 -14130 55142 -14096
rect 55494 -14098 55510 -14096
rect 55494 -14130 55506 -14098
rect 55130 -14136 55506 -14130
rect 53930 -14162 54730 -14156
rect 53930 -14196 53942 -14162
rect 54718 -14196 54730 -14162
rect 55020 -14182 55090 -14168
rect 53930 -14202 54730 -14196
rect 53940 -14208 54730 -14202
rect 54920 -14198 54980 -14188
rect 53940 -14248 54920 -14208
rect 53830 -14338 53920 -14328
rect 53830 -14448 53850 -14338
rect 53830 -14458 53920 -14448
rect 54320 -14748 54510 -14248
rect 54710 -14268 54920 -14248
rect 54910 -14278 54980 -14268
rect 55020 -14216 55046 -14182
rect 55080 -14216 55090 -14182
rect 55020 -14328 55090 -14216
rect 55142 -14262 55494 -14136
rect 55540 -14182 55620 -14168
rect 55540 -14216 55556 -14182
rect 55590 -14216 55620 -14182
rect 55130 -14268 55506 -14262
rect 55130 -14302 55142 -14268
rect 55494 -14302 55506 -14268
rect 55130 -14308 55506 -14302
rect 55000 -14338 55090 -14328
rect 55000 -14448 55090 -14438
rect 55540 -14328 55620 -14216
rect 55540 -14338 55630 -14328
rect 55630 -14438 55680 -14348
rect 55540 -14448 55680 -14438
rect 55274 -14538 55320 -14536
rect 55220 -14548 55320 -14538
rect 55220 -14724 55280 -14718
rect 55314 -14724 55320 -14548
rect 55220 -14728 55320 -14724
rect 55274 -14736 55320 -14728
rect 55362 -14548 55408 -14536
rect 55362 -14724 55368 -14548
rect 55402 -14558 55510 -14548
rect 55402 -14724 55410 -14558
rect 55362 -14728 55410 -14724
rect 55500 -14728 55510 -14558
rect 55362 -14736 55510 -14728
rect 55390 -14738 55510 -14736
rect 53636 -14788 53760 -14784
rect 53636 -14796 53682 -14788
rect 16408 -16182 16420 -16086
rect 16490 -14808 34630 -14802
rect 16490 -16086 16496 -14808
rect 16578 -14904 16987 -14892
rect 16578 -14912 16584 -14904
rect 16981 -14912 16987 -14904
rect 34160 -14904 34630 -14808
rect 16570 -16022 16580 -14912
rect 16990 -16022 17000 -14912
rect 34160 -16018 34171 -14904
rect 34568 -16018 34630 -14904
rect 16578 -16030 16987 -16022
rect 34160 -16086 34630 -16018
rect 16490 -16092 34630 -16086
rect 34720 -14808 34736 -14802
rect 53940 -14808 54020 -14768
rect 54080 -14782 54860 -14748
rect 55311 -14774 55371 -14768
rect 34720 -16086 34726 -14808
rect 53514 -14834 53626 -14828
rect 53514 -14838 53526 -14834
rect 53510 -14868 53526 -14838
rect 53614 -14838 53626 -14834
rect 53614 -14868 53630 -14838
rect 53510 -14928 53630 -14868
rect 53940 -14888 53950 -14808
rect 54010 -14838 54020 -14808
rect 54069 -14788 54869 -14782
rect 54069 -14822 54081 -14788
rect 54857 -14822 54869 -14788
rect 54069 -14828 54869 -14822
rect 54910 -14798 54980 -14788
rect 54010 -14850 54028 -14838
rect 54022 -14888 54028 -14850
rect 53940 -14900 54028 -14888
rect 53940 -14908 54020 -14900
rect 54910 -14908 54980 -14898
rect 55311 -14808 55324 -14774
rect 55358 -14808 55371 -14774
rect 54070 -14910 54870 -14908
rect 54069 -14916 54870 -14910
rect 54069 -14938 54081 -14916
rect 54041 -14950 54081 -14938
rect 54857 -14918 54870 -14916
rect 54857 -14950 54880 -14918
rect 55311 -14948 55371 -14808
rect 54041 -14958 54880 -14950
rect 55240 -14958 55371 -14948
rect 54041 -14968 55240 -14958
rect 53510 -15058 53630 -15048
rect 53961 -15008 55240 -14968
rect 53961 -15206 54031 -15008
rect 54730 -15068 54860 -15058
rect 54730 -15088 54740 -15068
rect 54080 -15138 54740 -15088
rect 54069 -15144 54740 -15138
rect 54850 -15138 54860 -15068
rect 54850 -15144 54869 -15138
rect 54069 -15178 54081 -15144
rect 54857 -15178 54869 -15144
rect 54069 -15184 54869 -15178
rect 54911 -15194 54981 -15008
rect 55370 -15008 55371 -14958
rect 55240 -15028 55370 -15018
rect 55410 -15048 55510 -14738
rect 55410 -15158 55510 -15138
rect 55570 -15068 55680 -14448
rect 55780 -14830 55820 -14078
rect 55854 -14830 55860 -14054
rect 55780 -14838 55860 -14830
rect 55814 -14842 55860 -14838
rect 55992 -14054 56300 -14042
rect 55992 -14830 55998 -14054
rect 56032 -14828 56300 -14054
rect 56410 -14098 56430 -13499
rect 56380 -14275 56430 -14098
rect 56464 -14275 56470 -13499
rect 56380 -14287 56470 -14275
rect 56552 -13499 56750 -13487
rect 56552 -14275 56558 -13499
rect 56592 -13638 56750 -13499
rect 57066 -13480 57098 -13450
rect 57368 -13450 57372 -13364
rect 58896 -13359 59076 -13350
rect 58896 -13360 59084 -13359
rect 59156 -13360 59202 -13359
rect 57368 -13480 57396 -13450
rect 57066 -13610 57086 -13480
rect 57376 -13610 57396 -13480
rect 56592 -14275 56610 -13638
rect 57066 -13640 57396 -13610
rect 56860 -13790 57060 -13778
rect 56860 -13818 57236 -13790
rect 56860 -13948 56900 -13818
rect 57020 -13948 57236 -13818
rect 56860 -13988 57236 -13948
rect 57036 -13990 57236 -13988
rect 58556 -13880 58756 -13860
rect 58556 -14040 58576 -13880
rect 58736 -14040 58756 -13880
rect 58556 -14060 58756 -14040
rect 56552 -14278 56610 -14275
rect 57036 -14140 57446 -14130
rect 56552 -14287 56598 -14278
rect 57036 -14280 57056 -14140
rect 57416 -14280 57446 -14140
rect 56380 -14558 56440 -14287
rect 57036 -14300 57098 -14280
rect 56480 -14328 56550 -14318
rect 56480 -14398 56550 -14388
rect 57096 -14414 57098 -14334
rect 57368 -14300 57446 -14280
rect 57368 -14414 57372 -14334
rect 57096 -14430 57372 -14414
rect 58896 -14490 58926 -13360
rect 58966 -13371 59086 -13360
rect 58966 -13747 59044 -13371
rect 59078 -13747 59086 -13371
rect 58966 -13770 59086 -13747
rect 59156 -13371 59256 -13360
rect 59756 -13370 59826 -13340
rect 59966 -13352 59976 -13322
rect 60316 -13322 60346 -13316
rect 61036 -13320 61466 -13310
rect 60316 -13352 60326 -13322
rect 59966 -13360 60326 -13352
rect 59156 -13747 59162 -13371
rect 59196 -13440 59256 -13371
rect 59236 -13520 59256 -13440
rect 59196 -13640 59256 -13520
rect 59236 -13720 59256 -13640
rect 59196 -13747 59256 -13720
rect 59156 -13760 59256 -13747
rect 58966 -14080 59036 -13770
rect 59066 -13806 59176 -13800
rect 59066 -13810 59103 -13806
rect 59137 -13810 59176 -13806
rect 59066 -13880 59076 -13810
rect 59166 -13880 59176 -13810
rect 59066 -13890 59176 -13880
rect 59206 -13960 59256 -13760
rect 59376 -13390 59826 -13370
rect 59376 -13430 59476 -13390
rect 59656 -13430 59826 -13390
rect 59376 -13440 59826 -13430
rect 59376 -13490 59436 -13440
rect 59376 -13850 59386 -13490
rect 59426 -13850 59436 -13490
rect 59526 -13498 59576 -13470
rect 59526 -13532 59546 -13498
rect 59636 -13530 59706 -13470
rect 59580 -13532 59706 -13530
rect 59526 -13540 59706 -13532
rect 59476 -13582 59546 -13570
rect 59476 -13650 59502 -13582
rect 59476 -13758 59502 -13720
rect 59536 -13758 59546 -13582
rect 59476 -13770 59546 -13758
rect 59576 -13582 59636 -13570
rect 59576 -13590 59590 -13582
rect 59624 -13590 59636 -13582
rect 59576 -13770 59636 -13760
rect 59534 -13808 59592 -13802
rect 59534 -13810 59546 -13808
rect 59066 -13970 59176 -13960
rect 59066 -14040 59076 -13970
rect 59166 -14040 59176 -13970
rect 59066 -14042 59103 -14040
rect 59137 -14042 59176 -14040
rect 59066 -14050 59176 -14042
rect 59206 -13970 59266 -13960
rect 59206 -14050 59266 -14040
rect 59376 -14000 59436 -13850
rect 59516 -13842 59546 -13810
rect 59580 -13810 59592 -13808
rect 59666 -13810 59706 -13540
rect 59580 -13842 59706 -13810
rect 59516 -13880 59706 -13842
rect 59746 -13498 59936 -13470
rect 59746 -13532 59862 -13498
rect 59896 -13532 59936 -13498
rect 59746 -13540 59936 -13532
rect 61036 -13500 61206 -13320
rect 61346 -13500 61466 -13320
rect 61036 -13540 61466 -13500
rect 59746 -13800 59776 -13540
rect 60286 -13550 60476 -13540
rect 59806 -13582 59866 -13570
rect 59806 -13600 59818 -13582
rect 59852 -13600 59866 -13582
rect 59806 -13758 59818 -13740
rect 59852 -13758 59866 -13740
rect 59806 -13770 59866 -13758
rect 59900 -13580 60016 -13570
rect 59900 -13582 59916 -13580
rect 59900 -13758 59906 -13582
rect 59900 -13760 59916 -13758
rect 60006 -13760 60016 -13580
rect 60286 -13690 60306 -13550
rect 60456 -13690 60476 -13550
rect 61176 -13600 61386 -13580
rect 60286 -13700 60476 -13690
rect 61026 -13620 61136 -13610
rect 59900 -13770 60016 -13760
rect 60076 -13757 60196 -13720
rect 60076 -13791 60127 -13757
rect 60161 -13791 60196 -13757
rect 59746 -13808 59926 -13800
rect 59746 -13810 59862 -13808
rect 59896 -13810 59926 -13808
rect 59746 -13880 59826 -13810
rect 59916 -13880 59926 -13810
rect 59746 -13890 59926 -13880
rect 60076 -13849 60196 -13791
rect 60336 -13760 60446 -13700
rect 60336 -13800 60366 -13760
rect 60406 -13800 60446 -13760
rect 60636 -13757 60816 -13720
rect 60636 -13791 60671 -13757
rect 60705 -13791 60747 -13757
rect 60781 -13791 60816 -13757
rect 60076 -13880 60127 -13849
rect 60161 -13880 60196 -13849
rect 59736 -13970 59936 -13960
rect 58966 -14101 59086 -14080
rect 58966 -14477 59044 -14101
rect 59078 -14477 59086 -14101
rect 58966 -14490 59086 -14477
rect 59156 -14090 59202 -14089
rect 59156 -14101 59236 -14090
rect 59156 -14477 59162 -14101
rect 59196 -14130 59236 -14101
rect 59226 -14210 59236 -14130
rect 59196 -14360 59236 -14210
rect 59226 -14440 59236 -14360
rect 59196 -14477 59236 -14440
rect 59376 -14370 59386 -14000
rect 59426 -14370 59436 -14000
rect 59516 -14011 59706 -13970
rect 59516 -14045 59545 -14011
rect 59579 -14045 59706 -14011
rect 59516 -14050 59706 -14045
rect 59533 -14051 59591 -14050
rect 59466 -14095 59546 -14080
rect 59586 -14083 59646 -14080
rect 59466 -14130 59501 -14095
rect 59466 -14271 59501 -14210
rect 59535 -14271 59546 -14095
rect 59466 -14280 59546 -14271
rect 59583 -14095 59646 -14083
rect 59583 -14110 59589 -14095
rect 59623 -14110 59646 -14095
rect 59583 -14250 59586 -14110
rect 59583 -14271 59589 -14250
rect 59623 -14271 59646 -14250
rect 59583 -14280 59646 -14271
rect 59495 -14283 59541 -14280
rect 59583 -14283 59629 -14280
rect 59533 -14320 59591 -14315
rect 59676 -14320 59706 -14050
rect 59376 -14410 59436 -14370
rect 59506 -14380 59516 -14320
rect 59596 -14380 59706 -14320
rect 59736 -14040 59826 -13970
rect 59926 -14040 59936 -13970
rect 59736 -14045 59861 -14040
rect 59895 -14045 59936 -14040
rect 59736 -14050 59936 -14045
rect 60076 -14040 60096 -13880
rect 60176 -14040 60196 -13880
rect 59736 -14320 59766 -14050
rect 59849 -14051 59907 -14050
rect 60076 -14067 60127 -14040
rect 60161 -14067 60196 -14040
rect 59796 -14083 59856 -14080
rect 59796 -14090 59857 -14083
rect 59856 -14270 59857 -14090
rect 59796 -14271 59817 -14270
rect 59851 -14271 59857 -14270
rect 59796 -14280 59857 -14271
rect 59811 -14283 59857 -14280
rect 59899 -14090 59945 -14083
rect 59899 -14095 59916 -14090
rect 59899 -14271 59905 -14095
rect 59899 -14280 59916 -14271
rect 60006 -14280 60016 -14090
rect 60076 -14125 60196 -14067
rect 60346 -13850 60426 -13800
rect 60346 -13890 60366 -13850
rect 60406 -13890 60426 -13850
rect 60346 -13940 60426 -13890
rect 60346 -13980 60366 -13940
rect 60406 -13980 60426 -13940
rect 60346 -14020 60426 -13980
rect 60346 -14060 60366 -14020
rect 60406 -14060 60426 -14020
rect 60346 -14070 60426 -14060
rect 60636 -13849 60816 -13791
rect 60636 -13883 60671 -13849
rect 60705 -13883 60747 -13849
rect 60781 -13883 60816 -13849
rect 60636 -13941 60816 -13883
rect 60636 -13975 60671 -13941
rect 60705 -13975 60747 -13941
rect 60781 -13975 60816 -13941
rect 60636 -14033 60816 -13975
rect 60636 -14067 60671 -14033
rect 60705 -14067 60747 -14033
rect 60781 -14067 60816 -14033
rect 60076 -14159 60127 -14125
rect 60161 -14159 60196 -14125
rect 60076 -14190 60196 -14159
rect 60276 -14110 60546 -14100
rect 60276 -14125 60476 -14110
rect 60276 -14159 60297 -14125
rect 60331 -14159 60369 -14125
rect 60405 -14159 60449 -14125
rect 60276 -14170 60476 -14159
rect 60536 -14170 60546 -14110
rect 60276 -14180 60546 -14170
rect 60636 -14125 60816 -14067
rect 61026 -13730 61036 -13620
rect 61126 -13730 61136 -13620
rect 61176 -13680 61196 -13600
rect 61366 -13680 61386 -13600
rect 61176 -13700 61386 -13680
rect 61026 -13760 61136 -13730
rect 61026 -13800 61046 -13760
rect 61086 -13800 61136 -13760
rect 61026 -13850 61136 -13800
rect 61026 -13890 61046 -13850
rect 61086 -13890 61136 -13850
rect 61026 -13940 61136 -13890
rect 61026 -13980 61046 -13940
rect 61086 -13980 61136 -13940
rect 61026 -14020 61136 -13980
rect 61026 -14060 61046 -14020
rect 61086 -14060 61136 -14020
rect 61026 -14080 61136 -14060
rect 61256 -13757 61366 -13700
rect 61256 -13791 61291 -13757
rect 61325 -13791 61366 -13757
rect 61256 -13849 61366 -13791
rect 61256 -13850 61291 -13849
rect 61325 -13850 61366 -13849
rect 61256 -14060 61276 -13850
rect 61356 -14060 61366 -13850
rect 61256 -14067 61291 -14060
rect 61325 -14067 61366 -14060
rect 60636 -14159 60671 -14125
rect 60705 -14159 60747 -14125
rect 60781 -14159 60816 -14125
rect 60636 -14240 60816 -14159
rect 60966 -14124 61177 -14110
rect 60966 -14125 61129 -14124
rect 60966 -14159 60980 -14125
rect 61015 -14159 61053 -14125
rect 61088 -14158 61129 -14125
rect 61164 -14158 61177 -14124
rect 61088 -14159 61177 -14158
rect 60966 -14190 61177 -14159
rect 61256 -14125 61366 -14067
rect 61256 -14159 61291 -14125
rect 61325 -14159 61366 -14125
rect 61256 -14190 61366 -14159
rect 60466 -14250 60546 -14240
rect 59899 -14283 59945 -14280
rect 60466 -14310 60476 -14250
rect 60536 -14310 60546 -14250
rect 59849 -14320 59907 -14315
rect 60466 -14320 60546 -14310
rect 60606 -14250 60826 -14240
rect 60606 -14310 60616 -14250
rect 60736 -14310 60756 -14250
rect 60816 -14310 60826 -14250
rect 60606 -14320 60826 -14310
rect 60886 -14250 60966 -14240
rect 60886 -14310 60896 -14250
rect 60956 -14310 60966 -14250
rect 60886 -14320 60966 -14310
rect 59736 -14321 59926 -14320
rect 59736 -14355 59861 -14321
rect 59895 -14355 59926 -14321
rect 59736 -14380 59926 -14355
rect 60636 -14370 60816 -14320
rect 59376 -14420 59826 -14410
rect 59376 -14460 59476 -14420
rect 59646 -14460 59826 -14420
rect 59376 -14470 59826 -14460
rect 59156 -14490 59236 -14477
rect 58896 -14500 59086 -14490
rect 56380 -14568 57000 -14558
rect 57356 -14564 57676 -14550
rect 56440 -14574 57000 -14568
rect 57314 -14570 57676 -14564
rect 56440 -14594 57178 -14574
rect 56440 -14644 57118 -14594
rect 57168 -14644 57178 -14594
rect 57314 -14610 57326 -14570
rect 57376 -14610 57676 -14570
rect 57314 -14616 57676 -14610
rect 57356 -14630 57676 -14616
rect 56440 -14654 57178 -14644
rect 56440 -14688 57000 -14654
rect 57112 -14656 57174 -14654
rect 56380 -14758 57000 -14688
rect 56032 -14830 56038 -14828
rect 55992 -14842 56038 -14830
rect 55880 -14874 55970 -14868
rect 55870 -14878 55982 -14874
rect 55870 -14920 55880 -14878
rect 55970 -14920 55982 -14878
rect 55880 -14968 55970 -14958
rect 56120 -14998 56300 -14828
rect 57096 -14909 57372 -14878
rect 57096 -14943 57125 -14909
rect 57159 -14943 57217 -14909
rect 57251 -14943 57309 -14909
rect 57343 -14920 57372 -14909
rect 57343 -14943 57376 -14920
rect 57096 -14980 57376 -14943
rect 57066 -14990 57376 -14980
rect 56426 -14998 57376 -14990
rect 56120 -15008 57376 -14998
rect 56014 -15058 56086 -15046
rect 55570 -15178 55830 -15068
rect 53961 -15244 53988 -15206
rect 54022 -15244 54031 -15206
rect 53961 -15258 54031 -15244
rect 54910 -15206 54981 -15194
rect 54910 -15244 54916 -15206
rect 54950 -15244 54981 -15206
rect 54910 -15256 54981 -15244
rect 54911 -15258 54981 -15256
rect 55220 -15218 55330 -15208
rect 54069 -15272 54869 -15266
rect 54069 -15306 54081 -15272
rect 54857 -15278 54869 -15272
rect 54857 -15306 54880 -15278
rect 54069 -15312 54880 -15306
rect 54090 -15388 54880 -15312
rect 55330 -15318 55380 -15218
rect 55330 -15328 55480 -15318
rect 55220 -15338 55480 -15328
rect 55280 -15352 55480 -15338
rect 55280 -15358 55488 -15352
rect 55280 -15378 55300 -15358
rect 54090 -15488 54150 -15388
rect 54840 -15488 54880 -15388
rect 55288 -15392 55300 -15378
rect 55476 -15392 55488 -15358
rect 55530 -15378 55610 -15368
rect 55288 -15398 55488 -15392
rect 55520 -15402 55530 -15390
rect 55520 -15436 55526 -15402
rect 55288 -15446 55488 -15440
rect 55288 -15480 55300 -15446
rect 55476 -15480 55488 -15446
rect 55520 -15448 55530 -15436
rect 55530 -15478 55610 -15468
rect 55288 -15486 55488 -15480
rect 54090 -15508 54140 -15488
rect 54100 -15748 54140 -15508
rect 54850 -15748 54880 -15488
rect 55300 -15528 55470 -15486
rect 55300 -15668 55320 -15528
rect 55470 -15614 55482 -15542
rect 55300 -15678 55470 -15668
rect 54100 -15788 54880 -15748
rect 55710 -15998 55830 -15178
rect 56014 -15208 56020 -15058
rect 56080 -15208 56086 -15058
rect 56014 -15220 56086 -15208
rect 56120 -15208 56170 -15008
rect 56390 -15060 57376 -15008
rect 56390 -15068 57156 -15060
rect 56390 -15208 56654 -15068
rect 56120 -15258 56654 -15208
rect 56306 -15286 56654 -15258
rect 56998 -15220 57156 -15068
rect 57316 -15220 57376 -15060
rect 56998 -15286 57376 -15220
rect 56306 -15700 57376 -15286
rect 57556 -15410 57676 -14630
rect 58896 -14660 58986 -14500
rect 59756 -14520 59826 -14470
rect 59066 -14536 59176 -14530
rect 59066 -14540 59103 -14536
rect 59137 -14540 59176 -14536
rect 59066 -14600 59076 -14540
rect 59166 -14600 59176 -14540
rect 59066 -14610 59176 -14600
rect 58896 -15030 58926 -14660
rect 58966 -15030 58986 -14730
rect 59116 -14660 59506 -14640
rect 59116 -14730 59146 -14660
rect 59226 -14730 59276 -14660
rect 59356 -14730 59396 -14660
rect 59476 -14730 59506 -14660
rect 59116 -14748 59506 -14730
rect 59646 -14660 59716 -14640
rect 59706 -14720 59716 -14660
rect 59646 -14730 59716 -14720
rect 59113 -14754 59513 -14748
rect 59113 -14788 59125 -14754
rect 59501 -14788 59513 -14754
rect 59113 -14794 59513 -14788
rect 59546 -14800 59616 -14790
rect 59246 -14856 59256 -14830
rect 59113 -14862 59256 -14856
rect 59366 -14856 59376 -14830
rect 59366 -14862 59513 -14856
rect 59016 -14900 59076 -14880
rect 59113 -14896 59125 -14862
rect 59501 -14896 59513 -14862
rect 59606 -14860 59616 -14800
rect 59546 -14870 59616 -14860
rect 59113 -14902 59513 -14896
rect 59016 -14990 59076 -14960
rect 59113 -14970 59513 -14964
rect 59113 -15004 59125 -14970
rect 59501 -15004 59513 -14970
rect 59113 -15010 59513 -15004
rect 58896 -15100 58906 -15030
rect 58896 -15120 58986 -15100
rect 59116 -15030 59516 -15010
rect 59116 -15100 59146 -15030
rect 59226 -15100 59276 -15030
rect 59356 -15100 59396 -15030
rect 59476 -15100 59516 -15030
rect 59116 -15120 59516 -15100
rect 59646 -15030 59656 -14730
rect 59706 -15030 59716 -14730
rect 59756 -14700 59766 -14520
rect 59806 -14700 59826 -14520
rect 59956 -14520 60336 -14510
rect 59956 -14534 59966 -14520
rect 59946 -14540 59966 -14534
rect 60326 -14534 60336 -14520
rect 60326 -14540 60346 -14534
rect 59856 -14580 59916 -14570
rect 59946 -14574 59958 -14540
rect 60334 -14574 60346 -14540
rect 61056 -14540 61176 -14190
rect 59946 -14580 59966 -14574
rect 60326 -14580 60346 -14574
rect 60376 -14580 60436 -14560
rect 59956 -14590 60336 -14580
rect 59856 -14660 59916 -14640
rect 59946 -14648 60346 -14642
rect 59756 -14740 59826 -14700
rect 59946 -14682 59958 -14648
rect 60334 -14682 60346 -14648
rect 60376 -14660 60436 -14640
rect 61126 -14640 61176 -14540
rect 61056 -14670 61176 -14640
rect 59946 -14688 60346 -14682
rect 59946 -14740 60336 -14688
rect 59756 -14760 60536 -14740
rect 59756 -14800 59866 -14760
rect 60426 -14800 60536 -14760
rect 59756 -14810 60536 -14800
rect 59796 -14920 59806 -14810
rect 59916 -14920 59926 -14810
rect 59796 -14930 59926 -14920
rect 60436 -14830 60536 -14810
rect 60436 -14950 60446 -14830
rect 60526 -14950 60536 -14830
rect 60436 -14960 60536 -14950
rect 59646 -15040 59716 -15030
rect 59706 -15100 59716 -15040
rect 59646 -15120 59716 -15100
rect 58806 -15410 59356 -15380
rect 59846 -15390 60256 -15380
rect 59846 -15400 59996 -15390
rect 57556 -15420 59356 -15410
rect 57556 -15560 58986 -15420
rect 59126 -15560 59356 -15420
rect 57556 -15610 59356 -15560
rect 58806 -15690 59356 -15610
rect 59700 -15500 59996 -15400
rect 60106 -15400 60256 -15390
rect 60106 -15500 60400 -15400
rect 59700 -15600 60400 -15500
rect 59700 -15900 59800 -15600
rect 60300 -15900 60400 -15600
rect 55710 -16000 55910 -15998
rect 59700 -16000 60400 -15900
rect 34720 -16092 34742 -16086
rect 34730 -16182 34742 -16092
rect 16408 -16188 34742 -16182
rect 55400 -16100 56100 -16000
rect 55400 -16500 55500 -16100
rect 56000 -16500 56100 -16100
rect 55400 -16600 56100 -16500
rect 55300 -17100 55800 -17000
rect 55300 -17400 55400 -17100
rect 55700 -17400 55800 -17100
rect 54090 -17538 54890 -17498
rect 55300 -17500 55800 -17400
rect 54090 -17668 54150 -17538
rect 53510 -17720 53800 -17718
rect 53480 -17740 53800 -17720
rect 53480 -17940 53500 -17740
rect 53780 -17940 53800 -17740
rect 54080 -17798 54150 -17668
rect 54860 -17778 54890 -17538
rect 54850 -17798 54890 -17778
rect 54080 -17866 54880 -17798
rect 54079 -17872 54880 -17866
rect 54079 -17906 54091 -17872
rect 54867 -17898 54880 -17872
rect 54867 -17906 54879 -17898
rect 54079 -17912 54879 -17906
rect 53480 -17960 53800 -17940
rect 53510 -18058 53800 -17960
rect 53002 -18220 53480 -18158
rect 53000 -18358 53480 -18220
rect 53510 -18168 53520 -18058
rect 53640 -18168 53800 -18058
rect 53510 -18288 53800 -18168
rect 53970 -17934 54040 -17918
rect 53970 -17972 53998 -17934
rect 54032 -17972 54040 -17934
rect 53970 -18168 54040 -17972
rect 54920 -17934 54990 -17918
rect 54920 -17972 54926 -17934
rect 54960 -17972 54990 -17934
rect 54079 -18000 54879 -17994
rect 54079 -18034 54091 -18000
rect 54867 -18034 54879 -18000
rect 54079 -18038 54879 -18034
rect 54079 -18040 54750 -18038
rect 54090 -18088 54750 -18040
rect 54740 -18118 54750 -18088
rect 54850 -18040 54879 -18038
rect 54850 -18108 54860 -18040
rect 54840 -18118 54860 -18108
rect 54750 -18128 54860 -18118
rect 54920 -18168 54990 -17972
rect 55430 -18018 55520 -18008
rect 55290 -18128 55390 -18118
rect 53970 -18198 55290 -18168
rect 55430 -18158 55520 -18088
rect 53970 -18208 55390 -18198
rect 54050 -18218 55380 -18208
rect 54050 -18228 54880 -18218
rect 54050 -18238 54091 -18228
rect 54079 -18262 54091 -18238
rect 54867 -18238 54880 -18228
rect 54867 -18262 54879 -18238
rect 54079 -18268 54879 -18262
rect 54920 -18278 54990 -18268
rect 53510 -18306 53630 -18288
rect 53510 -18338 53526 -18306
rect 53514 -18340 53526 -18338
rect 53614 -18338 53630 -18306
rect 53940 -18290 54038 -18278
rect 53940 -18298 53998 -18290
rect 53614 -18340 53626 -18338
rect 53514 -18346 53626 -18340
rect 53000 -20108 53050 -18358
rect 53250 -18368 53480 -18358
rect 53250 -19718 53330 -18368
rect 53400 -18378 53480 -18368
rect 53400 -18390 53504 -18378
rect 53400 -19166 53464 -18390
rect 53498 -19166 53504 -18390
rect 53400 -19178 53504 -19166
rect 53636 -18388 53682 -18378
rect 53636 -18390 53760 -18388
rect 53636 -19166 53642 -18390
rect 53676 -19166 53760 -18390
rect 53940 -18398 53950 -18298
rect 54032 -18328 54038 -18290
rect 54020 -18340 54038 -18328
rect 54020 -18398 54030 -18340
rect 54079 -18356 54879 -18350
rect 54079 -18390 54091 -18356
rect 54867 -18390 54879 -18356
rect 54920 -18378 54990 -18368
rect 55320 -18368 55380 -18218
rect 54079 -18396 54879 -18390
rect 53940 -18418 54030 -18398
rect 54090 -18428 54870 -18396
rect 55320 -18402 55334 -18368
rect 55368 -18402 55380 -18368
rect 55320 -18408 55380 -18402
rect 53840 -18728 53920 -18718
rect 53840 -18838 53860 -18728
rect 53840 -18848 53920 -18838
rect 53840 -19040 53900 -18848
rect 54320 -18928 54510 -18428
rect 55440 -18438 55520 -18158
rect 55410 -18440 55520 -18438
rect 55284 -18448 55330 -18440
rect 55230 -18452 55330 -18448
rect 55230 -18458 55290 -18452
rect 55324 -18628 55330 -18452
rect 55230 -18638 55330 -18628
rect 55284 -18640 55330 -18638
rect 55372 -18448 55520 -18440
rect 55372 -18452 55430 -18448
rect 55372 -18628 55378 -18452
rect 55412 -18618 55430 -18452
rect 55510 -18618 55520 -18448
rect 55412 -18628 55520 -18618
rect 55372 -18640 55418 -18628
rect 55580 -18728 55720 -17500
rect 58776 -17670 59306 -17550
rect 58776 -17680 58966 -17670
rect 56146 -17780 57366 -17730
rect 55954 -17928 56046 -17916
rect 56146 -17928 56506 -17780
rect 55954 -18098 55960 -17928
rect 56040 -18098 56046 -17928
rect 55954 -18110 56046 -18098
rect 56120 -17958 56506 -17928
rect 56120 -18168 56190 -17958
rect 56390 -18030 56506 -17958
rect 57016 -17934 57366 -17780
rect 57586 -17830 58966 -17680
rect 59126 -17830 59306 -17670
rect 57586 -17850 59306 -17830
rect 59946 -17700 60386 -17600
rect 57586 -17880 58986 -17850
rect 59946 -17860 59956 -17700
rect 60166 -17860 60386 -17700
rect 57016 -18030 57368 -17934
rect 56390 -18070 57368 -18030
rect 56390 -18168 57126 -18070
rect 56120 -18174 57126 -18168
rect 56120 -18178 56750 -18174
rect 55880 -18218 55970 -18208
rect 55870 -18296 55880 -18250
rect 55970 -18296 55982 -18250
rect 55880 -18308 55970 -18298
rect 55000 -18738 55090 -18728
rect 55000 -18848 55090 -18838
rect 54710 -18928 54960 -18908
rect 53940 -18968 54960 -18928
rect 53940 -18972 54730 -18968
rect 53930 -18978 54730 -18972
rect 53930 -19012 53942 -18978
rect 54718 -19012 54730 -18978
rect 53930 -19018 54730 -19012
rect 53840 -19128 53858 -19040
rect 53892 -19128 53900 -19040
rect 53840 -19148 53900 -19128
rect 54762 -19038 54850 -19028
rect 54762 -19040 54770 -19038
rect 54762 -19128 54768 -19040
rect 54840 -19128 54850 -19038
rect 54762 -19140 54850 -19128
rect 54770 -19148 54850 -19140
rect 53636 -19178 53760 -19166
rect 53400 -19396 53480 -19178
rect 53514 -19216 53626 -19210
rect 53514 -19218 53526 -19216
rect 53510 -19250 53526 -19218
rect 53614 -19218 53626 -19216
rect 53614 -19250 53630 -19218
rect 53510 -19324 53630 -19250
rect 53510 -19358 53526 -19324
rect 53614 -19358 53630 -19324
rect 53680 -19238 53760 -19178
rect 53930 -19156 54730 -19150
rect 53930 -19190 53942 -19156
rect 54718 -19190 54730 -19156
rect 53930 -19196 54730 -19190
rect 53940 -19228 54720 -19196
rect 53920 -19238 54720 -19228
rect 53680 -19328 54720 -19238
rect 53514 -19364 53626 -19358
rect 53680 -19396 53760 -19328
rect 53920 -19338 54720 -19328
rect 53940 -19378 54720 -19338
rect 54900 -19368 54960 -18968
rect 55010 -18960 55090 -18848
rect 55540 -18738 55720 -18728
rect 55630 -18838 55720 -18738
rect 55130 -18874 55506 -18868
rect 55130 -18908 55142 -18874
rect 55494 -18908 55506 -18874
rect 55130 -18914 55506 -18908
rect 55010 -18994 55046 -18960
rect 55080 -18994 55090 -18960
rect 55010 -19008 55090 -18994
rect 55142 -19040 55494 -18914
rect 55540 -18960 55720 -18838
rect 55540 -18994 55556 -18960
rect 55590 -18994 55720 -18960
rect 55540 -19008 55720 -18994
rect 55780 -18340 55860 -18328
rect 55130 -19046 55506 -19040
rect 55130 -19080 55142 -19046
rect 55494 -19078 55506 -19046
rect 55494 -19080 55510 -19078
rect 55130 -19086 55510 -19080
rect 55140 -19098 55510 -19086
rect 55780 -19098 55820 -18340
rect 55140 -19116 55820 -19098
rect 55854 -19116 55860 -18340
rect 55140 -19128 55860 -19116
rect 55992 -18340 56038 -18328
rect 55992 -19116 55998 -18340
rect 56032 -18348 56038 -18340
rect 56120 -18348 56300 -18178
rect 57098 -18200 57126 -18174
rect 57356 -18200 57368 -18070
rect 57098 -18214 57368 -18200
rect 57096 -18245 57372 -18214
rect 57096 -18279 57125 -18245
rect 57159 -18279 57217 -18245
rect 57251 -18279 57309 -18245
rect 57343 -18279 57372 -18245
rect 57096 -18310 57372 -18279
rect 56032 -18706 56300 -18348
rect 56590 -18468 56660 -18458
rect 56660 -18534 57000 -18468
rect 57586 -18530 57706 -17880
rect 59946 -17890 60386 -17860
rect 57366 -18534 57706 -18530
rect 56660 -18538 57188 -18534
rect 56660 -18544 57190 -18538
rect 56660 -18594 57118 -18544
rect 57178 -18594 57190 -18544
rect 57314 -18540 57706 -18534
rect 57314 -18580 57326 -18540
rect 57366 -18580 57706 -18540
rect 57314 -18586 57706 -18580
rect 57366 -18590 57706 -18586
rect 58896 -18170 58986 -18150
rect 58896 -18230 58906 -18170
rect 58896 -18520 58926 -18230
rect 58966 -18520 58986 -18170
rect 59106 -18170 59516 -18160
rect 59106 -18230 59216 -18170
rect 59276 -18230 59326 -18170
rect 59386 -18230 59436 -18170
rect 59496 -18230 59516 -18170
rect 59106 -18247 59516 -18230
rect 59626 -18170 59706 -18130
rect 59626 -18230 59636 -18170
rect 59626 -18240 59656 -18230
rect 59106 -18280 59125 -18247
rect 59113 -18281 59125 -18280
rect 59501 -18280 59516 -18247
rect 59501 -18281 59513 -18280
rect 59113 -18287 59513 -18281
rect 59546 -18290 59616 -18280
rect 59276 -18330 59356 -18320
rect 59276 -18349 59286 -18330
rect 59113 -18355 59286 -18349
rect 59346 -18349 59356 -18330
rect 59346 -18355 59513 -18349
rect 59113 -18389 59125 -18355
rect 59501 -18389 59513 -18355
rect 59606 -18350 59616 -18290
rect 59546 -18360 59616 -18350
rect 59113 -18390 59286 -18389
rect 59346 -18390 59513 -18389
rect 59016 -18400 59076 -18390
rect 59113 -18395 59513 -18390
rect 59276 -18400 59356 -18395
rect 59546 -18410 59616 -18400
rect 59016 -18470 59076 -18460
rect 59113 -18463 59513 -18457
rect 59113 -18497 59125 -18463
rect 59501 -18497 59513 -18463
rect 59606 -18470 59616 -18410
rect 59546 -18480 59616 -18470
rect 59113 -18500 59513 -18497
rect 59113 -18503 59516 -18500
rect 58896 -18530 58986 -18520
rect 58896 -18590 58906 -18530
rect 58966 -18590 58986 -18530
rect 58896 -18592 58986 -18590
rect 59116 -18520 59516 -18503
rect 59646 -18510 59656 -18240
rect 59116 -18580 59216 -18520
rect 59276 -18580 59336 -18520
rect 59396 -18580 59436 -18520
rect 59496 -18580 59516 -18520
rect 56660 -18598 57190 -18594
rect 56590 -18600 57190 -18598
rect 56590 -18604 57188 -18600
rect 56590 -18668 57000 -18604
rect 56032 -18718 56356 -18706
rect 56032 -19116 56280 -18718
rect 55992 -19128 56280 -19116
rect 55140 -19138 55200 -19128
rect 55450 -19158 55810 -19128
rect 55870 -19166 55982 -19160
rect 55870 -19200 55882 -19166
rect 55970 -19200 55982 -19166
rect 55870 -19206 55982 -19200
rect 55140 -19218 55200 -19208
rect 55024 -19248 55116 -19236
rect 55024 -19328 55030 -19248
rect 55110 -19328 55116 -19248
rect 55024 -19340 55116 -19328
rect 55734 -19248 55816 -19236
rect 55734 -19328 55740 -19248
rect 55810 -19328 55816 -19248
rect 55734 -19340 55816 -19328
rect 55880 -19238 55970 -19206
rect 55880 -19364 55970 -19328
rect 56060 -19348 56280 -19128
rect 56350 -19348 56356 -18718
rect 56480 -18788 56550 -18778
rect 56480 -18858 56550 -18848
rect 56590 -18887 56750 -18668
rect 58894 -18686 58988 -18592
rect 59116 -18600 59516 -18580
rect 59636 -18520 59656 -18510
rect 59696 -18520 59706 -18170
rect 59856 -18340 59976 -18330
rect 59856 -18430 59866 -18340
rect 59966 -18430 59976 -18340
rect 59856 -18440 59976 -18430
rect 60436 -18420 60446 -18320
rect 60526 -18420 60536 -18320
rect 60436 -18440 60536 -18420
rect 59636 -18530 59706 -18520
rect 59696 -18590 59706 -18530
rect 59636 -18610 59706 -18590
rect 59756 -18460 60536 -18440
rect 59756 -18500 59866 -18460
rect 60426 -18500 60536 -18460
rect 59756 -18510 60536 -18500
rect 59756 -18550 59826 -18510
rect 59066 -18640 59176 -18630
rect 58896 -18750 58986 -18686
rect 59066 -18710 59076 -18640
rect 59166 -18710 59176 -18640
rect 59066 -18712 59103 -18710
rect 59137 -18712 59176 -18710
rect 59066 -18720 59176 -18712
rect 59756 -18740 59766 -18550
rect 59806 -18740 59826 -18550
rect 59956 -18568 60046 -18540
rect 59946 -18574 60046 -18568
rect 60126 -18568 60336 -18540
rect 60126 -18574 60346 -18568
rect 59856 -18610 59916 -18600
rect 59946 -18608 59958 -18574
rect 60334 -18608 60346 -18574
rect 59946 -18614 60346 -18608
rect 60376 -18620 60446 -18610
rect 59856 -18690 59916 -18680
rect 59946 -18682 60346 -18676
rect 59946 -18716 59958 -18682
rect 60334 -18716 60346 -18682
rect 60376 -18690 60446 -18680
rect 59946 -18722 59976 -18716
rect 57098 -18758 57368 -18754
rect 57096 -18764 57372 -18758
rect 57096 -18850 57098 -18764
rect 56424 -18888 56470 -18887
rect 56060 -19360 56356 -19348
rect 56410 -18899 56470 -18888
rect 53400 -19408 53504 -19396
rect 53400 -19718 53464 -19408
rect 53250 -20108 53464 -19718
rect 53000 -20184 53464 -20108
rect 53498 -20184 53504 -19408
rect 53000 -20188 53504 -20184
rect 53458 -20196 53504 -20188
rect 53636 -19408 53760 -19396
rect 53636 -20184 53642 -19408
rect 53676 -20184 53760 -19408
rect 53930 -19384 54730 -19378
rect 53930 -19418 53942 -19384
rect 54718 -19418 54730 -19384
rect 53930 -19424 54730 -19418
rect 53830 -19446 53900 -19428
rect 53830 -19534 53858 -19446
rect 53892 -19534 53900 -19446
rect 53830 -19728 53900 -19534
rect 54760 -19446 54850 -19428
rect 54760 -19534 54768 -19446
rect 54802 -19448 54850 -19446
rect 54900 -19438 55200 -19368
rect 55870 -19370 55982 -19364
rect 55870 -19404 55882 -19370
rect 55970 -19404 55982 -19370
rect 55450 -19438 55810 -19408
rect 55870 -19410 55982 -19404
rect 56060 -19438 56300 -19360
rect 54900 -19442 55820 -19438
rect 56000 -19442 56300 -19438
rect 54900 -19448 55860 -19442
rect 54840 -19528 54850 -19448
rect 54802 -19534 54850 -19528
rect 54760 -19548 54850 -19534
rect 55130 -19454 55860 -19448
rect 55130 -19478 55820 -19454
rect 55130 -19496 55510 -19478
rect 55130 -19530 55142 -19496
rect 55494 -19498 55510 -19496
rect 55494 -19530 55506 -19498
rect 55130 -19536 55506 -19530
rect 53930 -19562 54730 -19556
rect 53930 -19596 53942 -19562
rect 54718 -19596 54730 -19562
rect 55020 -19582 55090 -19568
rect 53930 -19602 54730 -19596
rect 53940 -19608 54730 -19602
rect 54920 -19598 54980 -19588
rect 53940 -19648 54920 -19608
rect 53830 -19738 53920 -19728
rect 53830 -19848 53850 -19738
rect 53830 -19858 53920 -19848
rect 54320 -20148 54510 -19648
rect 54710 -19668 54920 -19648
rect 54910 -19678 54980 -19668
rect 55020 -19616 55046 -19582
rect 55080 -19616 55090 -19582
rect 55020 -19728 55090 -19616
rect 55142 -19662 55494 -19536
rect 55540 -19582 55620 -19568
rect 55540 -19616 55556 -19582
rect 55590 -19616 55620 -19582
rect 55130 -19668 55506 -19662
rect 55130 -19702 55142 -19668
rect 55494 -19702 55506 -19668
rect 55130 -19708 55506 -19702
rect 55000 -19738 55090 -19728
rect 55000 -19848 55090 -19838
rect 55540 -19728 55620 -19616
rect 55540 -19738 55630 -19728
rect 55630 -19838 55680 -19748
rect 55540 -19848 55680 -19838
rect 55274 -19938 55320 -19936
rect 55220 -19948 55320 -19938
rect 55220 -20124 55280 -20118
rect 55314 -20124 55320 -19948
rect 55220 -20128 55320 -20124
rect 55274 -20136 55320 -20128
rect 55362 -19948 55408 -19936
rect 55362 -20124 55368 -19948
rect 55402 -19958 55510 -19948
rect 55402 -20124 55410 -19958
rect 55362 -20128 55410 -20124
rect 55500 -20128 55510 -19958
rect 55362 -20136 55510 -20128
rect 55390 -20138 55510 -20136
rect 53636 -20188 53760 -20184
rect 53636 -20196 53682 -20188
rect 53940 -20208 54020 -20168
rect 54080 -20182 54860 -20148
rect 55311 -20174 55371 -20168
rect 53514 -20234 53626 -20228
rect 53514 -20238 53526 -20234
rect 53510 -20268 53526 -20238
rect 53614 -20238 53626 -20234
rect 53614 -20268 53630 -20238
rect 53510 -20328 53630 -20268
rect 53940 -20288 53950 -20208
rect 54010 -20238 54020 -20208
rect 54069 -20188 54869 -20182
rect 54069 -20222 54081 -20188
rect 54857 -20222 54869 -20188
rect 54069 -20228 54869 -20222
rect 54910 -20198 54980 -20188
rect 54010 -20250 54028 -20238
rect 54022 -20288 54028 -20250
rect 53940 -20300 54028 -20288
rect 53940 -20308 54020 -20300
rect 54910 -20308 54980 -20298
rect 55311 -20208 55324 -20174
rect 55358 -20208 55371 -20174
rect 54070 -20310 54870 -20308
rect 54069 -20316 54870 -20310
rect 54069 -20338 54081 -20316
rect 54041 -20350 54081 -20338
rect 54857 -20318 54870 -20316
rect 54857 -20350 54880 -20318
rect 55311 -20348 55371 -20208
rect 54041 -20358 54880 -20350
rect 55240 -20358 55371 -20348
rect 54041 -20368 55240 -20358
rect 53510 -20458 53630 -20448
rect 53961 -20408 55240 -20368
rect 53961 -20606 54031 -20408
rect 54730 -20468 54860 -20458
rect 54730 -20488 54740 -20468
rect 54080 -20538 54740 -20488
rect 54069 -20544 54740 -20538
rect 54850 -20538 54860 -20468
rect 54850 -20544 54869 -20538
rect 54069 -20578 54081 -20544
rect 54857 -20578 54869 -20544
rect 54069 -20584 54869 -20578
rect 54911 -20594 54981 -20408
rect 55370 -20408 55371 -20358
rect 55240 -20428 55370 -20418
rect 55410 -20448 55510 -20138
rect 55410 -20558 55510 -20538
rect 55570 -20468 55680 -19848
rect 55780 -20230 55820 -19478
rect 55854 -20230 55860 -19454
rect 55780 -20238 55860 -20230
rect 55814 -20242 55860 -20238
rect 55992 -19454 56300 -19442
rect 55992 -20230 55998 -19454
rect 56032 -20228 56300 -19454
rect 56410 -19498 56430 -18899
rect 56380 -19675 56430 -19498
rect 56464 -19675 56470 -18899
rect 56380 -19687 56470 -19675
rect 56552 -18899 56750 -18887
rect 56552 -19675 56558 -18899
rect 56592 -19038 56750 -18899
rect 57066 -18880 57098 -18850
rect 57368 -18850 57372 -18764
rect 58896 -18759 59076 -18750
rect 58896 -18760 59084 -18759
rect 59156 -18760 59202 -18759
rect 57368 -18880 57396 -18850
rect 57066 -19010 57086 -18880
rect 57376 -19010 57396 -18880
rect 56592 -19675 56610 -19038
rect 57066 -19040 57396 -19010
rect 56860 -19190 57060 -19178
rect 56860 -19218 57236 -19190
rect 56860 -19348 56900 -19218
rect 57020 -19348 57236 -19218
rect 56860 -19388 57236 -19348
rect 57036 -19390 57236 -19388
rect 58556 -19280 58756 -19260
rect 58556 -19440 58576 -19280
rect 58736 -19440 58756 -19280
rect 58556 -19460 58756 -19440
rect 56552 -19678 56610 -19675
rect 57036 -19540 57446 -19530
rect 56552 -19687 56598 -19678
rect 57036 -19680 57056 -19540
rect 57416 -19680 57446 -19540
rect 56380 -19958 56440 -19687
rect 57036 -19700 57098 -19680
rect 56480 -19728 56550 -19718
rect 56480 -19798 56550 -19788
rect 57096 -19814 57098 -19734
rect 57368 -19700 57446 -19680
rect 57368 -19814 57372 -19734
rect 57096 -19830 57372 -19814
rect 58896 -19890 58926 -18760
rect 58966 -18771 59086 -18760
rect 58966 -19147 59044 -18771
rect 59078 -19147 59086 -18771
rect 58966 -19170 59086 -19147
rect 59156 -18771 59256 -18760
rect 59756 -18770 59826 -18740
rect 59966 -18752 59976 -18722
rect 60316 -18722 60346 -18716
rect 61036 -18720 61466 -18710
rect 60316 -18752 60326 -18722
rect 59966 -18760 60326 -18752
rect 59156 -19147 59162 -18771
rect 59196 -18840 59256 -18771
rect 59236 -18920 59256 -18840
rect 59196 -19040 59256 -18920
rect 59236 -19120 59256 -19040
rect 59196 -19147 59256 -19120
rect 59156 -19160 59256 -19147
rect 58966 -19480 59036 -19170
rect 59066 -19206 59176 -19200
rect 59066 -19210 59103 -19206
rect 59137 -19210 59176 -19206
rect 59066 -19280 59076 -19210
rect 59166 -19280 59176 -19210
rect 59066 -19290 59176 -19280
rect 59206 -19360 59256 -19160
rect 59376 -18790 59826 -18770
rect 59376 -18830 59476 -18790
rect 59656 -18830 59826 -18790
rect 59376 -18840 59826 -18830
rect 59376 -18890 59436 -18840
rect 59376 -19250 59386 -18890
rect 59426 -19250 59436 -18890
rect 59526 -18898 59576 -18870
rect 59526 -18932 59546 -18898
rect 59636 -18930 59706 -18870
rect 59580 -18932 59706 -18930
rect 59526 -18940 59706 -18932
rect 59476 -18982 59546 -18970
rect 59476 -19050 59502 -18982
rect 59476 -19158 59502 -19120
rect 59536 -19158 59546 -18982
rect 59476 -19170 59546 -19158
rect 59576 -18982 59636 -18970
rect 59576 -18990 59590 -18982
rect 59624 -18990 59636 -18982
rect 59576 -19170 59636 -19160
rect 59534 -19208 59592 -19202
rect 59534 -19210 59546 -19208
rect 59066 -19370 59176 -19360
rect 59066 -19440 59076 -19370
rect 59166 -19440 59176 -19370
rect 59066 -19442 59103 -19440
rect 59137 -19442 59176 -19440
rect 59066 -19450 59176 -19442
rect 59206 -19370 59266 -19360
rect 59206 -19450 59266 -19440
rect 59376 -19400 59436 -19250
rect 59516 -19242 59546 -19210
rect 59580 -19210 59592 -19208
rect 59666 -19210 59706 -18940
rect 59580 -19242 59706 -19210
rect 59516 -19280 59706 -19242
rect 59746 -18898 59936 -18870
rect 59746 -18932 59862 -18898
rect 59896 -18932 59936 -18898
rect 59746 -18940 59936 -18932
rect 61036 -18900 61206 -18720
rect 61346 -18900 61466 -18720
rect 61036 -18940 61466 -18900
rect 59746 -19200 59776 -18940
rect 60286 -18950 60476 -18940
rect 59806 -18982 59866 -18970
rect 59806 -19000 59818 -18982
rect 59852 -19000 59866 -18982
rect 59806 -19158 59818 -19140
rect 59852 -19158 59866 -19140
rect 59806 -19170 59866 -19158
rect 59900 -18980 60016 -18970
rect 59900 -18982 59916 -18980
rect 59900 -19158 59906 -18982
rect 59900 -19160 59916 -19158
rect 60006 -19160 60016 -18980
rect 60286 -19090 60306 -18950
rect 60456 -19090 60476 -18950
rect 61176 -19000 61386 -18980
rect 60286 -19100 60476 -19090
rect 61026 -19020 61136 -19010
rect 59900 -19170 60016 -19160
rect 60076 -19157 60196 -19120
rect 60076 -19191 60127 -19157
rect 60161 -19191 60196 -19157
rect 59746 -19208 59926 -19200
rect 59746 -19210 59862 -19208
rect 59896 -19210 59926 -19208
rect 59746 -19280 59826 -19210
rect 59916 -19280 59926 -19210
rect 59746 -19290 59926 -19280
rect 60076 -19249 60196 -19191
rect 60336 -19160 60446 -19100
rect 60336 -19200 60366 -19160
rect 60406 -19200 60446 -19160
rect 60636 -19157 60816 -19120
rect 60636 -19191 60671 -19157
rect 60705 -19191 60747 -19157
rect 60781 -19191 60816 -19157
rect 60076 -19280 60127 -19249
rect 60161 -19280 60196 -19249
rect 59736 -19370 59936 -19360
rect 58966 -19501 59086 -19480
rect 58966 -19877 59044 -19501
rect 59078 -19877 59086 -19501
rect 58966 -19890 59086 -19877
rect 59156 -19490 59202 -19489
rect 59156 -19501 59236 -19490
rect 59156 -19877 59162 -19501
rect 59196 -19530 59236 -19501
rect 59226 -19610 59236 -19530
rect 59196 -19760 59236 -19610
rect 59226 -19840 59236 -19760
rect 59196 -19877 59236 -19840
rect 59376 -19770 59386 -19400
rect 59426 -19770 59436 -19400
rect 59516 -19411 59706 -19370
rect 59516 -19445 59545 -19411
rect 59579 -19445 59706 -19411
rect 59516 -19450 59706 -19445
rect 59533 -19451 59591 -19450
rect 59466 -19495 59546 -19480
rect 59586 -19483 59646 -19480
rect 59466 -19530 59501 -19495
rect 59466 -19671 59501 -19610
rect 59535 -19671 59546 -19495
rect 59466 -19680 59546 -19671
rect 59583 -19495 59646 -19483
rect 59583 -19510 59589 -19495
rect 59623 -19510 59646 -19495
rect 59583 -19650 59586 -19510
rect 59583 -19671 59589 -19650
rect 59623 -19671 59646 -19650
rect 59583 -19680 59646 -19671
rect 59495 -19683 59541 -19680
rect 59583 -19683 59629 -19680
rect 59533 -19720 59591 -19715
rect 59676 -19720 59706 -19450
rect 59376 -19810 59436 -19770
rect 59506 -19780 59516 -19720
rect 59596 -19780 59706 -19720
rect 59736 -19440 59826 -19370
rect 59926 -19440 59936 -19370
rect 59736 -19445 59861 -19440
rect 59895 -19445 59936 -19440
rect 59736 -19450 59936 -19445
rect 60076 -19440 60096 -19280
rect 60176 -19440 60196 -19280
rect 59736 -19720 59766 -19450
rect 59849 -19451 59907 -19450
rect 60076 -19467 60127 -19440
rect 60161 -19467 60196 -19440
rect 59796 -19483 59856 -19480
rect 59796 -19490 59857 -19483
rect 59856 -19670 59857 -19490
rect 59796 -19671 59817 -19670
rect 59851 -19671 59857 -19670
rect 59796 -19680 59857 -19671
rect 59811 -19683 59857 -19680
rect 59899 -19490 59945 -19483
rect 59899 -19495 59916 -19490
rect 59899 -19671 59905 -19495
rect 59899 -19680 59916 -19671
rect 60006 -19680 60016 -19490
rect 60076 -19525 60196 -19467
rect 60346 -19250 60426 -19200
rect 60346 -19290 60366 -19250
rect 60406 -19290 60426 -19250
rect 60346 -19340 60426 -19290
rect 60346 -19380 60366 -19340
rect 60406 -19380 60426 -19340
rect 60346 -19420 60426 -19380
rect 60346 -19460 60366 -19420
rect 60406 -19460 60426 -19420
rect 60346 -19470 60426 -19460
rect 60636 -19249 60816 -19191
rect 60636 -19283 60671 -19249
rect 60705 -19283 60747 -19249
rect 60781 -19283 60816 -19249
rect 60636 -19341 60816 -19283
rect 60636 -19375 60671 -19341
rect 60705 -19375 60747 -19341
rect 60781 -19375 60816 -19341
rect 60636 -19433 60816 -19375
rect 60636 -19467 60671 -19433
rect 60705 -19467 60747 -19433
rect 60781 -19467 60816 -19433
rect 60076 -19559 60127 -19525
rect 60161 -19559 60196 -19525
rect 60076 -19590 60196 -19559
rect 60276 -19510 60546 -19500
rect 60276 -19525 60476 -19510
rect 60276 -19559 60297 -19525
rect 60331 -19559 60369 -19525
rect 60405 -19559 60449 -19525
rect 60276 -19570 60476 -19559
rect 60536 -19570 60546 -19510
rect 60276 -19580 60546 -19570
rect 60636 -19525 60816 -19467
rect 61026 -19130 61036 -19020
rect 61126 -19130 61136 -19020
rect 61176 -19080 61196 -19000
rect 61366 -19080 61386 -19000
rect 61176 -19100 61386 -19080
rect 61026 -19160 61136 -19130
rect 61026 -19200 61046 -19160
rect 61086 -19200 61136 -19160
rect 61026 -19250 61136 -19200
rect 61026 -19290 61046 -19250
rect 61086 -19290 61136 -19250
rect 61026 -19340 61136 -19290
rect 61026 -19380 61046 -19340
rect 61086 -19380 61136 -19340
rect 61026 -19420 61136 -19380
rect 61026 -19460 61046 -19420
rect 61086 -19460 61136 -19420
rect 61026 -19480 61136 -19460
rect 61256 -19157 61366 -19100
rect 61256 -19191 61291 -19157
rect 61325 -19191 61366 -19157
rect 61256 -19249 61366 -19191
rect 61256 -19250 61291 -19249
rect 61325 -19250 61366 -19249
rect 61256 -19460 61276 -19250
rect 61356 -19460 61366 -19250
rect 61256 -19467 61291 -19460
rect 61325 -19467 61366 -19460
rect 60636 -19559 60671 -19525
rect 60705 -19559 60747 -19525
rect 60781 -19559 60816 -19525
rect 60636 -19640 60816 -19559
rect 60966 -19524 61177 -19510
rect 60966 -19525 61129 -19524
rect 60966 -19559 60980 -19525
rect 61015 -19559 61053 -19525
rect 61088 -19558 61129 -19525
rect 61164 -19558 61177 -19524
rect 61088 -19559 61177 -19558
rect 60966 -19590 61177 -19559
rect 61256 -19525 61366 -19467
rect 61256 -19559 61291 -19525
rect 61325 -19559 61366 -19525
rect 61256 -19590 61366 -19559
rect 60466 -19650 60546 -19640
rect 59899 -19683 59945 -19680
rect 60466 -19710 60476 -19650
rect 60536 -19710 60546 -19650
rect 59849 -19720 59907 -19715
rect 60466 -19720 60546 -19710
rect 60606 -19650 60826 -19640
rect 60606 -19710 60616 -19650
rect 60736 -19710 60756 -19650
rect 60816 -19710 60826 -19650
rect 60606 -19720 60826 -19710
rect 60886 -19650 60966 -19640
rect 60886 -19710 60896 -19650
rect 60956 -19710 60966 -19650
rect 60886 -19720 60966 -19710
rect 59736 -19721 59926 -19720
rect 59736 -19755 59861 -19721
rect 59895 -19755 59926 -19721
rect 59736 -19780 59926 -19755
rect 60636 -19770 60816 -19720
rect 59376 -19820 59826 -19810
rect 59376 -19860 59476 -19820
rect 59646 -19860 59826 -19820
rect 59376 -19870 59826 -19860
rect 59156 -19890 59236 -19877
rect 58896 -19900 59086 -19890
rect 56380 -19968 57000 -19958
rect 57356 -19964 57676 -19950
rect 56440 -19974 57000 -19968
rect 57314 -19970 57676 -19964
rect 56440 -19994 57178 -19974
rect 56440 -20044 57118 -19994
rect 57168 -20044 57178 -19994
rect 57314 -20010 57326 -19970
rect 57376 -20010 57676 -19970
rect 57314 -20016 57676 -20010
rect 57356 -20030 57676 -20016
rect 56440 -20054 57178 -20044
rect 56440 -20088 57000 -20054
rect 57112 -20056 57174 -20054
rect 56380 -20158 57000 -20088
rect 56032 -20230 56038 -20228
rect 55992 -20242 56038 -20230
rect 55880 -20274 55970 -20268
rect 55870 -20278 55982 -20274
rect 55870 -20320 55880 -20278
rect 55970 -20320 55982 -20278
rect 55880 -20368 55970 -20358
rect 56120 -20398 56300 -20228
rect 57096 -20309 57372 -20278
rect 57096 -20343 57125 -20309
rect 57159 -20343 57217 -20309
rect 57251 -20343 57309 -20309
rect 57343 -20320 57372 -20309
rect 57343 -20343 57376 -20320
rect 57096 -20380 57376 -20343
rect 57066 -20390 57376 -20380
rect 56426 -20398 57376 -20390
rect 56120 -20408 57376 -20398
rect 56014 -20458 56086 -20446
rect 55570 -20578 55830 -20468
rect 53961 -20644 53988 -20606
rect 54022 -20644 54031 -20606
rect 53961 -20658 54031 -20644
rect 54910 -20606 54981 -20594
rect 54910 -20644 54916 -20606
rect 54950 -20644 54981 -20606
rect 54910 -20656 54981 -20644
rect 54911 -20658 54981 -20656
rect 55220 -20618 55330 -20608
rect 54069 -20672 54869 -20666
rect 54069 -20706 54081 -20672
rect 54857 -20678 54869 -20672
rect 54857 -20706 54880 -20678
rect 54069 -20712 54880 -20706
rect 54090 -20788 54880 -20712
rect 55330 -20718 55380 -20618
rect 55330 -20728 55480 -20718
rect 55220 -20738 55480 -20728
rect 55280 -20752 55480 -20738
rect 55280 -20758 55488 -20752
rect 55280 -20778 55300 -20758
rect 54090 -20888 54150 -20788
rect 54840 -20888 54880 -20788
rect 55288 -20792 55300 -20778
rect 55476 -20792 55488 -20758
rect 55530 -20778 55610 -20768
rect 55288 -20798 55488 -20792
rect 55520 -20802 55530 -20790
rect 55520 -20836 55526 -20802
rect 55288 -20846 55488 -20840
rect 55288 -20880 55300 -20846
rect 55476 -20880 55488 -20846
rect 55520 -20848 55530 -20836
rect 55530 -20878 55610 -20868
rect 55288 -20886 55488 -20880
rect 54090 -20908 54140 -20888
rect 54100 -21148 54140 -20908
rect 54850 -21148 54880 -20888
rect 55300 -20928 55470 -20886
rect 55300 -21068 55320 -20928
rect 55470 -21014 55482 -20942
rect 55300 -21078 55470 -21068
rect 54100 -21188 54880 -21148
rect 55710 -21398 55830 -20578
rect 56014 -20608 56020 -20458
rect 56080 -20608 56086 -20458
rect 56014 -20620 56086 -20608
rect 56120 -20608 56170 -20408
rect 56390 -20460 57376 -20408
rect 56390 -20468 57156 -20460
rect 56390 -20608 56654 -20468
rect 56120 -20658 56654 -20608
rect 56306 -20686 56654 -20658
rect 56998 -20620 57156 -20468
rect 57316 -20620 57376 -20460
rect 56998 -20686 57376 -20620
rect 56306 -21100 57376 -20686
rect 57556 -20810 57676 -20030
rect 58896 -20060 58986 -19900
rect 59756 -19920 59826 -19870
rect 59066 -19936 59176 -19930
rect 59066 -19940 59103 -19936
rect 59137 -19940 59176 -19936
rect 59066 -20000 59076 -19940
rect 59166 -20000 59176 -19940
rect 59066 -20010 59176 -20000
rect 58896 -20430 58926 -20060
rect 58966 -20430 58986 -20130
rect 59116 -20060 59506 -20040
rect 59116 -20130 59146 -20060
rect 59226 -20130 59276 -20060
rect 59356 -20130 59396 -20060
rect 59476 -20130 59506 -20060
rect 59116 -20148 59506 -20130
rect 59646 -20060 59716 -20040
rect 59706 -20120 59716 -20060
rect 59646 -20130 59716 -20120
rect 59113 -20154 59513 -20148
rect 59113 -20188 59125 -20154
rect 59501 -20188 59513 -20154
rect 59113 -20194 59513 -20188
rect 59546 -20200 59616 -20190
rect 59246 -20256 59256 -20230
rect 59113 -20262 59256 -20256
rect 59366 -20256 59376 -20230
rect 59366 -20262 59513 -20256
rect 59016 -20300 59076 -20280
rect 59113 -20296 59125 -20262
rect 59501 -20296 59513 -20262
rect 59606 -20260 59616 -20200
rect 59546 -20270 59616 -20260
rect 59113 -20302 59513 -20296
rect 59016 -20390 59076 -20360
rect 59113 -20370 59513 -20364
rect 59113 -20404 59125 -20370
rect 59501 -20404 59513 -20370
rect 59113 -20410 59513 -20404
rect 58896 -20500 58906 -20430
rect 58896 -20520 58986 -20500
rect 59116 -20430 59516 -20410
rect 59116 -20500 59146 -20430
rect 59226 -20500 59276 -20430
rect 59356 -20500 59396 -20430
rect 59476 -20500 59516 -20430
rect 59116 -20520 59516 -20500
rect 59646 -20430 59656 -20130
rect 59706 -20430 59716 -20130
rect 59756 -20100 59766 -19920
rect 59806 -20100 59826 -19920
rect 59956 -19920 60336 -19910
rect 59956 -19934 59966 -19920
rect 59946 -19940 59966 -19934
rect 60326 -19934 60336 -19920
rect 60326 -19940 60346 -19934
rect 59856 -19980 59916 -19970
rect 59946 -19974 59958 -19940
rect 60334 -19974 60346 -19940
rect 61056 -19940 61176 -19590
rect 59946 -19980 59966 -19974
rect 60326 -19980 60346 -19974
rect 60376 -19980 60436 -19960
rect 59956 -19990 60336 -19980
rect 59856 -20060 59916 -20040
rect 59946 -20048 60346 -20042
rect 59756 -20140 59826 -20100
rect 59946 -20082 59958 -20048
rect 60334 -20082 60346 -20048
rect 60376 -20060 60436 -20040
rect 61126 -20040 61176 -19940
rect 61056 -20070 61176 -20040
rect 59946 -20088 60346 -20082
rect 59946 -20140 60336 -20088
rect 59756 -20160 60536 -20140
rect 59756 -20200 59866 -20160
rect 60426 -20200 60536 -20160
rect 59756 -20210 60536 -20200
rect 59796 -20320 59806 -20210
rect 59916 -20320 59926 -20210
rect 59796 -20330 59926 -20320
rect 60436 -20230 60536 -20210
rect 60436 -20350 60446 -20230
rect 60526 -20350 60536 -20230
rect 60436 -20360 60536 -20350
rect 59646 -20440 59716 -20430
rect 59706 -20500 59716 -20440
rect 59646 -20520 59716 -20500
rect 58806 -20810 59356 -20780
rect 59846 -20790 60256 -20780
rect 59846 -20800 59996 -20790
rect 57556 -20820 59356 -20810
rect 57556 -20960 58986 -20820
rect 59126 -20960 59356 -20820
rect 57556 -21010 59356 -20960
rect 58806 -21090 59356 -21010
rect 59700 -20900 59996 -20800
rect 60106 -20800 60256 -20790
rect 60106 -20900 60400 -20800
rect 59700 -21000 60400 -20900
rect 59700 -21300 59800 -21000
rect 60300 -21300 60400 -21000
rect 55710 -21400 55910 -21398
rect 59700 -21400 60400 -21300
rect 55400 -21500 56200 -21400
rect 55400 -21900 55500 -21500
rect 56100 -21900 56200 -21500
rect 55400 -22000 56200 -21900
rect 55360 -22480 55800 -22400
rect 55360 -22760 55440 -22480
rect 55720 -22760 55800 -22480
rect 55360 -22840 55800 -22760
rect 54090 -22938 54890 -22898
rect 54090 -23068 54150 -22938
rect 53510 -23120 53800 -23118
rect 53460 -23140 53800 -23120
rect 53460 -23340 53480 -23140
rect 53780 -23340 53800 -23140
rect 54080 -23198 54150 -23068
rect 54860 -23178 54890 -22938
rect 54850 -23198 54890 -23178
rect 54080 -23266 54880 -23198
rect 54079 -23272 54880 -23266
rect 54079 -23306 54091 -23272
rect 54867 -23298 54880 -23272
rect 54867 -23306 54879 -23298
rect 54079 -23312 54879 -23306
rect 53460 -23360 53800 -23340
rect 53510 -23458 53800 -23360
rect 53002 -23620 53480 -23558
rect 53000 -23758 53480 -23620
rect 53510 -23568 53520 -23458
rect 53640 -23568 53800 -23458
rect 53510 -23688 53800 -23568
rect 53970 -23334 54040 -23318
rect 53970 -23372 53998 -23334
rect 54032 -23372 54040 -23334
rect 53970 -23568 54040 -23372
rect 54920 -23334 54990 -23318
rect 54920 -23372 54926 -23334
rect 54960 -23372 54990 -23334
rect 54079 -23400 54879 -23394
rect 54079 -23434 54091 -23400
rect 54867 -23434 54879 -23400
rect 54079 -23438 54879 -23434
rect 54079 -23440 54750 -23438
rect 54090 -23488 54750 -23440
rect 54740 -23518 54750 -23488
rect 54850 -23440 54879 -23438
rect 54850 -23508 54860 -23440
rect 54840 -23518 54860 -23508
rect 54750 -23528 54860 -23518
rect 54920 -23568 54990 -23372
rect 55430 -23418 55520 -23408
rect 55290 -23528 55390 -23518
rect 53970 -23598 55290 -23568
rect 55430 -23558 55520 -23488
rect 53970 -23608 55390 -23598
rect 54050 -23618 55380 -23608
rect 54050 -23628 54880 -23618
rect 54050 -23638 54091 -23628
rect 54079 -23662 54091 -23638
rect 54867 -23638 54880 -23628
rect 54867 -23662 54879 -23638
rect 54079 -23668 54879 -23662
rect 54920 -23678 54990 -23668
rect 53510 -23706 53630 -23688
rect 53510 -23738 53526 -23706
rect 53514 -23740 53526 -23738
rect 53614 -23738 53630 -23706
rect 53940 -23690 54038 -23678
rect 53940 -23698 53998 -23690
rect 53614 -23740 53626 -23738
rect 53514 -23746 53626 -23740
rect 53000 -25508 53050 -23758
rect 53250 -23768 53480 -23758
rect 53250 -25118 53330 -23768
rect 53400 -23778 53480 -23768
rect 53400 -23790 53504 -23778
rect 53400 -24566 53464 -23790
rect 53498 -24566 53504 -23790
rect 53400 -24578 53504 -24566
rect 53636 -23788 53682 -23778
rect 53636 -23790 53760 -23788
rect 53636 -24566 53642 -23790
rect 53676 -24566 53760 -23790
rect 53940 -23798 53950 -23698
rect 54032 -23728 54038 -23690
rect 54020 -23740 54038 -23728
rect 54020 -23798 54030 -23740
rect 54079 -23756 54879 -23750
rect 54079 -23790 54091 -23756
rect 54867 -23790 54879 -23756
rect 54920 -23778 54990 -23768
rect 55320 -23768 55380 -23618
rect 54079 -23796 54879 -23790
rect 53940 -23818 54030 -23798
rect 54090 -23828 54870 -23796
rect 55320 -23802 55334 -23768
rect 55368 -23802 55380 -23768
rect 55320 -23808 55380 -23802
rect 53840 -24128 53920 -24118
rect 53840 -24238 53860 -24128
rect 53840 -24248 53920 -24238
rect 53840 -24440 53900 -24248
rect 54320 -24328 54510 -23828
rect 55440 -23838 55520 -23558
rect 55410 -23840 55520 -23838
rect 55284 -23848 55330 -23840
rect 55230 -23852 55330 -23848
rect 55230 -23858 55290 -23852
rect 55324 -24028 55330 -23852
rect 55230 -24038 55330 -24028
rect 55284 -24040 55330 -24038
rect 55372 -23848 55520 -23840
rect 55372 -23852 55430 -23848
rect 55372 -24028 55378 -23852
rect 55412 -24018 55430 -23852
rect 55510 -24018 55520 -23848
rect 55412 -24028 55520 -24018
rect 55372 -24040 55418 -24028
rect 55580 -24128 55720 -22840
rect 58776 -23070 59306 -22950
rect 58776 -23080 58966 -23070
rect 56146 -23180 57366 -23130
rect 55954 -23328 56046 -23316
rect 56146 -23328 56506 -23180
rect 55954 -23498 55960 -23328
rect 56040 -23498 56046 -23328
rect 55954 -23510 56046 -23498
rect 56120 -23358 56506 -23328
rect 56120 -23568 56190 -23358
rect 56390 -23430 56506 -23358
rect 57016 -23334 57366 -23180
rect 57586 -23230 58966 -23080
rect 59126 -23230 59306 -23070
rect 57586 -23250 59306 -23230
rect 59946 -23100 60386 -23000
rect 57586 -23280 58986 -23250
rect 59946 -23260 59956 -23100
rect 60166 -23260 60386 -23100
rect 57016 -23430 57368 -23334
rect 56390 -23470 57368 -23430
rect 56390 -23568 57126 -23470
rect 56120 -23574 57126 -23568
rect 56120 -23578 56750 -23574
rect 55880 -23618 55970 -23608
rect 55870 -23696 55880 -23650
rect 55970 -23696 55982 -23650
rect 55880 -23708 55970 -23698
rect 55000 -24138 55090 -24128
rect 55000 -24248 55090 -24238
rect 54710 -24328 54960 -24308
rect 53940 -24368 54960 -24328
rect 53940 -24372 54730 -24368
rect 53930 -24378 54730 -24372
rect 53930 -24412 53942 -24378
rect 54718 -24412 54730 -24378
rect 53930 -24418 54730 -24412
rect 53840 -24528 53858 -24440
rect 53892 -24528 53900 -24440
rect 53840 -24548 53900 -24528
rect 54762 -24438 54850 -24428
rect 54762 -24440 54770 -24438
rect 54762 -24528 54768 -24440
rect 54840 -24528 54850 -24438
rect 54762 -24540 54850 -24528
rect 54770 -24548 54850 -24540
rect 53636 -24578 53760 -24566
rect 53400 -24796 53480 -24578
rect 53514 -24616 53626 -24610
rect 53514 -24618 53526 -24616
rect 53510 -24650 53526 -24618
rect 53614 -24618 53626 -24616
rect 53614 -24650 53630 -24618
rect 53510 -24724 53630 -24650
rect 53510 -24758 53526 -24724
rect 53614 -24758 53630 -24724
rect 53680 -24638 53760 -24578
rect 53930 -24556 54730 -24550
rect 53930 -24590 53942 -24556
rect 54718 -24590 54730 -24556
rect 53930 -24596 54730 -24590
rect 53940 -24628 54720 -24596
rect 53920 -24638 54720 -24628
rect 53680 -24728 54720 -24638
rect 53514 -24764 53626 -24758
rect 53680 -24796 53760 -24728
rect 53920 -24738 54720 -24728
rect 53940 -24778 54720 -24738
rect 54900 -24768 54960 -24368
rect 55010 -24360 55090 -24248
rect 55540 -24138 55720 -24128
rect 55630 -24238 55720 -24138
rect 55130 -24274 55506 -24268
rect 55130 -24308 55142 -24274
rect 55494 -24308 55506 -24274
rect 55130 -24314 55506 -24308
rect 55010 -24394 55046 -24360
rect 55080 -24394 55090 -24360
rect 55010 -24408 55090 -24394
rect 55142 -24440 55494 -24314
rect 55540 -24360 55720 -24238
rect 55540 -24394 55556 -24360
rect 55590 -24394 55720 -24360
rect 55540 -24408 55720 -24394
rect 55780 -23740 55860 -23728
rect 55130 -24446 55506 -24440
rect 55130 -24480 55142 -24446
rect 55494 -24478 55506 -24446
rect 55494 -24480 55510 -24478
rect 55130 -24486 55510 -24480
rect 55140 -24498 55510 -24486
rect 55780 -24498 55820 -23740
rect 55140 -24516 55820 -24498
rect 55854 -24516 55860 -23740
rect 55140 -24528 55860 -24516
rect 55992 -23740 56038 -23728
rect 55992 -24516 55998 -23740
rect 56032 -23748 56038 -23740
rect 56120 -23748 56300 -23578
rect 57098 -23600 57126 -23574
rect 57356 -23600 57368 -23470
rect 57098 -23614 57368 -23600
rect 57096 -23645 57372 -23614
rect 57096 -23679 57125 -23645
rect 57159 -23679 57217 -23645
rect 57251 -23679 57309 -23645
rect 57343 -23679 57372 -23645
rect 57096 -23710 57372 -23679
rect 56032 -24106 56300 -23748
rect 56590 -23868 56660 -23858
rect 56660 -23934 57000 -23868
rect 57586 -23930 57706 -23280
rect 59946 -23290 60386 -23260
rect 57366 -23934 57706 -23930
rect 56660 -23938 57188 -23934
rect 56660 -23944 57190 -23938
rect 56660 -23994 57118 -23944
rect 57178 -23994 57190 -23944
rect 57314 -23940 57706 -23934
rect 57314 -23980 57326 -23940
rect 57366 -23980 57706 -23940
rect 57314 -23986 57706 -23980
rect 57366 -23990 57706 -23986
rect 58896 -23570 58986 -23550
rect 58896 -23630 58906 -23570
rect 58896 -23920 58926 -23630
rect 58966 -23920 58986 -23570
rect 59106 -23570 59516 -23560
rect 59106 -23630 59216 -23570
rect 59276 -23630 59326 -23570
rect 59386 -23630 59436 -23570
rect 59496 -23630 59516 -23570
rect 59106 -23647 59516 -23630
rect 59626 -23570 59706 -23530
rect 59626 -23630 59636 -23570
rect 59626 -23640 59656 -23630
rect 59106 -23680 59125 -23647
rect 59113 -23681 59125 -23680
rect 59501 -23680 59516 -23647
rect 59501 -23681 59513 -23680
rect 59113 -23687 59513 -23681
rect 59546 -23690 59616 -23680
rect 59276 -23730 59356 -23720
rect 59276 -23749 59286 -23730
rect 59113 -23755 59286 -23749
rect 59346 -23749 59356 -23730
rect 59346 -23755 59513 -23749
rect 59113 -23789 59125 -23755
rect 59501 -23789 59513 -23755
rect 59606 -23750 59616 -23690
rect 59546 -23760 59616 -23750
rect 59113 -23790 59286 -23789
rect 59346 -23790 59513 -23789
rect 59016 -23800 59076 -23790
rect 59113 -23795 59513 -23790
rect 59276 -23800 59356 -23795
rect 59546 -23810 59616 -23800
rect 59016 -23870 59076 -23860
rect 59113 -23863 59513 -23857
rect 59113 -23897 59125 -23863
rect 59501 -23897 59513 -23863
rect 59606 -23870 59616 -23810
rect 59546 -23880 59616 -23870
rect 59113 -23900 59513 -23897
rect 59113 -23903 59516 -23900
rect 58896 -23930 58986 -23920
rect 58896 -23990 58906 -23930
rect 58966 -23990 58986 -23930
rect 58896 -23992 58986 -23990
rect 59116 -23920 59516 -23903
rect 59646 -23910 59656 -23640
rect 59116 -23980 59216 -23920
rect 59276 -23980 59336 -23920
rect 59396 -23980 59436 -23920
rect 59496 -23980 59516 -23920
rect 56660 -23998 57190 -23994
rect 56590 -24000 57190 -23998
rect 56590 -24004 57188 -24000
rect 56590 -24068 57000 -24004
rect 56032 -24118 56356 -24106
rect 56032 -24516 56280 -24118
rect 55992 -24528 56280 -24516
rect 55140 -24538 55200 -24528
rect 55450 -24558 55810 -24528
rect 55870 -24566 55982 -24560
rect 55870 -24600 55882 -24566
rect 55970 -24600 55982 -24566
rect 55870 -24606 55982 -24600
rect 55140 -24618 55200 -24608
rect 55024 -24648 55116 -24636
rect 55024 -24728 55030 -24648
rect 55110 -24728 55116 -24648
rect 55024 -24740 55116 -24728
rect 55734 -24648 55816 -24636
rect 55734 -24728 55740 -24648
rect 55810 -24728 55816 -24648
rect 55734 -24740 55816 -24728
rect 55880 -24638 55970 -24606
rect 55880 -24764 55970 -24728
rect 56060 -24748 56280 -24528
rect 56350 -24748 56356 -24118
rect 56480 -24188 56550 -24178
rect 56480 -24258 56550 -24248
rect 56590 -24287 56750 -24068
rect 58894 -24086 58988 -23992
rect 59116 -24000 59516 -23980
rect 59636 -23920 59656 -23910
rect 59696 -23920 59706 -23570
rect 59856 -23740 59976 -23730
rect 59856 -23830 59866 -23740
rect 59966 -23830 59976 -23740
rect 59856 -23840 59976 -23830
rect 60436 -23820 60446 -23720
rect 60526 -23820 60536 -23720
rect 60436 -23840 60536 -23820
rect 59636 -23930 59706 -23920
rect 59696 -23990 59706 -23930
rect 59636 -24010 59706 -23990
rect 59756 -23860 60536 -23840
rect 59756 -23900 59866 -23860
rect 60426 -23900 60536 -23860
rect 59756 -23910 60536 -23900
rect 59756 -23950 59826 -23910
rect 59066 -24040 59176 -24030
rect 58896 -24150 58986 -24086
rect 59066 -24110 59076 -24040
rect 59166 -24110 59176 -24040
rect 59066 -24112 59103 -24110
rect 59137 -24112 59176 -24110
rect 59066 -24120 59176 -24112
rect 59756 -24140 59766 -23950
rect 59806 -24140 59826 -23950
rect 59956 -23968 60046 -23940
rect 59946 -23974 60046 -23968
rect 60126 -23968 60336 -23940
rect 60126 -23974 60346 -23968
rect 59856 -24010 59916 -24000
rect 59946 -24008 59958 -23974
rect 60334 -24008 60346 -23974
rect 59946 -24014 60346 -24008
rect 60376 -24020 60446 -24010
rect 59856 -24090 59916 -24080
rect 59946 -24082 60346 -24076
rect 59946 -24116 59958 -24082
rect 60334 -24116 60346 -24082
rect 60376 -24090 60446 -24080
rect 59946 -24122 59976 -24116
rect 57098 -24158 57368 -24154
rect 57096 -24164 57372 -24158
rect 57096 -24250 57098 -24164
rect 56424 -24288 56470 -24287
rect 56060 -24760 56356 -24748
rect 56410 -24299 56470 -24288
rect 53400 -24808 53504 -24796
rect 53400 -25118 53464 -24808
rect 53250 -25508 53464 -25118
rect 53000 -25584 53464 -25508
rect 53498 -25584 53504 -24808
rect 53000 -25588 53504 -25584
rect 53458 -25596 53504 -25588
rect 53636 -24808 53760 -24796
rect 53636 -25584 53642 -24808
rect 53676 -25584 53760 -24808
rect 53930 -24784 54730 -24778
rect 53930 -24818 53942 -24784
rect 54718 -24818 54730 -24784
rect 53930 -24824 54730 -24818
rect 53830 -24846 53900 -24828
rect 53830 -24934 53858 -24846
rect 53892 -24934 53900 -24846
rect 53830 -25128 53900 -24934
rect 54760 -24846 54850 -24828
rect 54760 -24934 54768 -24846
rect 54802 -24848 54850 -24846
rect 54900 -24838 55200 -24768
rect 55870 -24770 55982 -24764
rect 55870 -24804 55882 -24770
rect 55970 -24804 55982 -24770
rect 55450 -24838 55810 -24808
rect 55870 -24810 55982 -24804
rect 56060 -24838 56300 -24760
rect 54900 -24842 55820 -24838
rect 56000 -24842 56300 -24838
rect 54900 -24848 55860 -24842
rect 54840 -24928 54850 -24848
rect 54802 -24934 54850 -24928
rect 54760 -24948 54850 -24934
rect 55130 -24854 55860 -24848
rect 55130 -24878 55820 -24854
rect 55130 -24896 55510 -24878
rect 55130 -24930 55142 -24896
rect 55494 -24898 55510 -24896
rect 55494 -24930 55506 -24898
rect 55130 -24936 55506 -24930
rect 53930 -24962 54730 -24956
rect 53930 -24996 53942 -24962
rect 54718 -24996 54730 -24962
rect 55020 -24982 55090 -24968
rect 53930 -25002 54730 -24996
rect 53940 -25008 54730 -25002
rect 54920 -24998 54980 -24988
rect 53940 -25048 54920 -25008
rect 53830 -25138 53920 -25128
rect 53830 -25248 53850 -25138
rect 53830 -25258 53920 -25248
rect 54320 -25548 54510 -25048
rect 54710 -25068 54920 -25048
rect 54910 -25078 54980 -25068
rect 55020 -25016 55046 -24982
rect 55080 -25016 55090 -24982
rect 55020 -25128 55090 -25016
rect 55142 -25062 55494 -24936
rect 55540 -24982 55620 -24968
rect 55540 -25016 55556 -24982
rect 55590 -25016 55620 -24982
rect 55130 -25068 55506 -25062
rect 55130 -25102 55142 -25068
rect 55494 -25102 55506 -25068
rect 55130 -25108 55506 -25102
rect 55000 -25138 55090 -25128
rect 55000 -25248 55090 -25238
rect 55540 -25128 55620 -25016
rect 55540 -25138 55630 -25128
rect 55630 -25238 55680 -25148
rect 55540 -25248 55680 -25238
rect 55274 -25338 55320 -25336
rect 55220 -25348 55320 -25338
rect 55220 -25524 55280 -25518
rect 55314 -25524 55320 -25348
rect 55220 -25528 55320 -25524
rect 55274 -25536 55320 -25528
rect 55362 -25348 55408 -25336
rect 55362 -25524 55368 -25348
rect 55402 -25358 55510 -25348
rect 55402 -25524 55410 -25358
rect 55362 -25528 55410 -25524
rect 55500 -25528 55510 -25358
rect 55362 -25536 55510 -25528
rect 55390 -25538 55510 -25536
rect 53636 -25588 53760 -25584
rect 53636 -25596 53682 -25588
rect 53940 -25608 54020 -25568
rect 54080 -25582 54860 -25548
rect 55311 -25574 55371 -25568
rect 53514 -25634 53626 -25628
rect 53514 -25638 53526 -25634
rect 53510 -25668 53526 -25638
rect 53614 -25638 53626 -25634
rect 53614 -25668 53630 -25638
rect 53510 -25728 53630 -25668
rect 53940 -25688 53950 -25608
rect 54010 -25638 54020 -25608
rect 54069 -25588 54869 -25582
rect 54069 -25622 54081 -25588
rect 54857 -25622 54869 -25588
rect 54069 -25628 54869 -25622
rect 54910 -25598 54980 -25588
rect 54010 -25650 54028 -25638
rect 54022 -25688 54028 -25650
rect 53940 -25700 54028 -25688
rect 53940 -25708 54020 -25700
rect 54910 -25708 54980 -25698
rect 55311 -25608 55324 -25574
rect 55358 -25608 55371 -25574
rect 54070 -25710 54870 -25708
rect 14400 -26400 20000 -25800
rect 14400 -27200 15000 -26400
rect 10800 -30600 15000 -27200
rect 14400 -31200 15000 -30600
rect 19400 -31200 20000 -26400
rect 26000 -26400 35800 -25800
rect 54069 -25716 54870 -25710
rect 54069 -25738 54081 -25716
rect 54041 -25750 54081 -25738
rect 54857 -25718 54870 -25716
rect 54857 -25750 54880 -25718
rect 55311 -25748 55371 -25608
rect 54041 -25758 54880 -25750
rect 55240 -25758 55371 -25748
rect 54041 -25768 55240 -25758
rect 53510 -25858 53630 -25848
rect 53961 -25808 55240 -25768
rect 53961 -26006 54031 -25808
rect 54730 -25868 54860 -25858
rect 54730 -25888 54740 -25868
rect 54080 -25938 54740 -25888
rect 54069 -25944 54740 -25938
rect 54850 -25938 54860 -25868
rect 54850 -25944 54869 -25938
rect 54069 -25978 54081 -25944
rect 54857 -25978 54869 -25944
rect 54069 -25984 54869 -25978
rect 54911 -25994 54981 -25808
rect 55370 -25808 55371 -25758
rect 55240 -25828 55370 -25818
rect 55410 -25848 55510 -25538
rect 55410 -25958 55510 -25938
rect 55570 -25868 55680 -25248
rect 55780 -25630 55820 -24878
rect 55854 -25630 55860 -24854
rect 55780 -25638 55860 -25630
rect 55814 -25642 55860 -25638
rect 55992 -24854 56300 -24842
rect 55992 -25630 55998 -24854
rect 56032 -25628 56300 -24854
rect 56410 -24898 56430 -24299
rect 56380 -25075 56430 -24898
rect 56464 -25075 56470 -24299
rect 56380 -25087 56470 -25075
rect 56552 -24299 56750 -24287
rect 56552 -25075 56558 -24299
rect 56592 -24438 56750 -24299
rect 57066 -24280 57098 -24250
rect 57368 -24250 57372 -24164
rect 58896 -24159 59076 -24150
rect 58896 -24160 59084 -24159
rect 59156 -24160 59202 -24159
rect 57368 -24280 57396 -24250
rect 57066 -24410 57086 -24280
rect 57376 -24410 57396 -24280
rect 56592 -25075 56610 -24438
rect 57066 -24440 57396 -24410
rect 56860 -24590 57060 -24578
rect 56860 -24618 57236 -24590
rect 56860 -24748 56900 -24618
rect 57020 -24748 57236 -24618
rect 56860 -24788 57236 -24748
rect 57036 -24790 57236 -24788
rect 58556 -24680 58756 -24660
rect 58556 -24840 58576 -24680
rect 58736 -24840 58756 -24680
rect 58556 -24860 58756 -24840
rect 56552 -25078 56610 -25075
rect 57036 -24940 57446 -24930
rect 56552 -25087 56598 -25078
rect 57036 -25080 57056 -24940
rect 57416 -25080 57446 -24940
rect 56380 -25358 56440 -25087
rect 57036 -25100 57098 -25080
rect 56480 -25128 56550 -25118
rect 56480 -25198 56550 -25188
rect 57096 -25214 57098 -25134
rect 57368 -25100 57446 -25080
rect 57368 -25214 57372 -25134
rect 57096 -25230 57372 -25214
rect 58896 -25290 58926 -24160
rect 58966 -24171 59086 -24160
rect 58966 -24547 59044 -24171
rect 59078 -24547 59086 -24171
rect 58966 -24570 59086 -24547
rect 59156 -24171 59256 -24160
rect 59756 -24170 59826 -24140
rect 59966 -24152 59976 -24122
rect 60316 -24122 60346 -24116
rect 61036 -24120 61466 -24110
rect 60316 -24152 60326 -24122
rect 59966 -24160 60326 -24152
rect 59156 -24547 59162 -24171
rect 59196 -24240 59256 -24171
rect 59236 -24320 59256 -24240
rect 59196 -24440 59256 -24320
rect 59236 -24520 59256 -24440
rect 59196 -24547 59256 -24520
rect 59156 -24560 59256 -24547
rect 58966 -24880 59036 -24570
rect 59066 -24606 59176 -24600
rect 59066 -24610 59103 -24606
rect 59137 -24610 59176 -24606
rect 59066 -24680 59076 -24610
rect 59166 -24680 59176 -24610
rect 59066 -24690 59176 -24680
rect 59206 -24760 59256 -24560
rect 59376 -24190 59826 -24170
rect 59376 -24230 59476 -24190
rect 59656 -24230 59826 -24190
rect 59376 -24240 59826 -24230
rect 59376 -24290 59436 -24240
rect 59376 -24650 59386 -24290
rect 59426 -24650 59436 -24290
rect 59526 -24298 59576 -24270
rect 59526 -24332 59546 -24298
rect 59636 -24330 59706 -24270
rect 59580 -24332 59706 -24330
rect 59526 -24340 59706 -24332
rect 59476 -24382 59546 -24370
rect 59476 -24450 59502 -24382
rect 59476 -24558 59502 -24520
rect 59536 -24558 59546 -24382
rect 59476 -24570 59546 -24558
rect 59576 -24382 59636 -24370
rect 59576 -24390 59590 -24382
rect 59624 -24390 59636 -24382
rect 59576 -24570 59636 -24560
rect 59534 -24608 59592 -24602
rect 59534 -24610 59546 -24608
rect 59066 -24770 59176 -24760
rect 59066 -24840 59076 -24770
rect 59166 -24840 59176 -24770
rect 59066 -24842 59103 -24840
rect 59137 -24842 59176 -24840
rect 59066 -24850 59176 -24842
rect 59206 -24770 59266 -24760
rect 59206 -24850 59266 -24840
rect 59376 -24800 59436 -24650
rect 59516 -24642 59546 -24610
rect 59580 -24610 59592 -24608
rect 59666 -24610 59706 -24340
rect 59580 -24642 59706 -24610
rect 59516 -24680 59706 -24642
rect 59746 -24298 59936 -24270
rect 59746 -24332 59862 -24298
rect 59896 -24332 59936 -24298
rect 59746 -24340 59936 -24332
rect 61036 -24300 61206 -24120
rect 61346 -24300 61466 -24120
rect 61036 -24340 61466 -24300
rect 59746 -24600 59776 -24340
rect 60286 -24350 60476 -24340
rect 59806 -24382 59866 -24370
rect 59806 -24400 59818 -24382
rect 59852 -24400 59866 -24382
rect 59806 -24558 59818 -24540
rect 59852 -24558 59866 -24540
rect 59806 -24570 59866 -24558
rect 59900 -24380 60016 -24370
rect 59900 -24382 59916 -24380
rect 59900 -24558 59906 -24382
rect 59900 -24560 59916 -24558
rect 60006 -24560 60016 -24380
rect 60286 -24490 60306 -24350
rect 60456 -24490 60476 -24350
rect 61176 -24400 61386 -24380
rect 60286 -24500 60476 -24490
rect 61026 -24420 61136 -24410
rect 59900 -24570 60016 -24560
rect 60076 -24557 60196 -24520
rect 60076 -24591 60127 -24557
rect 60161 -24591 60196 -24557
rect 59746 -24608 59926 -24600
rect 59746 -24610 59862 -24608
rect 59896 -24610 59926 -24608
rect 59746 -24680 59826 -24610
rect 59916 -24680 59926 -24610
rect 59746 -24690 59926 -24680
rect 60076 -24649 60196 -24591
rect 60336 -24560 60446 -24500
rect 60336 -24600 60366 -24560
rect 60406 -24600 60446 -24560
rect 60636 -24557 60816 -24520
rect 60636 -24591 60671 -24557
rect 60705 -24591 60747 -24557
rect 60781 -24591 60816 -24557
rect 60076 -24680 60127 -24649
rect 60161 -24680 60196 -24649
rect 59736 -24770 59936 -24760
rect 58966 -24901 59086 -24880
rect 58966 -25277 59044 -24901
rect 59078 -25277 59086 -24901
rect 58966 -25290 59086 -25277
rect 59156 -24890 59202 -24889
rect 59156 -24901 59236 -24890
rect 59156 -25277 59162 -24901
rect 59196 -24930 59236 -24901
rect 59226 -25010 59236 -24930
rect 59196 -25160 59236 -25010
rect 59226 -25240 59236 -25160
rect 59196 -25277 59236 -25240
rect 59376 -25170 59386 -24800
rect 59426 -25170 59436 -24800
rect 59516 -24811 59706 -24770
rect 59516 -24845 59545 -24811
rect 59579 -24845 59706 -24811
rect 59516 -24850 59706 -24845
rect 59533 -24851 59591 -24850
rect 59466 -24895 59546 -24880
rect 59586 -24883 59646 -24880
rect 59466 -24930 59501 -24895
rect 59466 -25071 59501 -25010
rect 59535 -25071 59546 -24895
rect 59466 -25080 59546 -25071
rect 59583 -24895 59646 -24883
rect 59583 -24910 59589 -24895
rect 59623 -24910 59646 -24895
rect 59583 -25050 59586 -24910
rect 59583 -25071 59589 -25050
rect 59623 -25071 59646 -25050
rect 59583 -25080 59646 -25071
rect 59495 -25083 59541 -25080
rect 59583 -25083 59629 -25080
rect 59533 -25120 59591 -25115
rect 59676 -25120 59706 -24850
rect 59376 -25210 59436 -25170
rect 59506 -25180 59516 -25120
rect 59596 -25180 59706 -25120
rect 59736 -24840 59826 -24770
rect 59926 -24840 59936 -24770
rect 59736 -24845 59861 -24840
rect 59895 -24845 59936 -24840
rect 59736 -24850 59936 -24845
rect 60076 -24840 60096 -24680
rect 60176 -24840 60196 -24680
rect 59736 -25120 59766 -24850
rect 59849 -24851 59907 -24850
rect 60076 -24867 60127 -24840
rect 60161 -24867 60196 -24840
rect 59796 -24883 59856 -24880
rect 59796 -24890 59857 -24883
rect 59856 -25070 59857 -24890
rect 59796 -25071 59817 -25070
rect 59851 -25071 59857 -25070
rect 59796 -25080 59857 -25071
rect 59811 -25083 59857 -25080
rect 59899 -24890 59945 -24883
rect 59899 -24895 59916 -24890
rect 59899 -25071 59905 -24895
rect 59899 -25080 59916 -25071
rect 60006 -25080 60016 -24890
rect 60076 -24925 60196 -24867
rect 60346 -24650 60426 -24600
rect 60346 -24690 60366 -24650
rect 60406 -24690 60426 -24650
rect 60346 -24740 60426 -24690
rect 60346 -24780 60366 -24740
rect 60406 -24780 60426 -24740
rect 60346 -24820 60426 -24780
rect 60346 -24860 60366 -24820
rect 60406 -24860 60426 -24820
rect 60346 -24870 60426 -24860
rect 60636 -24649 60816 -24591
rect 60636 -24683 60671 -24649
rect 60705 -24683 60747 -24649
rect 60781 -24683 60816 -24649
rect 60636 -24741 60816 -24683
rect 60636 -24775 60671 -24741
rect 60705 -24775 60747 -24741
rect 60781 -24775 60816 -24741
rect 60636 -24833 60816 -24775
rect 60636 -24867 60671 -24833
rect 60705 -24867 60747 -24833
rect 60781 -24867 60816 -24833
rect 60076 -24959 60127 -24925
rect 60161 -24959 60196 -24925
rect 60076 -24990 60196 -24959
rect 60276 -24910 60546 -24900
rect 60276 -24925 60476 -24910
rect 60276 -24959 60297 -24925
rect 60331 -24959 60369 -24925
rect 60405 -24959 60449 -24925
rect 60276 -24970 60476 -24959
rect 60536 -24970 60546 -24910
rect 60276 -24980 60546 -24970
rect 60636 -24925 60816 -24867
rect 61026 -24530 61036 -24420
rect 61126 -24530 61136 -24420
rect 61176 -24480 61196 -24400
rect 61366 -24480 61386 -24400
rect 61176 -24500 61386 -24480
rect 61026 -24560 61136 -24530
rect 61026 -24600 61046 -24560
rect 61086 -24600 61136 -24560
rect 61026 -24650 61136 -24600
rect 61026 -24690 61046 -24650
rect 61086 -24690 61136 -24650
rect 61026 -24740 61136 -24690
rect 61026 -24780 61046 -24740
rect 61086 -24780 61136 -24740
rect 61026 -24820 61136 -24780
rect 61026 -24860 61046 -24820
rect 61086 -24860 61136 -24820
rect 61026 -24880 61136 -24860
rect 61256 -24557 61366 -24500
rect 61256 -24591 61291 -24557
rect 61325 -24591 61366 -24557
rect 61256 -24649 61366 -24591
rect 61256 -24650 61291 -24649
rect 61325 -24650 61366 -24649
rect 61256 -24860 61276 -24650
rect 61356 -24860 61366 -24650
rect 61256 -24867 61291 -24860
rect 61325 -24867 61366 -24860
rect 60636 -24959 60671 -24925
rect 60705 -24959 60747 -24925
rect 60781 -24959 60816 -24925
rect 60636 -25040 60816 -24959
rect 60966 -24924 61177 -24910
rect 60966 -24925 61129 -24924
rect 60966 -24959 60980 -24925
rect 61015 -24959 61053 -24925
rect 61088 -24958 61129 -24925
rect 61164 -24958 61177 -24924
rect 61088 -24959 61177 -24958
rect 60966 -24990 61177 -24959
rect 61256 -24925 61366 -24867
rect 61256 -24959 61291 -24925
rect 61325 -24959 61366 -24925
rect 61256 -24990 61366 -24959
rect 60466 -25050 60546 -25040
rect 59899 -25083 59945 -25080
rect 60466 -25110 60476 -25050
rect 60536 -25110 60546 -25050
rect 59849 -25120 59907 -25115
rect 60466 -25120 60546 -25110
rect 60606 -25050 60826 -25040
rect 60606 -25110 60616 -25050
rect 60736 -25110 60756 -25050
rect 60816 -25110 60826 -25050
rect 60606 -25120 60826 -25110
rect 60886 -25050 60966 -25040
rect 60886 -25110 60896 -25050
rect 60956 -25110 60966 -25050
rect 60886 -25120 60966 -25110
rect 59736 -25121 59926 -25120
rect 59736 -25155 59861 -25121
rect 59895 -25155 59926 -25121
rect 59736 -25180 59926 -25155
rect 60636 -25170 60816 -25120
rect 59376 -25220 59826 -25210
rect 59376 -25260 59476 -25220
rect 59646 -25260 59826 -25220
rect 59376 -25270 59826 -25260
rect 59156 -25290 59236 -25277
rect 58896 -25300 59086 -25290
rect 56380 -25368 57000 -25358
rect 57356 -25364 57676 -25350
rect 56440 -25374 57000 -25368
rect 57314 -25370 57676 -25364
rect 56440 -25394 57178 -25374
rect 56440 -25444 57118 -25394
rect 57168 -25444 57178 -25394
rect 57314 -25410 57326 -25370
rect 57376 -25410 57676 -25370
rect 57314 -25416 57676 -25410
rect 57356 -25430 57676 -25416
rect 56440 -25454 57178 -25444
rect 56440 -25488 57000 -25454
rect 57112 -25456 57174 -25454
rect 56380 -25558 57000 -25488
rect 56032 -25630 56038 -25628
rect 55992 -25642 56038 -25630
rect 55880 -25674 55970 -25668
rect 55870 -25678 55982 -25674
rect 55870 -25720 55880 -25678
rect 55970 -25720 55982 -25678
rect 55880 -25768 55970 -25758
rect 56120 -25798 56300 -25628
rect 57096 -25709 57372 -25678
rect 57096 -25743 57125 -25709
rect 57159 -25743 57217 -25709
rect 57251 -25743 57309 -25709
rect 57343 -25720 57372 -25709
rect 57343 -25743 57376 -25720
rect 57096 -25780 57376 -25743
rect 57066 -25790 57376 -25780
rect 56426 -25798 57376 -25790
rect 56120 -25808 57376 -25798
rect 56014 -25858 56086 -25846
rect 55570 -25978 55830 -25868
rect 53961 -26044 53988 -26006
rect 54022 -26044 54031 -26006
rect 53961 -26058 54031 -26044
rect 54910 -26006 54981 -25994
rect 54910 -26044 54916 -26006
rect 54950 -26044 54981 -26006
rect 54910 -26056 54981 -26044
rect 54911 -26058 54981 -26056
rect 55220 -26018 55330 -26008
rect 54069 -26072 54869 -26066
rect 54069 -26106 54081 -26072
rect 54857 -26078 54869 -26072
rect 54857 -26106 54880 -26078
rect 54069 -26112 54880 -26106
rect 54090 -26188 54880 -26112
rect 55330 -26118 55380 -26018
rect 55330 -26128 55480 -26118
rect 55220 -26138 55480 -26128
rect 55280 -26152 55480 -26138
rect 55280 -26158 55488 -26152
rect 55280 -26178 55300 -26158
rect 54090 -26288 54150 -26188
rect 54840 -26288 54880 -26188
rect 55288 -26192 55300 -26178
rect 55476 -26192 55488 -26158
rect 55530 -26178 55610 -26168
rect 55288 -26198 55488 -26192
rect 55520 -26202 55530 -26190
rect 55520 -26236 55526 -26202
rect 55288 -26246 55488 -26240
rect 55288 -26280 55300 -26246
rect 55476 -26280 55488 -26246
rect 55520 -26248 55530 -26236
rect 55530 -26278 55610 -26268
rect 55288 -26286 55488 -26280
rect 54090 -26308 54140 -26288
rect 26000 -30120 26600 -26400
rect 25860 -30400 26600 -30120
rect 35200 -30120 35800 -26400
rect 54100 -26548 54140 -26308
rect 54850 -26548 54880 -26288
rect 55300 -26328 55470 -26286
rect 55300 -26468 55320 -26328
rect 55470 -26414 55482 -26342
rect 55300 -26478 55470 -26468
rect 54100 -26588 54880 -26548
rect 55710 -26798 55830 -25978
rect 56014 -26008 56020 -25858
rect 56080 -26008 56086 -25858
rect 56014 -26020 56086 -26008
rect 56120 -26008 56170 -25808
rect 56390 -25860 57376 -25808
rect 56390 -25868 57156 -25860
rect 56390 -26008 56654 -25868
rect 56120 -26058 56654 -26008
rect 56306 -26086 56654 -26058
rect 56998 -26020 57156 -25868
rect 57316 -26020 57376 -25860
rect 56998 -26086 57376 -26020
rect 56306 -26500 57376 -26086
rect 57556 -26210 57676 -25430
rect 58896 -25460 58986 -25300
rect 59756 -25320 59826 -25270
rect 59066 -25336 59176 -25330
rect 59066 -25340 59103 -25336
rect 59137 -25340 59176 -25336
rect 59066 -25400 59076 -25340
rect 59166 -25400 59176 -25340
rect 59066 -25410 59176 -25400
rect 58896 -25830 58926 -25460
rect 58966 -25830 58986 -25530
rect 59116 -25460 59506 -25440
rect 59116 -25530 59146 -25460
rect 59226 -25530 59276 -25460
rect 59356 -25530 59396 -25460
rect 59476 -25530 59506 -25460
rect 59116 -25548 59506 -25530
rect 59646 -25460 59716 -25440
rect 59706 -25520 59716 -25460
rect 59646 -25530 59716 -25520
rect 59113 -25554 59513 -25548
rect 59113 -25588 59125 -25554
rect 59501 -25588 59513 -25554
rect 59113 -25594 59513 -25588
rect 59546 -25600 59616 -25590
rect 59246 -25656 59256 -25630
rect 59113 -25662 59256 -25656
rect 59366 -25656 59376 -25630
rect 59366 -25662 59513 -25656
rect 59016 -25700 59076 -25680
rect 59113 -25696 59125 -25662
rect 59501 -25696 59513 -25662
rect 59606 -25660 59616 -25600
rect 59546 -25670 59616 -25660
rect 59113 -25702 59513 -25696
rect 59016 -25790 59076 -25760
rect 59113 -25770 59513 -25764
rect 59113 -25804 59125 -25770
rect 59501 -25804 59513 -25770
rect 59113 -25810 59513 -25804
rect 58896 -25900 58906 -25830
rect 58896 -25920 58986 -25900
rect 59116 -25830 59516 -25810
rect 59116 -25900 59146 -25830
rect 59226 -25900 59276 -25830
rect 59356 -25900 59396 -25830
rect 59476 -25900 59516 -25830
rect 59116 -25920 59516 -25900
rect 59646 -25830 59656 -25530
rect 59706 -25830 59716 -25530
rect 59756 -25500 59766 -25320
rect 59806 -25500 59826 -25320
rect 59956 -25320 60336 -25310
rect 59956 -25334 59966 -25320
rect 59946 -25340 59966 -25334
rect 60326 -25334 60336 -25320
rect 60326 -25340 60346 -25334
rect 59856 -25380 59916 -25370
rect 59946 -25374 59958 -25340
rect 60334 -25374 60346 -25340
rect 61056 -25340 61176 -24990
rect 59946 -25380 59966 -25374
rect 60326 -25380 60346 -25374
rect 60376 -25380 60436 -25360
rect 59956 -25390 60336 -25380
rect 59856 -25460 59916 -25440
rect 59946 -25448 60346 -25442
rect 59756 -25540 59826 -25500
rect 59946 -25482 59958 -25448
rect 60334 -25482 60346 -25448
rect 60376 -25460 60436 -25440
rect 61126 -25440 61176 -25340
rect 61056 -25470 61176 -25440
rect 59946 -25488 60346 -25482
rect 59946 -25540 60336 -25488
rect 59756 -25560 60536 -25540
rect 59756 -25600 59866 -25560
rect 60426 -25600 60536 -25560
rect 59756 -25610 60536 -25600
rect 59796 -25720 59806 -25610
rect 59916 -25720 59926 -25610
rect 59796 -25730 59926 -25720
rect 60436 -25630 60536 -25610
rect 60436 -25750 60446 -25630
rect 60526 -25750 60536 -25630
rect 60436 -25760 60536 -25750
rect 59646 -25840 59716 -25830
rect 59706 -25900 59716 -25840
rect 59646 -25920 59716 -25900
rect 58806 -26210 59356 -26180
rect 59846 -26190 60256 -26180
rect 59846 -26200 59996 -26190
rect 57556 -26220 59356 -26210
rect 57556 -26360 58986 -26220
rect 59126 -26360 59356 -26220
rect 57556 -26410 59356 -26360
rect 58806 -26490 59356 -26410
rect 59600 -26300 59996 -26200
rect 60106 -26200 60256 -26190
rect 60106 -26300 60500 -26200
rect 59600 -26400 60500 -26300
rect 55710 -26800 55910 -26798
rect 59600 -26800 59700 -26400
rect 60400 -26800 60500 -26400
rect 55400 -26900 56200 -26800
rect 59600 -26900 60500 -26800
rect 55400 -27300 55500 -26900
rect 56100 -27300 56200 -26900
rect 55400 -27400 56200 -27300
rect 55380 -27880 55800 -27800
rect 55380 -28160 55460 -27880
rect 55720 -28160 55800 -27880
rect 55380 -28240 55800 -28160
rect 54090 -28338 54890 -28298
rect 54090 -28468 54150 -28338
rect 53510 -28520 53800 -28518
rect 53460 -28540 53800 -28520
rect 53460 -28740 53480 -28540
rect 53780 -28740 53800 -28540
rect 54080 -28598 54150 -28468
rect 54860 -28578 54890 -28338
rect 54850 -28598 54890 -28578
rect 54080 -28666 54880 -28598
rect 54079 -28672 54880 -28666
rect 54079 -28706 54091 -28672
rect 54867 -28698 54880 -28672
rect 54867 -28706 54879 -28698
rect 54079 -28712 54879 -28706
rect 53460 -28760 53800 -28740
rect 53510 -28858 53800 -28760
rect 53002 -29020 53480 -28958
rect 53000 -29158 53480 -29020
rect 53510 -28968 53520 -28858
rect 53640 -28968 53800 -28858
rect 53510 -29088 53800 -28968
rect 53970 -28734 54040 -28718
rect 53970 -28772 53998 -28734
rect 54032 -28772 54040 -28734
rect 53970 -28968 54040 -28772
rect 54920 -28734 54990 -28718
rect 54920 -28772 54926 -28734
rect 54960 -28772 54990 -28734
rect 54079 -28800 54879 -28794
rect 54079 -28834 54091 -28800
rect 54867 -28834 54879 -28800
rect 54079 -28838 54879 -28834
rect 54079 -28840 54750 -28838
rect 54090 -28888 54750 -28840
rect 54740 -28918 54750 -28888
rect 54850 -28840 54879 -28838
rect 54850 -28908 54860 -28840
rect 54840 -28918 54860 -28908
rect 54750 -28928 54860 -28918
rect 54920 -28968 54990 -28772
rect 55430 -28818 55520 -28808
rect 55290 -28928 55390 -28918
rect 53970 -28998 55290 -28968
rect 55430 -28958 55520 -28888
rect 53970 -29008 55390 -28998
rect 54050 -29018 55380 -29008
rect 54050 -29028 54880 -29018
rect 54050 -29038 54091 -29028
rect 54079 -29062 54091 -29038
rect 54867 -29038 54880 -29028
rect 54867 -29062 54879 -29038
rect 54079 -29068 54879 -29062
rect 54920 -29078 54990 -29068
rect 53510 -29106 53630 -29088
rect 53510 -29138 53526 -29106
rect 53514 -29140 53526 -29138
rect 53614 -29138 53630 -29106
rect 53940 -29090 54038 -29078
rect 53940 -29098 53998 -29090
rect 53614 -29140 53626 -29138
rect 53514 -29146 53626 -29140
rect 35200 -30400 35890 -30120
rect 14400 -31800 20000 -31200
rect 24380 -31020 25800 -30980
rect 24380 -33000 25700 -31020
rect 14000 -38000 25700 -33000
rect 14000 -49000 15000 -38000
rect 24000 -49000 25700 -38000
rect 14000 -55000 25700 -49000
rect 24380 -57980 25700 -55000
rect 25780 -57980 25800 -31020
rect 25860 -31146 35890 -30400
rect 53000 -30908 53050 -29158
rect 53250 -29168 53480 -29158
rect 53250 -30518 53330 -29168
rect 53400 -29178 53480 -29168
rect 53400 -29190 53504 -29178
rect 53400 -29966 53464 -29190
rect 53498 -29966 53504 -29190
rect 53400 -29978 53504 -29966
rect 53636 -29188 53682 -29178
rect 53636 -29190 53760 -29188
rect 53636 -29966 53642 -29190
rect 53676 -29966 53760 -29190
rect 53940 -29198 53950 -29098
rect 54032 -29128 54038 -29090
rect 54020 -29140 54038 -29128
rect 54020 -29198 54030 -29140
rect 54079 -29156 54879 -29150
rect 54079 -29190 54091 -29156
rect 54867 -29190 54879 -29156
rect 54920 -29178 54990 -29168
rect 55320 -29168 55380 -29018
rect 54079 -29196 54879 -29190
rect 53940 -29218 54030 -29198
rect 54090 -29228 54870 -29196
rect 55320 -29202 55334 -29168
rect 55368 -29202 55380 -29168
rect 55320 -29208 55380 -29202
rect 53840 -29528 53920 -29518
rect 53840 -29638 53860 -29528
rect 53840 -29648 53920 -29638
rect 53840 -29840 53900 -29648
rect 54320 -29728 54510 -29228
rect 55440 -29238 55520 -28958
rect 55410 -29240 55520 -29238
rect 55284 -29248 55330 -29240
rect 55230 -29252 55330 -29248
rect 55230 -29258 55290 -29252
rect 55324 -29428 55330 -29252
rect 55230 -29438 55330 -29428
rect 55284 -29440 55330 -29438
rect 55372 -29248 55520 -29240
rect 55372 -29252 55430 -29248
rect 55372 -29428 55378 -29252
rect 55412 -29418 55430 -29252
rect 55510 -29418 55520 -29248
rect 55412 -29428 55520 -29418
rect 55372 -29440 55418 -29428
rect 55580 -29528 55720 -28240
rect 58776 -28470 59306 -28350
rect 58776 -28480 58966 -28470
rect 56146 -28580 57366 -28530
rect 55954 -28728 56046 -28716
rect 56146 -28728 56506 -28580
rect 55954 -28898 55960 -28728
rect 56040 -28898 56046 -28728
rect 55954 -28910 56046 -28898
rect 56120 -28758 56506 -28728
rect 56120 -28968 56190 -28758
rect 56390 -28830 56506 -28758
rect 57016 -28734 57366 -28580
rect 57586 -28630 58966 -28480
rect 59126 -28630 59306 -28470
rect 57586 -28650 59306 -28630
rect 59946 -28500 60386 -28400
rect 57586 -28680 58986 -28650
rect 59946 -28660 59956 -28500
rect 60166 -28660 60386 -28500
rect 57016 -28830 57368 -28734
rect 56390 -28870 57368 -28830
rect 56390 -28968 57126 -28870
rect 56120 -28974 57126 -28968
rect 56120 -28978 56750 -28974
rect 55880 -29018 55970 -29008
rect 55870 -29096 55880 -29050
rect 55970 -29096 55982 -29050
rect 55880 -29108 55970 -29098
rect 55000 -29538 55090 -29528
rect 55000 -29648 55090 -29638
rect 54710 -29728 54960 -29708
rect 53940 -29768 54960 -29728
rect 53940 -29772 54730 -29768
rect 53930 -29778 54730 -29772
rect 53930 -29812 53942 -29778
rect 54718 -29812 54730 -29778
rect 53930 -29818 54730 -29812
rect 53840 -29928 53858 -29840
rect 53892 -29928 53900 -29840
rect 53840 -29948 53900 -29928
rect 54762 -29838 54850 -29828
rect 54762 -29840 54770 -29838
rect 54762 -29928 54768 -29840
rect 54840 -29928 54850 -29838
rect 54762 -29940 54850 -29928
rect 54770 -29948 54850 -29940
rect 53636 -29978 53760 -29966
rect 53400 -30196 53480 -29978
rect 53514 -30016 53626 -30010
rect 53514 -30018 53526 -30016
rect 53510 -30050 53526 -30018
rect 53614 -30018 53626 -30016
rect 53614 -30050 53630 -30018
rect 53510 -30124 53630 -30050
rect 53510 -30158 53526 -30124
rect 53614 -30158 53630 -30124
rect 53680 -30038 53760 -29978
rect 53930 -29956 54730 -29950
rect 53930 -29990 53942 -29956
rect 54718 -29990 54730 -29956
rect 53930 -29996 54730 -29990
rect 53940 -30028 54720 -29996
rect 53920 -30038 54720 -30028
rect 53680 -30128 54720 -30038
rect 53514 -30164 53626 -30158
rect 53680 -30196 53760 -30128
rect 53920 -30138 54720 -30128
rect 53940 -30178 54720 -30138
rect 54900 -30168 54960 -29768
rect 55010 -29760 55090 -29648
rect 55540 -29538 55720 -29528
rect 55630 -29638 55720 -29538
rect 55130 -29674 55506 -29668
rect 55130 -29708 55142 -29674
rect 55494 -29708 55506 -29674
rect 55130 -29714 55506 -29708
rect 55010 -29794 55046 -29760
rect 55080 -29794 55090 -29760
rect 55010 -29808 55090 -29794
rect 55142 -29840 55494 -29714
rect 55540 -29760 55720 -29638
rect 55540 -29794 55556 -29760
rect 55590 -29794 55720 -29760
rect 55540 -29808 55720 -29794
rect 55780 -29140 55860 -29128
rect 55130 -29846 55506 -29840
rect 55130 -29880 55142 -29846
rect 55494 -29878 55506 -29846
rect 55494 -29880 55510 -29878
rect 55130 -29886 55510 -29880
rect 55140 -29898 55510 -29886
rect 55780 -29898 55820 -29140
rect 55140 -29916 55820 -29898
rect 55854 -29916 55860 -29140
rect 55140 -29928 55860 -29916
rect 55992 -29140 56038 -29128
rect 55992 -29916 55998 -29140
rect 56032 -29148 56038 -29140
rect 56120 -29148 56300 -28978
rect 57098 -29000 57126 -28974
rect 57356 -29000 57368 -28870
rect 57098 -29014 57368 -29000
rect 57096 -29045 57372 -29014
rect 57096 -29079 57125 -29045
rect 57159 -29079 57217 -29045
rect 57251 -29079 57309 -29045
rect 57343 -29079 57372 -29045
rect 57096 -29110 57372 -29079
rect 56032 -29506 56300 -29148
rect 56590 -29268 56660 -29258
rect 56660 -29334 57000 -29268
rect 57586 -29330 57706 -28680
rect 59946 -28690 60386 -28660
rect 57366 -29334 57706 -29330
rect 56660 -29338 57188 -29334
rect 56660 -29344 57190 -29338
rect 56660 -29394 57118 -29344
rect 57178 -29394 57190 -29344
rect 57314 -29340 57706 -29334
rect 57314 -29380 57326 -29340
rect 57366 -29380 57706 -29340
rect 57314 -29386 57706 -29380
rect 57366 -29390 57706 -29386
rect 58896 -28970 58986 -28950
rect 58896 -29030 58906 -28970
rect 58896 -29320 58926 -29030
rect 58966 -29320 58986 -28970
rect 59106 -28970 59516 -28960
rect 59106 -29030 59216 -28970
rect 59276 -29030 59326 -28970
rect 59386 -29030 59436 -28970
rect 59496 -29030 59516 -28970
rect 59106 -29047 59516 -29030
rect 59626 -28970 59706 -28930
rect 59626 -29030 59636 -28970
rect 59626 -29040 59656 -29030
rect 59106 -29080 59125 -29047
rect 59113 -29081 59125 -29080
rect 59501 -29080 59516 -29047
rect 59501 -29081 59513 -29080
rect 59113 -29087 59513 -29081
rect 59546 -29090 59616 -29080
rect 59276 -29130 59356 -29120
rect 59276 -29149 59286 -29130
rect 59113 -29155 59286 -29149
rect 59346 -29149 59356 -29130
rect 59346 -29155 59513 -29149
rect 59113 -29189 59125 -29155
rect 59501 -29189 59513 -29155
rect 59606 -29150 59616 -29090
rect 59546 -29160 59616 -29150
rect 59113 -29190 59286 -29189
rect 59346 -29190 59513 -29189
rect 59016 -29200 59076 -29190
rect 59113 -29195 59513 -29190
rect 59276 -29200 59356 -29195
rect 59546 -29210 59616 -29200
rect 59016 -29270 59076 -29260
rect 59113 -29263 59513 -29257
rect 59113 -29297 59125 -29263
rect 59501 -29297 59513 -29263
rect 59606 -29270 59616 -29210
rect 59546 -29280 59616 -29270
rect 59113 -29300 59513 -29297
rect 59113 -29303 59516 -29300
rect 58896 -29330 58986 -29320
rect 58896 -29390 58906 -29330
rect 58966 -29390 58986 -29330
rect 58896 -29392 58986 -29390
rect 59116 -29320 59516 -29303
rect 59646 -29310 59656 -29040
rect 59116 -29380 59216 -29320
rect 59276 -29380 59336 -29320
rect 59396 -29380 59436 -29320
rect 59496 -29380 59516 -29320
rect 56660 -29398 57190 -29394
rect 56590 -29400 57190 -29398
rect 56590 -29404 57188 -29400
rect 56590 -29468 57000 -29404
rect 56032 -29518 56356 -29506
rect 56032 -29916 56280 -29518
rect 55992 -29928 56280 -29916
rect 55140 -29938 55200 -29928
rect 55450 -29958 55810 -29928
rect 55870 -29966 55982 -29960
rect 55870 -30000 55882 -29966
rect 55970 -30000 55982 -29966
rect 55870 -30006 55982 -30000
rect 55140 -30018 55200 -30008
rect 55024 -30048 55116 -30036
rect 55024 -30128 55030 -30048
rect 55110 -30128 55116 -30048
rect 55024 -30140 55116 -30128
rect 55734 -30048 55816 -30036
rect 55734 -30128 55740 -30048
rect 55810 -30128 55816 -30048
rect 55734 -30140 55816 -30128
rect 55880 -30038 55970 -30006
rect 55880 -30164 55970 -30128
rect 56060 -30148 56280 -29928
rect 56350 -30148 56356 -29518
rect 56480 -29588 56550 -29578
rect 56480 -29658 56550 -29648
rect 56590 -29687 56750 -29468
rect 58894 -29486 58988 -29392
rect 59116 -29400 59516 -29380
rect 59636 -29320 59656 -29310
rect 59696 -29320 59706 -28970
rect 59856 -29140 59976 -29130
rect 59856 -29230 59866 -29140
rect 59966 -29230 59976 -29140
rect 59856 -29240 59976 -29230
rect 60436 -29220 60446 -29120
rect 60526 -29220 60536 -29120
rect 60436 -29240 60536 -29220
rect 59636 -29330 59706 -29320
rect 59696 -29390 59706 -29330
rect 59636 -29410 59706 -29390
rect 59756 -29260 60536 -29240
rect 59756 -29300 59866 -29260
rect 60426 -29300 60536 -29260
rect 59756 -29310 60536 -29300
rect 59756 -29350 59826 -29310
rect 59066 -29440 59176 -29430
rect 58896 -29550 58986 -29486
rect 59066 -29510 59076 -29440
rect 59166 -29510 59176 -29440
rect 59066 -29512 59103 -29510
rect 59137 -29512 59176 -29510
rect 59066 -29520 59176 -29512
rect 59756 -29540 59766 -29350
rect 59806 -29540 59826 -29350
rect 59956 -29368 60046 -29340
rect 59946 -29374 60046 -29368
rect 60126 -29368 60336 -29340
rect 60126 -29374 60346 -29368
rect 59856 -29410 59916 -29400
rect 59946 -29408 59958 -29374
rect 60334 -29408 60346 -29374
rect 59946 -29414 60346 -29408
rect 60376 -29420 60446 -29410
rect 59856 -29490 59916 -29480
rect 59946 -29482 60346 -29476
rect 59946 -29516 59958 -29482
rect 60334 -29516 60346 -29482
rect 60376 -29490 60446 -29480
rect 59946 -29522 59976 -29516
rect 57098 -29558 57368 -29554
rect 57096 -29564 57372 -29558
rect 57096 -29650 57098 -29564
rect 56424 -29688 56470 -29687
rect 56060 -30160 56356 -30148
rect 56410 -29699 56470 -29688
rect 53400 -30208 53504 -30196
rect 53400 -30518 53464 -30208
rect 53250 -30908 53464 -30518
rect 53000 -30984 53464 -30908
rect 53498 -30984 53504 -30208
rect 53000 -30988 53504 -30984
rect 53458 -30996 53504 -30988
rect 53636 -30208 53760 -30196
rect 53636 -30984 53642 -30208
rect 53676 -30984 53760 -30208
rect 53930 -30184 54730 -30178
rect 53930 -30218 53942 -30184
rect 54718 -30218 54730 -30184
rect 53930 -30224 54730 -30218
rect 53830 -30246 53900 -30228
rect 53830 -30334 53858 -30246
rect 53892 -30334 53900 -30246
rect 53830 -30528 53900 -30334
rect 54760 -30246 54850 -30228
rect 54760 -30334 54768 -30246
rect 54802 -30248 54850 -30246
rect 54900 -30238 55200 -30168
rect 55870 -30170 55982 -30164
rect 55870 -30204 55882 -30170
rect 55970 -30204 55982 -30170
rect 55450 -30238 55810 -30208
rect 55870 -30210 55982 -30204
rect 56060 -30238 56300 -30160
rect 54900 -30242 55820 -30238
rect 56000 -30242 56300 -30238
rect 54900 -30248 55860 -30242
rect 54840 -30328 54850 -30248
rect 54802 -30334 54850 -30328
rect 54760 -30348 54850 -30334
rect 55130 -30254 55860 -30248
rect 55130 -30278 55820 -30254
rect 55130 -30296 55510 -30278
rect 55130 -30330 55142 -30296
rect 55494 -30298 55510 -30296
rect 55494 -30330 55506 -30298
rect 55130 -30336 55506 -30330
rect 53930 -30362 54730 -30356
rect 53930 -30396 53942 -30362
rect 54718 -30396 54730 -30362
rect 55020 -30382 55090 -30368
rect 53930 -30402 54730 -30396
rect 53940 -30408 54730 -30402
rect 54920 -30398 54980 -30388
rect 53940 -30448 54920 -30408
rect 53830 -30538 53920 -30528
rect 53830 -30648 53850 -30538
rect 53830 -30658 53920 -30648
rect 54320 -30948 54510 -30448
rect 54710 -30468 54920 -30448
rect 54910 -30478 54980 -30468
rect 55020 -30416 55046 -30382
rect 55080 -30416 55090 -30382
rect 55020 -30528 55090 -30416
rect 55142 -30462 55494 -30336
rect 55540 -30382 55620 -30368
rect 55540 -30416 55556 -30382
rect 55590 -30416 55620 -30382
rect 55130 -30468 55506 -30462
rect 55130 -30502 55142 -30468
rect 55494 -30502 55506 -30468
rect 55130 -30508 55506 -30502
rect 55000 -30538 55090 -30528
rect 55000 -30648 55090 -30638
rect 55540 -30528 55620 -30416
rect 55540 -30538 55630 -30528
rect 55630 -30638 55680 -30548
rect 55540 -30648 55680 -30638
rect 55274 -30738 55320 -30736
rect 55220 -30748 55320 -30738
rect 55220 -30924 55280 -30918
rect 55314 -30924 55320 -30748
rect 55220 -30928 55320 -30924
rect 55274 -30936 55320 -30928
rect 55362 -30748 55408 -30736
rect 55362 -30924 55368 -30748
rect 55402 -30758 55510 -30748
rect 55402 -30924 55410 -30758
rect 55362 -30928 55410 -30924
rect 55500 -30928 55510 -30758
rect 55362 -30936 55510 -30928
rect 55390 -30938 55510 -30936
rect 53636 -30988 53760 -30984
rect 53636 -30996 53682 -30988
rect 53940 -31008 54020 -30968
rect 54080 -30982 54860 -30948
rect 55311 -30974 55371 -30968
rect 53514 -31034 53626 -31028
rect 53514 -31038 53526 -31034
rect 25860 -31543 25884 -31146
rect 26998 -31543 27126 -31146
rect 28240 -31543 28368 -31146
rect 29482 -31543 29610 -31146
rect 30724 -31543 30852 -31146
rect 31966 -31543 32094 -31146
rect 33208 -31543 33336 -31146
rect 34450 -31543 34578 -31146
rect 35692 -31543 35890 -31146
rect 53510 -31068 53526 -31038
rect 53614 -31038 53626 -31034
rect 53614 -31068 53630 -31038
rect 53510 -31128 53630 -31068
rect 53940 -31088 53950 -31008
rect 54010 -31038 54020 -31008
rect 54069 -30988 54869 -30982
rect 54069 -31022 54081 -30988
rect 54857 -31022 54869 -30988
rect 54069 -31028 54869 -31022
rect 54910 -30998 54980 -30988
rect 54010 -31050 54028 -31038
rect 54022 -31088 54028 -31050
rect 53940 -31100 54028 -31088
rect 53940 -31108 54020 -31100
rect 54910 -31108 54980 -31098
rect 55311 -31008 55324 -30974
rect 55358 -31008 55371 -30974
rect 54070 -31110 54870 -31108
rect 54069 -31116 54870 -31110
rect 54069 -31138 54081 -31116
rect 54041 -31150 54081 -31138
rect 54857 -31118 54870 -31116
rect 54857 -31150 54880 -31118
rect 55311 -31148 55371 -31008
rect 54041 -31158 54880 -31150
rect 55240 -31158 55371 -31148
rect 54041 -31168 55240 -31158
rect 53510 -31258 53630 -31248
rect 53961 -31208 55240 -31168
rect 53961 -31406 54031 -31208
rect 54730 -31268 54860 -31258
rect 54730 -31288 54740 -31268
rect 54080 -31338 54740 -31288
rect 54069 -31344 54740 -31338
rect 54850 -31338 54860 -31268
rect 54850 -31344 54869 -31338
rect 54069 -31378 54081 -31344
rect 54857 -31378 54869 -31344
rect 54069 -31384 54869 -31378
rect 54911 -31394 54981 -31208
rect 55370 -31208 55371 -31158
rect 55240 -31228 55370 -31218
rect 55410 -31248 55510 -30938
rect 55410 -31358 55510 -31338
rect 55570 -31268 55680 -30648
rect 55780 -31030 55820 -30278
rect 55854 -31030 55860 -30254
rect 55780 -31038 55860 -31030
rect 55814 -31042 55860 -31038
rect 55992 -30254 56300 -30242
rect 55992 -31030 55998 -30254
rect 56032 -31028 56300 -30254
rect 56410 -30298 56430 -29699
rect 56380 -30475 56430 -30298
rect 56464 -30475 56470 -29699
rect 56380 -30487 56470 -30475
rect 56552 -29699 56750 -29687
rect 56552 -30475 56558 -29699
rect 56592 -29838 56750 -29699
rect 57066 -29680 57098 -29650
rect 57368 -29650 57372 -29564
rect 58896 -29559 59076 -29550
rect 58896 -29560 59084 -29559
rect 59156 -29560 59202 -29559
rect 57368 -29680 57396 -29650
rect 57066 -29810 57086 -29680
rect 57376 -29810 57396 -29680
rect 56592 -30475 56610 -29838
rect 57066 -29840 57396 -29810
rect 56860 -29990 57060 -29978
rect 56860 -30018 57236 -29990
rect 56860 -30148 56900 -30018
rect 57020 -30148 57236 -30018
rect 56860 -30188 57236 -30148
rect 57036 -30190 57236 -30188
rect 58556 -30080 58756 -30060
rect 58556 -30240 58576 -30080
rect 58736 -30240 58756 -30080
rect 58556 -30260 58756 -30240
rect 56552 -30478 56610 -30475
rect 57036 -30340 57446 -30330
rect 56552 -30487 56598 -30478
rect 57036 -30480 57056 -30340
rect 57416 -30480 57446 -30340
rect 56380 -30758 56440 -30487
rect 57036 -30500 57098 -30480
rect 56480 -30528 56550 -30518
rect 56480 -30598 56550 -30588
rect 57096 -30614 57098 -30534
rect 57368 -30500 57446 -30480
rect 57368 -30614 57372 -30534
rect 57096 -30630 57372 -30614
rect 58896 -30690 58926 -29560
rect 58966 -29571 59086 -29560
rect 58966 -29947 59044 -29571
rect 59078 -29947 59086 -29571
rect 58966 -29970 59086 -29947
rect 59156 -29571 59256 -29560
rect 59756 -29570 59826 -29540
rect 59966 -29552 59976 -29522
rect 60316 -29522 60346 -29516
rect 61036 -29520 61466 -29510
rect 60316 -29552 60326 -29522
rect 59966 -29560 60326 -29552
rect 59156 -29947 59162 -29571
rect 59196 -29640 59256 -29571
rect 59236 -29720 59256 -29640
rect 59196 -29840 59256 -29720
rect 59236 -29920 59256 -29840
rect 59196 -29947 59256 -29920
rect 59156 -29960 59256 -29947
rect 58966 -30280 59036 -29970
rect 59066 -30006 59176 -30000
rect 59066 -30010 59103 -30006
rect 59137 -30010 59176 -30006
rect 59066 -30080 59076 -30010
rect 59166 -30080 59176 -30010
rect 59066 -30090 59176 -30080
rect 59206 -30160 59256 -29960
rect 59376 -29590 59826 -29570
rect 59376 -29630 59476 -29590
rect 59656 -29630 59826 -29590
rect 59376 -29640 59826 -29630
rect 59376 -29690 59436 -29640
rect 59376 -30050 59386 -29690
rect 59426 -30050 59436 -29690
rect 59526 -29698 59576 -29670
rect 59526 -29732 59546 -29698
rect 59636 -29730 59706 -29670
rect 59580 -29732 59706 -29730
rect 59526 -29740 59706 -29732
rect 59476 -29782 59546 -29770
rect 59476 -29850 59502 -29782
rect 59476 -29958 59502 -29920
rect 59536 -29958 59546 -29782
rect 59476 -29970 59546 -29958
rect 59576 -29782 59636 -29770
rect 59576 -29790 59590 -29782
rect 59624 -29790 59636 -29782
rect 59576 -29970 59636 -29960
rect 59534 -30008 59592 -30002
rect 59534 -30010 59546 -30008
rect 59066 -30170 59176 -30160
rect 59066 -30240 59076 -30170
rect 59166 -30240 59176 -30170
rect 59066 -30242 59103 -30240
rect 59137 -30242 59176 -30240
rect 59066 -30250 59176 -30242
rect 59206 -30170 59266 -30160
rect 59206 -30250 59266 -30240
rect 59376 -30200 59436 -30050
rect 59516 -30042 59546 -30010
rect 59580 -30010 59592 -30008
rect 59666 -30010 59706 -29740
rect 59580 -30042 59706 -30010
rect 59516 -30080 59706 -30042
rect 59746 -29698 59936 -29670
rect 59746 -29732 59862 -29698
rect 59896 -29732 59936 -29698
rect 59746 -29740 59936 -29732
rect 61036 -29700 61206 -29520
rect 61346 -29700 61466 -29520
rect 61036 -29740 61466 -29700
rect 59746 -30000 59776 -29740
rect 60286 -29750 60476 -29740
rect 59806 -29782 59866 -29770
rect 59806 -29800 59818 -29782
rect 59852 -29800 59866 -29782
rect 59806 -29958 59818 -29940
rect 59852 -29958 59866 -29940
rect 59806 -29970 59866 -29958
rect 59900 -29780 60016 -29770
rect 59900 -29782 59916 -29780
rect 59900 -29958 59906 -29782
rect 59900 -29960 59916 -29958
rect 60006 -29960 60016 -29780
rect 60286 -29890 60306 -29750
rect 60456 -29890 60476 -29750
rect 61176 -29800 61386 -29780
rect 60286 -29900 60476 -29890
rect 61026 -29820 61136 -29810
rect 59900 -29970 60016 -29960
rect 60076 -29957 60196 -29920
rect 60076 -29991 60127 -29957
rect 60161 -29991 60196 -29957
rect 59746 -30008 59926 -30000
rect 59746 -30010 59862 -30008
rect 59896 -30010 59926 -30008
rect 59746 -30080 59826 -30010
rect 59916 -30080 59926 -30010
rect 59746 -30090 59926 -30080
rect 60076 -30049 60196 -29991
rect 60336 -29960 60446 -29900
rect 60336 -30000 60366 -29960
rect 60406 -30000 60446 -29960
rect 60636 -29957 60816 -29920
rect 60636 -29991 60671 -29957
rect 60705 -29991 60747 -29957
rect 60781 -29991 60816 -29957
rect 60076 -30080 60127 -30049
rect 60161 -30080 60196 -30049
rect 59736 -30170 59936 -30160
rect 58966 -30301 59086 -30280
rect 58966 -30677 59044 -30301
rect 59078 -30677 59086 -30301
rect 58966 -30690 59086 -30677
rect 59156 -30290 59202 -30289
rect 59156 -30301 59236 -30290
rect 59156 -30677 59162 -30301
rect 59196 -30330 59236 -30301
rect 59226 -30410 59236 -30330
rect 59196 -30560 59236 -30410
rect 59226 -30640 59236 -30560
rect 59196 -30677 59236 -30640
rect 59376 -30570 59386 -30200
rect 59426 -30570 59436 -30200
rect 59516 -30211 59706 -30170
rect 59516 -30245 59545 -30211
rect 59579 -30245 59706 -30211
rect 59516 -30250 59706 -30245
rect 59533 -30251 59591 -30250
rect 59466 -30295 59546 -30280
rect 59586 -30283 59646 -30280
rect 59466 -30330 59501 -30295
rect 59466 -30471 59501 -30410
rect 59535 -30471 59546 -30295
rect 59466 -30480 59546 -30471
rect 59583 -30295 59646 -30283
rect 59583 -30310 59589 -30295
rect 59623 -30310 59646 -30295
rect 59583 -30450 59586 -30310
rect 59583 -30471 59589 -30450
rect 59623 -30471 59646 -30450
rect 59583 -30480 59646 -30471
rect 59495 -30483 59541 -30480
rect 59583 -30483 59629 -30480
rect 59533 -30520 59591 -30515
rect 59676 -30520 59706 -30250
rect 59376 -30610 59436 -30570
rect 59506 -30580 59516 -30520
rect 59596 -30580 59706 -30520
rect 59736 -30240 59826 -30170
rect 59926 -30240 59936 -30170
rect 59736 -30245 59861 -30240
rect 59895 -30245 59936 -30240
rect 59736 -30250 59936 -30245
rect 60076 -30240 60096 -30080
rect 60176 -30240 60196 -30080
rect 59736 -30520 59766 -30250
rect 59849 -30251 59907 -30250
rect 60076 -30267 60127 -30240
rect 60161 -30267 60196 -30240
rect 59796 -30283 59856 -30280
rect 59796 -30290 59857 -30283
rect 59856 -30470 59857 -30290
rect 59796 -30471 59817 -30470
rect 59851 -30471 59857 -30470
rect 59796 -30480 59857 -30471
rect 59811 -30483 59857 -30480
rect 59899 -30290 59945 -30283
rect 59899 -30295 59916 -30290
rect 59899 -30471 59905 -30295
rect 59899 -30480 59916 -30471
rect 60006 -30480 60016 -30290
rect 60076 -30325 60196 -30267
rect 60346 -30050 60426 -30000
rect 60346 -30090 60366 -30050
rect 60406 -30090 60426 -30050
rect 60346 -30140 60426 -30090
rect 60346 -30180 60366 -30140
rect 60406 -30180 60426 -30140
rect 60346 -30220 60426 -30180
rect 60346 -30260 60366 -30220
rect 60406 -30260 60426 -30220
rect 60346 -30270 60426 -30260
rect 60636 -30049 60816 -29991
rect 60636 -30083 60671 -30049
rect 60705 -30083 60747 -30049
rect 60781 -30083 60816 -30049
rect 60636 -30141 60816 -30083
rect 60636 -30175 60671 -30141
rect 60705 -30175 60747 -30141
rect 60781 -30175 60816 -30141
rect 60636 -30233 60816 -30175
rect 60636 -30267 60671 -30233
rect 60705 -30267 60747 -30233
rect 60781 -30267 60816 -30233
rect 60076 -30359 60127 -30325
rect 60161 -30359 60196 -30325
rect 60076 -30390 60196 -30359
rect 60276 -30310 60546 -30300
rect 60276 -30325 60476 -30310
rect 60276 -30359 60297 -30325
rect 60331 -30359 60369 -30325
rect 60405 -30359 60449 -30325
rect 60276 -30370 60476 -30359
rect 60536 -30370 60546 -30310
rect 60276 -30380 60546 -30370
rect 60636 -30325 60816 -30267
rect 61026 -29930 61036 -29820
rect 61126 -29930 61136 -29820
rect 61176 -29880 61196 -29800
rect 61366 -29880 61386 -29800
rect 61176 -29900 61386 -29880
rect 61026 -29960 61136 -29930
rect 61026 -30000 61046 -29960
rect 61086 -30000 61136 -29960
rect 61026 -30050 61136 -30000
rect 61026 -30090 61046 -30050
rect 61086 -30090 61136 -30050
rect 61026 -30140 61136 -30090
rect 61026 -30180 61046 -30140
rect 61086 -30180 61136 -30140
rect 61026 -30220 61136 -30180
rect 61026 -30260 61046 -30220
rect 61086 -30260 61136 -30220
rect 61026 -30280 61136 -30260
rect 61256 -29957 61366 -29900
rect 61256 -29991 61291 -29957
rect 61325 -29991 61366 -29957
rect 61256 -30049 61366 -29991
rect 61256 -30050 61291 -30049
rect 61325 -30050 61366 -30049
rect 61256 -30260 61276 -30050
rect 61356 -30260 61366 -30050
rect 61256 -30267 61291 -30260
rect 61325 -30267 61366 -30260
rect 60636 -30359 60671 -30325
rect 60705 -30359 60747 -30325
rect 60781 -30359 60816 -30325
rect 60636 -30440 60816 -30359
rect 60966 -30324 61177 -30310
rect 60966 -30325 61129 -30324
rect 60966 -30359 60980 -30325
rect 61015 -30359 61053 -30325
rect 61088 -30358 61129 -30325
rect 61164 -30358 61177 -30324
rect 61088 -30359 61177 -30358
rect 60966 -30390 61177 -30359
rect 61256 -30325 61366 -30267
rect 61256 -30359 61291 -30325
rect 61325 -30359 61366 -30325
rect 61256 -30390 61366 -30359
rect 60466 -30450 60546 -30440
rect 59899 -30483 59945 -30480
rect 60466 -30510 60476 -30450
rect 60536 -30510 60546 -30450
rect 59849 -30520 59907 -30515
rect 60466 -30520 60546 -30510
rect 60606 -30450 60826 -30440
rect 60606 -30510 60616 -30450
rect 60736 -30510 60756 -30450
rect 60816 -30510 60826 -30450
rect 60606 -30520 60826 -30510
rect 60886 -30450 60966 -30440
rect 60886 -30510 60896 -30450
rect 60956 -30510 60966 -30450
rect 60886 -30520 60966 -30510
rect 59736 -30521 59926 -30520
rect 59736 -30555 59861 -30521
rect 59895 -30555 59926 -30521
rect 59736 -30580 59926 -30555
rect 60636 -30570 60816 -30520
rect 59376 -30620 59826 -30610
rect 59376 -30660 59476 -30620
rect 59646 -30660 59826 -30620
rect 59376 -30670 59826 -30660
rect 59156 -30690 59236 -30677
rect 58896 -30700 59086 -30690
rect 56380 -30768 57000 -30758
rect 57356 -30764 57676 -30750
rect 56440 -30774 57000 -30768
rect 57314 -30770 57676 -30764
rect 56440 -30794 57178 -30774
rect 56440 -30844 57118 -30794
rect 57168 -30844 57178 -30794
rect 57314 -30810 57326 -30770
rect 57376 -30810 57676 -30770
rect 57314 -30816 57676 -30810
rect 57356 -30830 57676 -30816
rect 56440 -30854 57178 -30844
rect 56440 -30888 57000 -30854
rect 57112 -30856 57174 -30854
rect 56380 -30958 57000 -30888
rect 56032 -31030 56038 -31028
rect 55992 -31042 56038 -31030
rect 55880 -31074 55970 -31068
rect 55870 -31078 55982 -31074
rect 55870 -31120 55880 -31078
rect 55970 -31120 55982 -31078
rect 55880 -31168 55970 -31158
rect 56120 -31198 56300 -31028
rect 57096 -31109 57372 -31078
rect 57096 -31143 57125 -31109
rect 57159 -31143 57217 -31109
rect 57251 -31143 57309 -31109
rect 57343 -31120 57372 -31109
rect 57343 -31143 57376 -31120
rect 57096 -31180 57376 -31143
rect 57066 -31190 57376 -31180
rect 56426 -31198 57376 -31190
rect 56120 -31208 57376 -31198
rect 56014 -31258 56086 -31246
rect 55570 -31378 55830 -31268
rect 53961 -31444 53988 -31406
rect 54022 -31444 54031 -31406
rect 53961 -31458 54031 -31444
rect 54910 -31406 54981 -31394
rect 54910 -31444 54916 -31406
rect 54950 -31444 54981 -31406
rect 54910 -31456 54981 -31444
rect 54911 -31458 54981 -31456
rect 55220 -31418 55330 -31408
rect 54069 -31472 54869 -31466
rect 54069 -31506 54081 -31472
rect 54857 -31478 54869 -31472
rect 54857 -31506 54880 -31478
rect 54069 -31512 54880 -31506
rect 25860 -31560 35890 -31543
rect 54090 -31588 54880 -31512
rect 55330 -31518 55380 -31418
rect 55330 -31528 55480 -31518
rect 55220 -31538 55480 -31528
rect 55280 -31552 55480 -31538
rect 55280 -31558 55488 -31552
rect 55280 -31578 55300 -31558
rect 54090 -31688 54150 -31588
rect 54840 -31688 54880 -31588
rect 55288 -31592 55300 -31578
rect 55476 -31592 55488 -31558
rect 55530 -31578 55610 -31568
rect 55288 -31598 55488 -31592
rect 55520 -31602 55530 -31590
rect 55520 -31636 55526 -31602
rect 55288 -31646 55488 -31640
rect 55288 -31680 55300 -31646
rect 55476 -31680 55488 -31646
rect 55520 -31648 55530 -31636
rect 55530 -31678 55610 -31668
rect 55288 -31686 55488 -31680
rect 54090 -31708 54140 -31688
rect 54100 -31948 54140 -31708
rect 54850 -31948 54880 -31688
rect 55300 -31728 55470 -31686
rect 55300 -31868 55320 -31728
rect 55470 -31814 55482 -31742
rect 55300 -31878 55470 -31868
rect 54100 -31988 54880 -31948
rect 36000 -32062 37000 -32000
rect 25862 -32081 37000 -32062
rect 25862 -32478 25884 -32081
rect 26998 -32478 27126 -32081
rect 28240 -32478 28368 -32081
rect 29482 -32478 29610 -32081
rect 30724 -32478 30852 -32081
rect 31966 -32478 32094 -32081
rect 33208 -32478 33336 -32081
rect 34450 -32478 34578 -32081
rect 35692 -32200 37000 -32081
rect 55710 -32198 55830 -31378
rect 56014 -31408 56020 -31258
rect 56080 -31408 56086 -31258
rect 56014 -31420 56086 -31408
rect 56120 -31408 56170 -31208
rect 56390 -31260 57376 -31208
rect 56390 -31268 57156 -31260
rect 56390 -31408 56654 -31268
rect 56120 -31458 56654 -31408
rect 56306 -31486 56654 -31458
rect 56998 -31420 57156 -31268
rect 57316 -31420 57376 -31260
rect 56998 -31486 57376 -31420
rect 56306 -31900 57376 -31486
rect 57556 -31610 57676 -30830
rect 58896 -30860 58986 -30700
rect 59756 -30720 59826 -30670
rect 59066 -30736 59176 -30730
rect 59066 -30740 59103 -30736
rect 59137 -30740 59176 -30736
rect 59066 -30800 59076 -30740
rect 59166 -30800 59176 -30740
rect 59066 -30810 59176 -30800
rect 58896 -31230 58926 -30860
rect 58966 -31230 58986 -30930
rect 59116 -30860 59506 -30840
rect 59116 -30930 59146 -30860
rect 59226 -30930 59276 -30860
rect 59356 -30930 59396 -30860
rect 59476 -30930 59506 -30860
rect 59116 -30948 59506 -30930
rect 59646 -30860 59716 -30840
rect 59706 -30920 59716 -30860
rect 59646 -30930 59716 -30920
rect 59113 -30954 59513 -30948
rect 59113 -30988 59125 -30954
rect 59501 -30988 59513 -30954
rect 59113 -30994 59513 -30988
rect 59546 -31000 59616 -30990
rect 59246 -31056 59256 -31030
rect 59113 -31062 59256 -31056
rect 59366 -31056 59376 -31030
rect 59366 -31062 59513 -31056
rect 59016 -31100 59076 -31080
rect 59113 -31096 59125 -31062
rect 59501 -31096 59513 -31062
rect 59606 -31060 59616 -31000
rect 59546 -31070 59616 -31060
rect 59113 -31102 59513 -31096
rect 59016 -31190 59076 -31160
rect 59113 -31170 59513 -31164
rect 59113 -31204 59125 -31170
rect 59501 -31204 59513 -31170
rect 59113 -31210 59513 -31204
rect 58896 -31300 58906 -31230
rect 58896 -31320 58986 -31300
rect 59116 -31230 59516 -31210
rect 59116 -31300 59146 -31230
rect 59226 -31300 59276 -31230
rect 59356 -31300 59396 -31230
rect 59476 -31300 59516 -31230
rect 59116 -31320 59516 -31300
rect 59646 -31230 59656 -30930
rect 59706 -31230 59716 -30930
rect 59756 -30900 59766 -30720
rect 59806 -30900 59826 -30720
rect 59956 -30720 60336 -30710
rect 59956 -30734 59966 -30720
rect 59946 -30740 59966 -30734
rect 60326 -30734 60336 -30720
rect 60326 -30740 60346 -30734
rect 59856 -30780 59916 -30770
rect 59946 -30774 59958 -30740
rect 60334 -30774 60346 -30740
rect 61056 -30740 61176 -30390
rect 59946 -30780 59966 -30774
rect 60326 -30780 60346 -30774
rect 60376 -30780 60436 -30760
rect 59956 -30790 60336 -30780
rect 59856 -30860 59916 -30840
rect 59946 -30848 60346 -30842
rect 59756 -30940 59826 -30900
rect 59946 -30882 59958 -30848
rect 60334 -30882 60346 -30848
rect 60376 -30860 60436 -30840
rect 61126 -30840 61176 -30740
rect 61056 -30870 61176 -30840
rect 59946 -30888 60346 -30882
rect 59946 -30940 60336 -30888
rect 59756 -30960 60536 -30940
rect 59756 -31000 59866 -30960
rect 60426 -31000 60536 -30960
rect 59756 -31010 60536 -31000
rect 59796 -31120 59806 -31010
rect 59916 -31120 59926 -31010
rect 59796 -31130 59926 -31120
rect 60436 -31030 60536 -31010
rect 60436 -31150 60446 -31030
rect 60526 -31150 60536 -31030
rect 60436 -31160 60536 -31150
rect 59646 -31240 59716 -31230
rect 59706 -31300 59716 -31240
rect 59646 -31320 59716 -31300
rect 58806 -31610 59356 -31580
rect 59846 -31590 60256 -31580
rect 59846 -31600 59996 -31590
rect 57556 -31620 59356 -31610
rect 57556 -31760 58986 -31620
rect 59126 -31760 59356 -31620
rect 57556 -31810 59356 -31760
rect 58806 -31890 59356 -31810
rect 59700 -31700 59996 -31600
rect 60106 -31600 60256 -31590
rect 60106 -31700 60400 -31600
rect 59700 -31800 60400 -31700
rect 59700 -32100 59800 -31800
rect 60300 -32100 60400 -31800
rect 55710 -32200 55910 -32198
rect 59700 -32200 60400 -32100
rect 35692 -32478 36200 -32200
rect 25862 -32744 36200 -32478
rect 25862 -33141 25882 -32744
rect 26996 -33141 27124 -32744
rect 28238 -33141 28366 -32744
rect 29480 -33141 29608 -32744
rect 30722 -33141 30850 -32744
rect 31964 -33141 32092 -32744
rect 33206 -33141 33334 -32744
rect 34448 -33141 34576 -32744
rect 35690 -33000 36200 -32744
rect 36800 -33000 37000 -32200
rect 55400 -32300 56200 -32200
rect 55400 -32700 55500 -32300
rect 56100 -32700 56200 -32300
rect 55400 -32800 56200 -32700
rect 35690 -33141 37000 -33000
rect 25862 -33162 37000 -33141
rect 36000 -33200 37000 -33162
rect 55380 -33280 55800 -33200
rect 55380 -33560 55460 -33280
rect 55720 -33560 55800 -33280
rect 35900 -33660 38200 -33600
rect 55380 -33640 55800 -33560
rect 25860 -33679 38200 -33660
rect 25860 -34076 25882 -33679
rect 26996 -34076 27124 -33679
rect 28238 -34076 28366 -33679
rect 29480 -34076 29608 -33679
rect 30722 -34076 30850 -33679
rect 31964 -34076 32092 -33679
rect 33206 -34076 33334 -33679
rect 34448 -34076 34576 -33679
rect 35690 -33700 38200 -33679
rect 35690 -34076 36000 -33700
rect 25860 -34342 36000 -34076
rect 25860 -34739 25882 -34342
rect 26996 -34739 27124 -34342
rect 28238 -34739 28366 -34342
rect 29480 -34739 29608 -34342
rect 30722 -34739 30850 -34342
rect 31964 -34739 32092 -34342
rect 33206 -34739 33334 -34342
rect 34448 -34739 34576 -34342
rect 35690 -34700 36000 -34342
rect 38100 -34700 38200 -33700
rect 54090 -33738 54890 -33698
rect 54090 -33868 54150 -33738
rect 53510 -33920 53800 -33918
rect 53460 -33940 53800 -33920
rect 53460 -34140 53480 -33940
rect 53780 -34140 53800 -33940
rect 54080 -33998 54150 -33868
rect 54860 -33978 54890 -33738
rect 54850 -33998 54890 -33978
rect 54080 -34066 54880 -33998
rect 54079 -34072 54880 -34066
rect 54079 -34106 54091 -34072
rect 54867 -34098 54880 -34072
rect 54867 -34106 54879 -34098
rect 54079 -34112 54879 -34106
rect 53460 -34160 53800 -34140
rect 53510 -34258 53800 -34160
rect 53002 -34420 53480 -34358
rect 35690 -34739 38200 -34700
rect 25860 -34760 38200 -34739
rect 35900 -34800 38200 -34760
rect 53000 -34558 53480 -34420
rect 53510 -34368 53520 -34258
rect 53640 -34368 53800 -34258
rect 53510 -34488 53800 -34368
rect 53970 -34134 54040 -34118
rect 53970 -34172 53998 -34134
rect 54032 -34172 54040 -34134
rect 53970 -34368 54040 -34172
rect 54920 -34134 54990 -34118
rect 54920 -34172 54926 -34134
rect 54960 -34172 54990 -34134
rect 54079 -34200 54879 -34194
rect 54079 -34234 54091 -34200
rect 54867 -34234 54879 -34200
rect 54079 -34238 54879 -34234
rect 54079 -34240 54750 -34238
rect 54090 -34288 54750 -34240
rect 54740 -34318 54750 -34288
rect 54850 -34240 54879 -34238
rect 54850 -34308 54860 -34240
rect 54840 -34318 54860 -34308
rect 54750 -34328 54860 -34318
rect 54920 -34368 54990 -34172
rect 55430 -34218 55520 -34208
rect 55290 -34328 55390 -34318
rect 53970 -34398 55290 -34368
rect 55430 -34358 55520 -34288
rect 53970 -34408 55390 -34398
rect 54050 -34418 55380 -34408
rect 54050 -34428 54880 -34418
rect 54050 -34438 54091 -34428
rect 54079 -34462 54091 -34438
rect 54867 -34438 54880 -34428
rect 54867 -34462 54879 -34438
rect 54079 -34468 54879 -34462
rect 54920 -34478 54990 -34468
rect 53510 -34506 53630 -34488
rect 53510 -34538 53526 -34506
rect 53514 -34540 53526 -34538
rect 53614 -34538 53630 -34506
rect 53940 -34490 54038 -34478
rect 53940 -34498 53998 -34490
rect 53614 -34540 53626 -34538
rect 53514 -34546 53626 -34540
rect 35900 -35258 39100 -35200
rect 25860 -35277 39100 -35258
rect 25860 -35674 25882 -35277
rect 26996 -35674 27124 -35277
rect 28238 -35674 28366 -35277
rect 29480 -35674 29608 -35277
rect 30722 -35674 30850 -35277
rect 31964 -35674 32092 -35277
rect 33206 -35674 33334 -35277
rect 34448 -35674 34576 -35277
rect 35690 -35300 39100 -35277
rect 35690 -35674 36000 -35300
rect 25860 -35944 36000 -35674
rect 25860 -36341 25882 -35944
rect 26996 -36341 27124 -35944
rect 28238 -36341 28366 -35944
rect 29480 -36341 29608 -35944
rect 30722 -36341 30850 -35944
rect 31964 -36341 32092 -35944
rect 33206 -36341 33334 -35944
rect 34448 -36341 34576 -35944
rect 35690 -36300 36000 -35944
rect 39000 -36300 39100 -35300
rect 35690 -36341 39100 -36300
rect 25860 -36358 39100 -36341
rect 35900 -36400 39100 -36358
rect 53000 -36308 53050 -34558
rect 53250 -34568 53480 -34558
rect 53250 -35918 53330 -34568
rect 53400 -34578 53480 -34568
rect 53400 -34590 53504 -34578
rect 53400 -35366 53464 -34590
rect 53498 -35366 53504 -34590
rect 53400 -35378 53504 -35366
rect 53636 -34588 53682 -34578
rect 53636 -34590 53760 -34588
rect 53636 -35366 53642 -34590
rect 53676 -35366 53760 -34590
rect 53940 -34598 53950 -34498
rect 54032 -34528 54038 -34490
rect 54020 -34540 54038 -34528
rect 54020 -34598 54030 -34540
rect 54079 -34556 54879 -34550
rect 54079 -34590 54091 -34556
rect 54867 -34590 54879 -34556
rect 54920 -34578 54990 -34568
rect 55320 -34568 55380 -34418
rect 54079 -34596 54879 -34590
rect 53940 -34618 54030 -34598
rect 54090 -34628 54870 -34596
rect 55320 -34602 55334 -34568
rect 55368 -34602 55380 -34568
rect 55320 -34608 55380 -34602
rect 53840 -34928 53920 -34918
rect 53840 -35038 53860 -34928
rect 53840 -35048 53920 -35038
rect 53840 -35240 53900 -35048
rect 54320 -35128 54510 -34628
rect 55440 -34638 55520 -34358
rect 55410 -34640 55520 -34638
rect 55284 -34648 55330 -34640
rect 55230 -34652 55330 -34648
rect 55230 -34658 55290 -34652
rect 55324 -34828 55330 -34652
rect 55230 -34838 55330 -34828
rect 55284 -34840 55330 -34838
rect 55372 -34648 55520 -34640
rect 55372 -34652 55430 -34648
rect 55372 -34828 55378 -34652
rect 55412 -34818 55430 -34652
rect 55510 -34818 55520 -34648
rect 55412 -34828 55520 -34818
rect 55372 -34840 55418 -34828
rect 55580 -34928 55720 -33640
rect 58776 -33870 59306 -33750
rect 58776 -33880 58966 -33870
rect 56146 -33980 57366 -33930
rect 55954 -34128 56046 -34116
rect 56146 -34128 56506 -33980
rect 55954 -34298 55960 -34128
rect 56040 -34298 56046 -34128
rect 55954 -34310 56046 -34298
rect 56120 -34158 56506 -34128
rect 56120 -34368 56190 -34158
rect 56390 -34230 56506 -34158
rect 57016 -34134 57366 -33980
rect 57586 -34030 58966 -33880
rect 59126 -34030 59306 -33870
rect 57586 -34050 59306 -34030
rect 59946 -33900 60386 -33800
rect 57586 -34080 58986 -34050
rect 59946 -34060 59956 -33900
rect 60166 -34060 60386 -33900
rect 57016 -34230 57368 -34134
rect 56390 -34270 57368 -34230
rect 56390 -34368 57126 -34270
rect 56120 -34374 57126 -34368
rect 56120 -34378 56750 -34374
rect 55880 -34418 55970 -34408
rect 55870 -34496 55880 -34450
rect 55970 -34496 55982 -34450
rect 55880 -34508 55970 -34498
rect 55000 -34938 55090 -34928
rect 55000 -35048 55090 -35038
rect 54710 -35128 54960 -35108
rect 53940 -35168 54960 -35128
rect 53940 -35172 54730 -35168
rect 53930 -35178 54730 -35172
rect 53930 -35212 53942 -35178
rect 54718 -35212 54730 -35178
rect 53930 -35218 54730 -35212
rect 53840 -35328 53858 -35240
rect 53892 -35328 53900 -35240
rect 53840 -35348 53900 -35328
rect 54762 -35238 54850 -35228
rect 54762 -35240 54770 -35238
rect 54762 -35328 54768 -35240
rect 54840 -35328 54850 -35238
rect 54762 -35340 54850 -35328
rect 54770 -35348 54850 -35340
rect 53636 -35378 53760 -35366
rect 53400 -35596 53480 -35378
rect 53514 -35416 53626 -35410
rect 53514 -35418 53526 -35416
rect 53510 -35450 53526 -35418
rect 53614 -35418 53626 -35416
rect 53614 -35450 53630 -35418
rect 53510 -35524 53630 -35450
rect 53510 -35558 53526 -35524
rect 53614 -35558 53630 -35524
rect 53680 -35438 53760 -35378
rect 53930 -35356 54730 -35350
rect 53930 -35390 53942 -35356
rect 54718 -35390 54730 -35356
rect 53930 -35396 54730 -35390
rect 53940 -35428 54720 -35396
rect 53920 -35438 54720 -35428
rect 53680 -35528 54720 -35438
rect 53514 -35564 53626 -35558
rect 53680 -35596 53760 -35528
rect 53920 -35538 54720 -35528
rect 53940 -35578 54720 -35538
rect 54900 -35568 54960 -35168
rect 55010 -35160 55090 -35048
rect 55540 -34938 55720 -34928
rect 55630 -35038 55720 -34938
rect 55130 -35074 55506 -35068
rect 55130 -35108 55142 -35074
rect 55494 -35108 55506 -35074
rect 55130 -35114 55506 -35108
rect 55010 -35194 55046 -35160
rect 55080 -35194 55090 -35160
rect 55010 -35208 55090 -35194
rect 55142 -35240 55494 -35114
rect 55540 -35160 55720 -35038
rect 55540 -35194 55556 -35160
rect 55590 -35194 55720 -35160
rect 55540 -35208 55720 -35194
rect 55780 -34540 55860 -34528
rect 55130 -35246 55506 -35240
rect 55130 -35280 55142 -35246
rect 55494 -35278 55506 -35246
rect 55494 -35280 55510 -35278
rect 55130 -35286 55510 -35280
rect 55140 -35298 55510 -35286
rect 55780 -35298 55820 -34540
rect 55140 -35316 55820 -35298
rect 55854 -35316 55860 -34540
rect 55140 -35328 55860 -35316
rect 55992 -34540 56038 -34528
rect 55992 -35316 55998 -34540
rect 56032 -34548 56038 -34540
rect 56120 -34548 56300 -34378
rect 57098 -34400 57126 -34374
rect 57356 -34400 57368 -34270
rect 57098 -34414 57368 -34400
rect 57096 -34445 57372 -34414
rect 57096 -34479 57125 -34445
rect 57159 -34479 57217 -34445
rect 57251 -34479 57309 -34445
rect 57343 -34479 57372 -34445
rect 57096 -34510 57372 -34479
rect 56032 -34906 56300 -34548
rect 56590 -34668 56660 -34658
rect 56660 -34734 57000 -34668
rect 57586 -34730 57706 -34080
rect 59946 -34090 60386 -34060
rect 71900 -34100 74100 -34000
rect 57366 -34734 57706 -34730
rect 56660 -34738 57188 -34734
rect 56660 -34744 57190 -34738
rect 56660 -34794 57118 -34744
rect 57178 -34794 57190 -34744
rect 57314 -34740 57706 -34734
rect 57314 -34780 57326 -34740
rect 57366 -34780 57706 -34740
rect 57314 -34786 57706 -34780
rect 57366 -34790 57706 -34786
rect 58896 -34370 58986 -34350
rect 58896 -34430 58906 -34370
rect 58896 -34720 58926 -34430
rect 58966 -34720 58986 -34370
rect 59106 -34370 59516 -34360
rect 59106 -34430 59216 -34370
rect 59276 -34430 59326 -34370
rect 59386 -34430 59436 -34370
rect 59496 -34430 59516 -34370
rect 59106 -34447 59516 -34430
rect 59626 -34370 59706 -34330
rect 59626 -34430 59636 -34370
rect 59626 -34440 59656 -34430
rect 59106 -34480 59125 -34447
rect 59113 -34481 59125 -34480
rect 59501 -34480 59516 -34447
rect 59501 -34481 59513 -34480
rect 59113 -34487 59513 -34481
rect 59546 -34490 59616 -34480
rect 59276 -34530 59356 -34520
rect 59276 -34549 59286 -34530
rect 59113 -34555 59286 -34549
rect 59346 -34549 59356 -34530
rect 59346 -34555 59513 -34549
rect 59113 -34589 59125 -34555
rect 59501 -34589 59513 -34555
rect 59606 -34550 59616 -34490
rect 59546 -34560 59616 -34550
rect 59113 -34590 59286 -34589
rect 59346 -34590 59513 -34589
rect 59016 -34600 59076 -34590
rect 59113 -34595 59513 -34590
rect 59276 -34600 59356 -34595
rect 59546 -34610 59616 -34600
rect 59016 -34670 59076 -34660
rect 59113 -34663 59513 -34657
rect 59113 -34697 59125 -34663
rect 59501 -34697 59513 -34663
rect 59606 -34670 59616 -34610
rect 59546 -34680 59616 -34670
rect 59113 -34700 59513 -34697
rect 59113 -34703 59516 -34700
rect 58896 -34730 58986 -34720
rect 58896 -34790 58906 -34730
rect 58966 -34790 58986 -34730
rect 58896 -34792 58986 -34790
rect 59116 -34720 59516 -34703
rect 59646 -34710 59656 -34440
rect 59116 -34780 59216 -34720
rect 59276 -34780 59336 -34720
rect 59396 -34780 59436 -34720
rect 59496 -34780 59516 -34720
rect 56660 -34798 57190 -34794
rect 56590 -34800 57190 -34798
rect 56590 -34804 57188 -34800
rect 56590 -34868 57000 -34804
rect 56032 -34918 56356 -34906
rect 56032 -35316 56280 -34918
rect 55992 -35328 56280 -35316
rect 55140 -35338 55200 -35328
rect 55450 -35358 55810 -35328
rect 55870 -35366 55982 -35360
rect 55870 -35400 55882 -35366
rect 55970 -35400 55982 -35366
rect 55870 -35406 55982 -35400
rect 55140 -35418 55200 -35408
rect 55024 -35448 55116 -35436
rect 55024 -35528 55030 -35448
rect 55110 -35528 55116 -35448
rect 55024 -35540 55116 -35528
rect 55734 -35448 55816 -35436
rect 55734 -35528 55740 -35448
rect 55810 -35528 55816 -35448
rect 55734 -35540 55816 -35528
rect 55880 -35438 55970 -35406
rect 55880 -35564 55970 -35528
rect 56060 -35548 56280 -35328
rect 56350 -35548 56356 -34918
rect 56480 -34988 56550 -34978
rect 56480 -35058 56550 -35048
rect 56590 -35087 56750 -34868
rect 58894 -34886 58988 -34792
rect 59116 -34800 59516 -34780
rect 59636 -34720 59656 -34710
rect 59696 -34720 59706 -34370
rect 59856 -34540 59976 -34530
rect 59856 -34630 59866 -34540
rect 59966 -34630 59976 -34540
rect 59856 -34640 59976 -34630
rect 60436 -34620 60446 -34520
rect 60526 -34620 60536 -34520
rect 60436 -34640 60536 -34620
rect 59636 -34730 59706 -34720
rect 59696 -34790 59706 -34730
rect 59636 -34810 59706 -34790
rect 59756 -34660 60536 -34640
rect 59756 -34700 59866 -34660
rect 60426 -34700 60536 -34660
rect 59756 -34710 60536 -34700
rect 59756 -34750 59826 -34710
rect 59066 -34840 59176 -34830
rect 58896 -34950 58986 -34886
rect 59066 -34910 59076 -34840
rect 59166 -34910 59176 -34840
rect 59066 -34912 59103 -34910
rect 59137 -34912 59176 -34910
rect 59066 -34920 59176 -34912
rect 59756 -34940 59766 -34750
rect 59806 -34940 59826 -34750
rect 59956 -34768 60046 -34740
rect 59946 -34774 60046 -34768
rect 60126 -34768 60336 -34740
rect 60126 -34774 60346 -34768
rect 59856 -34810 59916 -34800
rect 59946 -34808 59958 -34774
rect 60334 -34808 60346 -34774
rect 59946 -34814 60346 -34808
rect 60376 -34820 60446 -34810
rect 59856 -34890 59916 -34880
rect 59946 -34882 60346 -34876
rect 59946 -34916 59958 -34882
rect 60334 -34916 60346 -34882
rect 60376 -34890 60446 -34880
rect 59946 -34922 59976 -34916
rect 57098 -34958 57368 -34954
rect 57096 -34964 57372 -34958
rect 57096 -35050 57098 -34964
rect 56424 -35088 56470 -35087
rect 56060 -35560 56356 -35548
rect 56410 -35099 56470 -35088
rect 53400 -35608 53504 -35596
rect 53400 -35918 53464 -35608
rect 53250 -36308 53464 -35918
rect 53000 -36384 53464 -36308
rect 53498 -36384 53504 -35608
rect 53000 -36388 53504 -36384
rect 53458 -36396 53504 -36388
rect 53636 -35608 53760 -35596
rect 53636 -36384 53642 -35608
rect 53676 -36384 53760 -35608
rect 53930 -35584 54730 -35578
rect 53930 -35618 53942 -35584
rect 54718 -35618 54730 -35584
rect 53930 -35624 54730 -35618
rect 53830 -35646 53900 -35628
rect 53830 -35734 53858 -35646
rect 53892 -35734 53900 -35646
rect 53830 -35928 53900 -35734
rect 54760 -35646 54850 -35628
rect 54760 -35734 54768 -35646
rect 54802 -35648 54850 -35646
rect 54900 -35638 55200 -35568
rect 55870 -35570 55982 -35564
rect 55870 -35604 55882 -35570
rect 55970 -35604 55982 -35570
rect 55450 -35638 55810 -35608
rect 55870 -35610 55982 -35604
rect 56060 -35638 56300 -35560
rect 54900 -35642 55820 -35638
rect 56000 -35642 56300 -35638
rect 54900 -35648 55860 -35642
rect 54840 -35728 54850 -35648
rect 54802 -35734 54850 -35728
rect 54760 -35748 54850 -35734
rect 55130 -35654 55860 -35648
rect 55130 -35678 55820 -35654
rect 55130 -35696 55510 -35678
rect 55130 -35730 55142 -35696
rect 55494 -35698 55510 -35696
rect 55494 -35730 55506 -35698
rect 55130 -35736 55506 -35730
rect 53930 -35762 54730 -35756
rect 53930 -35796 53942 -35762
rect 54718 -35796 54730 -35762
rect 55020 -35782 55090 -35768
rect 53930 -35802 54730 -35796
rect 53940 -35808 54730 -35802
rect 54920 -35798 54980 -35788
rect 53940 -35848 54920 -35808
rect 53830 -35938 53920 -35928
rect 53830 -36048 53850 -35938
rect 53830 -36058 53920 -36048
rect 54320 -36348 54510 -35848
rect 54710 -35868 54920 -35848
rect 54910 -35878 54980 -35868
rect 55020 -35816 55046 -35782
rect 55080 -35816 55090 -35782
rect 55020 -35928 55090 -35816
rect 55142 -35862 55494 -35736
rect 55540 -35782 55620 -35768
rect 55540 -35816 55556 -35782
rect 55590 -35816 55620 -35782
rect 55130 -35868 55506 -35862
rect 55130 -35902 55142 -35868
rect 55494 -35902 55506 -35868
rect 55130 -35908 55506 -35902
rect 55000 -35938 55090 -35928
rect 55000 -36048 55090 -36038
rect 55540 -35928 55620 -35816
rect 55540 -35938 55630 -35928
rect 55630 -36038 55680 -35948
rect 55540 -36048 55680 -36038
rect 55274 -36138 55320 -36136
rect 55220 -36148 55320 -36138
rect 55220 -36324 55280 -36318
rect 55314 -36324 55320 -36148
rect 55220 -36328 55320 -36324
rect 55274 -36336 55320 -36328
rect 55362 -36148 55408 -36136
rect 55362 -36324 55368 -36148
rect 55402 -36158 55510 -36148
rect 55402 -36324 55410 -36158
rect 55362 -36328 55410 -36324
rect 55500 -36328 55510 -36158
rect 55362 -36336 55510 -36328
rect 55390 -36338 55510 -36336
rect 53636 -36388 53760 -36384
rect 53636 -36396 53682 -36388
rect 53940 -36408 54020 -36368
rect 54080 -36382 54860 -36348
rect 55311 -36374 55371 -36368
rect 53514 -36434 53626 -36428
rect 53514 -36438 53526 -36434
rect 53510 -36468 53526 -36438
rect 53614 -36438 53626 -36434
rect 53614 -36468 53630 -36438
rect 53510 -36528 53630 -36468
rect 53940 -36488 53950 -36408
rect 54010 -36438 54020 -36408
rect 54069 -36388 54869 -36382
rect 54069 -36422 54081 -36388
rect 54857 -36422 54869 -36388
rect 54069 -36428 54869 -36422
rect 54910 -36398 54980 -36388
rect 54010 -36450 54028 -36438
rect 54022 -36488 54028 -36450
rect 53940 -36500 54028 -36488
rect 53940 -36508 54020 -36500
rect 54910 -36508 54980 -36498
rect 55311 -36408 55324 -36374
rect 55358 -36408 55371 -36374
rect 54070 -36510 54870 -36508
rect 54069 -36516 54870 -36510
rect 54069 -36538 54081 -36516
rect 54041 -36550 54081 -36538
rect 54857 -36518 54870 -36516
rect 54857 -36550 54880 -36518
rect 55311 -36548 55371 -36408
rect 54041 -36558 54880 -36550
rect 55240 -36558 55371 -36548
rect 54041 -36568 55240 -36558
rect 53510 -36658 53630 -36648
rect 53961 -36608 55240 -36568
rect 35900 -36860 40100 -36800
rect 53961 -36806 54031 -36608
rect 54730 -36668 54860 -36658
rect 54730 -36688 54740 -36668
rect 54080 -36738 54740 -36688
rect 54069 -36744 54740 -36738
rect 54850 -36738 54860 -36668
rect 54850 -36744 54869 -36738
rect 54069 -36778 54081 -36744
rect 54857 -36778 54869 -36744
rect 54069 -36784 54869 -36778
rect 54911 -36794 54981 -36608
rect 55370 -36608 55371 -36558
rect 55240 -36628 55370 -36618
rect 55410 -36648 55510 -36338
rect 55410 -36758 55510 -36738
rect 55570 -36668 55680 -36048
rect 55780 -36430 55820 -35678
rect 55854 -36430 55860 -35654
rect 55780 -36438 55860 -36430
rect 55814 -36442 55860 -36438
rect 55992 -35654 56300 -35642
rect 55992 -36430 55998 -35654
rect 56032 -36428 56300 -35654
rect 56410 -35698 56430 -35099
rect 56380 -35875 56430 -35698
rect 56464 -35875 56470 -35099
rect 56380 -35887 56470 -35875
rect 56552 -35099 56750 -35087
rect 56552 -35875 56558 -35099
rect 56592 -35238 56750 -35099
rect 57066 -35080 57098 -35050
rect 57368 -35050 57372 -34964
rect 58896 -34959 59076 -34950
rect 58896 -34960 59084 -34959
rect 59156 -34960 59202 -34959
rect 57368 -35080 57396 -35050
rect 57066 -35210 57086 -35080
rect 57376 -35210 57396 -35080
rect 56592 -35875 56610 -35238
rect 57066 -35240 57396 -35210
rect 56860 -35390 57060 -35378
rect 56860 -35418 57236 -35390
rect 56860 -35548 56900 -35418
rect 57020 -35548 57236 -35418
rect 56860 -35588 57236 -35548
rect 57036 -35590 57236 -35588
rect 58556 -35480 58756 -35460
rect 58556 -35640 58576 -35480
rect 58736 -35640 58756 -35480
rect 58556 -35660 58756 -35640
rect 56552 -35878 56610 -35875
rect 57036 -35740 57446 -35730
rect 56552 -35887 56598 -35878
rect 57036 -35880 57056 -35740
rect 57416 -35880 57446 -35740
rect 56380 -36158 56440 -35887
rect 57036 -35900 57098 -35880
rect 56480 -35928 56550 -35918
rect 56480 -35998 56550 -35988
rect 57096 -36014 57098 -35934
rect 57368 -35900 57446 -35880
rect 57368 -36014 57372 -35934
rect 57096 -36030 57372 -36014
rect 58896 -36090 58926 -34960
rect 58966 -34971 59086 -34960
rect 58966 -35347 59044 -34971
rect 59078 -35347 59086 -34971
rect 58966 -35370 59086 -35347
rect 59156 -34971 59256 -34960
rect 59756 -34970 59826 -34940
rect 59966 -34952 59976 -34922
rect 60316 -34922 60346 -34916
rect 61036 -34920 61466 -34910
rect 60316 -34952 60326 -34922
rect 59966 -34960 60326 -34952
rect 59156 -35347 59162 -34971
rect 59196 -35040 59256 -34971
rect 59236 -35120 59256 -35040
rect 59196 -35240 59256 -35120
rect 59236 -35320 59256 -35240
rect 59196 -35347 59256 -35320
rect 59156 -35360 59256 -35347
rect 58966 -35680 59036 -35370
rect 59066 -35406 59176 -35400
rect 59066 -35410 59103 -35406
rect 59137 -35410 59176 -35406
rect 59066 -35480 59076 -35410
rect 59166 -35480 59176 -35410
rect 59066 -35490 59176 -35480
rect 59206 -35560 59256 -35360
rect 59376 -34990 59826 -34970
rect 59376 -35030 59476 -34990
rect 59656 -35030 59826 -34990
rect 59376 -35040 59826 -35030
rect 59376 -35090 59436 -35040
rect 59376 -35450 59386 -35090
rect 59426 -35450 59436 -35090
rect 59526 -35098 59576 -35070
rect 59526 -35132 59546 -35098
rect 59636 -35130 59706 -35070
rect 59580 -35132 59706 -35130
rect 59526 -35140 59706 -35132
rect 59476 -35182 59546 -35170
rect 59476 -35250 59502 -35182
rect 59476 -35358 59502 -35320
rect 59536 -35358 59546 -35182
rect 59476 -35370 59546 -35358
rect 59576 -35182 59636 -35170
rect 59576 -35190 59590 -35182
rect 59624 -35190 59636 -35182
rect 59576 -35370 59636 -35360
rect 59534 -35408 59592 -35402
rect 59534 -35410 59546 -35408
rect 59066 -35570 59176 -35560
rect 59066 -35640 59076 -35570
rect 59166 -35640 59176 -35570
rect 59066 -35642 59103 -35640
rect 59137 -35642 59176 -35640
rect 59066 -35650 59176 -35642
rect 59206 -35570 59266 -35560
rect 59206 -35650 59266 -35640
rect 59376 -35600 59436 -35450
rect 59516 -35442 59546 -35410
rect 59580 -35410 59592 -35408
rect 59666 -35410 59706 -35140
rect 59580 -35442 59706 -35410
rect 59516 -35480 59706 -35442
rect 59746 -35098 59936 -35070
rect 59746 -35132 59862 -35098
rect 59896 -35132 59936 -35098
rect 59746 -35140 59936 -35132
rect 61036 -35100 61206 -34920
rect 61346 -35100 61466 -34920
rect 61036 -35140 61466 -35100
rect 59746 -35400 59776 -35140
rect 60286 -35150 60476 -35140
rect 59806 -35182 59866 -35170
rect 59806 -35200 59818 -35182
rect 59852 -35200 59866 -35182
rect 59806 -35358 59818 -35340
rect 59852 -35358 59866 -35340
rect 59806 -35370 59866 -35358
rect 59900 -35180 60016 -35170
rect 59900 -35182 59916 -35180
rect 59900 -35358 59906 -35182
rect 59900 -35360 59916 -35358
rect 60006 -35360 60016 -35180
rect 60286 -35290 60306 -35150
rect 60456 -35290 60476 -35150
rect 61176 -35200 61386 -35180
rect 60286 -35300 60476 -35290
rect 61026 -35220 61136 -35210
rect 59900 -35370 60016 -35360
rect 60076 -35357 60196 -35320
rect 60076 -35391 60127 -35357
rect 60161 -35391 60196 -35357
rect 59746 -35408 59926 -35400
rect 59746 -35410 59862 -35408
rect 59896 -35410 59926 -35408
rect 59746 -35480 59826 -35410
rect 59916 -35480 59926 -35410
rect 59746 -35490 59926 -35480
rect 60076 -35449 60196 -35391
rect 60336 -35360 60446 -35300
rect 60336 -35400 60366 -35360
rect 60406 -35400 60446 -35360
rect 60636 -35357 60816 -35320
rect 60636 -35391 60671 -35357
rect 60705 -35391 60747 -35357
rect 60781 -35391 60816 -35357
rect 60076 -35480 60127 -35449
rect 60161 -35480 60196 -35449
rect 59736 -35570 59936 -35560
rect 58966 -35701 59086 -35680
rect 58966 -36077 59044 -35701
rect 59078 -36077 59086 -35701
rect 58966 -36090 59086 -36077
rect 59156 -35690 59202 -35689
rect 59156 -35701 59236 -35690
rect 59156 -36077 59162 -35701
rect 59196 -35730 59236 -35701
rect 59226 -35810 59236 -35730
rect 59196 -35960 59236 -35810
rect 59226 -36040 59236 -35960
rect 59196 -36077 59236 -36040
rect 59376 -35970 59386 -35600
rect 59426 -35970 59436 -35600
rect 59516 -35611 59706 -35570
rect 59516 -35645 59545 -35611
rect 59579 -35645 59706 -35611
rect 59516 -35650 59706 -35645
rect 59533 -35651 59591 -35650
rect 59466 -35695 59546 -35680
rect 59586 -35683 59646 -35680
rect 59466 -35730 59501 -35695
rect 59466 -35871 59501 -35810
rect 59535 -35871 59546 -35695
rect 59466 -35880 59546 -35871
rect 59583 -35695 59646 -35683
rect 59583 -35710 59589 -35695
rect 59623 -35710 59646 -35695
rect 59583 -35850 59586 -35710
rect 59583 -35871 59589 -35850
rect 59623 -35871 59646 -35850
rect 59583 -35880 59646 -35871
rect 59495 -35883 59541 -35880
rect 59583 -35883 59629 -35880
rect 59533 -35920 59591 -35915
rect 59676 -35920 59706 -35650
rect 59376 -36010 59436 -35970
rect 59506 -35980 59516 -35920
rect 59596 -35980 59706 -35920
rect 59736 -35640 59826 -35570
rect 59926 -35640 59936 -35570
rect 59736 -35645 59861 -35640
rect 59895 -35645 59936 -35640
rect 59736 -35650 59936 -35645
rect 60076 -35640 60096 -35480
rect 60176 -35640 60196 -35480
rect 59736 -35920 59766 -35650
rect 59849 -35651 59907 -35650
rect 60076 -35667 60127 -35640
rect 60161 -35667 60196 -35640
rect 59796 -35683 59856 -35680
rect 59796 -35690 59857 -35683
rect 59856 -35870 59857 -35690
rect 59796 -35871 59817 -35870
rect 59851 -35871 59857 -35870
rect 59796 -35880 59857 -35871
rect 59811 -35883 59857 -35880
rect 59899 -35690 59945 -35683
rect 59899 -35695 59916 -35690
rect 59899 -35871 59905 -35695
rect 59899 -35880 59916 -35871
rect 60006 -35880 60016 -35690
rect 60076 -35725 60196 -35667
rect 60346 -35450 60426 -35400
rect 60346 -35490 60366 -35450
rect 60406 -35490 60426 -35450
rect 60346 -35540 60426 -35490
rect 60346 -35580 60366 -35540
rect 60406 -35580 60426 -35540
rect 60346 -35620 60426 -35580
rect 60346 -35660 60366 -35620
rect 60406 -35660 60426 -35620
rect 60346 -35670 60426 -35660
rect 60636 -35449 60816 -35391
rect 60636 -35483 60671 -35449
rect 60705 -35483 60747 -35449
rect 60781 -35483 60816 -35449
rect 60636 -35541 60816 -35483
rect 60636 -35575 60671 -35541
rect 60705 -35575 60747 -35541
rect 60781 -35575 60816 -35541
rect 60636 -35633 60816 -35575
rect 60636 -35667 60671 -35633
rect 60705 -35667 60747 -35633
rect 60781 -35667 60816 -35633
rect 60076 -35759 60127 -35725
rect 60161 -35759 60196 -35725
rect 60076 -35790 60196 -35759
rect 60276 -35710 60546 -35700
rect 60276 -35725 60476 -35710
rect 60276 -35759 60297 -35725
rect 60331 -35759 60369 -35725
rect 60405 -35759 60449 -35725
rect 60276 -35770 60476 -35759
rect 60536 -35770 60546 -35710
rect 60276 -35780 60546 -35770
rect 60636 -35725 60816 -35667
rect 61026 -35330 61036 -35220
rect 61126 -35330 61136 -35220
rect 61176 -35280 61196 -35200
rect 61366 -35280 61386 -35200
rect 61176 -35300 61386 -35280
rect 61026 -35360 61136 -35330
rect 61026 -35400 61046 -35360
rect 61086 -35400 61136 -35360
rect 61026 -35450 61136 -35400
rect 61026 -35490 61046 -35450
rect 61086 -35490 61136 -35450
rect 61026 -35540 61136 -35490
rect 61026 -35580 61046 -35540
rect 61086 -35580 61136 -35540
rect 61026 -35620 61136 -35580
rect 61026 -35660 61046 -35620
rect 61086 -35660 61136 -35620
rect 61026 -35680 61136 -35660
rect 61256 -35357 61366 -35300
rect 61256 -35391 61291 -35357
rect 61325 -35391 61366 -35357
rect 61256 -35449 61366 -35391
rect 61256 -35450 61291 -35449
rect 61325 -35450 61366 -35449
rect 61256 -35660 61276 -35450
rect 61356 -35660 61366 -35450
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 61256 -35667 61291 -35660
rect 61325 -35667 61366 -35660
rect 60636 -35759 60671 -35725
rect 60705 -35759 60747 -35725
rect 60781 -35759 60816 -35725
rect 60636 -35840 60816 -35759
rect 60966 -35724 61177 -35710
rect 60966 -35725 61129 -35724
rect 60966 -35759 60980 -35725
rect 61015 -35759 61053 -35725
rect 61088 -35758 61129 -35725
rect 61164 -35758 61177 -35724
rect 61088 -35759 61177 -35758
rect 60966 -35790 61177 -35759
rect 61256 -35725 61366 -35667
rect 61256 -35759 61291 -35725
rect 61325 -35759 61366 -35725
rect 61256 -35790 61366 -35759
rect 60466 -35850 60546 -35840
rect 59899 -35883 59945 -35880
rect 60466 -35910 60476 -35850
rect 60536 -35910 60546 -35850
rect 59849 -35920 59907 -35915
rect 60466 -35920 60546 -35910
rect 60606 -35850 60826 -35840
rect 60606 -35910 60616 -35850
rect 60736 -35910 60756 -35850
rect 60816 -35910 60826 -35850
rect 60606 -35920 60826 -35910
rect 60886 -35850 60966 -35840
rect 60886 -35910 60896 -35850
rect 60956 -35910 60966 -35850
rect 60886 -35920 60966 -35910
rect 59736 -35921 59926 -35920
rect 59736 -35955 59861 -35921
rect 59895 -35955 59926 -35921
rect 59736 -35980 59926 -35955
rect 60636 -35970 60816 -35920
rect 59376 -36020 59826 -36010
rect 59376 -36060 59476 -36020
rect 59646 -36060 59826 -36020
rect 59376 -36070 59826 -36060
rect 59156 -36090 59236 -36077
rect 58896 -36100 59086 -36090
rect 56380 -36168 57000 -36158
rect 57356 -36164 57676 -36150
rect 56440 -36174 57000 -36168
rect 57314 -36170 57676 -36164
rect 56440 -36194 57178 -36174
rect 56440 -36244 57118 -36194
rect 57168 -36244 57178 -36194
rect 57314 -36210 57326 -36170
rect 57376 -36210 57676 -36170
rect 57314 -36216 57676 -36210
rect 57356 -36230 57676 -36216
rect 56440 -36254 57178 -36244
rect 56440 -36288 57000 -36254
rect 57112 -36256 57174 -36254
rect 56380 -36358 57000 -36288
rect 56032 -36430 56038 -36428
rect 55992 -36442 56038 -36430
rect 55880 -36474 55970 -36468
rect 55870 -36478 55982 -36474
rect 55870 -36520 55880 -36478
rect 55970 -36520 55982 -36478
rect 55880 -36568 55970 -36558
rect 56120 -36598 56300 -36428
rect 57096 -36509 57372 -36478
rect 57096 -36543 57125 -36509
rect 57159 -36543 57217 -36509
rect 57251 -36543 57309 -36509
rect 57343 -36520 57372 -36509
rect 57343 -36543 57376 -36520
rect 57096 -36580 57376 -36543
rect 57066 -36590 57376 -36580
rect 56426 -36598 57376 -36590
rect 56120 -36608 57376 -36598
rect 56014 -36658 56086 -36646
rect 55570 -36778 55830 -36668
rect 53961 -36844 53988 -36806
rect 54022 -36844 54031 -36806
rect 53961 -36858 54031 -36844
rect 54910 -36806 54981 -36794
rect 54910 -36844 54916 -36806
rect 54950 -36844 54981 -36806
rect 54910 -36856 54981 -36844
rect 54911 -36858 54981 -36856
rect 55220 -36818 55330 -36808
rect 25862 -36879 40100 -36860
rect 25862 -37276 25882 -36879
rect 26996 -37276 27124 -36879
rect 28238 -37276 28366 -36879
rect 29480 -37276 29608 -36879
rect 30722 -37276 30850 -36879
rect 31964 -37276 32092 -36879
rect 33206 -37276 33334 -36879
rect 34448 -37276 34576 -36879
rect 35690 -36900 40100 -36879
rect 35690 -37276 36000 -36900
rect 25862 -37544 36000 -37276
rect 25862 -37941 25882 -37544
rect 26996 -37941 27124 -37544
rect 28238 -37941 28366 -37544
rect 29480 -37941 29608 -37544
rect 30722 -37941 30850 -37544
rect 31964 -37941 32092 -37544
rect 33206 -37941 33334 -37544
rect 34448 -37941 34576 -37544
rect 35690 -37900 36000 -37544
rect 40000 -37900 40100 -36900
rect 54069 -36872 54869 -36866
rect 54069 -36906 54081 -36872
rect 54857 -36878 54869 -36872
rect 54857 -36906 54880 -36878
rect 54069 -36912 54880 -36906
rect 54090 -36988 54880 -36912
rect 55330 -36918 55380 -36818
rect 55330 -36928 55480 -36918
rect 55220 -36938 55480 -36928
rect 55280 -36952 55480 -36938
rect 55280 -36958 55488 -36952
rect 55280 -36978 55300 -36958
rect 54090 -37088 54150 -36988
rect 54840 -37088 54880 -36988
rect 55288 -36992 55300 -36978
rect 55476 -36992 55488 -36958
rect 55530 -36978 55610 -36968
rect 55288 -36998 55488 -36992
rect 55520 -37002 55530 -36990
rect 55520 -37036 55526 -37002
rect 55288 -37046 55488 -37040
rect 55288 -37080 55300 -37046
rect 55476 -37080 55488 -37046
rect 55520 -37048 55530 -37036
rect 55530 -37078 55610 -37068
rect 55288 -37086 55488 -37080
rect 54090 -37108 54140 -37088
rect 54100 -37348 54140 -37108
rect 54850 -37348 54880 -37088
rect 55300 -37128 55470 -37086
rect 55300 -37268 55320 -37128
rect 55470 -37214 55482 -37142
rect 55300 -37278 55470 -37268
rect 54100 -37388 54880 -37348
rect 55710 -37598 55830 -36778
rect 56014 -36808 56020 -36658
rect 56080 -36808 56086 -36658
rect 56014 -36820 56086 -36808
rect 56120 -36808 56170 -36608
rect 56390 -36660 57376 -36608
rect 56390 -36668 57156 -36660
rect 56390 -36808 56654 -36668
rect 56120 -36858 56654 -36808
rect 56306 -36886 56654 -36858
rect 56998 -36820 57156 -36668
rect 57316 -36820 57376 -36660
rect 56998 -36886 57376 -36820
rect 56306 -37300 57376 -36886
rect 57556 -37010 57676 -36230
rect 58896 -36260 58986 -36100
rect 59756 -36120 59826 -36070
rect 59066 -36136 59176 -36130
rect 59066 -36140 59103 -36136
rect 59137 -36140 59176 -36136
rect 59066 -36200 59076 -36140
rect 59166 -36200 59176 -36140
rect 59066 -36210 59176 -36200
rect 58896 -36630 58926 -36260
rect 58966 -36630 58986 -36330
rect 59116 -36260 59506 -36240
rect 59116 -36330 59146 -36260
rect 59226 -36330 59276 -36260
rect 59356 -36330 59396 -36260
rect 59476 -36330 59506 -36260
rect 59116 -36348 59506 -36330
rect 59646 -36260 59716 -36240
rect 59706 -36320 59716 -36260
rect 59646 -36330 59716 -36320
rect 59113 -36354 59513 -36348
rect 59113 -36388 59125 -36354
rect 59501 -36388 59513 -36354
rect 59113 -36394 59513 -36388
rect 59546 -36400 59616 -36390
rect 59246 -36456 59256 -36430
rect 59113 -36462 59256 -36456
rect 59366 -36456 59376 -36430
rect 59366 -36462 59513 -36456
rect 59016 -36500 59076 -36480
rect 59113 -36496 59125 -36462
rect 59501 -36496 59513 -36462
rect 59606 -36460 59616 -36400
rect 59546 -36470 59616 -36460
rect 59113 -36502 59513 -36496
rect 59016 -36590 59076 -36560
rect 59113 -36570 59513 -36564
rect 59113 -36604 59125 -36570
rect 59501 -36604 59513 -36570
rect 59113 -36610 59513 -36604
rect 58896 -36700 58906 -36630
rect 58896 -36720 58986 -36700
rect 59116 -36630 59516 -36610
rect 59116 -36700 59146 -36630
rect 59226 -36700 59276 -36630
rect 59356 -36700 59396 -36630
rect 59476 -36700 59516 -36630
rect 59116 -36720 59516 -36700
rect 59646 -36630 59656 -36330
rect 59706 -36630 59716 -36330
rect 59756 -36300 59766 -36120
rect 59806 -36300 59826 -36120
rect 59956 -36120 60336 -36110
rect 59956 -36134 59966 -36120
rect 59946 -36140 59966 -36134
rect 60326 -36134 60336 -36120
rect 60326 -36140 60346 -36134
rect 59856 -36180 59916 -36170
rect 59946 -36174 59958 -36140
rect 60334 -36174 60346 -36140
rect 61056 -36140 61176 -35790
rect 59946 -36180 59966 -36174
rect 60326 -36180 60346 -36174
rect 60376 -36180 60436 -36160
rect 59956 -36190 60336 -36180
rect 59856 -36260 59916 -36240
rect 59946 -36248 60346 -36242
rect 59756 -36340 59826 -36300
rect 59946 -36282 59958 -36248
rect 60334 -36282 60346 -36248
rect 60376 -36260 60436 -36240
rect 61126 -36240 61176 -36140
rect 61056 -36270 61176 -36240
rect 59946 -36288 60346 -36282
rect 59946 -36340 60336 -36288
rect 59756 -36360 60536 -36340
rect 59756 -36400 59866 -36360
rect 60426 -36400 60536 -36360
rect 59756 -36410 60536 -36400
rect 59796 -36520 59806 -36410
rect 59916 -36520 59926 -36410
rect 59796 -36530 59926 -36520
rect 60436 -36430 60536 -36410
rect 60436 -36550 60446 -36430
rect 60526 -36550 60536 -36430
rect 60436 -36560 60536 -36550
rect 59646 -36640 59716 -36630
rect 59706 -36700 59716 -36640
rect 59646 -36720 59716 -36700
rect 58806 -37010 59356 -36980
rect 59846 -36990 60256 -36980
rect 59846 -37000 59996 -36990
rect 57556 -37020 59356 -37010
rect 57556 -37160 58986 -37020
rect 59126 -37160 59356 -37020
rect 57556 -37210 59356 -37160
rect 58806 -37290 59356 -37210
rect 59800 -37100 59996 -37000
rect 60106 -37000 60256 -36990
rect 60106 -37100 60300 -37000
rect 59800 -37200 60300 -37100
rect 59800 -37400 59900 -37200
rect 60200 -37400 60300 -37200
rect 59800 -37500 60300 -37400
rect 55710 -37600 55910 -37598
rect 35690 -37941 40100 -37900
rect 25862 -37960 40100 -37941
rect 35900 -38000 40100 -37960
rect 55300 -37700 56200 -37600
rect 55300 -38100 55400 -37700
rect 56100 -38100 56200 -37700
rect 55300 -38200 56200 -38100
rect 84700 -38050 85660 -37780
rect 73180 -38360 73380 -38140
rect 35900 -38460 41100 -38400
rect 25860 -38479 41100 -38460
rect 25860 -38876 25882 -38479
rect 26996 -38876 27124 -38479
rect 28238 -38876 28366 -38479
rect 29480 -38876 29608 -38479
rect 30722 -38876 30850 -38479
rect 31964 -38876 32092 -38479
rect 33206 -38876 33334 -38479
rect 34448 -38876 34576 -38479
rect 35690 -38500 41100 -38479
rect 35690 -38876 36000 -38500
rect 25860 -39146 36000 -38876
rect 25860 -39543 25884 -39146
rect 26998 -39543 27126 -39146
rect 28240 -39543 28368 -39146
rect 29482 -39543 29610 -39146
rect 30724 -39543 30852 -39146
rect 31966 -39543 32094 -39146
rect 33208 -39543 33336 -39146
rect 34450 -39543 34578 -39146
rect 35692 -39500 36000 -39146
rect 41000 -39500 41100 -38500
rect 73180 -38550 73220 -38360
rect 73340 -38550 73380 -38360
rect 73180 -38560 73380 -38550
rect 73430 -38360 73630 -38140
rect 73430 -38550 73470 -38360
rect 73590 -38550 73630 -38360
rect 73430 -38560 73630 -38550
rect 73680 -38360 73880 -38140
rect 73680 -38550 73720 -38360
rect 73840 -38550 73880 -38360
rect 73680 -38560 73880 -38550
rect 73930 -38360 74130 -38140
rect 73930 -38550 73970 -38360
rect 74090 -38550 74130 -38360
rect 73930 -38560 74130 -38550
rect 74180 -38360 74380 -38140
rect 74180 -38550 74220 -38360
rect 74340 -38550 74380 -38360
rect 74180 -38560 74380 -38550
rect 74430 -38360 74630 -38140
rect 74430 -38550 74470 -38360
rect 74590 -38550 74630 -38360
rect 74430 -38560 74630 -38550
rect 74680 -38360 74880 -38140
rect 74680 -38550 74720 -38360
rect 74840 -38550 74880 -38360
rect 74680 -38560 74880 -38550
rect 74930 -38360 75130 -38140
rect 74930 -38550 74970 -38360
rect 75090 -38550 75130 -38360
rect 74930 -38560 75130 -38550
rect 75180 -38150 75560 -38140
rect 75180 -38270 75390 -38150
rect 75550 -38270 75560 -38150
rect 75180 -38280 75560 -38270
rect 75180 -38360 75380 -38280
rect 76880 -38340 77260 -38336
rect 75180 -38550 75220 -38360
rect 75340 -38550 75380 -38360
rect 75500 -38350 77260 -38340
rect 75500 -38371 77110 -38350
rect 75500 -38405 75535 -38371
rect 75569 -38405 75627 -38371
rect 75661 -38405 75719 -38371
rect 75753 -38405 75811 -38371
rect 75845 -38405 75903 -38371
rect 75937 -38405 75995 -38371
rect 76029 -38405 76085 -38371
rect 76119 -38405 76177 -38371
rect 76211 -38405 76269 -38371
rect 76303 -38405 76361 -38371
rect 76395 -38405 76453 -38371
rect 76487 -38405 76545 -38371
rect 76579 -38405 76637 -38371
rect 76671 -38405 76729 -38371
rect 76763 -38405 76821 -38371
rect 76855 -38405 77110 -38371
rect 75500 -38410 77110 -38405
rect 75500 -38440 76920 -38410
rect 75661 -38500 75728 -38494
rect 75180 -38560 75380 -38550
rect 75660 -38517 75728 -38500
rect 75660 -38551 75670 -38517
rect 75704 -38551 75728 -38517
rect 75660 -38570 75728 -38551
rect 75933 -38520 76011 -38492
rect 76765 -38498 76817 -38492
rect 75933 -38554 75942 -38520
rect 75976 -38554 76011 -38520
rect 75933 -38570 76011 -38554
rect 76204 -38519 76268 -38503
rect 76204 -38553 76217 -38519
rect 76251 -38553 76268 -38519
rect 76204 -38570 76268 -38553
rect 76483 -38519 76549 -38506
rect 76483 -38553 76492 -38519
rect 76526 -38553 76549 -38519
rect 75400 -38590 75480 -38580
rect 75660 -38583 75764 -38570
rect 75390 -38596 75410 -38590
rect 55380 -38680 55800 -38600
rect 73710 -38648 73723 -38596
rect 73840 -38648 75410 -38596
rect 75400 -38650 75410 -38648
rect 75470 -38596 75490 -38590
rect 75560 -38596 75630 -38590
rect 75470 -38610 75630 -38596
rect 75470 -38648 75580 -38610
rect 75470 -38650 75480 -38648
rect 75400 -38660 75480 -38650
rect 75560 -38650 75580 -38648
rect 75620 -38650 75630 -38610
rect 75560 -38670 75630 -38650
rect 75660 -38609 75673 -38583
rect 75660 -38643 75670 -38609
rect 75660 -38661 75673 -38643
rect 75751 -38661 75764 -38583
rect 55380 -38960 55460 -38680
rect 55720 -38960 55800 -38680
rect 75660 -38674 75764 -38661
rect 75840 -38582 75900 -38581
rect 75840 -38603 75902 -38582
rect 75840 -38637 75862 -38603
rect 75896 -38637 75902 -38603
rect 75840 -38663 75902 -38637
rect 75933 -38583 76037 -38570
rect 75933 -38661 75946 -38583
rect 76024 -38661 76037 -38583
rect 75660 -38698 75730 -38674
rect 72610 -38740 73050 -38730
rect 72610 -38920 72820 -38740
rect 73040 -38920 73050 -38740
rect 75660 -38732 75670 -38698
rect 75704 -38732 75730 -38698
rect 74210 -38760 75440 -38750
rect 75660 -38760 75730 -38732
rect 74210 -38840 74220 -38760
rect 74340 -38790 75440 -38760
rect 75840 -38790 75900 -38663
rect 75933 -38674 76037 -38661
rect 76102 -38583 76167 -38570
rect 76204 -38583 76323 -38570
rect 76483 -38583 76549 -38553
rect 76759 -38521 76817 -38498
rect 76759 -38555 76768 -38521
rect 76802 -38555 76817 -38521
rect 76759 -38583 76817 -38555
rect 76882 -38530 76920 -38440
rect 77060 -38530 77110 -38410
rect 76882 -38570 77110 -38530
rect 77220 -38570 77260 -38350
rect 76882 -38580 77260 -38570
rect 84700 -38480 84960 -38050
rect 85400 -38480 85660 -38050
rect 76167 -38661 76168 -38596
rect 76204 -38610 76232 -38583
rect 76204 -38644 76224 -38610
rect 76204 -38661 76232 -38644
rect 76310 -38661 76323 -38583
rect 76102 -38674 76167 -38661
rect 76204 -38674 76323 -38661
rect 76362 -38594 76453 -38583
rect 76362 -38600 76455 -38594
rect 76362 -38660 76380 -38600
rect 76440 -38660 76455 -38600
rect 76362 -38663 76455 -38660
rect 76483 -38596 76596 -38583
rect 76483 -38609 76505 -38596
rect 76483 -38643 76497 -38609
rect 76483 -38661 76505 -38643
rect 76583 -38661 76596 -38596
rect 76362 -38674 76453 -38663
rect 76483 -38674 76596 -38661
rect 76635 -38596 76726 -38583
rect 76635 -38674 76648 -38596
rect 75933 -38703 76011 -38674
rect 75933 -38737 75943 -38703
rect 75977 -38737 76011 -38703
rect 75933 -38778 76011 -38737
rect 76204 -38704 76268 -38674
rect 76370 -38680 76450 -38674
rect 76204 -38738 76215 -38704
rect 76249 -38738 76268 -38704
rect 76204 -38776 76268 -38738
rect 76483 -38703 76549 -38674
rect 76635 -38687 76726 -38674
rect 76759 -38596 76843 -38583
rect 76759 -38610 76791 -38596
rect 76759 -38644 76772 -38610
rect 76759 -38674 76791 -38644
rect 76759 -38687 76843 -38674
rect 76483 -38737 76492 -38703
rect 76526 -38737 76549 -38703
rect 76483 -38754 76549 -38737
rect 76759 -38703 76817 -38687
rect 84700 -38690 85660 -38480
rect 87880 -38390 88840 -38140
rect 87880 -38690 88150 -38390
rect 76759 -38737 76768 -38703
rect 76802 -38737 76817 -38703
rect 76759 -38756 76817 -38737
rect 74340 -38830 75900 -38790
rect 76204 -38810 76218 -38776
rect 76252 -38810 76268 -38776
rect 76204 -38823 76268 -38810
rect 76765 -38830 76817 -38756
rect 76850 -38790 79050 -38760
rect 76850 -38800 77170 -38790
rect 74340 -38840 75440 -38830
rect 74210 -38850 75440 -38840
rect 76850 -38880 76930 -38800
rect 72610 -38930 73050 -38920
rect 75500 -38915 76930 -38880
rect 55380 -39040 55800 -38960
rect 75500 -38949 75535 -38915
rect 75569 -38949 75627 -38915
rect 75661 -38949 75719 -38915
rect 75753 -38949 75811 -38915
rect 75845 -38949 75903 -38915
rect 75937 -38949 75995 -38915
rect 76029 -38949 76085 -38915
rect 76119 -38949 76177 -38915
rect 76211 -38949 76269 -38915
rect 76303 -38949 76361 -38915
rect 76395 -38949 76453 -38915
rect 76487 -38949 76545 -38915
rect 76579 -38949 76637 -38915
rect 76671 -38949 76729 -38915
rect 76763 -38949 76821 -38915
rect 76855 -38949 76930 -38915
rect 75500 -38980 76930 -38949
rect 76850 -39040 76930 -38980
rect 77040 -39040 77170 -38800
rect 77430 -39040 79050 -38790
rect 54090 -39138 54890 -39098
rect 54090 -39268 54150 -39138
rect 53510 -39320 53800 -39318
rect 35692 -39543 41100 -39500
rect 25860 -39560 41100 -39543
rect 53460 -39340 53800 -39320
rect 53460 -39540 53480 -39340
rect 53780 -39540 53800 -39340
rect 54080 -39398 54150 -39268
rect 54860 -39378 54890 -39138
rect 54850 -39398 54890 -39378
rect 54080 -39466 54880 -39398
rect 54079 -39472 54880 -39466
rect 54079 -39506 54091 -39472
rect 54867 -39498 54880 -39472
rect 54867 -39506 54879 -39498
rect 54079 -39512 54879 -39506
rect 53460 -39560 53800 -39540
rect 35900 -39600 41100 -39560
rect 53510 -39658 53800 -39560
rect 53002 -39820 53480 -39758
rect 53000 -39958 53480 -39820
rect 53510 -39768 53520 -39658
rect 53640 -39768 53800 -39658
rect 53510 -39888 53800 -39768
rect 53970 -39534 54040 -39518
rect 53970 -39572 53998 -39534
rect 54032 -39572 54040 -39534
rect 53970 -39768 54040 -39572
rect 54920 -39534 54990 -39518
rect 54920 -39572 54926 -39534
rect 54960 -39572 54990 -39534
rect 54079 -39600 54879 -39594
rect 54079 -39634 54091 -39600
rect 54867 -39634 54879 -39600
rect 54079 -39638 54879 -39634
rect 54079 -39640 54750 -39638
rect 54090 -39688 54750 -39640
rect 54740 -39718 54750 -39688
rect 54850 -39640 54879 -39638
rect 54850 -39708 54860 -39640
rect 54840 -39718 54860 -39708
rect 54750 -39728 54860 -39718
rect 54920 -39768 54990 -39572
rect 55430 -39618 55520 -39608
rect 55290 -39728 55390 -39718
rect 53970 -39798 55290 -39768
rect 55430 -39758 55520 -39688
rect 53970 -39808 55390 -39798
rect 54050 -39818 55380 -39808
rect 54050 -39828 54880 -39818
rect 54050 -39838 54091 -39828
rect 54079 -39862 54091 -39838
rect 54867 -39838 54880 -39828
rect 54867 -39862 54879 -39838
rect 54079 -39868 54879 -39862
rect 54920 -39878 54990 -39868
rect 53510 -39906 53630 -39888
rect 53510 -39938 53526 -39906
rect 53514 -39940 53526 -39938
rect 53614 -39938 53630 -39906
rect 53940 -39890 54038 -39878
rect 53940 -39898 53998 -39890
rect 53614 -39940 53626 -39938
rect 53514 -39946 53626 -39940
rect 35900 -40062 42200 -40000
rect 25862 -40081 42200 -40062
rect 25862 -40478 25884 -40081
rect 26998 -40478 27126 -40081
rect 28240 -40478 28368 -40081
rect 29482 -40478 29610 -40081
rect 30724 -40478 30852 -40081
rect 31966 -40478 32094 -40081
rect 33208 -40478 33336 -40081
rect 34450 -40478 34578 -40081
rect 35692 -40100 42200 -40081
rect 35692 -40478 36000 -40100
rect 25862 -40744 36000 -40478
rect 25862 -41141 25882 -40744
rect 26996 -41141 27124 -40744
rect 28238 -41141 28366 -40744
rect 29480 -41141 29608 -40744
rect 30722 -41141 30850 -40744
rect 31964 -41141 32092 -40744
rect 33206 -41141 33334 -40744
rect 34448 -41141 34576 -40744
rect 35690 -41100 36000 -40744
rect 42100 -41100 42200 -40100
rect 35690 -41141 42200 -41100
rect 25862 -41162 42200 -41141
rect 35900 -41200 42200 -41162
rect 35900 -41660 43200 -41600
rect 25860 -41679 43200 -41660
rect 25860 -42076 25882 -41679
rect 26996 -42076 27124 -41679
rect 28238 -42076 28366 -41679
rect 29480 -42076 29608 -41679
rect 30722 -42076 30850 -41679
rect 31964 -42076 32092 -41679
rect 33206 -42076 33334 -41679
rect 34448 -42076 34576 -41679
rect 35690 -41700 43200 -41679
rect 35690 -42076 36000 -41700
rect 25860 -42342 36000 -42076
rect 25860 -42739 25882 -42342
rect 26996 -42739 27124 -42342
rect 28238 -42739 28366 -42342
rect 29480 -42739 29608 -42342
rect 30722 -42739 30850 -42342
rect 31964 -42739 32092 -42342
rect 33206 -42739 33334 -42342
rect 34448 -42739 34576 -42342
rect 35690 -42700 36000 -42342
rect 43100 -42700 43200 -41700
rect 53000 -41708 53050 -39958
rect 53250 -39968 53480 -39958
rect 53250 -41318 53330 -39968
rect 53400 -39978 53480 -39968
rect 53400 -39990 53504 -39978
rect 53400 -40766 53464 -39990
rect 53498 -40766 53504 -39990
rect 53400 -40778 53504 -40766
rect 53636 -39988 53682 -39978
rect 53636 -39990 53760 -39988
rect 53636 -40766 53642 -39990
rect 53676 -40766 53760 -39990
rect 53940 -39998 53950 -39898
rect 54032 -39928 54038 -39890
rect 54020 -39940 54038 -39928
rect 54020 -39998 54030 -39940
rect 54079 -39956 54879 -39950
rect 54079 -39990 54091 -39956
rect 54867 -39990 54879 -39956
rect 54920 -39978 54990 -39968
rect 55320 -39968 55380 -39818
rect 54079 -39996 54879 -39990
rect 53940 -40018 54030 -39998
rect 54090 -40028 54870 -39996
rect 55320 -40002 55334 -39968
rect 55368 -40002 55380 -39968
rect 55320 -40008 55380 -40002
rect 53840 -40328 53920 -40318
rect 53840 -40438 53860 -40328
rect 53840 -40448 53920 -40438
rect 53840 -40640 53900 -40448
rect 54320 -40528 54510 -40028
rect 55440 -40038 55520 -39758
rect 55410 -40040 55520 -40038
rect 55284 -40048 55330 -40040
rect 55230 -40052 55330 -40048
rect 55230 -40058 55290 -40052
rect 55324 -40228 55330 -40052
rect 55230 -40238 55330 -40228
rect 55284 -40240 55330 -40238
rect 55372 -40048 55520 -40040
rect 55372 -40052 55430 -40048
rect 55372 -40228 55378 -40052
rect 55412 -40218 55430 -40052
rect 55510 -40218 55520 -40048
rect 55412 -40228 55520 -40218
rect 55372 -40240 55418 -40228
rect 55580 -40328 55720 -39040
rect 76850 -39041 79050 -39040
rect 72610 -39070 73050 -39060
rect 58776 -39270 59306 -39150
rect 58776 -39280 58966 -39270
rect 56146 -39380 57366 -39330
rect 55954 -39528 56046 -39516
rect 56146 -39528 56506 -39380
rect 55954 -39698 55960 -39528
rect 56040 -39698 56046 -39528
rect 55954 -39710 56046 -39698
rect 56120 -39558 56506 -39528
rect 56120 -39768 56190 -39558
rect 56390 -39630 56506 -39558
rect 57016 -39534 57366 -39380
rect 57586 -39430 58966 -39280
rect 59126 -39430 59306 -39270
rect 57586 -39450 59306 -39430
rect 59946 -39300 60386 -39200
rect 72610 -39250 72820 -39070
rect 73040 -39250 73050 -39070
rect 76850 -39075 77607 -39041
rect 77641 -39075 77699 -39041
rect 77733 -39075 77791 -39041
rect 77825 -39075 77883 -39041
rect 77917 -39075 77975 -39041
rect 78009 -39075 78067 -39041
rect 78101 -39075 78159 -39041
rect 78193 -39075 78251 -39041
rect 78285 -39075 78343 -39041
rect 78377 -39075 78435 -39041
rect 78469 -39075 78527 -39041
rect 78561 -39075 78619 -39041
rect 78653 -39075 78711 -39041
rect 78745 -39075 78803 -39041
rect 78837 -39075 78895 -39041
rect 78929 -39075 78987 -39041
rect 79021 -39075 79050 -39041
rect 76850 -39080 79050 -39075
rect 77578 -39106 79050 -39080
rect 73460 -39180 73480 -39120
rect 73580 -39130 77540 -39120
rect 73580 -39170 77430 -39130
rect 77520 -39170 77540 -39130
rect 78600 -39140 79050 -39106
rect 80730 -38790 88150 -38690
rect 80730 -38960 80890 -38790
rect 81070 -38960 81500 -38790
rect 81680 -38800 88150 -38790
rect 81680 -38960 82110 -38800
rect 80730 -38970 82110 -38960
rect 82290 -38810 83470 -38800
rect 82290 -38970 82760 -38810
rect 80730 -38980 82760 -38970
rect 82940 -38970 83470 -38810
rect 83650 -38970 84190 -38800
rect 84370 -38820 88150 -38800
rect 88590 -38820 88840 -38390
rect 84370 -38970 85840 -38820
rect 82940 -38980 85840 -38970
rect 80730 -38990 85840 -38980
rect 86020 -38830 88840 -38820
rect 86020 -38990 87280 -38830
rect 80730 -39000 87280 -38990
rect 87460 -39000 88840 -38830
rect 80730 -39091 88840 -39000
rect 80730 -39125 80767 -39091
rect 80801 -39125 80859 -39091
rect 80893 -39125 80951 -39091
rect 80985 -39125 81043 -39091
rect 81077 -39125 81135 -39091
rect 81169 -39125 81227 -39091
rect 81261 -39125 81319 -39091
rect 81353 -39125 81411 -39091
rect 81445 -39125 81503 -39091
rect 81537 -39125 81595 -39091
rect 81629 -39125 81687 -39091
rect 81721 -39125 81779 -39091
rect 81813 -39125 81871 -39091
rect 81905 -39125 81963 -39091
rect 81997 -39125 82055 -39091
rect 82089 -39125 82147 -39091
rect 82181 -39125 82239 -39091
rect 82273 -39125 82331 -39091
rect 82365 -39125 82423 -39091
rect 82457 -39125 82515 -39091
rect 82549 -39125 82607 -39091
rect 82641 -39125 82699 -39091
rect 82733 -39125 82791 -39091
rect 82825 -39125 82883 -39091
rect 82917 -39125 82975 -39091
rect 83009 -39125 83067 -39091
rect 83101 -39125 83159 -39091
rect 83193 -39125 83251 -39091
rect 83285 -39125 83343 -39091
rect 83377 -39125 83435 -39091
rect 83469 -39125 83527 -39091
rect 83561 -39125 83619 -39091
rect 83653 -39125 83711 -39091
rect 83745 -39125 83803 -39091
rect 83837 -39125 83895 -39091
rect 83929 -39125 83987 -39091
rect 84021 -39125 84079 -39091
rect 84113 -39125 84171 -39091
rect 84205 -39125 84263 -39091
rect 84297 -39125 84355 -39091
rect 84389 -39125 84447 -39091
rect 84481 -39125 84539 -39091
rect 84573 -39125 84631 -39091
rect 84665 -39125 84723 -39091
rect 84757 -39125 84815 -39091
rect 84849 -39125 84907 -39091
rect 84941 -39125 84999 -39091
rect 85033 -39125 85091 -39091
rect 85125 -39125 85183 -39091
rect 85217 -39125 85275 -39091
rect 85309 -39125 85367 -39091
rect 85401 -39125 85459 -39091
rect 85493 -39125 85551 -39091
rect 85585 -39125 85643 -39091
rect 85677 -39125 85735 -39091
rect 85769 -39125 85827 -39091
rect 85861 -39125 85919 -39091
rect 85953 -39125 86011 -39091
rect 86045 -39125 86103 -39091
rect 86137 -39125 86195 -39091
rect 86229 -39125 86287 -39091
rect 86321 -39125 86379 -39091
rect 86413 -39125 86471 -39091
rect 86505 -39125 86563 -39091
rect 86597 -39125 86655 -39091
rect 86689 -39125 86747 -39091
rect 86781 -39125 86839 -39091
rect 86873 -39125 86931 -39091
rect 86965 -39125 87023 -39091
rect 87057 -39125 87115 -39091
rect 87149 -39125 87207 -39091
rect 87241 -39125 87299 -39091
rect 87333 -39125 87391 -39091
rect 87425 -39125 87483 -39091
rect 87517 -39125 87575 -39091
rect 87609 -39125 87667 -39091
rect 87701 -39125 87759 -39091
rect 87793 -39125 87851 -39091
rect 87885 -39125 87943 -39091
rect 87977 -39125 88035 -39091
rect 88069 -39125 88127 -39091
rect 88161 -39125 88219 -39091
rect 88253 -39125 88311 -39091
rect 88345 -39125 88403 -39091
rect 88437 -39125 88495 -39091
rect 88529 -39125 88587 -39091
rect 88621 -39125 88679 -39091
rect 88713 -39125 88771 -39091
rect 88805 -39125 88840 -39091
rect 80730 -39160 88840 -39125
rect 73580 -39180 77540 -39170
rect 72610 -39260 73050 -39250
rect 73710 -39290 73730 -39230
rect 73830 -39270 77690 -39230
rect 82760 -39240 82910 -39230
rect 87170 -39240 87270 -39230
rect 80050 -39270 80460 -39240
rect 73830 -39280 77840 -39270
rect 73830 -39290 77780 -39280
rect 57586 -39480 58986 -39450
rect 59946 -39460 59956 -39300
rect 60166 -39460 60386 -39300
rect 77580 -39320 77780 -39290
rect 77820 -39320 77840 -39280
rect 77580 -39330 77840 -39320
rect 78570 -39320 78650 -39310
rect 73210 -39340 77510 -39330
rect 73210 -39400 73230 -39340
rect 73330 -39360 77510 -39340
rect 77870 -39350 77970 -39330
rect 77860 -39360 77900 -39350
rect 73330 -39390 77900 -39360
rect 77940 -39390 77970 -39350
rect 73330 -39400 77970 -39390
rect 73210 -39410 77970 -39400
rect 78140 -39340 78220 -39330
rect 78270 -39340 78350 -39330
rect 78140 -39400 78150 -39340
rect 78210 -39400 78220 -39340
rect 78140 -39410 78220 -39400
rect 78250 -39400 78280 -39340
rect 78340 -39350 78430 -39340
rect 78340 -39390 78370 -39350
rect 78410 -39390 78430 -39350
rect 78570 -39380 78580 -39320
rect 78640 -39380 78650 -39320
rect 78570 -39390 78650 -39380
rect 78790 -39330 78860 -39320
rect 78790 -39390 78800 -39330
rect 78340 -39400 78430 -39390
rect 78790 -39400 78860 -39390
rect 79060 -39340 79270 -39330
rect 78250 -39403 78410 -39400
rect 78270 -39410 78350 -39403
rect 57016 -39630 57368 -39534
rect 56390 -39670 57368 -39630
rect 56390 -39768 57126 -39670
rect 56120 -39774 57126 -39768
rect 56120 -39778 56750 -39774
rect 55880 -39818 55970 -39808
rect 55870 -39896 55880 -39850
rect 55970 -39896 55982 -39850
rect 55880 -39908 55970 -39898
rect 55000 -40338 55090 -40328
rect 55000 -40448 55090 -40438
rect 54710 -40528 54960 -40508
rect 53940 -40568 54960 -40528
rect 53940 -40572 54730 -40568
rect 53930 -40578 54730 -40572
rect 53930 -40612 53942 -40578
rect 54718 -40612 54730 -40578
rect 53930 -40618 54730 -40612
rect 53840 -40728 53858 -40640
rect 53892 -40728 53900 -40640
rect 53840 -40748 53900 -40728
rect 54762 -40638 54850 -40628
rect 54762 -40640 54770 -40638
rect 54762 -40728 54768 -40640
rect 54840 -40728 54850 -40638
rect 54762 -40740 54850 -40728
rect 54770 -40748 54850 -40740
rect 53636 -40778 53760 -40766
rect 53400 -40996 53480 -40778
rect 53514 -40816 53626 -40810
rect 53514 -40818 53526 -40816
rect 53510 -40850 53526 -40818
rect 53614 -40818 53626 -40816
rect 53614 -40850 53630 -40818
rect 53510 -40924 53630 -40850
rect 53510 -40958 53526 -40924
rect 53614 -40958 53630 -40924
rect 53680 -40838 53760 -40778
rect 53930 -40756 54730 -40750
rect 53930 -40790 53942 -40756
rect 54718 -40790 54730 -40756
rect 53930 -40796 54730 -40790
rect 53940 -40828 54720 -40796
rect 53920 -40838 54720 -40828
rect 53680 -40928 54720 -40838
rect 53514 -40964 53626 -40958
rect 53680 -40996 53760 -40928
rect 53920 -40938 54720 -40928
rect 53940 -40978 54720 -40938
rect 54900 -40968 54960 -40568
rect 55010 -40560 55090 -40448
rect 55540 -40338 55720 -40328
rect 55630 -40438 55720 -40338
rect 55130 -40474 55506 -40468
rect 55130 -40508 55142 -40474
rect 55494 -40508 55506 -40474
rect 55130 -40514 55506 -40508
rect 55010 -40594 55046 -40560
rect 55080 -40594 55090 -40560
rect 55010 -40608 55090 -40594
rect 55142 -40640 55494 -40514
rect 55540 -40560 55720 -40438
rect 55540 -40594 55556 -40560
rect 55590 -40594 55720 -40560
rect 55540 -40608 55720 -40594
rect 55780 -39940 55860 -39928
rect 55130 -40646 55506 -40640
rect 55130 -40680 55142 -40646
rect 55494 -40678 55506 -40646
rect 55494 -40680 55510 -40678
rect 55130 -40686 55510 -40680
rect 55140 -40698 55510 -40686
rect 55780 -40698 55820 -39940
rect 55140 -40716 55820 -40698
rect 55854 -40716 55860 -39940
rect 55140 -40728 55860 -40716
rect 55992 -39940 56038 -39928
rect 55992 -40716 55998 -39940
rect 56032 -39948 56038 -39940
rect 56120 -39948 56300 -39778
rect 57098 -39800 57126 -39774
rect 57356 -39800 57368 -39670
rect 57098 -39814 57368 -39800
rect 57096 -39845 57372 -39814
rect 57096 -39879 57125 -39845
rect 57159 -39879 57217 -39845
rect 57251 -39879 57309 -39845
rect 57343 -39879 57372 -39845
rect 57096 -39910 57372 -39879
rect 56032 -40306 56300 -39948
rect 56590 -40068 56660 -40058
rect 56660 -40134 57000 -40068
rect 57586 -40130 57706 -39480
rect 59946 -39490 60386 -39460
rect 77220 -39500 77230 -39440
rect 77310 -39500 77320 -39440
rect 77220 -39510 77320 -39500
rect 77400 -39460 77560 -39440
rect 77400 -39550 77420 -39460
rect 72610 -39560 73050 -39550
rect 57366 -40134 57706 -40130
rect 56660 -40138 57188 -40134
rect 56660 -40144 57190 -40138
rect 56660 -40194 57118 -40144
rect 57178 -40194 57190 -40144
rect 57314 -40140 57706 -40134
rect 57314 -40180 57326 -40140
rect 57366 -40180 57706 -40140
rect 57314 -40186 57706 -40180
rect 57366 -40190 57706 -40186
rect 58896 -39770 58986 -39750
rect 58896 -39830 58906 -39770
rect 58896 -40120 58926 -39830
rect 58966 -40120 58986 -39770
rect 59106 -39770 59516 -39760
rect 59106 -39830 59216 -39770
rect 59276 -39830 59326 -39770
rect 59386 -39830 59436 -39770
rect 59496 -39830 59516 -39770
rect 59106 -39847 59516 -39830
rect 59626 -39770 59706 -39730
rect 72610 -39740 72820 -39560
rect 73040 -39740 73050 -39560
rect 76900 -39570 77420 -39550
rect 76900 -39720 76920 -39570
rect 77060 -39580 77420 -39570
rect 77540 -39550 77560 -39460
rect 79060 -39510 79080 -39340
rect 79140 -39350 79270 -39340
rect 79250 -39510 79270 -39350
rect 79060 -39520 79270 -39510
rect 77540 -39580 79050 -39550
rect 77060 -39585 79050 -39580
rect 77060 -39619 77607 -39585
rect 77641 -39619 77699 -39585
rect 77733 -39619 77791 -39585
rect 77825 -39619 77883 -39585
rect 77917 -39619 77975 -39585
rect 78009 -39619 78067 -39585
rect 78101 -39619 78159 -39585
rect 78193 -39619 78251 -39585
rect 78285 -39619 78343 -39585
rect 78377 -39619 78435 -39585
rect 78469 -39619 78527 -39585
rect 78561 -39619 78619 -39585
rect 78653 -39619 78711 -39585
rect 78745 -39619 78803 -39585
rect 78837 -39619 78895 -39585
rect 78929 -39619 78987 -39585
rect 79021 -39619 79050 -39585
rect 80050 -39580 80080 -39270
rect 80430 -39330 80460 -39270
rect 80430 -39350 80660 -39330
rect 80430 -39510 80480 -39350
rect 80640 -39510 80660 -39350
rect 80430 -39530 80660 -39510
rect 82760 -39530 82780 -39240
rect 82820 -39270 82910 -39240
rect 82890 -39520 82910 -39270
rect 84220 -39250 84320 -39240
rect 83350 -39380 83790 -39370
rect 83350 -39394 83370 -39380
rect 83770 -39394 83790 -39380
rect 83350 -39434 83368 -39394
rect 83773 -39434 83790 -39394
rect 83350 -39450 83370 -39434
rect 83770 -39450 83790 -39434
rect 83350 -39460 83790 -39450
rect 82820 -39530 82910 -39520
rect 80430 -39580 80460 -39530
rect 82760 -39560 82910 -39530
rect 84220 -39540 84230 -39250
rect 84310 -39540 84320 -39250
rect 85700 -39260 85800 -39240
rect 84850 -39380 85260 -39370
rect 84850 -39450 84870 -39380
rect 85240 -39450 85260 -39380
rect 84850 -39460 85260 -39450
rect 84220 -39550 84320 -39540
rect 85700 -39550 85710 -39260
rect 85790 -39550 85800 -39260
rect 86310 -39380 86720 -39370
rect 86310 -39450 86320 -39380
rect 86710 -39450 86720 -39380
rect 86310 -39460 86720 -39450
rect 87170 -39510 87180 -39240
rect 87260 -39510 87270 -39240
rect 88640 -39250 88740 -39240
rect 87440 -39380 87770 -39370
rect 87440 -39450 87450 -39380
rect 87760 -39450 87770 -39380
rect 87440 -39460 87770 -39450
rect 87170 -39520 87270 -39510
rect 88640 -39540 88650 -39250
rect 88730 -39540 88740 -39250
rect 92000 -39550 95800 -38600
rect 85700 -39560 85800 -39550
rect 80050 -39610 80460 -39580
rect 91750 -39580 95800 -39550
rect 77060 -39660 79050 -39619
rect 80730 -39635 88840 -39600
rect 77060 -39720 77420 -39660
rect 76900 -39740 77420 -39720
rect 72610 -39750 73050 -39740
rect 59626 -39830 59636 -39770
rect 59626 -39840 59656 -39830
rect 59106 -39880 59125 -39847
rect 59113 -39881 59125 -39880
rect 59501 -39880 59516 -39847
rect 59501 -39881 59513 -39880
rect 59113 -39887 59513 -39881
rect 59546 -39890 59616 -39880
rect 59276 -39930 59356 -39920
rect 59276 -39949 59286 -39930
rect 59113 -39955 59286 -39949
rect 59346 -39949 59356 -39930
rect 59346 -39955 59513 -39949
rect 59113 -39989 59125 -39955
rect 59501 -39989 59513 -39955
rect 59606 -39950 59616 -39890
rect 59546 -39960 59616 -39950
rect 59113 -39990 59286 -39989
rect 59346 -39990 59513 -39989
rect 59016 -40000 59076 -39990
rect 59113 -39995 59513 -39990
rect 59276 -40000 59356 -39995
rect 59546 -40010 59616 -40000
rect 59016 -40070 59076 -40060
rect 59113 -40063 59513 -40057
rect 59113 -40097 59125 -40063
rect 59501 -40097 59513 -40063
rect 59606 -40070 59616 -40010
rect 59546 -40080 59616 -40070
rect 59113 -40100 59513 -40097
rect 59113 -40103 59516 -40100
rect 58896 -40130 58986 -40120
rect 58896 -40190 58906 -40130
rect 58966 -40190 58986 -40130
rect 58896 -40192 58986 -40190
rect 59116 -40120 59516 -40103
rect 59646 -40110 59656 -39840
rect 59116 -40180 59216 -40120
rect 59276 -40180 59336 -40120
rect 59396 -40180 59436 -40120
rect 59496 -40180 59516 -40120
rect 56660 -40198 57190 -40194
rect 56590 -40200 57190 -40198
rect 56590 -40204 57188 -40200
rect 56590 -40268 57000 -40204
rect 56032 -40318 56356 -40306
rect 56032 -40716 56280 -40318
rect 55992 -40728 56280 -40716
rect 55140 -40738 55200 -40728
rect 55450 -40758 55810 -40728
rect 55870 -40766 55982 -40760
rect 55870 -40800 55882 -40766
rect 55970 -40800 55982 -40766
rect 55870 -40806 55982 -40800
rect 55140 -40818 55200 -40808
rect 55024 -40848 55116 -40836
rect 55024 -40928 55030 -40848
rect 55110 -40928 55116 -40848
rect 55024 -40940 55116 -40928
rect 55734 -40848 55816 -40836
rect 55734 -40928 55740 -40848
rect 55810 -40928 55816 -40848
rect 55734 -40940 55816 -40928
rect 55880 -40838 55970 -40806
rect 55880 -40964 55970 -40928
rect 56060 -40948 56280 -40728
rect 56350 -40948 56356 -40318
rect 56480 -40388 56550 -40378
rect 56480 -40458 56550 -40448
rect 56590 -40487 56750 -40268
rect 58894 -40286 58988 -40192
rect 59116 -40200 59516 -40180
rect 59636 -40120 59656 -40110
rect 59696 -40120 59706 -39770
rect 77160 -39780 77270 -39770
rect 72610 -39840 73050 -39830
rect 59856 -39940 59976 -39930
rect 59856 -40030 59866 -39940
rect 59966 -40030 59976 -39940
rect 59856 -40040 59976 -40030
rect 60436 -40020 60446 -39920
rect 60526 -40020 60536 -39920
rect 60436 -40040 60536 -40020
rect 72610 -40020 72820 -39840
rect 73040 -40020 73050 -39840
rect 77160 -39850 77170 -39780
rect 77260 -39850 77270 -39780
rect 77400 -39780 77420 -39740
rect 77540 -39671 79050 -39660
rect 77540 -39705 77607 -39671
rect 77641 -39705 77699 -39671
rect 77733 -39705 77791 -39671
rect 77825 -39705 77883 -39671
rect 77917 -39705 77975 -39671
rect 78009 -39705 78067 -39671
rect 78101 -39705 79050 -39671
rect 77540 -39740 79050 -39705
rect 80050 -39680 80460 -39650
rect 77540 -39780 77560 -39740
rect 77400 -39800 77560 -39780
rect 78140 -39790 78220 -39770
rect 77160 -39860 77270 -39850
rect 77690 -39890 77960 -39880
rect 74210 -39950 74230 -39890
rect 74330 -39900 77960 -39890
rect 74330 -39920 77900 -39900
rect 74330 -39950 77700 -39920
rect 77860 -39940 77900 -39920
rect 77940 -39940 77960 -39900
rect 77860 -39950 77960 -39940
rect 77750 -39960 77830 -39950
rect 77750 -39980 77770 -39960
rect 72610 -40030 73050 -40020
rect 74710 -40040 74730 -39980
rect 74830 -40000 77770 -39980
rect 77810 -40000 77830 -39960
rect 74830 -40040 77830 -40000
rect 59636 -40130 59706 -40120
rect 59696 -40190 59706 -40130
rect 59636 -40210 59706 -40190
rect 59756 -40060 60536 -40040
rect 59756 -40100 59866 -40060
rect 60426 -40100 60536 -40060
rect 78140 -40080 78150 -39790
rect 78210 -40080 78220 -39790
rect 78140 -40100 78220 -40080
rect 80050 -40060 80080 -39680
rect 80430 -39780 80460 -39680
rect 80730 -39669 80767 -39635
rect 80801 -39669 80859 -39635
rect 80893 -39669 80951 -39635
rect 80985 -39669 81043 -39635
rect 81077 -39669 81135 -39635
rect 81169 -39669 81227 -39635
rect 81261 -39669 81319 -39635
rect 81353 -39669 81411 -39635
rect 81445 -39669 81503 -39635
rect 81537 -39669 81595 -39635
rect 81629 -39669 81687 -39635
rect 81721 -39669 81779 -39635
rect 81813 -39669 81871 -39635
rect 81905 -39669 81963 -39635
rect 81997 -39669 82055 -39635
rect 82089 -39669 82147 -39635
rect 82181 -39669 82239 -39635
rect 82273 -39669 82331 -39635
rect 82365 -39669 82423 -39635
rect 82457 -39669 82515 -39635
rect 82549 -39669 82607 -39635
rect 82641 -39669 82699 -39635
rect 82733 -39669 82791 -39635
rect 82825 -39669 82883 -39635
rect 82917 -39669 82975 -39635
rect 83009 -39669 83067 -39635
rect 83101 -39669 83159 -39635
rect 83193 -39669 83251 -39635
rect 83285 -39669 83343 -39635
rect 83377 -39669 83435 -39635
rect 83469 -39669 83527 -39635
rect 83561 -39669 83619 -39635
rect 83653 -39669 83711 -39635
rect 83745 -39669 83803 -39635
rect 83837 -39669 83895 -39635
rect 83929 -39669 83987 -39635
rect 84021 -39669 84079 -39635
rect 84113 -39669 84171 -39635
rect 84205 -39669 84263 -39635
rect 84297 -39669 84355 -39635
rect 84389 -39669 84447 -39635
rect 84481 -39669 84539 -39635
rect 84573 -39669 84631 -39635
rect 84665 -39669 84723 -39635
rect 84757 -39669 84815 -39635
rect 84849 -39669 84907 -39635
rect 84941 -39669 84999 -39635
rect 85033 -39669 85091 -39635
rect 85125 -39669 85183 -39635
rect 85217 -39669 85275 -39635
rect 85309 -39669 85367 -39635
rect 85401 -39669 85459 -39635
rect 85493 -39669 85551 -39635
rect 85585 -39669 85643 -39635
rect 85677 -39669 85735 -39635
rect 85769 -39669 85827 -39635
rect 85861 -39669 85919 -39635
rect 85953 -39669 86011 -39635
rect 86045 -39669 86103 -39635
rect 86137 -39669 86195 -39635
rect 86229 -39669 86287 -39635
rect 86321 -39669 86379 -39635
rect 86413 -39669 86471 -39635
rect 86505 -39669 86563 -39635
rect 86597 -39669 86655 -39635
rect 86689 -39669 86747 -39635
rect 86781 -39669 86839 -39635
rect 86873 -39669 86931 -39635
rect 86965 -39669 87023 -39635
rect 87057 -39669 87115 -39635
rect 87149 -39669 87207 -39635
rect 87241 -39669 87299 -39635
rect 87333 -39669 87391 -39635
rect 87425 -39669 87483 -39635
rect 87517 -39669 87575 -39635
rect 87609 -39669 87667 -39635
rect 87701 -39669 87759 -39635
rect 87793 -39669 87851 -39635
rect 87885 -39669 87943 -39635
rect 87977 -39669 88035 -39635
rect 88069 -39669 88127 -39635
rect 88161 -39669 88219 -39635
rect 88253 -39669 88311 -39635
rect 88345 -39669 88403 -39635
rect 88437 -39669 88495 -39635
rect 88529 -39669 88587 -39635
rect 88621 -39669 88679 -39635
rect 88713 -39669 88771 -39635
rect 88805 -39669 88840 -39635
rect 80730 -39711 88840 -39669
rect 80730 -39745 80817 -39711
rect 80851 -39745 80909 -39711
rect 80943 -39745 81001 -39711
rect 81035 -39730 88840 -39711
rect 81035 -39740 88500 -39730
rect 81035 -39745 82490 -39740
rect 80730 -39770 82490 -39745
rect 80730 -39780 81590 -39770
rect 80430 -39800 80660 -39780
rect 80430 -39960 80480 -39800
rect 80640 -39960 80660 -39800
rect 80430 -39980 80660 -39960
rect 81480 -39940 81590 -39780
rect 81760 -39910 82490 -39770
rect 82660 -39750 85160 -39740
rect 82660 -39830 83750 -39750
rect 82660 -39910 83150 -39830
rect 81760 -39940 83150 -39910
rect 81480 -39980 83150 -39940
rect 80430 -40060 80460 -39980
rect 80050 -40090 80460 -40060
rect 80510 -40050 81000 -40030
rect 59756 -40110 60536 -40100
rect 77400 -40110 77490 -40100
rect 59756 -40150 59826 -40110
rect 59066 -40240 59176 -40230
rect 58896 -40350 58986 -40286
rect 59066 -40310 59076 -40240
rect 59166 -40310 59176 -40240
rect 59066 -40312 59103 -40310
rect 59137 -40312 59176 -40310
rect 59066 -40320 59176 -40312
rect 59756 -40340 59766 -40150
rect 59806 -40340 59826 -40150
rect 59956 -40168 60046 -40140
rect 59946 -40174 60046 -40168
rect 60126 -40168 60336 -40140
rect 60126 -40174 60346 -40168
rect 59856 -40210 59916 -40200
rect 59946 -40208 59958 -40174
rect 60334 -40208 60346 -40174
rect 77400 -40180 77410 -40110
rect 77480 -40180 77490 -40110
rect 80510 -40120 80940 -40050
rect 79380 -40150 79710 -40120
rect 79380 -40180 79410 -40150
rect 77400 -40190 77490 -40180
rect 59946 -40214 60346 -40208
rect 60376 -40220 60446 -40210
rect 59856 -40290 59916 -40280
rect 59946 -40282 60346 -40276
rect 59946 -40316 59958 -40282
rect 60334 -40316 60346 -40282
rect 60376 -40290 60446 -40280
rect 77570 -40215 79410 -40180
rect 77570 -40249 77607 -40215
rect 77641 -40249 77699 -40215
rect 77733 -40249 77791 -40215
rect 77825 -40249 77883 -40215
rect 77917 -40249 77975 -40215
rect 78009 -40249 78067 -40215
rect 78101 -40220 79410 -40215
rect 78101 -40249 78250 -40220
rect 72610 -40300 73050 -40290
rect 59946 -40322 59976 -40316
rect 57098 -40358 57368 -40354
rect 57096 -40364 57372 -40358
rect 57096 -40450 57098 -40364
rect 56424 -40488 56470 -40487
rect 56060 -40960 56356 -40948
rect 56410 -40499 56470 -40488
rect 53400 -41008 53504 -40996
rect 53400 -41318 53464 -41008
rect 53250 -41708 53464 -41318
rect 53000 -41784 53464 -41708
rect 53498 -41784 53504 -41008
rect 53000 -41788 53504 -41784
rect 53458 -41796 53504 -41788
rect 53636 -41008 53760 -40996
rect 53636 -41784 53642 -41008
rect 53676 -41784 53760 -41008
rect 53930 -40984 54730 -40978
rect 53930 -41018 53942 -40984
rect 54718 -41018 54730 -40984
rect 53930 -41024 54730 -41018
rect 53830 -41046 53900 -41028
rect 53830 -41134 53858 -41046
rect 53892 -41134 53900 -41046
rect 53830 -41328 53900 -41134
rect 54760 -41046 54850 -41028
rect 54760 -41134 54768 -41046
rect 54802 -41048 54850 -41046
rect 54900 -41038 55200 -40968
rect 55870 -40970 55982 -40964
rect 55870 -41004 55882 -40970
rect 55970 -41004 55982 -40970
rect 55450 -41038 55810 -41008
rect 55870 -41010 55982 -41004
rect 56060 -41038 56300 -40960
rect 54900 -41042 55820 -41038
rect 56000 -41042 56300 -41038
rect 54900 -41048 55860 -41042
rect 54840 -41128 54850 -41048
rect 54802 -41134 54850 -41128
rect 54760 -41148 54850 -41134
rect 55130 -41054 55860 -41048
rect 55130 -41078 55820 -41054
rect 55130 -41096 55510 -41078
rect 55130 -41130 55142 -41096
rect 55494 -41098 55510 -41096
rect 55494 -41130 55506 -41098
rect 55130 -41136 55506 -41130
rect 53930 -41162 54730 -41156
rect 53930 -41196 53942 -41162
rect 54718 -41196 54730 -41162
rect 55020 -41182 55090 -41168
rect 53930 -41202 54730 -41196
rect 53940 -41208 54730 -41202
rect 54920 -41198 54980 -41188
rect 53940 -41248 54920 -41208
rect 53830 -41338 53920 -41328
rect 53830 -41448 53850 -41338
rect 53830 -41458 53920 -41448
rect 54320 -41748 54510 -41248
rect 54710 -41268 54920 -41248
rect 54910 -41278 54980 -41268
rect 55020 -41216 55046 -41182
rect 55080 -41216 55090 -41182
rect 55020 -41328 55090 -41216
rect 55142 -41262 55494 -41136
rect 55540 -41182 55620 -41168
rect 55540 -41216 55556 -41182
rect 55590 -41216 55620 -41182
rect 55130 -41268 55506 -41262
rect 55130 -41302 55142 -41268
rect 55494 -41302 55506 -41268
rect 55130 -41308 55506 -41302
rect 55000 -41338 55090 -41328
rect 55000 -41448 55090 -41438
rect 55540 -41328 55620 -41216
rect 55540 -41338 55630 -41328
rect 55630 -41438 55680 -41348
rect 55540 -41448 55680 -41438
rect 55274 -41538 55320 -41536
rect 55220 -41548 55320 -41538
rect 55220 -41724 55280 -41718
rect 55314 -41724 55320 -41548
rect 55220 -41728 55320 -41724
rect 55274 -41736 55320 -41728
rect 55362 -41548 55408 -41536
rect 55362 -41724 55368 -41548
rect 55402 -41558 55510 -41548
rect 55402 -41724 55410 -41558
rect 55362 -41728 55410 -41724
rect 55500 -41728 55510 -41558
rect 55362 -41736 55510 -41728
rect 55390 -41738 55510 -41736
rect 53636 -41788 53760 -41784
rect 53636 -41796 53682 -41788
rect 53940 -41808 54020 -41768
rect 54080 -41782 54860 -41748
rect 55311 -41774 55371 -41768
rect 53514 -41834 53626 -41828
rect 53514 -41838 53526 -41834
rect 53510 -41868 53526 -41838
rect 53614 -41838 53626 -41834
rect 53614 -41868 53630 -41838
rect 53510 -41928 53630 -41868
rect 53940 -41888 53950 -41808
rect 54010 -41838 54020 -41808
rect 54069 -41788 54869 -41782
rect 54069 -41822 54081 -41788
rect 54857 -41822 54869 -41788
rect 54069 -41828 54869 -41822
rect 54910 -41798 54980 -41788
rect 54010 -41850 54028 -41838
rect 54022 -41888 54028 -41850
rect 53940 -41900 54028 -41888
rect 53940 -41908 54020 -41900
rect 54910 -41908 54980 -41898
rect 55311 -41808 55324 -41774
rect 55358 -41808 55371 -41774
rect 54070 -41910 54870 -41908
rect 54069 -41916 54870 -41910
rect 54069 -41938 54081 -41916
rect 54041 -41950 54081 -41938
rect 54857 -41918 54870 -41916
rect 54857 -41950 54880 -41918
rect 55311 -41948 55371 -41808
rect 54041 -41958 54880 -41950
rect 55240 -41958 55371 -41948
rect 54041 -41968 55240 -41958
rect 53510 -42058 53630 -42048
rect 53961 -42008 55240 -41968
rect 53961 -42206 54031 -42008
rect 54730 -42068 54860 -42058
rect 54730 -42088 54740 -42068
rect 54080 -42138 54740 -42088
rect 54069 -42144 54740 -42138
rect 54850 -42138 54860 -42068
rect 54850 -42144 54869 -42138
rect 54069 -42178 54081 -42144
rect 54857 -42178 54869 -42144
rect 54069 -42184 54869 -42178
rect 54911 -42194 54981 -42008
rect 55370 -42008 55371 -41958
rect 55240 -42028 55370 -42018
rect 55410 -42048 55510 -41738
rect 55410 -42158 55510 -42138
rect 55570 -42068 55680 -41448
rect 55780 -41830 55820 -41078
rect 55854 -41830 55860 -41054
rect 55780 -41838 55860 -41830
rect 55814 -41842 55860 -41838
rect 55992 -41054 56300 -41042
rect 55992 -41830 55998 -41054
rect 56032 -41828 56300 -41054
rect 56410 -41098 56430 -40499
rect 56380 -41275 56430 -41098
rect 56464 -41275 56470 -40499
rect 56380 -41287 56470 -41275
rect 56552 -40499 56750 -40487
rect 56552 -41275 56558 -40499
rect 56592 -40638 56750 -40499
rect 57066 -40480 57098 -40450
rect 57368 -40450 57372 -40364
rect 58896 -40359 59076 -40350
rect 58896 -40360 59084 -40359
rect 59156 -40360 59202 -40359
rect 57368 -40480 57396 -40450
rect 57066 -40610 57086 -40480
rect 57376 -40610 57396 -40480
rect 56592 -41275 56610 -40638
rect 57066 -40640 57396 -40610
rect 56860 -40790 57060 -40778
rect 56860 -40818 57236 -40790
rect 56860 -40948 56900 -40818
rect 57020 -40948 57236 -40818
rect 56860 -40988 57236 -40948
rect 57036 -40990 57236 -40988
rect 58556 -40880 58756 -40860
rect 58556 -41040 58576 -40880
rect 58736 -41040 58756 -40880
rect 58556 -41060 58756 -41040
rect 56552 -41278 56610 -41275
rect 57036 -41140 57446 -41130
rect 56552 -41287 56598 -41278
rect 57036 -41280 57056 -41140
rect 57416 -41280 57446 -41140
rect 56380 -41558 56440 -41287
rect 57036 -41300 57098 -41280
rect 56480 -41328 56550 -41318
rect 56480 -41398 56550 -41388
rect 57096 -41414 57098 -41334
rect 57368 -41300 57446 -41280
rect 57368 -41414 57372 -41334
rect 57096 -41430 57372 -41414
rect 58896 -41490 58926 -40360
rect 58966 -40371 59086 -40360
rect 58966 -40747 59044 -40371
rect 59078 -40747 59086 -40371
rect 58966 -40770 59086 -40747
rect 59156 -40371 59256 -40360
rect 59756 -40370 59826 -40340
rect 59966 -40352 59976 -40322
rect 60316 -40322 60346 -40316
rect 61036 -40320 61466 -40310
rect 60316 -40352 60326 -40322
rect 59966 -40360 60326 -40352
rect 59156 -40747 59162 -40371
rect 59196 -40440 59256 -40371
rect 59236 -40520 59256 -40440
rect 59196 -40640 59256 -40520
rect 59236 -40720 59256 -40640
rect 59196 -40747 59256 -40720
rect 59156 -40760 59256 -40747
rect 58966 -41080 59036 -40770
rect 59066 -40806 59176 -40800
rect 59066 -40810 59103 -40806
rect 59137 -40810 59176 -40806
rect 59066 -40880 59076 -40810
rect 59166 -40880 59176 -40810
rect 59066 -40890 59176 -40880
rect 59206 -40960 59256 -40760
rect 59376 -40390 59826 -40370
rect 59376 -40430 59476 -40390
rect 59656 -40430 59826 -40390
rect 59376 -40440 59826 -40430
rect 59376 -40490 59436 -40440
rect 59376 -40850 59386 -40490
rect 59426 -40850 59436 -40490
rect 59526 -40498 59576 -40470
rect 59526 -40532 59546 -40498
rect 59636 -40530 59706 -40470
rect 59580 -40532 59706 -40530
rect 59526 -40540 59706 -40532
rect 59476 -40582 59546 -40570
rect 59476 -40650 59502 -40582
rect 59476 -40758 59502 -40720
rect 59536 -40758 59546 -40582
rect 59476 -40770 59546 -40758
rect 59576 -40582 59636 -40570
rect 59576 -40590 59590 -40582
rect 59624 -40590 59636 -40582
rect 59576 -40770 59636 -40760
rect 59534 -40808 59592 -40802
rect 59534 -40810 59546 -40808
rect 59066 -40970 59176 -40960
rect 59066 -41040 59076 -40970
rect 59166 -41040 59176 -40970
rect 59066 -41042 59103 -41040
rect 59137 -41042 59176 -41040
rect 59066 -41050 59176 -41042
rect 59206 -40970 59266 -40960
rect 59206 -41050 59266 -41040
rect 59376 -41000 59436 -40850
rect 59516 -40842 59546 -40810
rect 59580 -40810 59592 -40808
rect 59666 -40810 59706 -40540
rect 59580 -40842 59706 -40810
rect 59516 -40880 59706 -40842
rect 59746 -40498 59936 -40470
rect 59746 -40532 59862 -40498
rect 59896 -40532 59936 -40498
rect 59746 -40540 59936 -40532
rect 61036 -40500 61206 -40320
rect 61346 -40500 61466 -40320
rect 72610 -40480 72820 -40300
rect 73040 -40480 73050 -40300
rect 77570 -40291 78250 -40249
rect 77570 -40325 77607 -40291
rect 77641 -40325 77699 -40291
rect 77733 -40325 77791 -40291
rect 77825 -40325 77883 -40291
rect 77917 -40325 77975 -40291
rect 78009 -40325 78250 -40291
rect 77570 -40330 78250 -40325
rect 78360 -40330 78560 -40220
rect 78670 -40330 78800 -40220
rect 78910 -40330 79060 -40220
rect 79170 -40330 79410 -40220
rect 77570 -40360 79410 -40330
rect 79380 -40390 79410 -40360
rect 79680 -40390 79710 -40150
rect 79770 -40130 80940 -40120
rect 79770 -40370 79780 -40130
rect 79910 -40160 80940 -40130
rect 80990 -40160 81000 -40050
rect 79910 -40180 81000 -40160
rect 83000 -40180 83150 -39980
rect 83510 -39920 83750 -39830
rect 83920 -39910 85160 -39750
rect 85330 -39750 87390 -39740
rect 85330 -39910 86320 -39750
rect 83920 -39920 86320 -39910
rect 86490 -39910 87390 -39750
rect 87560 -39900 88500 -39740
rect 88670 -39900 88840 -39730
rect 87560 -39910 88840 -39900
rect 86490 -39920 88840 -39910
rect 83510 -39980 88840 -39920
rect 83510 -40180 83640 -39980
rect 79910 -40370 80690 -40180
rect 79770 -40380 80690 -40370
rect 80730 -40250 81600 -40220
rect 80730 -40255 81140 -40250
rect 80730 -40289 80817 -40255
rect 80851 -40289 80909 -40255
rect 80943 -40289 81001 -40255
rect 81035 -40289 81140 -40255
rect 80730 -40330 81140 -40289
rect 79380 -40410 79710 -40390
rect 72610 -40490 73050 -40480
rect 61036 -40540 61466 -40500
rect 80730 -40500 80850 -40330
rect 81020 -40500 81140 -40330
rect 80730 -40510 81140 -40500
rect 81570 -40510 81600 -40250
rect 83000 -40290 83640 -40180
rect 87520 -40240 88840 -39980
rect 91750 -39960 91780 -39580
rect 92130 -39960 95800 -39580
rect 91750 -39990 95800 -39960
rect 77980 -40530 78420 -40510
rect 77440 -40540 77530 -40530
rect 59746 -40800 59776 -40540
rect 60286 -40550 60476 -40540
rect 59806 -40582 59866 -40570
rect 59806 -40600 59818 -40582
rect 59852 -40600 59866 -40582
rect 59806 -40758 59818 -40740
rect 59852 -40758 59866 -40740
rect 59806 -40770 59866 -40758
rect 59900 -40580 60016 -40570
rect 59900 -40582 59916 -40580
rect 59900 -40758 59906 -40582
rect 59900 -40760 59916 -40758
rect 60006 -40760 60016 -40580
rect 60286 -40690 60306 -40550
rect 60456 -40690 60476 -40550
rect 61176 -40600 61386 -40580
rect 60286 -40700 60476 -40690
rect 61026 -40620 61136 -40610
rect 59900 -40770 60016 -40760
rect 60076 -40757 60196 -40720
rect 60076 -40791 60127 -40757
rect 60161 -40791 60196 -40757
rect 59746 -40808 59926 -40800
rect 59746 -40810 59862 -40808
rect 59896 -40810 59926 -40808
rect 59746 -40880 59826 -40810
rect 59916 -40880 59926 -40810
rect 59746 -40890 59926 -40880
rect 60076 -40849 60196 -40791
rect 60336 -40760 60446 -40700
rect 60336 -40800 60366 -40760
rect 60406 -40800 60446 -40760
rect 60636 -40757 60816 -40720
rect 60636 -40791 60671 -40757
rect 60705 -40791 60747 -40757
rect 60781 -40791 60816 -40757
rect 60076 -40880 60127 -40849
rect 60161 -40880 60196 -40849
rect 59736 -40970 59936 -40960
rect 58966 -41101 59086 -41080
rect 58966 -41477 59044 -41101
rect 59078 -41477 59086 -41101
rect 58966 -41490 59086 -41477
rect 59156 -41090 59202 -41089
rect 59156 -41101 59236 -41090
rect 59156 -41477 59162 -41101
rect 59196 -41130 59236 -41101
rect 59226 -41210 59236 -41130
rect 59196 -41360 59236 -41210
rect 59226 -41440 59236 -41360
rect 59196 -41477 59236 -41440
rect 59376 -41370 59386 -41000
rect 59426 -41370 59436 -41000
rect 59516 -41011 59706 -40970
rect 59516 -41045 59545 -41011
rect 59579 -41045 59706 -41011
rect 59516 -41050 59706 -41045
rect 59533 -41051 59591 -41050
rect 59466 -41095 59546 -41080
rect 59586 -41083 59646 -41080
rect 59466 -41130 59501 -41095
rect 59466 -41271 59501 -41210
rect 59535 -41271 59546 -41095
rect 59466 -41280 59546 -41271
rect 59583 -41095 59646 -41083
rect 59583 -41110 59589 -41095
rect 59623 -41110 59646 -41095
rect 59583 -41250 59586 -41110
rect 59583 -41271 59589 -41250
rect 59623 -41271 59646 -41250
rect 59583 -41280 59646 -41271
rect 59495 -41283 59541 -41280
rect 59583 -41283 59629 -41280
rect 59533 -41320 59591 -41315
rect 59676 -41320 59706 -41050
rect 59376 -41410 59436 -41370
rect 59506 -41380 59516 -41320
rect 59596 -41380 59706 -41320
rect 59736 -41040 59826 -40970
rect 59926 -41040 59936 -40970
rect 59736 -41045 59861 -41040
rect 59895 -41045 59936 -41040
rect 59736 -41050 59936 -41045
rect 60076 -41040 60096 -40880
rect 60176 -41040 60196 -40880
rect 59736 -41320 59766 -41050
rect 59849 -41051 59907 -41050
rect 60076 -41067 60127 -41040
rect 60161 -41067 60196 -41040
rect 59796 -41083 59856 -41080
rect 59796 -41090 59857 -41083
rect 59856 -41270 59857 -41090
rect 59796 -41271 59817 -41270
rect 59851 -41271 59857 -41270
rect 59796 -41280 59857 -41271
rect 59811 -41283 59857 -41280
rect 59899 -41090 59945 -41083
rect 59899 -41095 59916 -41090
rect 59899 -41271 59905 -41095
rect 59899 -41280 59916 -41271
rect 60006 -41280 60016 -41090
rect 60076 -41125 60196 -41067
rect 60346 -40850 60426 -40800
rect 60346 -40890 60366 -40850
rect 60406 -40890 60426 -40850
rect 60346 -40940 60426 -40890
rect 60346 -40980 60366 -40940
rect 60406 -40980 60426 -40940
rect 60346 -41020 60426 -40980
rect 60346 -41060 60366 -41020
rect 60406 -41060 60426 -41020
rect 60346 -41070 60426 -41060
rect 60636 -40849 60816 -40791
rect 60636 -40883 60671 -40849
rect 60705 -40883 60747 -40849
rect 60781 -40883 60816 -40849
rect 60636 -40941 60816 -40883
rect 60636 -40975 60671 -40941
rect 60705 -40975 60747 -40941
rect 60781 -40975 60816 -40941
rect 60636 -41033 60816 -40975
rect 60636 -41067 60671 -41033
rect 60705 -41067 60747 -41033
rect 60781 -41067 60816 -41033
rect 60076 -41159 60127 -41125
rect 60161 -41159 60196 -41125
rect 60076 -41190 60196 -41159
rect 60276 -41110 60546 -41100
rect 60276 -41125 60476 -41110
rect 60276 -41159 60297 -41125
rect 60331 -41159 60369 -41125
rect 60405 -41159 60449 -41125
rect 60276 -41170 60476 -41159
rect 60536 -41170 60546 -41110
rect 60276 -41180 60546 -41170
rect 60636 -41125 60816 -41067
rect 61026 -40730 61036 -40620
rect 61126 -40730 61136 -40620
rect 61176 -40680 61196 -40600
rect 61366 -40680 61386 -40600
rect 77440 -40610 77450 -40540
rect 77520 -40610 77530 -40540
rect 77980 -40570 78000 -40530
rect 78040 -40570 78420 -40530
rect 80730 -40540 81600 -40510
rect 77440 -40620 77530 -40610
rect 77770 -40630 77780 -40570
rect 77840 -40630 77850 -40570
rect 77770 -40640 77850 -40630
rect 77980 -40620 78420 -40570
rect 61176 -40700 61386 -40680
rect 72610 -40660 73050 -40650
rect 61026 -40760 61136 -40730
rect 61026 -40800 61046 -40760
rect 61086 -40800 61136 -40760
rect 61026 -40850 61136 -40800
rect 61026 -40890 61046 -40850
rect 61086 -40890 61136 -40850
rect 61026 -40940 61136 -40890
rect 61026 -40980 61046 -40940
rect 61086 -40980 61136 -40940
rect 61026 -41020 61136 -40980
rect 61026 -41060 61046 -41020
rect 61086 -41060 61136 -41020
rect 61026 -41080 61136 -41060
rect 61256 -40757 61366 -40700
rect 61256 -40791 61291 -40757
rect 61325 -40791 61366 -40757
rect 61256 -40849 61366 -40791
rect 61256 -40850 61291 -40849
rect 61325 -40850 61366 -40849
rect 72610 -40840 72820 -40660
rect 73040 -40840 73050 -40660
rect 77980 -40660 78000 -40620
rect 78040 -40650 78420 -40620
rect 78040 -40660 78310 -40650
rect 77380 -40700 77540 -40680
rect 77380 -40800 77400 -40700
rect 72610 -40850 73050 -40840
rect 76900 -40820 77400 -40800
rect 77520 -40800 77540 -40700
rect 77980 -40700 78310 -40660
rect 77980 -40740 78000 -40700
rect 78040 -40740 78310 -40700
rect 77980 -40760 78310 -40740
rect 78410 -40760 78420 -40650
rect 77980 -40770 78420 -40760
rect 87520 -40590 87830 -40240
rect 88190 -40270 88840 -40240
rect 88190 -40590 88480 -40270
rect 77520 -40820 78590 -40800
rect 61256 -41060 61276 -40850
rect 61356 -41060 61366 -40850
rect 76900 -40960 76920 -40820
rect 77060 -40835 78590 -40820
rect 77060 -40869 77607 -40835
rect 77641 -40869 77699 -40835
rect 77733 -40869 77791 -40835
rect 77825 -40869 77883 -40835
rect 77917 -40869 77975 -40835
rect 78009 -40869 78590 -40835
rect 77060 -40911 78590 -40869
rect 77060 -40945 77607 -40911
rect 77641 -40945 77699 -40911
rect 77733 -40945 77791 -40911
rect 77825 -40945 77883 -40911
rect 77917 -40945 77975 -40911
rect 78009 -40945 78067 -40911
rect 78101 -40945 78159 -40911
rect 78193 -40945 78251 -40911
rect 78285 -40945 78343 -40911
rect 78377 -40945 78435 -40911
rect 78469 -40945 78527 -40911
rect 78561 -40945 78590 -40911
rect 77060 -40950 78590 -40945
rect 77060 -40960 77400 -40950
rect 76900 -40980 77400 -40960
rect 61256 -41067 61291 -41060
rect 61325 -41067 61366 -41060
rect 60636 -41159 60671 -41125
rect 60705 -41159 60747 -41125
rect 60781 -41159 60816 -41125
rect 60636 -41240 60816 -41159
rect 60966 -41124 61177 -41110
rect 60966 -41125 61129 -41124
rect 60966 -41159 60980 -41125
rect 61015 -41159 61053 -41125
rect 61088 -41158 61129 -41125
rect 61164 -41158 61177 -41124
rect 61088 -41159 61177 -41158
rect 60966 -41190 61177 -41159
rect 61256 -41125 61366 -41067
rect 61256 -41159 61291 -41125
rect 61325 -41159 61366 -41125
rect 61256 -41190 61366 -41159
rect 72610 -41060 73050 -41050
rect 60466 -41250 60546 -41240
rect 59899 -41283 59945 -41280
rect 60466 -41310 60476 -41250
rect 60536 -41310 60546 -41250
rect 59849 -41320 59907 -41315
rect 60466 -41320 60546 -41310
rect 60606 -41250 60826 -41240
rect 60606 -41310 60616 -41250
rect 60736 -41310 60756 -41250
rect 60816 -41310 60826 -41250
rect 60606 -41320 60826 -41310
rect 60886 -41250 60966 -41240
rect 60886 -41310 60896 -41250
rect 60956 -41310 60966 -41250
rect 60886 -41320 60966 -41310
rect 59736 -41321 59926 -41320
rect 59736 -41355 59861 -41321
rect 59895 -41355 59926 -41321
rect 59736 -41380 59926 -41355
rect 60636 -41370 60816 -41320
rect 59376 -41420 59826 -41410
rect 59376 -41460 59476 -41420
rect 59646 -41460 59826 -41420
rect 59376 -41470 59826 -41460
rect 59156 -41490 59236 -41477
rect 58896 -41500 59086 -41490
rect 56380 -41568 57000 -41558
rect 57356 -41564 57676 -41550
rect 56440 -41574 57000 -41568
rect 57314 -41570 57676 -41564
rect 56440 -41594 57178 -41574
rect 56440 -41644 57118 -41594
rect 57168 -41644 57178 -41594
rect 57314 -41610 57326 -41570
rect 57376 -41610 57676 -41570
rect 57314 -41616 57676 -41610
rect 57356 -41630 57676 -41616
rect 56440 -41654 57178 -41644
rect 56440 -41688 57000 -41654
rect 57112 -41656 57174 -41654
rect 56380 -41758 57000 -41688
rect 56032 -41830 56038 -41828
rect 55992 -41842 56038 -41830
rect 55880 -41874 55970 -41868
rect 55870 -41878 55982 -41874
rect 55870 -41920 55880 -41878
rect 55970 -41920 55982 -41878
rect 55880 -41968 55970 -41958
rect 56120 -41998 56300 -41828
rect 57096 -41909 57372 -41878
rect 57096 -41943 57125 -41909
rect 57159 -41943 57217 -41909
rect 57251 -41943 57309 -41909
rect 57343 -41920 57372 -41909
rect 57343 -41943 57376 -41920
rect 57096 -41980 57376 -41943
rect 57066 -41990 57376 -41980
rect 56426 -41998 57376 -41990
rect 56120 -42008 57376 -41998
rect 56014 -42058 56086 -42046
rect 55570 -42178 55830 -42068
rect 53961 -42244 53988 -42206
rect 54022 -42244 54031 -42206
rect 53961 -42258 54031 -42244
rect 54910 -42206 54981 -42194
rect 54910 -42244 54916 -42206
rect 54950 -42244 54981 -42206
rect 54910 -42256 54981 -42244
rect 54911 -42258 54981 -42256
rect 55220 -42218 55330 -42208
rect 54069 -42272 54869 -42266
rect 54069 -42306 54081 -42272
rect 54857 -42278 54869 -42272
rect 54857 -42306 54880 -42278
rect 54069 -42312 54880 -42306
rect 54090 -42388 54880 -42312
rect 55330 -42318 55380 -42218
rect 55330 -42328 55480 -42318
rect 55220 -42338 55480 -42328
rect 55280 -42352 55480 -42338
rect 55280 -42358 55488 -42352
rect 55280 -42378 55300 -42358
rect 54090 -42488 54150 -42388
rect 54840 -42488 54880 -42388
rect 55288 -42392 55300 -42378
rect 55476 -42392 55488 -42358
rect 55530 -42378 55610 -42368
rect 55288 -42398 55488 -42392
rect 55520 -42402 55530 -42390
rect 55520 -42436 55526 -42402
rect 55288 -42446 55488 -42440
rect 55288 -42480 55300 -42446
rect 55476 -42480 55488 -42446
rect 55520 -42448 55530 -42436
rect 55530 -42478 55610 -42468
rect 55288 -42486 55488 -42480
rect 54090 -42508 54140 -42488
rect 35690 -42739 43200 -42700
rect 25860 -42760 43200 -42739
rect 35900 -42800 43200 -42760
rect 54100 -42748 54140 -42508
rect 54850 -42748 54880 -42488
rect 55300 -42528 55470 -42486
rect 55300 -42668 55320 -42528
rect 55470 -42614 55482 -42542
rect 55300 -42678 55470 -42668
rect 54100 -42788 54880 -42748
rect 55710 -42998 55830 -42178
rect 56014 -42208 56020 -42058
rect 56080 -42208 56086 -42058
rect 56014 -42220 56086 -42208
rect 56120 -42208 56170 -42008
rect 56390 -42060 57376 -42008
rect 56390 -42068 57156 -42060
rect 56390 -42208 56654 -42068
rect 56120 -42258 56654 -42208
rect 56306 -42286 56654 -42258
rect 56998 -42220 57156 -42068
rect 57316 -42220 57376 -42060
rect 56998 -42286 57376 -42220
rect 56306 -42700 57376 -42286
rect 57556 -42410 57676 -41630
rect 58896 -41660 58986 -41500
rect 59756 -41520 59826 -41470
rect 59066 -41536 59176 -41530
rect 59066 -41540 59103 -41536
rect 59137 -41540 59176 -41536
rect 59066 -41600 59076 -41540
rect 59166 -41600 59176 -41540
rect 59066 -41610 59176 -41600
rect 58896 -42030 58926 -41660
rect 58966 -42030 58986 -41730
rect 59116 -41660 59506 -41640
rect 59116 -41730 59146 -41660
rect 59226 -41730 59276 -41660
rect 59356 -41730 59396 -41660
rect 59476 -41730 59506 -41660
rect 59116 -41748 59506 -41730
rect 59646 -41660 59716 -41640
rect 59706 -41720 59716 -41660
rect 59646 -41730 59716 -41720
rect 59113 -41754 59513 -41748
rect 59113 -41788 59125 -41754
rect 59501 -41788 59513 -41754
rect 59113 -41794 59513 -41788
rect 59546 -41800 59616 -41790
rect 59246 -41856 59256 -41830
rect 59113 -41862 59256 -41856
rect 59366 -41856 59376 -41830
rect 59366 -41862 59513 -41856
rect 59016 -41900 59076 -41880
rect 59113 -41896 59125 -41862
rect 59501 -41896 59513 -41862
rect 59606 -41860 59616 -41800
rect 59546 -41870 59616 -41860
rect 59113 -41902 59513 -41896
rect 59016 -41990 59076 -41960
rect 59113 -41970 59513 -41964
rect 59113 -42004 59125 -41970
rect 59501 -42004 59513 -41970
rect 59113 -42010 59513 -42004
rect 58896 -42100 58906 -42030
rect 58896 -42120 58986 -42100
rect 59116 -42030 59516 -42010
rect 59116 -42100 59146 -42030
rect 59226 -42100 59276 -42030
rect 59356 -42100 59396 -42030
rect 59476 -42100 59516 -42030
rect 59116 -42120 59516 -42100
rect 59646 -42030 59656 -41730
rect 59706 -42030 59716 -41730
rect 59756 -41700 59766 -41520
rect 59806 -41700 59826 -41520
rect 59956 -41520 60336 -41510
rect 59956 -41534 59966 -41520
rect 59946 -41540 59966 -41534
rect 60326 -41534 60336 -41520
rect 60326 -41540 60346 -41534
rect 59856 -41580 59916 -41570
rect 59946 -41574 59958 -41540
rect 60334 -41574 60346 -41540
rect 61056 -41540 61176 -41190
rect 72610 -41240 72820 -41060
rect 73040 -41240 73050 -41060
rect 77380 -41070 77400 -40980
rect 77520 -40980 78590 -40950
rect 80050 -40910 80460 -40880
rect 87520 -40890 88480 -40590
rect 92000 -40800 95800 -39990
rect 77520 -41070 77540 -40980
rect 77380 -41090 77540 -41070
rect 78550 -41030 78790 -41020
rect 78050 -41090 78130 -41080
rect 77770 -41140 77850 -41130
rect 72610 -41250 73050 -41240
rect 77440 -41160 77540 -41150
rect 77440 -41240 77450 -41160
rect 77530 -41240 77540 -41160
rect 77770 -41200 77780 -41140
rect 77840 -41200 77850 -41140
rect 78050 -41180 78060 -41090
rect 78120 -41180 78130 -41090
rect 78550 -41100 78570 -41030
rect 78640 -41100 78670 -41030
rect 78350 -41130 78410 -41120
rect 78050 -41190 78130 -41180
rect 78170 -41140 78300 -41130
rect 77770 -41210 77850 -41200
rect 77440 -41250 77540 -41240
rect 78170 -41240 78180 -41140
rect 78290 -41240 78300 -41140
rect 78350 -41200 78410 -41190
rect 78550 -41170 78670 -41100
rect 78170 -41250 78300 -41240
rect 78550 -41240 78570 -41170
rect 78640 -41240 78670 -41170
rect 78550 -41310 78670 -41240
rect 78550 -41380 78570 -41310
rect 78640 -41380 78670 -41310
rect 78780 -41380 78790 -41030
rect 80050 -41290 80080 -40910
rect 80430 -41000 80460 -40910
rect 80430 -41200 80660 -41000
rect 80430 -41290 80460 -41200
rect 80050 -41320 80460 -41290
rect 78550 -41390 78790 -41380
rect 79380 -41380 79710 -41350
rect 79380 -41420 79410 -41380
rect 77570 -41455 79410 -41420
rect 77570 -41489 77607 -41455
rect 77641 -41489 77699 -41455
rect 77733 -41489 77791 -41455
rect 77825 -41489 77883 -41455
rect 77917 -41489 77975 -41455
rect 78009 -41489 78067 -41455
rect 78101 -41489 78159 -41455
rect 78193 -41489 78251 -41455
rect 78285 -41489 78343 -41455
rect 78377 -41489 78435 -41455
rect 78469 -41489 78527 -41455
rect 78561 -41460 79410 -41455
rect 78561 -41489 78630 -41460
rect 59946 -41580 59966 -41574
rect 60326 -41580 60346 -41574
rect 60376 -41580 60436 -41560
rect 59956 -41590 60336 -41580
rect 59856 -41660 59916 -41640
rect 59946 -41648 60346 -41642
rect 59756 -41740 59826 -41700
rect 59946 -41682 59958 -41648
rect 60334 -41682 60346 -41648
rect 60376 -41660 60436 -41640
rect 61126 -41640 61176 -41540
rect 61056 -41670 61176 -41640
rect 72610 -41510 73050 -41500
rect 59946 -41688 60346 -41682
rect 59946 -41740 60336 -41688
rect 72610 -41690 72820 -41510
rect 73040 -41690 73050 -41510
rect 77570 -41531 78630 -41489
rect 77570 -41565 77607 -41531
rect 77641 -41565 77699 -41531
rect 77733 -41565 77791 -41531
rect 77825 -41565 77883 -41531
rect 77917 -41565 77975 -41531
rect 78009 -41565 78630 -41531
rect 77570 -41570 78630 -41565
rect 78740 -41570 78850 -41460
rect 78960 -41570 79090 -41460
rect 79200 -41570 79410 -41460
rect 77570 -41600 79410 -41570
rect 79380 -41620 79410 -41600
rect 79680 -41620 79710 -41380
rect 79380 -41650 79710 -41620
rect 72610 -41700 73050 -41690
rect 77960 -41730 78600 -41720
rect 77960 -41740 78170 -41730
rect 59756 -41760 60536 -41740
rect 59756 -41800 59866 -41760
rect 60426 -41800 60536 -41760
rect 59756 -41810 60536 -41800
rect 59796 -41920 59806 -41810
rect 59916 -41920 59926 -41810
rect 59796 -41930 59926 -41920
rect 60436 -41830 60536 -41810
rect 60436 -41950 60446 -41830
rect 60526 -41950 60536 -41830
rect 77480 -41770 77590 -41760
rect 77480 -41860 77490 -41770
rect 77580 -41860 77590 -41770
rect 77960 -41780 77980 -41740
rect 78020 -41780 78170 -41740
rect 77480 -41870 77590 -41860
rect 77770 -41870 77780 -41810
rect 77840 -41870 77850 -41810
rect 60436 -41960 60536 -41950
rect 72610 -41880 73050 -41870
rect 77770 -41880 77850 -41870
rect 77960 -41860 78170 -41780
rect 59646 -42040 59716 -42030
rect 59706 -42100 59716 -42040
rect 72610 -42060 72820 -41880
rect 73040 -42060 73050 -41880
rect 77960 -41900 77980 -41860
rect 78020 -41900 78170 -41860
rect 77400 -41960 77560 -41940
rect 77400 -42040 77420 -41960
rect 72610 -42070 73050 -42060
rect 76900 -42060 77420 -42040
rect 59646 -42120 59716 -42100
rect 76900 -42220 76920 -42060
rect 77060 -42220 77420 -42060
rect 76900 -42240 77420 -42220
rect 77400 -42250 77420 -42240
rect 77540 -42040 77560 -41960
rect 77960 -41960 78170 -41900
rect 77960 -42000 77980 -41960
rect 78020 -42000 78170 -41960
rect 78290 -42000 78530 -41730
rect 78590 -42000 78600 -41730
rect 77960 -42010 78600 -42000
rect 77540 -42075 78040 -42040
rect 77540 -42109 77607 -42075
rect 77641 -42109 77699 -42075
rect 77733 -42109 77791 -42075
rect 77825 -42109 77883 -42075
rect 77917 -42109 77975 -42075
rect 78009 -42109 78040 -42075
rect 77540 -42165 78040 -42109
rect 77540 -42199 77609 -42165
rect 77643 -42199 77701 -42165
rect 77735 -42199 77793 -42165
rect 77827 -42199 77885 -42165
rect 77919 -42199 77977 -42165
rect 78011 -42199 78040 -42165
rect 77540 -42240 78040 -42199
rect 77540 -42250 77560 -42240
rect 77400 -42270 77560 -42250
rect 77960 -42340 78310 -42330
rect 77960 -42380 77980 -42340
rect 78020 -42380 78060 -42340
rect 58806 -42410 59356 -42380
rect 59846 -42390 60256 -42380
rect 59846 -42400 59996 -42390
rect 57556 -42420 59356 -42410
rect 57556 -42560 58986 -42420
rect 59126 -42560 59356 -42420
rect 57556 -42610 59356 -42560
rect 58806 -42690 59356 -42610
rect 59600 -42500 59996 -42400
rect 60106 -42400 60256 -42390
rect 60106 -42500 60600 -42400
rect 59600 -42800 60600 -42500
rect 77460 -42410 77570 -42400
rect 77460 -42500 77470 -42410
rect 77560 -42500 77570 -42410
rect 77770 -42440 77780 -42380
rect 77840 -42440 77850 -42380
rect 77770 -42450 77850 -42440
rect 77960 -42420 78060 -42380
rect 77460 -42510 77570 -42500
rect 77960 -42460 77980 -42420
rect 78020 -42460 78060 -42420
rect 77960 -42520 78060 -42460
rect 77960 -42560 77980 -42520
rect 78020 -42560 78060 -42520
rect 77960 -42600 78060 -42560
rect 77960 -42640 77980 -42600
rect 78020 -42640 78060 -42600
rect 78120 -42640 78310 -42340
rect 77960 -42650 78310 -42640
rect 79380 -42640 79710 -42610
rect 77580 -42680 78040 -42678
rect 79380 -42680 79410 -42640
rect 55710 -43000 55910 -42998
rect 43100 -43200 44400 -43000
rect 35900 -43258 44400 -43200
rect 25860 -43277 44400 -43258
rect 25860 -43674 25882 -43277
rect 26996 -43674 27124 -43277
rect 28238 -43674 28366 -43277
rect 29480 -43674 29608 -43277
rect 30722 -43674 30850 -43277
rect 31964 -43674 32092 -43277
rect 33206 -43674 33334 -43277
rect 34448 -43674 34576 -43277
rect 35690 -43300 44400 -43277
rect 35690 -43674 36000 -43300
rect 25860 -43944 36000 -43674
rect 25860 -44341 25882 -43944
rect 26996 -44341 27124 -43944
rect 28238 -44341 28366 -43944
rect 29480 -44341 29608 -43944
rect 30722 -44341 30850 -43944
rect 31964 -44341 32092 -43944
rect 33206 -44341 33334 -43944
rect 34448 -44341 34576 -43944
rect 35690 -44300 36000 -43944
rect 44300 -44300 44400 -43300
rect 55400 -43100 56200 -43000
rect 55400 -43500 55500 -43100
rect 56100 -43500 56200 -43100
rect 55400 -43600 56200 -43500
rect 59600 -43400 59800 -42800
rect 60400 -43400 60600 -42800
rect 77570 -42709 79410 -42680
rect 77570 -42743 77609 -42709
rect 77643 -42743 77701 -42709
rect 77735 -42743 77793 -42709
rect 77827 -42743 77885 -42709
rect 77919 -42743 77977 -42709
rect 78011 -42710 79410 -42709
rect 78011 -42743 78940 -42710
rect 77570 -42781 78940 -42743
rect 77570 -42815 77607 -42781
rect 77641 -42815 77699 -42781
rect 77733 -42815 77791 -42781
rect 77825 -42815 77883 -42781
rect 77917 -42815 77975 -42781
rect 78009 -42815 78067 -42781
rect 78101 -42815 78159 -42781
rect 78193 -42815 78351 -42781
rect 78385 -42815 78443 -42781
rect 78477 -42815 78535 -42781
rect 78569 -42815 78627 -42781
rect 78661 -42815 78719 -42781
rect 78753 -42815 78811 -42781
rect 78845 -42815 78940 -42781
rect 77570 -42820 78940 -42815
rect 79050 -42820 79130 -42710
rect 79240 -42820 79410 -42710
rect 77570 -42830 79410 -42820
rect 77570 -42846 78222 -42830
rect 78320 -42840 79410 -42830
rect 78322 -42846 79410 -42840
rect 77570 -42850 78210 -42846
rect 78589 -42850 79410 -42846
rect 78238 -42880 78310 -42877
rect 77460 -42930 77640 -42920
rect 77460 -43000 77470 -42930
rect 77540 -42940 77640 -42930
rect 77540 -42990 77580 -42940
rect 77630 -42990 77640 -42940
rect 78230 -42940 78240 -42880
rect 78300 -42940 78310 -42880
rect 79380 -42880 79410 -42850
rect 79680 -42880 79710 -42640
rect 82790 -42740 91440 -42710
rect 78830 -42920 79000 -42900
rect 79380 -42910 79710 -42880
rect 79980 -42910 80390 -42880
rect 78230 -42950 78300 -42940
rect 78830 -42970 78850 -42920
rect 77540 -43000 77640 -42990
rect 77460 -43010 77640 -43000
rect 78160 -43010 78230 -42990
rect 77860 -43050 77920 -43040
rect 77190 -43080 77270 -43070
rect 75920 -43140 75940 -43080
rect 76050 -43140 77200 -43080
rect 77260 -43090 77830 -43080
rect 77260 -43130 77770 -43090
rect 77810 -43130 77830 -43090
rect 77260 -43140 77830 -43130
rect 77860 -43120 77920 -43110
rect 77190 -43150 77270 -43140
rect 77860 -43160 77870 -43120
rect 77910 -43160 77920 -43120
rect 77390 -43210 77550 -43190
rect 77390 -43290 77410 -43210
rect 59600 -43600 60600 -43400
rect 76900 -43310 77410 -43290
rect 76900 -43450 76920 -43310
rect 77060 -43330 77410 -43310
rect 77530 -43290 77550 -43210
rect 77860 -43200 77920 -43160
rect 78160 -43180 78170 -43010
rect 78220 -43020 78230 -43010
rect 78220 -43040 78580 -43020
rect 78220 -43090 78470 -43040
rect 78560 -43090 78580 -43040
rect 78830 -43040 78860 -42970
rect 78220 -43100 78580 -43090
rect 78620 -43080 78710 -43070
rect 78220 -43180 78230 -43100
rect 78340 -43140 78410 -43130
rect 78620 -43140 78630 -43080
rect 78700 -43140 78710 -43080
rect 77860 -43240 77870 -43200
rect 77910 -43240 77920 -43200
rect 77860 -43260 77920 -43240
rect 77950 -43190 78030 -43180
rect 77950 -43250 77960 -43190
rect 78020 -43250 78030 -43190
rect 78160 -43200 78230 -43180
rect 78330 -43200 78340 -43140
rect 78410 -43200 78420 -43140
rect 78620 -43150 78710 -43140
rect 78830 -43090 78850 -43040
rect 78830 -43160 78860 -43090
rect 78830 -43210 78850 -43160
rect 78980 -43210 79000 -42920
rect 78830 -43230 79000 -43210
rect 77950 -43260 78030 -43250
rect 79980 -43290 80010 -42910
rect 80360 -42990 80390 -42910
rect 80360 -43190 80590 -42990
rect 80360 -43290 80390 -43190
rect 77530 -43325 78880 -43290
rect 79980 -43320 80390 -43290
rect 82790 -43310 82820 -42740
rect 91410 -43310 91440 -42740
rect 77530 -43330 77607 -43325
rect 77060 -43359 77607 -43330
rect 77641 -43359 77699 -43325
rect 77733 -43359 77791 -43325
rect 77825 -43359 77883 -43325
rect 77917 -43359 77975 -43325
rect 78009 -43359 78067 -43325
rect 78101 -43359 78159 -43325
rect 78193 -43359 78351 -43325
rect 78385 -43359 78443 -43325
rect 78477 -43359 78535 -43325
rect 78569 -43359 78627 -43325
rect 78661 -43359 78719 -43325
rect 78753 -43359 78811 -43325
rect 78845 -43359 78880 -43325
rect 77060 -43390 78880 -43359
rect 77060 -43450 77410 -43390
rect 76900 -43470 77410 -43450
rect 77390 -43510 77410 -43470
rect 77530 -43397 78880 -43390
rect 77530 -43431 77607 -43397
rect 77641 -43431 77699 -43397
rect 77733 -43431 77791 -43397
rect 77825 -43431 77883 -43397
rect 77917 -43431 77975 -43397
rect 78009 -43431 78067 -43397
rect 78101 -43431 78159 -43397
rect 78193 -43431 78880 -43397
rect 77530 -43470 78880 -43431
rect 82790 -43380 91440 -43310
rect 77530 -43510 77550 -43470
rect 77190 -43530 77270 -43520
rect 77390 -43530 77550 -43510
rect 77760 -43520 77820 -43500
rect 77190 -43590 77200 -43530
rect 77260 -43560 77270 -43530
rect 77760 -43560 77770 -43520
rect 77810 -43560 77820 -43520
rect 77260 -43590 77820 -43560
rect 77190 -43600 77820 -43590
rect 77760 -43610 77820 -43600
rect 77760 -43650 77770 -43610
rect 77810 -43650 77820 -43610
rect 77760 -43670 77820 -43650
rect 77850 -43670 77860 -43500
rect 77920 -43670 77930 -43500
rect 78170 -43510 78240 -43500
rect 78170 -43560 78200 -43510
rect 77850 -43680 77930 -43670
rect 77960 -43620 78030 -43610
rect 77960 -43680 77970 -43620
rect 77960 -43690 78030 -43680
rect 78170 -43650 78240 -43560
rect 78170 -43700 78200 -43650
rect 77420 -43760 77510 -43750
rect 77420 -43830 77430 -43760
rect 77500 -43830 77510 -43760
rect 77420 -43840 77510 -43830
rect 78170 -43790 78240 -43700
rect 78170 -43840 78200 -43790
rect 78170 -43870 78240 -43840
rect 78300 -43870 78310 -43500
rect 82790 -43550 83450 -43380
rect 83620 -43550 85150 -43380
rect 85320 -43550 86530 -43380
rect 86700 -43550 87820 -43380
rect 87990 -43550 89340 -43380
rect 89510 -43550 90750 -43380
rect 90920 -43550 91440 -43380
rect 82790 -43591 91440 -43550
rect 82790 -43625 82867 -43591
rect 82901 -43625 82959 -43591
rect 82993 -43625 83051 -43591
rect 83085 -43625 83143 -43591
rect 83177 -43625 83235 -43591
rect 83269 -43625 83327 -43591
rect 83361 -43625 83419 -43591
rect 83453 -43625 83511 -43591
rect 83545 -43625 83603 -43591
rect 83637 -43625 83695 -43591
rect 83729 -43625 83787 -43591
rect 83821 -43625 83879 -43591
rect 83913 -43625 83971 -43591
rect 84005 -43625 84063 -43591
rect 84097 -43625 84155 -43591
rect 84189 -43625 84247 -43591
rect 84281 -43625 84339 -43591
rect 84373 -43625 84431 -43591
rect 84465 -43625 84523 -43591
rect 84557 -43625 84615 -43591
rect 84649 -43625 84707 -43591
rect 84741 -43625 84799 -43591
rect 84833 -43625 84891 -43591
rect 84925 -43625 84983 -43591
rect 85017 -43625 85075 -43591
rect 85109 -43625 85167 -43591
rect 85201 -43625 85259 -43591
rect 85293 -43625 85351 -43591
rect 85385 -43625 85443 -43591
rect 85477 -43625 85535 -43591
rect 85569 -43625 85627 -43591
rect 85661 -43625 85719 -43591
rect 85753 -43625 85811 -43591
rect 85845 -43625 85903 -43591
rect 85937 -43625 85995 -43591
rect 86029 -43625 86087 -43591
rect 86121 -43625 86179 -43591
rect 86213 -43625 86271 -43591
rect 86305 -43625 86363 -43591
rect 86397 -43625 86455 -43591
rect 86489 -43625 86547 -43591
rect 86581 -43625 86639 -43591
rect 86673 -43625 86731 -43591
rect 86765 -43625 86823 -43591
rect 86857 -43625 86915 -43591
rect 86949 -43625 87007 -43591
rect 87041 -43625 87099 -43591
rect 87133 -43625 87191 -43591
rect 87225 -43625 87283 -43591
rect 87317 -43625 87375 -43591
rect 87409 -43625 87467 -43591
rect 87501 -43625 87559 -43591
rect 87593 -43625 87651 -43591
rect 87685 -43625 87743 -43591
rect 87777 -43625 87835 -43591
rect 87869 -43625 87927 -43591
rect 87961 -43625 88019 -43591
rect 88053 -43625 88111 -43591
rect 88145 -43625 88203 -43591
rect 88237 -43625 88295 -43591
rect 88329 -43625 88387 -43591
rect 88421 -43625 88479 -43591
rect 88513 -43625 88571 -43591
rect 88605 -43625 88663 -43591
rect 88697 -43625 88755 -43591
rect 88789 -43625 88847 -43591
rect 88881 -43625 88939 -43591
rect 88973 -43625 89031 -43591
rect 89065 -43625 89123 -43591
rect 89157 -43625 89215 -43591
rect 89249 -43625 89307 -43591
rect 89341 -43625 89399 -43591
rect 89433 -43625 89491 -43591
rect 89525 -43625 89583 -43591
rect 89617 -43625 89675 -43591
rect 89709 -43625 89767 -43591
rect 89801 -43625 89859 -43591
rect 89893 -43625 89951 -43591
rect 89985 -43625 90043 -43591
rect 90077 -43625 90135 -43591
rect 90169 -43625 90227 -43591
rect 90261 -43625 90319 -43591
rect 90353 -43625 90411 -43591
rect 90445 -43625 90503 -43591
rect 90537 -43625 90595 -43591
rect 90629 -43625 90687 -43591
rect 90721 -43625 90779 -43591
rect 90813 -43625 90871 -43591
rect 90905 -43625 90963 -43591
rect 90997 -43625 91055 -43591
rect 91089 -43625 91147 -43591
rect 91181 -43625 91239 -43591
rect 91273 -43625 91331 -43591
rect 91365 -43625 91440 -43591
rect 82790 -43660 91440 -43625
rect 86790 -43790 86880 -43780
rect 85310 -43810 85400 -43800
rect 78230 -43880 78310 -43870
rect 79380 -43860 79710 -43830
rect 79380 -43910 79410 -43860
rect 77570 -43940 79410 -43910
rect 77570 -43941 78280 -43940
rect 77570 -43975 77607 -43941
rect 77641 -43975 77699 -43941
rect 77733 -43975 77791 -43941
rect 77825 -43975 77883 -43941
rect 77917 -43975 77975 -43941
rect 78009 -43975 78067 -43941
rect 78101 -43975 78159 -43941
rect 78193 -43975 78280 -43941
rect 35690 -44341 44400 -44300
rect 25860 -44358 44400 -44341
rect 35900 -44400 44400 -44358
rect 55420 -44080 55800 -44000
rect 77570 -44013 78280 -43975
rect 77570 -44047 77607 -44013
rect 77641 -44047 77699 -44013
rect 77733 -44047 77791 -44013
rect 77825 -44047 77883 -44013
rect 77917 -44047 77975 -44013
rect 78009 -44047 78067 -44013
rect 78101 -44047 78159 -44013
rect 78193 -44047 78280 -44013
rect 77570 -44050 78280 -44047
rect 78390 -44050 78580 -43940
rect 78690 -44050 78880 -43940
rect 78990 -44050 79410 -43940
rect 77570 -44080 79410 -44050
rect 55420 -44360 55500 -44080
rect 55720 -44360 55800 -44080
rect 79380 -44100 79410 -44080
rect 79680 -44100 79710 -43860
rect 82460 -43890 82950 -43880
rect 82460 -44000 82470 -43890
rect 82550 -43900 82950 -43890
rect 82550 -43990 82880 -43900
rect 82930 -43990 82950 -43900
rect 82550 -44000 82950 -43990
rect 82460 -44010 82950 -44000
rect 83030 -43890 83110 -43880
rect 83030 -44000 83040 -43890
rect 83100 -44000 83110 -43890
rect 83030 -44010 83110 -44000
rect 85310 -44000 85320 -43810
rect 85390 -44000 85400 -43810
rect 85580 -43870 86490 -43860
rect 85580 -43950 85590 -43870
rect 86480 -43950 86490 -43870
rect 85580 -43960 86490 -43950
rect 85310 -44010 85400 -44000
rect 86790 -44000 86800 -43790
rect 86870 -44000 86880 -43790
rect 88260 -43800 88350 -43790
rect 87030 -43870 87930 -43860
rect 87030 -43950 87040 -43870
rect 87920 -43950 87930 -43870
rect 87030 -43960 87930 -43950
rect 86790 -44010 86880 -44000
rect 88260 -44000 88270 -43800
rect 88340 -44000 88350 -43800
rect 89730 -43800 89820 -43790
rect 88500 -43880 89400 -43870
rect 88500 -43950 88510 -43880
rect 89390 -43950 89400 -43880
rect 88500 -43960 89400 -43950
rect 88260 -44010 88350 -44000
rect 89730 -44010 89740 -43800
rect 89810 -44010 89820 -43800
rect 91200 -43800 91290 -43790
rect 89970 -43879 90770 -43870
rect 89970 -43897 89982 -43879
rect 89970 -43899 89980 -43897
rect 89970 -43933 89978 -43899
rect 89970 -43951 89982 -43933
rect 90762 -43951 90770 -43879
rect 89970 -43960 90770 -43951
rect 89730 -44020 89820 -44010
rect 91200 -44010 91210 -43800
rect 91280 -44010 91290 -43800
rect 91200 -44020 91290 -44010
rect 92000 -44050 95800 -43200
rect 91750 -44080 95800 -44050
rect 78160 -44130 78310 -44120
rect 79380 -44130 79710 -44100
rect 75920 -44240 75940 -44150
rect 76050 -44170 77530 -44150
rect 76050 -44220 77470 -44170
rect 77510 -44220 77530 -44170
rect 76050 -44240 77530 -44220
rect 75640 -44330 75660 -44270
rect 75760 -44300 77640 -44270
rect 75760 -44320 77920 -44300
rect 75760 -44330 77870 -44320
rect 77570 -44360 77870 -44330
rect 77910 -44360 77920 -44320
rect 55420 -44440 55800 -44360
rect 77380 -44380 77540 -44360
rect 77570 -44380 77920 -44360
rect 54090 -44538 54890 -44498
rect 54090 -44668 54150 -44538
rect 53510 -44720 53800 -44718
rect 53460 -44740 53800 -44720
rect 35900 -44860 44400 -44800
rect 25862 -44879 44400 -44860
rect 25862 -45276 25882 -44879
rect 26996 -45276 27124 -44879
rect 28238 -45276 28366 -44879
rect 29480 -45276 29608 -44879
rect 30722 -45276 30850 -44879
rect 31964 -45276 32092 -44879
rect 33206 -45276 33334 -44879
rect 34448 -45276 34576 -44879
rect 35690 -44900 44400 -44879
rect 35690 -45276 36000 -44900
rect 25862 -45542 36000 -45276
rect 25862 -45939 25882 -45542
rect 26996 -45939 27124 -45542
rect 28238 -45939 28366 -45542
rect 29480 -45939 29608 -45542
rect 30722 -45939 30850 -45542
rect 31964 -45939 32092 -45542
rect 33206 -45939 33334 -45542
rect 34448 -45939 34576 -45542
rect 35690 -45900 36000 -45542
rect 44300 -45900 44400 -44900
rect 53460 -44940 53480 -44740
rect 53780 -44940 53800 -44740
rect 54080 -44798 54150 -44668
rect 54860 -44778 54890 -44538
rect 54850 -44798 54890 -44778
rect 54080 -44866 54880 -44798
rect 54079 -44872 54880 -44866
rect 54079 -44906 54091 -44872
rect 54867 -44898 54880 -44872
rect 54867 -44906 54879 -44898
rect 54079 -44912 54879 -44906
rect 53460 -44960 53800 -44940
rect 53510 -45058 53800 -44960
rect 53002 -45220 53480 -45158
rect 35690 -45939 44400 -45900
rect 25862 -45960 44400 -45939
rect 35900 -46000 44400 -45960
rect 53000 -45358 53480 -45220
rect 53510 -45168 53520 -45058
rect 53640 -45168 53800 -45058
rect 53510 -45288 53800 -45168
rect 53970 -44934 54040 -44918
rect 53970 -44972 53998 -44934
rect 54032 -44972 54040 -44934
rect 53970 -45168 54040 -44972
rect 54920 -44934 54990 -44918
rect 54920 -44972 54926 -44934
rect 54960 -44972 54990 -44934
rect 54079 -45000 54879 -44994
rect 54079 -45034 54091 -45000
rect 54867 -45034 54879 -45000
rect 54079 -45038 54879 -45034
rect 54079 -45040 54750 -45038
rect 54090 -45088 54750 -45040
rect 54740 -45118 54750 -45088
rect 54850 -45040 54879 -45038
rect 54850 -45108 54860 -45040
rect 54840 -45118 54860 -45108
rect 54750 -45128 54860 -45118
rect 54920 -45168 54990 -44972
rect 55430 -45018 55520 -45008
rect 55290 -45128 55390 -45118
rect 53970 -45198 55290 -45168
rect 55430 -45158 55520 -45088
rect 53970 -45208 55390 -45198
rect 54050 -45218 55380 -45208
rect 54050 -45228 54880 -45218
rect 54050 -45238 54091 -45228
rect 54079 -45262 54091 -45238
rect 54867 -45238 54880 -45228
rect 54867 -45262 54879 -45238
rect 54079 -45268 54879 -45262
rect 54920 -45278 54990 -45268
rect 53510 -45306 53630 -45288
rect 53510 -45338 53526 -45306
rect 53514 -45340 53526 -45338
rect 53614 -45338 53630 -45306
rect 53940 -45290 54038 -45278
rect 53940 -45298 53998 -45290
rect 53614 -45340 53626 -45338
rect 53514 -45346 53626 -45340
rect 35900 -46458 43500 -46400
rect 25860 -46477 43500 -46458
rect 25860 -46874 25882 -46477
rect 26996 -46874 27124 -46477
rect 28238 -46874 28366 -46477
rect 29480 -46874 29608 -46477
rect 30722 -46874 30850 -46477
rect 31964 -46874 32092 -46477
rect 33206 -46874 33334 -46477
rect 34448 -46874 34576 -46477
rect 35690 -46500 43500 -46477
rect 35690 -46874 36000 -46500
rect 25860 -47136 36000 -46874
rect 25860 -47533 25882 -47136
rect 26996 -47533 27124 -47136
rect 28238 -47533 28366 -47136
rect 29480 -47533 29608 -47136
rect 30722 -47533 30850 -47136
rect 31964 -47533 32092 -47136
rect 33206 -47533 33334 -47136
rect 34448 -47533 34576 -47136
rect 35690 -47500 36000 -47136
rect 43400 -47500 43500 -46500
rect 53000 -47108 53050 -45358
rect 53250 -45368 53480 -45358
rect 53250 -46718 53330 -45368
rect 53400 -45378 53480 -45368
rect 53400 -45390 53504 -45378
rect 53400 -46166 53464 -45390
rect 53498 -46166 53504 -45390
rect 53400 -46178 53504 -46166
rect 53636 -45388 53682 -45378
rect 53636 -45390 53760 -45388
rect 53636 -46166 53642 -45390
rect 53676 -46166 53760 -45390
rect 53940 -45398 53950 -45298
rect 54032 -45328 54038 -45290
rect 54020 -45340 54038 -45328
rect 54020 -45398 54030 -45340
rect 54079 -45356 54879 -45350
rect 54079 -45390 54091 -45356
rect 54867 -45390 54879 -45356
rect 54920 -45378 54990 -45368
rect 55320 -45368 55380 -45218
rect 54079 -45396 54879 -45390
rect 53940 -45418 54030 -45398
rect 54090 -45428 54870 -45396
rect 55320 -45402 55334 -45368
rect 55368 -45402 55380 -45368
rect 55320 -45408 55380 -45402
rect 53840 -45728 53920 -45718
rect 53840 -45838 53860 -45728
rect 53840 -45848 53920 -45838
rect 53840 -46040 53900 -45848
rect 54320 -45928 54510 -45428
rect 55440 -45438 55520 -45158
rect 55410 -45440 55520 -45438
rect 55284 -45448 55330 -45440
rect 55230 -45452 55330 -45448
rect 55230 -45458 55290 -45452
rect 55324 -45628 55330 -45452
rect 55230 -45638 55330 -45628
rect 55284 -45640 55330 -45638
rect 55372 -45448 55520 -45440
rect 55372 -45452 55430 -45448
rect 55372 -45628 55378 -45452
rect 55412 -45618 55430 -45452
rect 55510 -45618 55520 -45448
rect 55412 -45628 55520 -45618
rect 55372 -45640 55418 -45628
rect 55580 -45728 55720 -44440
rect 77380 -44500 77400 -44380
rect 77520 -44500 77540 -44380
rect 77860 -44410 77920 -44380
rect 77750 -44420 77830 -44410
rect 77750 -44480 77760 -44420
rect 77820 -44480 77830 -44420
rect 77750 -44490 77830 -44480
rect 77860 -44470 77870 -44410
rect 77910 -44470 77920 -44410
rect 77860 -44490 77920 -44470
rect 77960 -44350 78040 -44340
rect 77960 -44470 77970 -44350
rect 78030 -44470 78040 -44350
rect 77960 -44480 78040 -44470
rect 78160 -44470 78180 -44130
rect 78300 -44470 78310 -44130
rect 78160 -44480 78310 -44470
rect 82790 -44135 91440 -44100
rect 82790 -44169 82867 -44135
rect 82901 -44169 82959 -44135
rect 82993 -44169 83051 -44135
rect 83085 -44169 83143 -44135
rect 83177 -44169 83235 -44135
rect 83269 -44169 83327 -44135
rect 83361 -44169 83419 -44135
rect 83453 -44169 83511 -44135
rect 83545 -44169 83603 -44135
rect 83637 -44169 83695 -44135
rect 83729 -44169 83787 -44135
rect 83821 -44169 83879 -44135
rect 83913 -44169 83971 -44135
rect 84005 -44169 84063 -44135
rect 84097 -44169 84155 -44135
rect 84189 -44169 84247 -44135
rect 84281 -44169 84339 -44135
rect 84373 -44169 84431 -44135
rect 84465 -44169 84523 -44135
rect 84557 -44169 84615 -44135
rect 84649 -44169 84707 -44135
rect 84741 -44169 84799 -44135
rect 84833 -44169 84891 -44135
rect 84925 -44169 84983 -44135
rect 85017 -44169 85075 -44135
rect 85109 -44169 85167 -44135
rect 85201 -44169 85259 -44135
rect 85293 -44169 85351 -44135
rect 85385 -44169 85443 -44135
rect 85477 -44169 85535 -44135
rect 85569 -44169 85627 -44135
rect 85661 -44169 85719 -44135
rect 85753 -44169 85811 -44135
rect 85845 -44169 85903 -44135
rect 85937 -44169 85995 -44135
rect 86029 -44169 86087 -44135
rect 86121 -44169 86179 -44135
rect 86213 -44169 86271 -44135
rect 86305 -44169 86363 -44135
rect 86397 -44169 86455 -44135
rect 86489 -44169 86547 -44135
rect 86581 -44169 86639 -44135
rect 86673 -44169 86731 -44135
rect 86765 -44169 86823 -44135
rect 86857 -44169 86915 -44135
rect 86949 -44169 87007 -44135
rect 87041 -44169 87099 -44135
rect 87133 -44169 87191 -44135
rect 87225 -44169 87283 -44135
rect 87317 -44169 87375 -44135
rect 87409 -44169 87467 -44135
rect 87501 -44169 87559 -44135
rect 87593 -44169 87651 -44135
rect 87685 -44169 87743 -44135
rect 87777 -44169 87835 -44135
rect 87869 -44169 87927 -44135
rect 87961 -44169 88019 -44135
rect 88053 -44169 88111 -44135
rect 88145 -44169 88203 -44135
rect 88237 -44169 88295 -44135
rect 88329 -44169 88387 -44135
rect 88421 -44169 88479 -44135
rect 88513 -44169 88571 -44135
rect 88605 -44169 88663 -44135
rect 88697 -44169 88755 -44135
rect 88789 -44169 88847 -44135
rect 88881 -44169 88939 -44135
rect 88973 -44169 89031 -44135
rect 89065 -44169 89123 -44135
rect 89157 -44169 89215 -44135
rect 89249 -44169 89307 -44135
rect 89341 -44169 89399 -44135
rect 89433 -44169 89491 -44135
rect 89525 -44169 89583 -44135
rect 89617 -44169 89675 -44135
rect 89709 -44169 89767 -44135
rect 89801 -44169 89859 -44135
rect 89893 -44169 89951 -44135
rect 89985 -44169 90043 -44135
rect 90077 -44169 90135 -44135
rect 90169 -44169 90227 -44135
rect 90261 -44169 90319 -44135
rect 90353 -44169 90411 -44135
rect 90445 -44169 90503 -44135
rect 90537 -44169 90595 -44135
rect 90629 -44169 90687 -44135
rect 90721 -44169 90779 -44135
rect 90813 -44169 90871 -44135
rect 90905 -44169 90963 -44135
rect 90997 -44169 91055 -44135
rect 91089 -44169 91147 -44135
rect 91181 -44169 91239 -44135
rect 91273 -44169 91331 -44135
rect 91365 -44169 91440 -44135
rect 82790 -44210 91440 -44169
rect 82790 -44380 83480 -44210
rect 83650 -44220 86530 -44210
rect 83650 -44380 85120 -44220
rect 82790 -44390 85120 -44380
rect 85290 -44380 86530 -44220
rect 86700 -44380 87910 -44210
rect 88080 -44220 91440 -44210
rect 88080 -44380 89450 -44220
rect 85290 -44390 89450 -44380
rect 89620 -44390 90730 -44220
rect 90900 -44390 91440 -44220
rect 82790 -44440 91440 -44390
rect 76900 -44520 77540 -44500
rect 58776 -44670 59306 -44550
rect 58776 -44680 58966 -44670
rect 56146 -44780 57366 -44730
rect 55954 -44928 56046 -44916
rect 56146 -44928 56506 -44780
rect 55954 -45098 55960 -44928
rect 56040 -45098 56046 -44928
rect 55954 -45110 56046 -45098
rect 56120 -44958 56506 -44928
rect 56120 -45168 56190 -44958
rect 56390 -45030 56506 -44958
rect 57016 -44934 57366 -44780
rect 57586 -44830 58966 -44680
rect 59126 -44830 59306 -44670
rect 57586 -44850 59306 -44830
rect 59946 -44700 60386 -44600
rect 76900 -44610 76920 -44520
rect 77060 -44557 78230 -44520
rect 77060 -44591 77607 -44557
rect 77641 -44591 77699 -44557
rect 77733 -44591 77791 -44557
rect 77825 -44591 77883 -44557
rect 77917 -44591 77975 -44557
rect 78009 -44591 78067 -44557
rect 78101 -44591 78159 -44557
rect 78193 -44591 78230 -44557
rect 77060 -44610 78230 -44591
rect 76900 -44630 78230 -44610
rect 57586 -44880 58986 -44850
rect 59946 -44860 59956 -44700
rect 60166 -44860 60386 -44700
rect 77380 -44750 77400 -44630
rect 77520 -44631 78230 -44630
rect 77520 -44665 77607 -44631
rect 77641 -44665 77699 -44631
rect 77733 -44665 77791 -44631
rect 77825 -44665 77883 -44631
rect 77917 -44665 77975 -44631
rect 78009 -44665 78067 -44631
rect 78101 -44665 78159 -44631
rect 78193 -44665 78230 -44631
rect 77520 -44700 78230 -44665
rect 77520 -44750 77540 -44700
rect 77380 -44770 77540 -44750
rect 77750 -44740 77830 -44730
rect 77750 -44800 77760 -44740
rect 77820 -44800 77830 -44740
rect 77750 -44810 77830 -44800
rect 77860 -44840 77920 -44830
rect 57016 -45030 57368 -44934
rect 56390 -45070 57368 -45030
rect 56390 -45168 57126 -45070
rect 56120 -45174 57126 -45168
rect 56120 -45178 56750 -45174
rect 55880 -45218 55970 -45208
rect 55870 -45296 55880 -45250
rect 55970 -45296 55982 -45250
rect 55880 -45308 55970 -45298
rect 55000 -45738 55090 -45728
rect 55000 -45848 55090 -45838
rect 54710 -45928 54960 -45908
rect 53940 -45968 54960 -45928
rect 53940 -45972 54730 -45968
rect 53930 -45978 54730 -45972
rect 53930 -46012 53942 -45978
rect 54718 -46012 54730 -45978
rect 53930 -46018 54730 -46012
rect 53840 -46128 53858 -46040
rect 53892 -46128 53900 -46040
rect 53840 -46148 53900 -46128
rect 54762 -46038 54850 -46028
rect 54762 -46040 54770 -46038
rect 54762 -46128 54768 -46040
rect 54840 -46128 54850 -46038
rect 54762 -46140 54850 -46128
rect 54770 -46148 54850 -46140
rect 53636 -46178 53760 -46166
rect 53400 -46396 53480 -46178
rect 53514 -46216 53626 -46210
rect 53514 -46218 53526 -46216
rect 53510 -46250 53526 -46218
rect 53614 -46218 53626 -46216
rect 53614 -46250 53630 -46218
rect 53510 -46324 53630 -46250
rect 53510 -46358 53526 -46324
rect 53614 -46358 53630 -46324
rect 53680 -46238 53760 -46178
rect 53930 -46156 54730 -46150
rect 53930 -46190 53942 -46156
rect 54718 -46190 54730 -46156
rect 53930 -46196 54730 -46190
rect 53940 -46228 54720 -46196
rect 53920 -46238 54720 -46228
rect 53680 -46328 54720 -46238
rect 53514 -46364 53626 -46358
rect 53680 -46396 53760 -46328
rect 53920 -46338 54720 -46328
rect 53940 -46378 54720 -46338
rect 54900 -46368 54960 -45968
rect 55010 -45960 55090 -45848
rect 55540 -45738 55720 -45728
rect 55630 -45838 55720 -45738
rect 55130 -45874 55506 -45868
rect 55130 -45908 55142 -45874
rect 55494 -45908 55506 -45874
rect 55130 -45914 55506 -45908
rect 55010 -45994 55046 -45960
rect 55080 -45994 55090 -45960
rect 55010 -46008 55090 -45994
rect 55142 -46040 55494 -45914
rect 55540 -45960 55720 -45838
rect 55540 -45994 55556 -45960
rect 55590 -45994 55720 -45960
rect 55540 -46008 55720 -45994
rect 55780 -45340 55860 -45328
rect 55130 -46046 55506 -46040
rect 55130 -46080 55142 -46046
rect 55494 -46078 55506 -46046
rect 55494 -46080 55510 -46078
rect 55130 -46086 55510 -46080
rect 55140 -46098 55510 -46086
rect 55780 -46098 55820 -45340
rect 55140 -46116 55820 -46098
rect 55854 -46116 55860 -45340
rect 55140 -46128 55860 -46116
rect 55992 -45340 56038 -45328
rect 55992 -46116 55998 -45340
rect 56032 -45348 56038 -45340
rect 56120 -45348 56300 -45178
rect 57098 -45200 57126 -45174
rect 57356 -45200 57368 -45070
rect 57098 -45214 57368 -45200
rect 57096 -45245 57372 -45214
rect 57096 -45279 57125 -45245
rect 57159 -45279 57217 -45245
rect 57251 -45279 57309 -45245
rect 57343 -45279 57372 -45245
rect 57096 -45310 57372 -45279
rect 56032 -45706 56300 -45348
rect 56590 -45468 56660 -45458
rect 56660 -45534 57000 -45468
rect 57586 -45530 57706 -44880
rect 59946 -44890 60386 -44860
rect 75920 -44900 75940 -44840
rect 76050 -44850 77920 -44840
rect 76050 -44890 77870 -44850
rect 77910 -44890 77920 -44850
rect 76050 -44900 77920 -44890
rect 77860 -44910 77920 -44900
rect 77950 -44850 78030 -44840
rect 77950 -44920 77960 -44850
rect 78020 -44920 78030 -44850
rect 77950 -44930 78030 -44920
rect 77560 -44950 77640 -44930
rect 77560 -44970 77580 -44950
rect 75210 -45060 75230 -44970
rect 75330 -45040 77580 -44970
rect 77630 -45040 77640 -44950
rect 75330 -45060 77640 -45040
rect 78170 -44950 78760 -44940
rect 78170 -45080 78190 -44950
rect 78260 -45080 78640 -44950
rect 78170 -45090 78640 -45080
rect 78750 -45090 78760 -44950
rect 82790 -45010 82820 -44440
rect 91410 -45010 91440 -44440
rect 91750 -44460 91780 -44080
rect 92130 -44460 95800 -44080
rect 91750 -44490 95800 -44460
rect 82790 -45040 91440 -45010
rect 78170 -45100 78760 -45090
rect 79380 -45120 79710 -45090
rect 57366 -45534 57706 -45530
rect 56660 -45538 57188 -45534
rect 56660 -45544 57190 -45538
rect 56660 -45594 57118 -45544
rect 57178 -45594 57190 -45544
rect 57314 -45540 57706 -45534
rect 57314 -45580 57326 -45540
rect 57366 -45580 57706 -45540
rect 57314 -45586 57706 -45580
rect 57366 -45590 57706 -45586
rect 58896 -45170 58986 -45150
rect 58896 -45230 58906 -45170
rect 58896 -45520 58926 -45230
rect 58966 -45520 58986 -45170
rect 59106 -45170 59516 -45160
rect 59106 -45230 59216 -45170
rect 59276 -45230 59326 -45170
rect 59386 -45230 59436 -45170
rect 59496 -45230 59516 -45170
rect 59106 -45247 59516 -45230
rect 59626 -45170 59706 -45130
rect 79380 -45140 79410 -45120
rect 59626 -45230 59636 -45170
rect 59626 -45240 59656 -45230
rect 59106 -45280 59125 -45247
rect 59113 -45281 59125 -45280
rect 59501 -45280 59516 -45247
rect 59501 -45281 59513 -45280
rect 59113 -45287 59513 -45281
rect 59546 -45290 59616 -45280
rect 59276 -45330 59356 -45320
rect 59276 -45349 59286 -45330
rect 59113 -45355 59286 -45349
rect 59346 -45349 59356 -45330
rect 59346 -45355 59513 -45349
rect 59113 -45389 59125 -45355
rect 59501 -45389 59513 -45355
rect 59606 -45350 59616 -45290
rect 59546 -45360 59616 -45350
rect 59113 -45390 59286 -45389
rect 59346 -45390 59513 -45389
rect 59016 -45400 59076 -45390
rect 59113 -45395 59513 -45390
rect 59276 -45400 59356 -45395
rect 59546 -45410 59616 -45400
rect 59016 -45470 59076 -45460
rect 59113 -45463 59513 -45457
rect 59113 -45497 59125 -45463
rect 59501 -45497 59513 -45463
rect 59606 -45470 59616 -45410
rect 59546 -45480 59616 -45470
rect 59113 -45500 59513 -45497
rect 59113 -45503 59516 -45500
rect 58896 -45530 58986 -45520
rect 58896 -45590 58906 -45530
rect 58966 -45590 58986 -45530
rect 58896 -45592 58986 -45590
rect 59116 -45520 59516 -45503
rect 59646 -45510 59656 -45240
rect 59116 -45580 59216 -45520
rect 59276 -45580 59336 -45520
rect 59396 -45580 59436 -45520
rect 59496 -45580 59516 -45520
rect 56660 -45598 57190 -45594
rect 56590 -45600 57190 -45598
rect 56590 -45604 57188 -45600
rect 56590 -45668 57000 -45604
rect 56032 -45718 56356 -45706
rect 56032 -46116 56280 -45718
rect 55992 -46128 56280 -46116
rect 55140 -46138 55200 -46128
rect 55450 -46158 55810 -46128
rect 55870 -46166 55982 -46160
rect 55870 -46200 55882 -46166
rect 55970 -46200 55982 -46166
rect 55870 -46206 55982 -46200
rect 55140 -46218 55200 -46208
rect 55024 -46248 55116 -46236
rect 55024 -46328 55030 -46248
rect 55110 -46328 55116 -46248
rect 55024 -46340 55116 -46328
rect 55734 -46248 55816 -46236
rect 55734 -46328 55740 -46248
rect 55810 -46328 55816 -46248
rect 55734 -46340 55816 -46328
rect 55880 -46238 55970 -46206
rect 55880 -46364 55970 -46328
rect 56060 -46348 56280 -46128
rect 56350 -46348 56356 -45718
rect 56480 -45788 56550 -45778
rect 56480 -45858 56550 -45848
rect 56590 -45887 56750 -45668
rect 58894 -45686 58988 -45592
rect 59116 -45600 59516 -45580
rect 59636 -45520 59656 -45510
rect 59696 -45520 59706 -45170
rect 77570 -45175 79410 -45140
rect 77570 -45209 77607 -45175
rect 77641 -45209 77699 -45175
rect 77733 -45209 77791 -45175
rect 77825 -45209 77883 -45175
rect 77917 -45209 77975 -45175
rect 78009 -45209 78067 -45175
rect 78101 -45209 78159 -45175
rect 78193 -45180 79410 -45175
rect 78193 -45209 79120 -45180
rect 77570 -45251 79120 -45209
rect 77570 -45285 77607 -45251
rect 77641 -45285 77699 -45251
rect 77733 -45285 77791 -45251
rect 77825 -45285 77883 -45251
rect 77917 -45285 77975 -45251
rect 78009 -45285 78067 -45251
rect 78101 -45285 78159 -45251
rect 78193 -45285 78251 -45251
rect 78285 -45285 78343 -45251
rect 78377 -45285 78435 -45251
rect 78469 -45285 78527 -45251
rect 78561 -45285 78619 -45251
rect 78653 -45285 78711 -45251
rect 78745 -45285 78803 -45251
rect 78837 -45285 78895 -45251
rect 78929 -45285 78987 -45251
rect 79021 -45285 79120 -45251
rect 77570 -45290 79120 -45285
rect 79230 -45290 79410 -45180
rect 77570 -45316 79410 -45290
rect 77570 -45320 77720 -45316
rect 77880 -45320 79410 -45316
rect 59856 -45340 59976 -45330
rect 59856 -45430 59866 -45340
rect 59966 -45430 59976 -45340
rect 59856 -45440 59976 -45430
rect 60436 -45420 60446 -45320
rect 60526 -45420 60536 -45320
rect 77750 -45350 77850 -45345
rect 76480 -45420 76500 -45350
rect 76600 -45352 77850 -45350
rect 76600 -45392 77770 -45352
rect 77830 -45392 77850 -45352
rect 79380 -45360 79410 -45320
rect 79680 -45360 79710 -45120
rect 76600 -45400 77850 -45392
rect 76600 -45420 77580 -45400
rect 77750 -45401 77850 -45400
rect 79000 -45370 79210 -45360
rect 60436 -45440 60536 -45420
rect 59636 -45530 59706 -45520
rect 59696 -45590 59706 -45530
rect 59636 -45610 59706 -45590
rect 59756 -45460 60536 -45440
rect 59756 -45500 59866 -45460
rect 60426 -45500 60536 -45460
rect 78060 -45480 78150 -45470
rect 59756 -45510 60536 -45500
rect 59756 -45550 59826 -45510
rect 59066 -45640 59176 -45630
rect 58896 -45750 58986 -45686
rect 59066 -45710 59076 -45640
rect 59166 -45710 59176 -45640
rect 59066 -45712 59103 -45710
rect 59137 -45712 59176 -45710
rect 59066 -45720 59176 -45712
rect 59756 -45740 59766 -45550
rect 59806 -45740 59826 -45550
rect 59956 -45568 60046 -45540
rect 59946 -45574 60046 -45568
rect 60126 -45568 60336 -45540
rect 60126 -45574 60346 -45568
rect 75210 -45570 75230 -45500
rect 75330 -45570 77880 -45500
rect 59856 -45610 59916 -45600
rect 59946 -45608 59958 -45574
rect 60334 -45608 60346 -45574
rect 77800 -45590 77880 -45570
rect 59946 -45614 60346 -45608
rect 77590 -45610 77720 -45600
rect 60376 -45620 60446 -45610
rect 77380 -45620 77520 -45610
rect 59856 -45690 59916 -45680
rect 59946 -45682 60346 -45676
rect 59946 -45716 59958 -45682
rect 60334 -45716 60346 -45682
rect 60376 -45690 60446 -45680
rect 76900 -45630 77520 -45620
rect 76900 -45640 77390 -45630
rect 59946 -45722 59976 -45716
rect 57098 -45758 57368 -45754
rect 57096 -45764 57372 -45758
rect 57096 -45850 57098 -45764
rect 56424 -45888 56470 -45887
rect 56060 -46360 56356 -46348
rect 56410 -45899 56470 -45888
rect 53400 -46408 53504 -46396
rect 53400 -46718 53464 -46408
rect 53250 -47108 53464 -46718
rect 53000 -47184 53464 -47108
rect 53498 -47184 53504 -46408
rect 53000 -47188 53504 -47184
rect 53458 -47196 53504 -47188
rect 53636 -46408 53760 -46396
rect 53636 -47184 53642 -46408
rect 53676 -47184 53760 -46408
rect 53930 -46384 54730 -46378
rect 53930 -46418 53942 -46384
rect 54718 -46418 54730 -46384
rect 53930 -46424 54730 -46418
rect 53830 -46446 53900 -46428
rect 53830 -46534 53858 -46446
rect 53892 -46534 53900 -46446
rect 53830 -46728 53900 -46534
rect 54760 -46446 54850 -46428
rect 54760 -46534 54768 -46446
rect 54802 -46448 54850 -46446
rect 54900 -46438 55200 -46368
rect 55870 -46370 55982 -46364
rect 55870 -46404 55882 -46370
rect 55970 -46404 55982 -46370
rect 55450 -46438 55810 -46408
rect 55870 -46410 55982 -46404
rect 56060 -46438 56300 -46360
rect 54900 -46442 55820 -46438
rect 56000 -46442 56300 -46438
rect 54900 -46448 55860 -46442
rect 54840 -46528 54850 -46448
rect 54802 -46534 54850 -46528
rect 54760 -46548 54850 -46534
rect 55130 -46454 55860 -46448
rect 55130 -46478 55820 -46454
rect 55130 -46496 55510 -46478
rect 55130 -46530 55142 -46496
rect 55494 -46498 55510 -46496
rect 55494 -46530 55506 -46498
rect 55130 -46536 55506 -46530
rect 53930 -46562 54730 -46556
rect 53930 -46596 53942 -46562
rect 54718 -46596 54730 -46562
rect 55020 -46582 55090 -46568
rect 53930 -46602 54730 -46596
rect 53940 -46608 54730 -46602
rect 54920 -46598 54980 -46588
rect 53940 -46648 54920 -46608
rect 53830 -46738 53920 -46728
rect 53830 -46848 53850 -46738
rect 53830 -46858 53920 -46848
rect 54320 -47148 54510 -46648
rect 54710 -46668 54920 -46648
rect 54910 -46678 54980 -46668
rect 55020 -46616 55046 -46582
rect 55080 -46616 55090 -46582
rect 55020 -46728 55090 -46616
rect 55142 -46662 55494 -46536
rect 55540 -46582 55620 -46568
rect 55540 -46616 55556 -46582
rect 55590 -46616 55620 -46582
rect 55130 -46668 55506 -46662
rect 55130 -46702 55142 -46668
rect 55494 -46702 55506 -46668
rect 55130 -46708 55506 -46702
rect 55000 -46738 55090 -46728
rect 55000 -46848 55090 -46838
rect 55540 -46728 55620 -46616
rect 55540 -46738 55630 -46728
rect 55630 -46838 55680 -46748
rect 55540 -46848 55680 -46838
rect 55274 -46938 55320 -46936
rect 55220 -46948 55320 -46938
rect 55220 -47124 55280 -47118
rect 55314 -47124 55320 -46948
rect 55220 -47128 55320 -47124
rect 55274 -47136 55320 -47128
rect 55362 -46948 55408 -46936
rect 55362 -47124 55368 -46948
rect 55402 -46958 55510 -46948
rect 55402 -47124 55410 -46958
rect 55362 -47128 55410 -47124
rect 55500 -47128 55510 -46958
rect 55362 -47136 55510 -47128
rect 55390 -47138 55510 -47136
rect 53636 -47188 53760 -47184
rect 53636 -47196 53682 -47188
rect 53940 -47208 54020 -47168
rect 54080 -47182 54860 -47148
rect 55311 -47174 55371 -47168
rect 53514 -47234 53626 -47228
rect 53514 -47238 53526 -47234
rect 53510 -47268 53526 -47238
rect 53614 -47238 53626 -47234
rect 53614 -47268 53630 -47238
rect 53510 -47328 53630 -47268
rect 53940 -47288 53950 -47208
rect 54010 -47238 54020 -47208
rect 54069 -47188 54869 -47182
rect 54069 -47222 54081 -47188
rect 54857 -47222 54869 -47188
rect 54069 -47228 54869 -47222
rect 54910 -47198 54980 -47188
rect 54010 -47250 54028 -47238
rect 54022 -47288 54028 -47250
rect 53940 -47300 54028 -47288
rect 53940 -47308 54020 -47300
rect 54910 -47308 54980 -47298
rect 55311 -47208 55324 -47174
rect 55358 -47208 55371 -47174
rect 54070 -47310 54870 -47308
rect 54069 -47316 54870 -47310
rect 54069 -47338 54081 -47316
rect 54041 -47350 54081 -47338
rect 54857 -47318 54870 -47316
rect 54857 -47350 54880 -47318
rect 55311 -47348 55371 -47208
rect 54041 -47358 54880 -47350
rect 55240 -47358 55371 -47348
rect 54041 -47368 55240 -47358
rect 53510 -47458 53630 -47448
rect 53961 -47408 55240 -47368
rect 35690 -47533 43500 -47500
rect 25860 -47558 43500 -47533
rect 35900 -47600 43500 -47558
rect 53961 -47606 54031 -47408
rect 54730 -47468 54860 -47458
rect 54730 -47488 54740 -47468
rect 54080 -47538 54740 -47488
rect 54069 -47544 54740 -47538
rect 54850 -47538 54860 -47468
rect 54850 -47544 54869 -47538
rect 54069 -47578 54081 -47544
rect 54857 -47578 54869 -47544
rect 54069 -47584 54869 -47578
rect 54911 -47594 54981 -47408
rect 55370 -47408 55371 -47358
rect 55240 -47428 55370 -47418
rect 55410 -47448 55510 -47138
rect 55410 -47558 55510 -47538
rect 55570 -47468 55680 -46848
rect 55780 -47230 55820 -46478
rect 55854 -47230 55860 -46454
rect 55780 -47238 55860 -47230
rect 55814 -47242 55860 -47238
rect 55992 -46454 56300 -46442
rect 55992 -47230 55998 -46454
rect 56032 -47228 56300 -46454
rect 56410 -46498 56430 -45899
rect 56380 -46675 56430 -46498
rect 56464 -46675 56470 -45899
rect 56380 -46687 56470 -46675
rect 56552 -45899 56750 -45887
rect 56552 -46675 56558 -45899
rect 56592 -46038 56750 -45899
rect 57066 -45880 57098 -45850
rect 57368 -45850 57372 -45764
rect 58896 -45759 59076 -45750
rect 58896 -45760 59084 -45759
rect 59156 -45760 59202 -45759
rect 57368 -45880 57396 -45850
rect 57066 -46010 57086 -45880
rect 57376 -46010 57396 -45880
rect 56592 -46675 56610 -46038
rect 57066 -46040 57396 -46010
rect 56860 -46190 57060 -46178
rect 56860 -46218 57236 -46190
rect 56860 -46348 56900 -46218
rect 57020 -46348 57236 -46218
rect 56860 -46388 57236 -46348
rect 57036 -46390 57236 -46388
rect 58556 -46280 58756 -46260
rect 58556 -46440 58576 -46280
rect 58736 -46440 58756 -46280
rect 58556 -46460 58756 -46440
rect 56552 -46678 56610 -46675
rect 57036 -46540 57446 -46530
rect 56552 -46687 56598 -46678
rect 57036 -46680 57056 -46540
rect 57416 -46680 57446 -46540
rect 56380 -46958 56440 -46687
rect 57036 -46700 57098 -46680
rect 56480 -46728 56550 -46718
rect 56480 -46798 56550 -46788
rect 57096 -46814 57098 -46734
rect 57368 -46700 57446 -46680
rect 57368 -46814 57372 -46734
rect 57096 -46830 57372 -46814
rect 58896 -46890 58926 -45760
rect 58966 -45771 59086 -45760
rect 58966 -46147 59044 -45771
rect 59078 -46147 59086 -45771
rect 58966 -46170 59086 -46147
rect 59156 -45771 59256 -45760
rect 59756 -45770 59826 -45740
rect 59966 -45752 59976 -45722
rect 60316 -45722 60346 -45716
rect 61036 -45720 61466 -45710
rect 60316 -45752 60326 -45722
rect 59966 -45760 60326 -45752
rect 59156 -46147 59162 -45771
rect 59196 -45840 59256 -45771
rect 59236 -45920 59256 -45840
rect 59196 -46040 59256 -45920
rect 59236 -46120 59256 -46040
rect 59196 -46147 59256 -46120
rect 59156 -46160 59256 -46147
rect 58966 -46480 59036 -46170
rect 59066 -46206 59176 -46200
rect 59066 -46210 59103 -46206
rect 59137 -46210 59176 -46206
rect 59066 -46280 59076 -46210
rect 59166 -46280 59176 -46210
rect 59066 -46290 59176 -46280
rect 59206 -46360 59256 -46160
rect 59376 -45790 59826 -45770
rect 59376 -45830 59476 -45790
rect 59656 -45830 59826 -45790
rect 59376 -45840 59826 -45830
rect 59376 -45890 59436 -45840
rect 59376 -46250 59386 -45890
rect 59426 -46250 59436 -45890
rect 59526 -45898 59576 -45870
rect 59526 -45932 59546 -45898
rect 59636 -45930 59706 -45870
rect 59580 -45932 59706 -45930
rect 59526 -45940 59706 -45932
rect 59476 -45982 59546 -45970
rect 59476 -46050 59502 -45982
rect 59476 -46158 59502 -46120
rect 59536 -46158 59546 -45982
rect 59476 -46170 59546 -46158
rect 59576 -45982 59636 -45970
rect 59576 -45990 59590 -45982
rect 59624 -45990 59636 -45982
rect 59576 -46170 59636 -46160
rect 59534 -46208 59592 -46202
rect 59534 -46210 59546 -46208
rect 59066 -46370 59176 -46360
rect 59066 -46440 59076 -46370
rect 59166 -46440 59176 -46370
rect 59066 -46442 59103 -46440
rect 59137 -46442 59176 -46440
rect 59066 -46450 59176 -46442
rect 59206 -46370 59266 -46360
rect 59206 -46450 59266 -46440
rect 59376 -46400 59436 -46250
rect 59516 -46242 59546 -46210
rect 59580 -46210 59592 -46208
rect 59666 -46210 59706 -45940
rect 59580 -46242 59706 -46210
rect 59516 -46280 59706 -46242
rect 59746 -45898 59936 -45870
rect 59746 -45932 59862 -45898
rect 59896 -45932 59936 -45898
rect 59746 -45940 59936 -45932
rect 61036 -45900 61206 -45720
rect 61346 -45900 61466 -45720
rect 76900 -45740 76920 -45640
rect 77060 -45740 77390 -45640
rect 76900 -45750 77390 -45740
rect 77510 -45750 77520 -45630
rect 77590 -45680 77600 -45610
rect 77710 -45680 77720 -45610
rect 77800 -45640 77820 -45590
rect 77860 -45640 77880 -45590
rect 78060 -45590 78070 -45480
rect 78140 -45590 78150 -45480
rect 78630 -45510 78750 -45500
rect 78060 -45600 78150 -45590
rect 78230 -45530 78310 -45520
rect 78230 -45590 78240 -45530
rect 78300 -45590 78310 -45530
rect 78230 -45600 78310 -45590
rect 78510 -45560 78590 -45540
rect 77800 -45650 77880 -45640
rect 78510 -45640 78530 -45560
rect 78570 -45640 78590 -45560
rect 78630 -45600 78640 -45510
rect 78740 -45600 78750 -45510
rect 78630 -45610 78750 -45600
rect 78800 -45550 78880 -45540
rect 78800 -45610 78810 -45550
rect 78870 -45610 78880 -45550
rect 78800 -45620 78880 -45610
rect 78510 -45670 78590 -45640
rect 77590 -45690 77720 -45680
rect 77970 -45680 78590 -45670
rect 77970 -45720 77990 -45680
rect 78030 -45720 78590 -45680
rect 79000 -45680 79020 -45370
rect 79070 -45380 79210 -45370
rect 79070 -45680 79080 -45380
rect 79190 -45680 79210 -45380
rect 79380 -45390 79710 -45360
rect 92000 -45400 95800 -44490
rect 79000 -45700 79210 -45680
rect 79980 -45430 80390 -45400
rect 77970 -45730 78590 -45720
rect 76900 -45760 77520 -45750
rect 77380 -45795 79060 -45760
rect 77380 -45829 77607 -45795
rect 77641 -45829 77699 -45795
rect 77733 -45829 77791 -45795
rect 77825 -45829 77883 -45795
rect 77917 -45829 77975 -45795
rect 78009 -45829 78067 -45795
rect 78101 -45829 78159 -45795
rect 78193 -45829 78251 -45795
rect 78285 -45829 78343 -45795
rect 78377 -45829 78435 -45795
rect 78469 -45829 78527 -45795
rect 78561 -45829 78619 -45795
rect 78653 -45829 78711 -45795
rect 78745 -45829 78803 -45795
rect 78837 -45829 78895 -45795
rect 78929 -45829 78987 -45795
rect 79021 -45829 79060 -45795
rect 77380 -45880 79060 -45829
rect 79980 -45810 80010 -45430
rect 80360 -45530 80390 -45430
rect 80360 -45730 80590 -45530
rect 80360 -45810 80390 -45730
rect 79980 -45840 80390 -45810
rect 61036 -45940 61466 -45900
rect 59746 -46200 59776 -45940
rect 60286 -45950 60476 -45940
rect 59806 -45982 59866 -45970
rect 59806 -46000 59818 -45982
rect 59852 -46000 59866 -45982
rect 59806 -46158 59818 -46140
rect 59852 -46158 59866 -46140
rect 59806 -46170 59866 -46158
rect 59900 -45980 60016 -45970
rect 59900 -45982 59916 -45980
rect 59900 -46158 59906 -45982
rect 59900 -46160 59916 -46158
rect 60006 -46160 60016 -45980
rect 60286 -46090 60306 -45950
rect 60456 -46090 60476 -45950
rect 61176 -46000 61386 -45980
rect 60286 -46100 60476 -46090
rect 61026 -46020 61136 -46010
rect 59900 -46170 60016 -46160
rect 60076 -46157 60196 -46120
rect 60076 -46191 60127 -46157
rect 60161 -46191 60196 -46157
rect 59746 -46208 59926 -46200
rect 59746 -46210 59862 -46208
rect 59896 -46210 59926 -46208
rect 59746 -46280 59826 -46210
rect 59916 -46280 59926 -46210
rect 59746 -46290 59926 -46280
rect 60076 -46249 60196 -46191
rect 60336 -46160 60446 -46100
rect 60336 -46200 60366 -46160
rect 60406 -46200 60446 -46160
rect 60636 -46157 60816 -46120
rect 60636 -46191 60671 -46157
rect 60705 -46191 60747 -46157
rect 60781 -46191 60816 -46157
rect 60076 -46280 60127 -46249
rect 60161 -46280 60196 -46249
rect 59736 -46370 59936 -46360
rect 58966 -46501 59086 -46480
rect 58966 -46877 59044 -46501
rect 59078 -46877 59086 -46501
rect 58966 -46890 59086 -46877
rect 59156 -46490 59202 -46489
rect 59156 -46501 59236 -46490
rect 59156 -46877 59162 -46501
rect 59196 -46530 59236 -46501
rect 59226 -46610 59236 -46530
rect 59196 -46760 59236 -46610
rect 59226 -46840 59236 -46760
rect 59196 -46877 59236 -46840
rect 59376 -46770 59386 -46400
rect 59426 -46770 59436 -46400
rect 59516 -46411 59706 -46370
rect 59516 -46445 59545 -46411
rect 59579 -46445 59706 -46411
rect 59516 -46450 59706 -46445
rect 59533 -46451 59591 -46450
rect 59466 -46495 59546 -46480
rect 59586 -46483 59646 -46480
rect 59466 -46530 59501 -46495
rect 59466 -46671 59501 -46610
rect 59535 -46671 59546 -46495
rect 59466 -46680 59546 -46671
rect 59583 -46495 59646 -46483
rect 59583 -46510 59589 -46495
rect 59623 -46510 59646 -46495
rect 59583 -46650 59586 -46510
rect 59583 -46671 59589 -46650
rect 59623 -46671 59646 -46650
rect 59583 -46680 59646 -46671
rect 59495 -46683 59541 -46680
rect 59583 -46683 59629 -46680
rect 59533 -46720 59591 -46715
rect 59676 -46720 59706 -46450
rect 59376 -46810 59436 -46770
rect 59506 -46780 59516 -46720
rect 59596 -46780 59706 -46720
rect 59736 -46440 59826 -46370
rect 59926 -46440 59936 -46370
rect 59736 -46445 59861 -46440
rect 59895 -46445 59936 -46440
rect 59736 -46450 59936 -46445
rect 60076 -46440 60096 -46280
rect 60176 -46440 60196 -46280
rect 59736 -46720 59766 -46450
rect 59849 -46451 59907 -46450
rect 60076 -46467 60127 -46440
rect 60161 -46467 60196 -46440
rect 59796 -46483 59856 -46480
rect 59796 -46490 59857 -46483
rect 59856 -46670 59857 -46490
rect 59796 -46671 59817 -46670
rect 59851 -46671 59857 -46670
rect 59796 -46680 59857 -46671
rect 59811 -46683 59857 -46680
rect 59899 -46490 59945 -46483
rect 59899 -46495 59916 -46490
rect 59899 -46671 59905 -46495
rect 59899 -46680 59916 -46671
rect 60006 -46680 60016 -46490
rect 60076 -46525 60196 -46467
rect 60346 -46250 60426 -46200
rect 60346 -46290 60366 -46250
rect 60406 -46290 60426 -46250
rect 60346 -46340 60426 -46290
rect 60346 -46380 60366 -46340
rect 60406 -46380 60426 -46340
rect 60346 -46420 60426 -46380
rect 60346 -46460 60366 -46420
rect 60406 -46460 60426 -46420
rect 60346 -46470 60426 -46460
rect 60636 -46249 60816 -46191
rect 60636 -46283 60671 -46249
rect 60705 -46283 60747 -46249
rect 60781 -46283 60816 -46249
rect 60636 -46341 60816 -46283
rect 60636 -46375 60671 -46341
rect 60705 -46375 60747 -46341
rect 60781 -46375 60816 -46341
rect 60636 -46433 60816 -46375
rect 60636 -46467 60671 -46433
rect 60705 -46467 60747 -46433
rect 60781 -46467 60816 -46433
rect 60076 -46559 60127 -46525
rect 60161 -46559 60196 -46525
rect 60076 -46590 60196 -46559
rect 60276 -46510 60546 -46500
rect 60276 -46525 60476 -46510
rect 60276 -46559 60297 -46525
rect 60331 -46559 60369 -46525
rect 60405 -46559 60449 -46525
rect 60276 -46570 60476 -46559
rect 60536 -46570 60546 -46510
rect 60276 -46580 60546 -46570
rect 60636 -46525 60816 -46467
rect 61026 -46130 61036 -46020
rect 61126 -46130 61136 -46020
rect 61176 -46080 61196 -46000
rect 61366 -46080 61386 -46000
rect 61176 -46100 61386 -46080
rect 61026 -46160 61136 -46130
rect 61026 -46200 61046 -46160
rect 61086 -46200 61136 -46160
rect 61026 -46250 61136 -46200
rect 61026 -46290 61046 -46250
rect 61086 -46290 61136 -46250
rect 61026 -46340 61136 -46290
rect 61026 -46380 61046 -46340
rect 61086 -46380 61136 -46340
rect 61026 -46420 61136 -46380
rect 61026 -46460 61046 -46420
rect 61086 -46460 61136 -46420
rect 61026 -46480 61136 -46460
rect 61256 -46157 61366 -46100
rect 61256 -46191 61291 -46157
rect 61325 -46191 61366 -46157
rect 61256 -46249 61366 -46191
rect 61256 -46250 61291 -46249
rect 61325 -46250 61366 -46249
rect 61256 -46460 61276 -46250
rect 61356 -46460 61366 -46250
rect 61256 -46467 61291 -46460
rect 61325 -46467 61366 -46460
rect 60636 -46559 60671 -46525
rect 60705 -46559 60747 -46525
rect 60781 -46559 60816 -46525
rect 60636 -46640 60816 -46559
rect 60966 -46524 61177 -46510
rect 60966 -46525 61129 -46524
rect 60966 -46559 60980 -46525
rect 61015 -46559 61053 -46525
rect 61088 -46558 61129 -46525
rect 61164 -46558 61177 -46524
rect 61088 -46559 61177 -46558
rect 60966 -46590 61177 -46559
rect 61256 -46525 61366 -46467
rect 61256 -46559 61291 -46525
rect 61325 -46559 61366 -46525
rect 61256 -46590 61366 -46559
rect 73180 -46400 73380 -46180
rect 73180 -46590 73220 -46400
rect 73340 -46590 73380 -46400
rect 60466 -46650 60546 -46640
rect 59899 -46683 59945 -46680
rect 60466 -46710 60476 -46650
rect 60536 -46710 60546 -46650
rect 59849 -46720 59907 -46715
rect 60466 -46720 60546 -46710
rect 60606 -46650 60826 -46640
rect 60606 -46710 60616 -46650
rect 60736 -46710 60756 -46650
rect 60816 -46710 60826 -46650
rect 60606 -46720 60826 -46710
rect 60886 -46650 60966 -46640
rect 60886 -46710 60896 -46650
rect 60956 -46710 60966 -46650
rect 60886 -46720 60966 -46710
rect 59736 -46721 59926 -46720
rect 59736 -46755 59861 -46721
rect 59895 -46755 59926 -46721
rect 59736 -46780 59926 -46755
rect 60636 -46770 60816 -46720
rect 59376 -46820 59826 -46810
rect 59376 -46860 59476 -46820
rect 59646 -46860 59826 -46820
rect 59376 -46870 59826 -46860
rect 59156 -46890 59236 -46877
rect 58896 -46900 59086 -46890
rect 56380 -46968 57000 -46958
rect 57356 -46964 57676 -46950
rect 56440 -46974 57000 -46968
rect 57314 -46970 57676 -46964
rect 56440 -46994 57178 -46974
rect 56440 -47044 57118 -46994
rect 57168 -47044 57178 -46994
rect 57314 -47010 57326 -46970
rect 57376 -47010 57676 -46970
rect 57314 -47016 57676 -47010
rect 57356 -47030 57676 -47016
rect 56440 -47054 57178 -47044
rect 56440 -47088 57000 -47054
rect 57112 -47056 57174 -47054
rect 56380 -47158 57000 -47088
rect 56032 -47230 56038 -47228
rect 55992 -47242 56038 -47230
rect 55880 -47274 55970 -47268
rect 55870 -47278 55982 -47274
rect 55870 -47320 55880 -47278
rect 55970 -47320 55982 -47278
rect 55880 -47368 55970 -47358
rect 56120 -47398 56300 -47228
rect 57096 -47309 57372 -47278
rect 57096 -47343 57125 -47309
rect 57159 -47343 57217 -47309
rect 57251 -47343 57309 -47309
rect 57343 -47320 57372 -47309
rect 57343 -47343 57376 -47320
rect 57096 -47380 57376 -47343
rect 57066 -47390 57376 -47380
rect 56426 -47398 57376 -47390
rect 56120 -47408 57376 -47398
rect 56014 -47458 56086 -47446
rect 55570 -47578 55830 -47468
rect 53961 -47644 53988 -47606
rect 54022 -47644 54031 -47606
rect 53961 -47658 54031 -47644
rect 54910 -47606 54981 -47594
rect 54910 -47644 54916 -47606
rect 54950 -47644 54981 -47606
rect 54910 -47656 54981 -47644
rect 54911 -47658 54981 -47656
rect 55220 -47618 55330 -47608
rect 54069 -47672 54869 -47666
rect 54069 -47706 54081 -47672
rect 54857 -47678 54869 -47672
rect 54857 -47706 54880 -47678
rect 54069 -47712 54880 -47706
rect 54090 -47788 54880 -47712
rect 55330 -47718 55380 -47618
rect 55330 -47728 55480 -47718
rect 55220 -47738 55480 -47728
rect 55280 -47752 55480 -47738
rect 55280 -47758 55488 -47752
rect 55280 -47778 55300 -47758
rect 54090 -47888 54150 -47788
rect 54840 -47888 54880 -47788
rect 55288 -47792 55300 -47778
rect 55476 -47792 55488 -47758
rect 55530 -47778 55610 -47768
rect 55288 -47798 55488 -47792
rect 55520 -47802 55530 -47790
rect 55520 -47836 55526 -47802
rect 55288 -47846 55488 -47840
rect 55288 -47880 55300 -47846
rect 55476 -47880 55488 -47846
rect 55520 -47848 55530 -47836
rect 55530 -47878 55610 -47868
rect 55288 -47886 55488 -47880
rect 54090 -47908 54140 -47888
rect 35900 -48052 42600 -48000
rect 25860 -48071 42600 -48052
rect 25860 -48468 25882 -48071
rect 26996 -48468 27124 -48071
rect 28238 -48468 28366 -48071
rect 29480 -48468 29608 -48071
rect 30722 -48468 30850 -48071
rect 31964 -48468 32092 -48071
rect 33206 -48468 33334 -48071
rect 34448 -48468 34576 -48071
rect 35690 -48100 42600 -48071
rect 35690 -48468 36000 -48100
rect 25860 -48734 36000 -48468
rect 25860 -49131 25882 -48734
rect 26996 -49131 27124 -48734
rect 28238 -49131 28366 -48734
rect 29480 -49131 29608 -48734
rect 30722 -49131 30850 -48734
rect 31964 -49131 32092 -48734
rect 33206 -49131 33334 -48734
rect 34448 -49131 34576 -48734
rect 35690 -49100 36000 -48734
rect 42500 -49100 42600 -48100
rect 54100 -48148 54140 -47908
rect 54850 -48148 54880 -47888
rect 55300 -47928 55470 -47886
rect 55300 -48068 55320 -47928
rect 55470 -48014 55482 -47942
rect 55300 -48078 55470 -48068
rect 54100 -48188 54880 -48148
rect 55710 -48398 55830 -47578
rect 56014 -47608 56020 -47458
rect 56080 -47608 56086 -47458
rect 56014 -47620 56086 -47608
rect 56120 -47608 56170 -47408
rect 56390 -47460 57376 -47408
rect 56390 -47468 57156 -47460
rect 56390 -47608 56654 -47468
rect 56120 -47658 56654 -47608
rect 56306 -47686 56654 -47658
rect 56998 -47620 57156 -47468
rect 57316 -47620 57376 -47460
rect 56998 -47686 57376 -47620
rect 56306 -48100 57376 -47686
rect 57556 -47810 57676 -47030
rect 58896 -47060 58986 -46900
rect 59756 -46920 59826 -46870
rect 59066 -46936 59176 -46930
rect 59066 -46940 59103 -46936
rect 59137 -46940 59176 -46936
rect 59066 -47000 59076 -46940
rect 59166 -47000 59176 -46940
rect 59066 -47010 59176 -47000
rect 58896 -47430 58926 -47060
rect 58966 -47430 58986 -47130
rect 59116 -47060 59506 -47040
rect 59116 -47130 59146 -47060
rect 59226 -47130 59276 -47060
rect 59356 -47130 59396 -47060
rect 59476 -47130 59506 -47060
rect 59116 -47148 59506 -47130
rect 59646 -47060 59716 -47040
rect 59706 -47120 59716 -47060
rect 59646 -47130 59716 -47120
rect 59113 -47154 59513 -47148
rect 59113 -47188 59125 -47154
rect 59501 -47188 59513 -47154
rect 59113 -47194 59513 -47188
rect 59546 -47200 59616 -47190
rect 59246 -47256 59256 -47230
rect 59113 -47262 59256 -47256
rect 59366 -47256 59376 -47230
rect 59366 -47262 59513 -47256
rect 59016 -47300 59076 -47280
rect 59113 -47296 59125 -47262
rect 59501 -47296 59513 -47262
rect 59606 -47260 59616 -47200
rect 59546 -47270 59616 -47260
rect 59113 -47302 59513 -47296
rect 59016 -47390 59076 -47360
rect 59113 -47370 59513 -47364
rect 59113 -47404 59125 -47370
rect 59501 -47404 59513 -47370
rect 59113 -47410 59513 -47404
rect 58896 -47500 58906 -47430
rect 58896 -47520 58986 -47500
rect 59116 -47430 59516 -47410
rect 59116 -47500 59146 -47430
rect 59226 -47500 59276 -47430
rect 59356 -47500 59396 -47430
rect 59476 -47500 59516 -47430
rect 59116 -47520 59516 -47500
rect 59646 -47430 59656 -47130
rect 59706 -47430 59716 -47130
rect 59756 -47100 59766 -46920
rect 59806 -47100 59826 -46920
rect 59956 -46920 60336 -46910
rect 59956 -46934 59966 -46920
rect 59946 -46940 59966 -46934
rect 60326 -46934 60336 -46920
rect 60326 -46940 60346 -46934
rect 59856 -46980 59916 -46970
rect 59946 -46974 59958 -46940
rect 60334 -46974 60346 -46940
rect 61056 -46940 61176 -46590
rect 73180 -46600 73380 -46590
rect 73430 -46400 73630 -46180
rect 73430 -46590 73470 -46400
rect 73590 -46590 73630 -46400
rect 73430 -46600 73630 -46590
rect 73680 -46400 73880 -46180
rect 73680 -46590 73720 -46400
rect 73840 -46590 73880 -46400
rect 73680 -46600 73880 -46590
rect 73930 -46400 74130 -46180
rect 73930 -46590 73970 -46400
rect 74090 -46590 74130 -46400
rect 73930 -46600 74130 -46590
rect 74180 -46400 74380 -46180
rect 74180 -46590 74220 -46400
rect 74340 -46590 74380 -46400
rect 74180 -46600 74380 -46590
rect 74430 -46400 74630 -46180
rect 74430 -46590 74470 -46400
rect 74590 -46590 74630 -46400
rect 74430 -46600 74630 -46590
rect 74680 -46400 74880 -46180
rect 74680 -46590 74720 -46400
rect 74840 -46590 74880 -46400
rect 74680 -46600 74880 -46590
rect 74930 -46400 75130 -46180
rect 74930 -46590 74970 -46400
rect 75090 -46590 75130 -46400
rect 74930 -46600 75130 -46590
rect 75180 -46190 75560 -46180
rect 75180 -46310 75390 -46190
rect 75550 -46310 75560 -46190
rect 75180 -46320 75560 -46310
rect 75180 -46400 75380 -46320
rect 76880 -46380 77260 -46376
rect 75180 -46590 75220 -46400
rect 75340 -46590 75380 -46400
rect 75500 -46390 77260 -46380
rect 75500 -46411 77110 -46390
rect 75500 -46445 75535 -46411
rect 75569 -46445 75627 -46411
rect 75661 -46445 75719 -46411
rect 75753 -46445 75811 -46411
rect 75845 -46445 75903 -46411
rect 75937 -46445 75995 -46411
rect 76029 -46445 76085 -46411
rect 76119 -46445 76177 -46411
rect 76211 -46445 76269 -46411
rect 76303 -46445 76361 -46411
rect 76395 -46445 76453 -46411
rect 76487 -46445 76545 -46411
rect 76579 -46445 76637 -46411
rect 76671 -46445 76729 -46411
rect 76763 -46445 76821 -46411
rect 76855 -46445 77110 -46411
rect 75500 -46450 77110 -46445
rect 75500 -46480 76920 -46450
rect 75661 -46540 75728 -46534
rect 75180 -46600 75380 -46590
rect 75660 -46557 75728 -46540
rect 75660 -46591 75670 -46557
rect 75704 -46591 75728 -46557
rect 75660 -46610 75728 -46591
rect 75933 -46560 76011 -46532
rect 76765 -46538 76817 -46532
rect 75933 -46594 75942 -46560
rect 75976 -46594 76011 -46560
rect 75933 -46610 76011 -46594
rect 76204 -46559 76268 -46543
rect 76204 -46593 76217 -46559
rect 76251 -46593 76268 -46559
rect 76204 -46610 76268 -46593
rect 76483 -46559 76549 -46546
rect 76483 -46593 76492 -46559
rect 76526 -46593 76549 -46559
rect 75400 -46630 75480 -46620
rect 75660 -46623 75764 -46610
rect 75390 -46636 75410 -46630
rect 73710 -46688 73723 -46636
rect 73840 -46688 75410 -46636
rect 75400 -46690 75410 -46688
rect 75470 -46636 75490 -46630
rect 75560 -46636 75630 -46630
rect 75470 -46650 75630 -46636
rect 75470 -46688 75580 -46650
rect 75470 -46690 75480 -46688
rect 75400 -46700 75480 -46690
rect 75560 -46690 75580 -46688
rect 75620 -46690 75630 -46650
rect 75560 -46710 75630 -46690
rect 75660 -46649 75673 -46623
rect 75660 -46683 75670 -46649
rect 75660 -46701 75673 -46683
rect 75751 -46701 75764 -46623
rect 75660 -46714 75764 -46701
rect 75840 -46622 75900 -46621
rect 75840 -46643 75902 -46622
rect 75840 -46677 75862 -46643
rect 75896 -46677 75902 -46643
rect 75840 -46703 75902 -46677
rect 75933 -46623 76037 -46610
rect 75933 -46701 75946 -46623
rect 76024 -46701 76037 -46623
rect 75660 -46738 75730 -46714
rect 75660 -46772 75670 -46738
rect 75704 -46772 75730 -46738
rect 74210 -46800 75440 -46790
rect 75660 -46800 75730 -46772
rect 74210 -46880 74220 -46800
rect 74340 -46830 75440 -46800
rect 75840 -46830 75900 -46703
rect 75933 -46714 76037 -46701
rect 76102 -46623 76167 -46610
rect 76204 -46623 76323 -46610
rect 76483 -46623 76549 -46593
rect 76759 -46561 76817 -46538
rect 76759 -46595 76768 -46561
rect 76802 -46595 76817 -46561
rect 76759 -46623 76817 -46595
rect 76882 -46570 76920 -46480
rect 77060 -46570 77110 -46450
rect 76882 -46610 77110 -46570
rect 77220 -46610 77260 -46390
rect 76882 -46620 77260 -46610
rect 76167 -46701 76168 -46636
rect 76204 -46650 76232 -46623
rect 76204 -46684 76224 -46650
rect 76204 -46701 76232 -46684
rect 76310 -46701 76323 -46623
rect 76102 -46714 76167 -46701
rect 76204 -46714 76323 -46701
rect 76362 -46634 76453 -46623
rect 76362 -46640 76455 -46634
rect 76362 -46700 76380 -46640
rect 76440 -46700 76455 -46640
rect 76362 -46703 76455 -46700
rect 76483 -46636 76596 -46623
rect 76483 -46649 76505 -46636
rect 76483 -46683 76497 -46649
rect 76483 -46701 76505 -46683
rect 76583 -46701 76596 -46636
rect 76362 -46714 76453 -46703
rect 76483 -46714 76596 -46701
rect 76635 -46636 76726 -46623
rect 76635 -46714 76648 -46636
rect 75933 -46743 76011 -46714
rect 75933 -46777 75943 -46743
rect 75977 -46777 76011 -46743
rect 75933 -46818 76011 -46777
rect 76204 -46744 76268 -46714
rect 76370 -46720 76450 -46714
rect 76204 -46778 76215 -46744
rect 76249 -46778 76268 -46744
rect 76204 -46816 76268 -46778
rect 76483 -46743 76549 -46714
rect 76635 -46727 76726 -46714
rect 76759 -46636 76843 -46623
rect 76759 -46650 76791 -46636
rect 76759 -46684 76772 -46650
rect 76759 -46714 76791 -46684
rect 76759 -46727 76843 -46714
rect 76483 -46777 76492 -46743
rect 76526 -46777 76549 -46743
rect 76483 -46794 76549 -46777
rect 76759 -46743 76817 -46727
rect 76759 -46777 76768 -46743
rect 76802 -46777 76817 -46743
rect 76759 -46796 76817 -46777
rect 74340 -46870 75900 -46830
rect 76204 -46850 76218 -46816
rect 76252 -46850 76268 -46816
rect 76204 -46863 76268 -46850
rect 76765 -46870 76817 -46796
rect 76850 -46830 79050 -46800
rect 76850 -46840 77170 -46830
rect 74340 -46880 75440 -46870
rect 74210 -46890 75440 -46880
rect 59946 -46980 59966 -46974
rect 60326 -46980 60346 -46974
rect 60376 -46980 60436 -46960
rect 59956 -46990 60336 -46980
rect 59856 -47060 59916 -47040
rect 59946 -47048 60346 -47042
rect 59756 -47140 59826 -47100
rect 59946 -47082 59958 -47048
rect 60334 -47082 60346 -47048
rect 60376 -47060 60436 -47040
rect 61126 -47040 61176 -46940
rect 61056 -47070 61176 -47040
rect 72810 -46900 73050 -46890
rect 59946 -47088 60346 -47082
rect 72810 -47080 72820 -46900
rect 73040 -47080 73050 -46900
rect 76850 -46920 76930 -46840
rect 75500 -46955 76930 -46920
rect 75500 -46989 75535 -46955
rect 75569 -46989 75627 -46955
rect 75661 -46989 75719 -46955
rect 75753 -46989 75811 -46955
rect 75845 -46989 75903 -46955
rect 75937 -46989 75995 -46955
rect 76029 -46989 76085 -46955
rect 76119 -46989 76177 -46955
rect 76211 -46989 76269 -46955
rect 76303 -46989 76361 -46955
rect 76395 -46989 76453 -46955
rect 76487 -46989 76545 -46955
rect 76579 -46989 76637 -46955
rect 76671 -46989 76729 -46955
rect 76763 -46989 76821 -46955
rect 76855 -46989 76930 -46955
rect 75500 -47020 76930 -46989
rect 59946 -47140 60336 -47088
rect 72810 -47090 73050 -47080
rect 76850 -47080 76930 -47020
rect 77040 -47080 77170 -46840
rect 77430 -47080 79050 -46830
rect 76850 -47081 79050 -47080
rect 76850 -47115 77607 -47081
rect 77641 -47115 77699 -47081
rect 77733 -47115 77791 -47081
rect 77825 -47115 77883 -47081
rect 77917 -47115 77975 -47081
rect 78009 -47115 78067 -47081
rect 78101 -47115 78159 -47081
rect 78193 -47115 78251 -47081
rect 78285 -47115 78343 -47081
rect 78377 -47115 78435 -47081
rect 78469 -47115 78527 -47081
rect 78561 -47115 78619 -47081
rect 78653 -47115 78711 -47081
rect 78745 -47115 78803 -47081
rect 78837 -47115 78895 -47081
rect 78929 -47115 78987 -47081
rect 79021 -47115 79050 -47081
rect 76850 -47120 79050 -47115
rect 59756 -47160 60536 -47140
rect 77578 -47146 79050 -47120
rect 59756 -47200 59866 -47160
rect 60426 -47200 60536 -47160
rect 59756 -47210 60536 -47200
rect 59796 -47320 59806 -47210
rect 59916 -47320 59926 -47210
rect 59796 -47330 59926 -47320
rect 60436 -47230 60536 -47210
rect 73460 -47220 73480 -47160
rect 73580 -47170 77540 -47160
rect 73580 -47210 77430 -47170
rect 77520 -47210 77540 -47170
rect 78600 -47180 79050 -47146
rect 82794 -46878 91444 -46848
rect 73580 -47220 77540 -47210
rect 60436 -47350 60446 -47230
rect 60526 -47350 60536 -47230
rect 60436 -47360 60536 -47350
rect 72600 -47230 73050 -47220
rect 72600 -47410 72820 -47230
rect 73040 -47410 73050 -47230
rect 73710 -47330 73730 -47270
rect 73830 -47310 77690 -47270
rect 80050 -47310 80460 -47280
rect 73830 -47320 77840 -47310
rect 73830 -47330 77780 -47320
rect 77580 -47360 77780 -47330
rect 77820 -47360 77840 -47320
rect 77580 -47370 77840 -47360
rect 78570 -47360 78650 -47350
rect 72600 -47420 73050 -47410
rect 73210 -47380 77510 -47370
rect 59646 -47440 59716 -47430
rect 59706 -47500 59716 -47440
rect 73210 -47440 73230 -47380
rect 73330 -47400 77510 -47380
rect 77870 -47390 77970 -47370
rect 77860 -47400 77900 -47390
rect 73330 -47430 77900 -47400
rect 77940 -47430 77970 -47390
rect 73330 -47440 77970 -47430
rect 73210 -47450 77970 -47440
rect 78140 -47380 78220 -47370
rect 78270 -47380 78350 -47370
rect 78140 -47440 78150 -47380
rect 78210 -47440 78220 -47380
rect 78140 -47450 78220 -47440
rect 78250 -47440 78280 -47380
rect 78340 -47390 78430 -47380
rect 78340 -47430 78370 -47390
rect 78410 -47430 78430 -47390
rect 78570 -47420 78580 -47360
rect 78640 -47420 78650 -47360
rect 78570 -47430 78650 -47420
rect 78790 -47370 78860 -47360
rect 78790 -47430 78800 -47370
rect 78340 -47440 78430 -47430
rect 78790 -47440 78860 -47430
rect 79060 -47380 79270 -47370
rect 78250 -47443 78410 -47440
rect 78270 -47450 78350 -47443
rect 59646 -47520 59716 -47500
rect 77220 -47540 77230 -47480
rect 77310 -47540 77320 -47480
rect 77220 -47550 77320 -47540
rect 77400 -47500 77560 -47480
rect 77400 -47590 77420 -47500
rect 76900 -47610 77420 -47590
rect 72600 -47720 73050 -47710
rect 58806 -47810 59356 -47780
rect 57556 -47820 59356 -47810
rect 57556 -47960 58986 -47820
rect 59126 -47960 59356 -47820
rect 59846 -47790 60256 -47780
rect 59846 -47900 59996 -47790
rect 60106 -47900 60256 -47790
rect 72600 -47900 72820 -47720
rect 73040 -47900 73050 -47720
rect 76900 -47760 76920 -47610
rect 77060 -47620 77420 -47610
rect 77540 -47590 77560 -47500
rect 79060 -47550 79080 -47380
rect 79140 -47390 79270 -47380
rect 79250 -47550 79270 -47390
rect 79060 -47560 79270 -47550
rect 77540 -47620 79050 -47590
rect 77060 -47625 79050 -47620
rect 77060 -47659 77607 -47625
rect 77641 -47659 77699 -47625
rect 77733 -47659 77791 -47625
rect 77825 -47659 77883 -47625
rect 77917 -47659 77975 -47625
rect 78009 -47659 78067 -47625
rect 78101 -47659 78159 -47625
rect 78193 -47659 78251 -47625
rect 78285 -47659 78343 -47625
rect 78377 -47659 78435 -47625
rect 78469 -47659 78527 -47625
rect 78561 -47659 78619 -47625
rect 78653 -47659 78711 -47625
rect 78745 -47659 78803 -47625
rect 78837 -47659 78895 -47625
rect 78929 -47659 78987 -47625
rect 79021 -47659 79050 -47625
rect 80050 -47620 80080 -47310
rect 80430 -47370 80460 -47310
rect 80430 -47570 80660 -47370
rect 82794 -47448 82824 -46878
rect 91414 -47448 91444 -46878
rect 82794 -47518 91444 -47448
rect 80430 -47620 80460 -47570
rect 80050 -47650 80460 -47620
rect 77060 -47700 79050 -47659
rect 82794 -47688 83454 -47518
rect 83624 -47688 85154 -47518
rect 85324 -47688 86534 -47518
rect 86704 -47688 87824 -47518
rect 87994 -47688 89344 -47518
rect 89514 -47688 90754 -47518
rect 90924 -47688 91444 -47518
rect 77060 -47760 77420 -47700
rect 76900 -47780 77420 -47760
rect 77160 -47820 77270 -47810
rect 77160 -47890 77170 -47820
rect 77260 -47890 77270 -47820
rect 77400 -47820 77420 -47780
rect 77540 -47711 79050 -47700
rect 77540 -47745 77607 -47711
rect 77641 -47745 77699 -47711
rect 77733 -47745 77791 -47711
rect 77825 -47745 77883 -47711
rect 77917 -47745 77975 -47711
rect 78009 -47745 78067 -47711
rect 78101 -47745 79050 -47711
rect 77540 -47780 79050 -47745
rect 80050 -47720 80460 -47690
rect 77540 -47820 77560 -47780
rect 77400 -47840 77560 -47820
rect 78140 -47830 78220 -47810
rect 77160 -47900 77270 -47890
rect 57556 -48010 59356 -47960
rect 58806 -48090 59356 -48010
rect 55710 -48400 55910 -48398
rect 55400 -48500 56200 -48400
rect 59600 -48500 60500 -47900
rect 72600 -47910 73050 -47900
rect 77690 -47930 77960 -47920
rect 74210 -47990 74230 -47930
rect 74330 -47940 77960 -47930
rect 74330 -47960 77900 -47940
rect 74330 -47990 77700 -47960
rect 77860 -47980 77900 -47960
rect 77940 -47980 77960 -47940
rect 77860 -47990 77960 -47980
rect 72600 -48000 73050 -47990
rect 72600 -48180 72820 -48000
rect 73040 -48180 73050 -48000
rect 77750 -48000 77830 -47990
rect 77750 -48020 77770 -48000
rect 74710 -48080 74730 -48020
rect 74830 -48040 77770 -48020
rect 77810 -48040 77830 -48000
rect 74830 -48080 77830 -48040
rect 78140 -48120 78150 -47830
rect 78210 -48120 78220 -47830
rect 78140 -48140 78220 -48120
rect 80050 -48100 80080 -47720
rect 80430 -47820 80460 -47720
rect 82794 -47731 91444 -47688
rect 82794 -47765 82867 -47731
rect 82901 -47765 82959 -47731
rect 82993 -47765 83051 -47731
rect 83085 -47765 83143 -47731
rect 83177 -47765 83235 -47731
rect 83269 -47765 83327 -47731
rect 83361 -47765 83419 -47731
rect 83453 -47765 83511 -47731
rect 83545 -47765 83603 -47731
rect 83637 -47765 83695 -47731
rect 83729 -47765 83787 -47731
rect 83821 -47765 83879 -47731
rect 83913 -47765 83971 -47731
rect 84005 -47765 84063 -47731
rect 84097 -47765 84155 -47731
rect 84189 -47765 84247 -47731
rect 84281 -47765 84339 -47731
rect 84373 -47765 84431 -47731
rect 84465 -47765 84523 -47731
rect 84557 -47765 84615 -47731
rect 84649 -47765 84707 -47731
rect 84741 -47765 84799 -47731
rect 84833 -47765 84891 -47731
rect 84925 -47765 84983 -47731
rect 85017 -47765 85075 -47731
rect 85109 -47765 85167 -47731
rect 85201 -47765 85259 -47731
rect 85293 -47765 85351 -47731
rect 85385 -47765 85443 -47731
rect 85477 -47765 85535 -47731
rect 85569 -47765 85627 -47731
rect 85661 -47765 85719 -47731
rect 85753 -47765 85811 -47731
rect 85845 -47765 85903 -47731
rect 85937 -47765 85995 -47731
rect 86029 -47765 86087 -47731
rect 86121 -47765 86179 -47731
rect 86213 -47765 86271 -47731
rect 86305 -47765 86363 -47731
rect 86397 -47765 86455 -47731
rect 86489 -47765 86547 -47731
rect 86581 -47765 86639 -47731
rect 86673 -47765 86731 -47731
rect 86765 -47765 86823 -47731
rect 86857 -47765 86915 -47731
rect 86949 -47765 87007 -47731
rect 87041 -47765 87099 -47731
rect 87133 -47765 87191 -47731
rect 87225 -47765 87283 -47731
rect 87317 -47765 87375 -47731
rect 87409 -47765 87467 -47731
rect 87501 -47765 87559 -47731
rect 87593 -47765 87651 -47731
rect 87685 -47765 87743 -47731
rect 87777 -47765 87835 -47731
rect 87869 -47765 87927 -47731
rect 87961 -47765 88019 -47731
rect 88053 -47765 88111 -47731
rect 88145 -47765 88203 -47731
rect 88237 -47765 88295 -47731
rect 88329 -47765 88387 -47731
rect 88421 -47765 88479 -47731
rect 88513 -47765 88571 -47731
rect 88605 -47765 88663 -47731
rect 88697 -47765 88755 -47731
rect 88789 -47765 88847 -47731
rect 88881 -47765 88939 -47731
rect 88973 -47765 89031 -47731
rect 89065 -47765 89123 -47731
rect 89157 -47765 89215 -47731
rect 89249 -47765 89307 -47731
rect 89341 -47765 89399 -47731
rect 89433 -47765 89491 -47731
rect 89525 -47765 89583 -47731
rect 89617 -47765 89675 -47731
rect 89709 -47765 89767 -47731
rect 89801 -47765 89859 -47731
rect 89893 -47765 89951 -47731
rect 89985 -47765 90043 -47731
rect 90077 -47765 90135 -47731
rect 90169 -47765 90227 -47731
rect 90261 -47765 90319 -47731
rect 90353 -47765 90411 -47731
rect 90445 -47765 90503 -47731
rect 90537 -47765 90595 -47731
rect 90629 -47765 90687 -47731
rect 90721 -47765 90779 -47731
rect 90813 -47765 90871 -47731
rect 90905 -47765 90963 -47731
rect 90997 -47765 91055 -47731
rect 91089 -47765 91147 -47731
rect 91181 -47765 91239 -47731
rect 91273 -47765 91331 -47731
rect 91365 -47765 91444 -47731
rect 82794 -47798 91444 -47765
rect 80430 -48020 80660 -47820
rect 86794 -47928 86884 -47918
rect 85314 -47948 85404 -47938
rect 81940 -48020 82950 -48010
rect 80430 -48100 80460 -48020
rect 80050 -48130 80460 -48100
rect 81940 -48140 81950 -48020
rect 82070 -48040 82950 -48020
rect 82070 -48130 82870 -48040
rect 82930 -48130 82950 -48040
rect 82070 -48140 82950 -48130
rect 72600 -48190 73050 -48180
rect 77400 -48150 77490 -48140
rect 81940 -48150 82950 -48140
rect 83030 -48020 83110 -48010
rect 83030 -48140 83040 -48020
rect 83100 -48140 83110 -48020
rect 83030 -48150 83110 -48140
rect 85314 -48138 85324 -47948
rect 85394 -48138 85404 -47948
rect 85584 -48008 86494 -47998
rect 85584 -48088 85594 -48008
rect 86484 -48088 86494 -48008
rect 85584 -48098 86494 -48088
rect 85314 -48148 85404 -48138
rect 86794 -48138 86804 -47928
rect 86874 -48138 86884 -47928
rect 88264 -47938 88354 -47928
rect 87034 -48008 87934 -47998
rect 87034 -48088 87044 -48008
rect 87924 -48088 87934 -48008
rect 87034 -48098 87934 -48088
rect 86794 -48148 86884 -48138
rect 88264 -48138 88274 -47938
rect 88344 -48138 88354 -47938
rect 89734 -47938 89824 -47928
rect 88504 -48018 89404 -48008
rect 88504 -48088 88514 -48018
rect 89394 -48088 89404 -48018
rect 88504 -48098 89404 -48088
rect 88264 -48148 88354 -48138
rect 89734 -48148 89744 -47938
rect 89814 -48148 89824 -47938
rect 91204 -47938 91294 -47928
rect 89974 -48017 90774 -48008
rect 89974 -48035 89986 -48017
rect 89974 -48037 89984 -48035
rect 89974 -48071 89982 -48037
rect 89974 -48089 89986 -48071
rect 90766 -48089 90774 -48017
rect 89974 -48098 90774 -48089
rect 77400 -48220 77410 -48150
rect 77480 -48220 77490 -48150
rect 89734 -48158 89824 -48148
rect 91204 -48148 91214 -47938
rect 91284 -48148 91294 -47938
rect 91204 -48158 91294 -48148
rect 79380 -48190 79710 -48160
rect 79380 -48220 79410 -48190
rect 77400 -48230 77490 -48220
rect 77570 -48255 79410 -48220
rect 77570 -48289 77607 -48255
rect 77641 -48289 77699 -48255
rect 77733 -48289 77791 -48255
rect 77825 -48289 77883 -48255
rect 77917 -48289 77975 -48255
rect 78009 -48289 78067 -48255
rect 78101 -48260 79410 -48255
rect 78101 -48289 78250 -48260
rect 77570 -48331 78250 -48289
rect 77570 -48365 77607 -48331
rect 77641 -48365 77699 -48331
rect 77733 -48365 77791 -48331
rect 77825 -48365 77883 -48331
rect 77917 -48365 77975 -48331
rect 78009 -48365 78250 -48331
rect 77570 -48370 78250 -48365
rect 78360 -48370 78560 -48260
rect 78670 -48370 78800 -48260
rect 78910 -48370 79060 -48260
rect 79170 -48370 79410 -48260
rect 77570 -48400 79410 -48370
rect 79380 -48430 79410 -48400
rect 79680 -48430 79710 -48190
rect 92000 -48210 95800 -47200
rect 79380 -48450 79710 -48430
rect 82794 -48275 91444 -48238
rect 82794 -48309 82867 -48275
rect 82901 -48309 82959 -48275
rect 82993 -48309 83051 -48275
rect 83085 -48309 83143 -48275
rect 83177 -48309 83235 -48275
rect 83269 -48309 83327 -48275
rect 83361 -48309 83419 -48275
rect 83453 -48309 83511 -48275
rect 83545 -48309 83603 -48275
rect 83637 -48309 83695 -48275
rect 83729 -48309 83787 -48275
rect 83821 -48309 83879 -48275
rect 83913 -48309 83971 -48275
rect 84005 -48309 84063 -48275
rect 84097 -48309 84155 -48275
rect 84189 -48309 84247 -48275
rect 84281 -48309 84339 -48275
rect 84373 -48309 84431 -48275
rect 84465 -48309 84523 -48275
rect 84557 -48309 84615 -48275
rect 84649 -48309 84707 -48275
rect 84741 -48309 84799 -48275
rect 84833 -48309 84891 -48275
rect 84925 -48309 84983 -48275
rect 85017 -48309 85075 -48275
rect 85109 -48309 85167 -48275
rect 85201 -48309 85259 -48275
rect 85293 -48309 85351 -48275
rect 85385 -48309 85443 -48275
rect 85477 -48309 85535 -48275
rect 85569 -48309 85627 -48275
rect 85661 -48309 85719 -48275
rect 85753 -48309 85811 -48275
rect 85845 -48309 85903 -48275
rect 85937 -48309 85995 -48275
rect 86029 -48309 86087 -48275
rect 86121 -48309 86179 -48275
rect 86213 -48309 86271 -48275
rect 86305 -48309 86363 -48275
rect 86397 -48309 86455 -48275
rect 86489 -48309 86547 -48275
rect 86581 -48309 86639 -48275
rect 86673 -48309 86731 -48275
rect 86765 -48309 86823 -48275
rect 86857 -48309 86915 -48275
rect 86949 -48309 87007 -48275
rect 87041 -48309 87099 -48275
rect 87133 -48309 87191 -48275
rect 87225 -48309 87283 -48275
rect 87317 -48309 87375 -48275
rect 87409 -48309 87467 -48275
rect 87501 -48309 87559 -48275
rect 87593 -48309 87651 -48275
rect 87685 -48309 87743 -48275
rect 87777 -48309 87835 -48275
rect 87869 -48309 87927 -48275
rect 87961 -48309 88019 -48275
rect 88053 -48309 88111 -48275
rect 88145 -48309 88203 -48275
rect 88237 -48309 88295 -48275
rect 88329 -48309 88387 -48275
rect 88421 -48309 88479 -48275
rect 88513 -48309 88571 -48275
rect 88605 -48309 88663 -48275
rect 88697 -48309 88755 -48275
rect 88789 -48309 88847 -48275
rect 88881 -48309 88939 -48275
rect 88973 -48309 89031 -48275
rect 89065 -48309 89123 -48275
rect 89157 -48309 89215 -48275
rect 89249 -48309 89307 -48275
rect 89341 -48309 89399 -48275
rect 89433 -48309 89491 -48275
rect 89525 -48309 89583 -48275
rect 89617 -48309 89675 -48275
rect 89709 -48309 89767 -48275
rect 89801 -48309 89859 -48275
rect 89893 -48309 89951 -48275
rect 89985 -48309 90043 -48275
rect 90077 -48309 90135 -48275
rect 90169 -48309 90227 -48275
rect 90261 -48309 90319 -48275
rect 90353 -48309 90411 -48275
rect 90445 -48309 90503 -48275
rect 90537 -48309 90595 -48275
rect 90629 -48309 90687 -48275
rect 90721 -48309 90779 -48275
rect 90813 -48309 90871 -48275
rect 90905 -48309 90963 -48275
rect 90997 -48309 91055 -48275
rect 91089 -48309 91147 -48275
rect 91181 -48309 91239 -48275
rect 91273 -48309 91331 -48275
rect 91365 -48309 91444 -48275
rect 82794 -48348 91444 -48309
rect 72600 -48460 73050 -48450
rect 55400 -48900 55500 -48500
rect 56100 -48900 56200 -48500
rect 72600 -48640 72820 -48460
rect 73040 -48640 73050 -48460
rect 82794 -48518 83484 -48348
rect 83654 -48358 86534 -48348
rect 83654 -48518 85124 -48358
rect 82794 -48528 85124 -48518
rect 85294 -48518 86534 -48358
rect 86704 -48518 87914 -48348
rect 88084 -48358 91444 -48348
rect 88084 -48518 89454 -48358
rect 85294 -48528 89454 -48518
rect 89624 -48528 90734 -48358
rect 90904 -48528 91444 -48358
rect 77980 -48570 78420 -48550
rect 72600 -48650 73050 -48640
rect 77440 -48580 77530 -48570
rect 77440 -48650 77450 -48580
rect 77520 -48650 77530 -48580
rect 77980 -48610 78000 -48570
rect 78040 -48610 78420 -48570
rect 77440 -48660 77530 -48650
rect 77770 -48670 77780 -48610
rect 77840 -48670 77850 -48610
rect 77770 -48680 77850 -48670
rect 77980 -48660 78420 -48610
rect 77980 -48700 78000 -48660
rect 78040 -48690 78420 -48660
rect 78040 -48700 78310 -48690
rect 77380 -48740 77540 -48720
rect 55400 -49000 56200 -48900
rect 72600 -48820 73050 -48810
rect 72600 -49000 72820 -48820
rect 73040 -49000 73050 -48820
rect 77380 -48840 77400 -48740
rect 72600 -49010 73050 -49000
rect 76900 -48860 77400 -48840
rect 77520 -48840 77540 -48740
rect 77980 -48740 78310 -48700
rect 77980 -48780 78000 -48740
rect 78040 -48780 78310 -48740
rect 77980 -48800 78310 -48780
rect 78410 -48800 78420 -48690
rect 77980 -48810 78420 -48800
rect 82794 -48578 91444 -48528
rect 77520 -48860 78590 -48840
rect 76900 -49000 76920 -48860
rect 77060 -48875 78590 -48860
rect 77060 -48909 77607 -48875
rect 77641 -48909 77699 -48875
rect 77733 -48909 77791 -48875
rect 77825 -48909 77883 -48875
rect 77917 -48909 77975 -48875
rect 78009 -48909 78590 -48875
rect 77060 -48951 78590 -48909
rect 77060 -48985 77607 -48951
rect 77641 -48985 77699 -48951
rect 77733 -48985 77791 -48951
rect 77825 -48985 77883 -48951
rect 77917 -48985 77975 -48951
rect 78009 -48985 78067 -48951
rect 78101 -48985 78159 -48951
rect 78193 -48985 78251 -48951
rect 78285 -48985 78343 -48951
rect 78377 -48985 78435 -48951
rect 78469 -48985 78527 -48951
rect 78561 -48985 78590 -48951
rect 77060 -48990 78590 -48985
rect 77060 -49000 77400 -48990
rect 76900 -49020 77400 -49000
rect 35690 -49131 42600 -49100
rect 77380 -49110 77400 -49020
rect 77520 -49020 78590 -48990
rect 80050 -48950 80460 -48920
rect 77520 -49110 77540 -49020
rect 77380 -49130 77540 -49110
rect 78550 -49070 78790 -49060
rect 78050 -49130 78130 -49120
rect 25860 -49152 42600 -49131
rect 35900 -49200 42600 -49152
rect 77770 -49180 77850 -49170
rect 77440 -49200 77540 -49190
rect 72600 -49220 73050 -49210
rect 72600 -49400 72820 -49220
rect 73040 -49400 73050 -49220
rect 77440 -49280 77450 -49200
rect 77530 -49280 77540 -49200
rect 77770 -49240 77780 -49180
rect 77840 -49240 77850 -49180
rect 78050 -49220 78060 -49130
rect 78120 -49220 78130 -49130
rect 78550 -49140 78570 -49070
rect 78640 -49140 78670 -49070
rect 78350 -49170 78410 -49160
rect 78050 -49230 78130 -49220
rect 78170 -49180 78300 -49170
rect 77770 -49250 77850 -49240
rect 77440 -49290 77540 -49280
rect 78170 -49280 78180 -49180
rect 78290 -49280 78300 -49180
rect 78350 -49240 78410 -49230
rect 78550 -49210 78670 -49140
rect 78170 -49290 78300 -49280
rect 78550 -49280 78570 -49210
rect 78640 -49280 78670 -49210
rect 55380 -49480 55800 -49400
rect 72600 -49410 73050 -49400
rect 78550 -49350 78670 -49280
rect 78550 -49420 78570 -49350
rect 78640 -49420 78670 -49350
rect 78780 -49420 78790 -49070
rect 80050 -49330 80080 -48950
rect 80430 -49040 80460 -48950
rect 80430 -49240 80660 -49040
rect 82794 -49148 82824 -48578
rect 91414 -49148 91444 -48578
rect 91750 -48240 95800 -48210
rect 91750 -48620 91780 -48240
rect 92130 -48620 95800 -48240
rect 91750 -48650 95800 -48620
rect 82794 -49178 91444 -49148
rect 80430 -49330 80460 -49240
rect 80050 -49360 80460 -49330
rect 78550 -49430 78790 -49420
rect 79380 -49420 79710 -49390
rect 92000 -49400 95800 -48650
rect 79380 -49460 79410 -49420
rect 35900 -49654 41700 -49600
rect 25862 -49669 41700 -49654
rect 25862 -50066 25882 -49669
rect 26996 -50066 27124 -49669
rect 28238 -50066 28366 -49669
rect 29480 -50066 29608 -49669
rect 30722 -50066 30850 -49669
rect 31964 -50066 32092 -49669
rect 33206 -50066 33334 -49669
rect 34448 -50066 34576 -49669
rect 35690 -49700 41700 -49669
rect 35690 -50066 36000 -49700
rect 25862 -50336 36000 -50066
rect 25862 -50733 25882 -50336
rect 26996 -50733 27124 -50336
rect 28238 -50733 28366 -50336
rect 29480 -50733 29608 -50336
rect 30722 -50733 30850 -50336
rect 31964 -50733 32092 -50336
rect 33206 -50733 33334 -50336
rect 34448 -50733 34576 -50336
rect 35690 -50700 36000 -50336
rect 41600 -50700 41700 -49700
rect 55380 -49760 55460 -49480
rect 55720 -49760 55800 -49480
rect 77570 -49495 79410 -49460
rect 77570 -49529 77607 -49495
rect 77641 -49529 77699 -49495
rect 77733 -49529 77791 -49495
rect 77825 -49529 77883 -49495
rect 77917 -49529 77975 -49495
rect 78009 -49529 78067 -49495
rect 78101 -49529 78159 -49495
rect 78193 -49529 78251 -49495
rect 78285 -49529 78343 -49495
rect 78377 -49529 78435 -49495
rect 78469 -49529 78527 -49495
rect 78561 -49500 79410 -49495
rect 78561 -49529 78630 -49500
rect 77570 -49571 78630 -49529
rect 77570 -49605 77607 -49571
rect 77641 -49605 77699 -49571
rect 77733 -49605 77791 -49571
rect 77825 -49605 77883 -49571
rect 77917 -49605 77975 -49571
rect 78009 -49605 78630 -49571
rect 77570 -49610 78630 -49605
rect 78740 -49610 78850 -49500
rect 78960 -49610 79090 -49500
rect 79200 -49610 79410 -49500
rect 77570 -49640 79410 -49610
rect 79380 -49660 79410 -49640
rect 79680 -49660 79710 -49420
rect 55380 -49840 55800 -49760
rect 72600 -49670 73050 -49660
rect 54090 -49938 54890 -49898
rect 54090 -50068 54150 -49938
rect 53510 -50120 53800 -50118
rect 53440 -50140 53800 -50120
rect 53440 -50340 53460 -50140
rect 53780 -50340 53800 -50140
rect 54080 -50198 54150 -50068
rect 54860 -50178 54890 -49938
rect 54850 -50198 54890 -50178
rect 54080 -50266 54880 -50198
rect 54079 -50272 54880 -50266
rect 54079 -50306 54091 -50272
rect 54867 -50298 54880 -50272
rect 54867 -50306 54879 -50298
rect 54079 -50312 54879 -50306
rect 53440 -50360 53800 -50340
rect 53510 -50458 53800 -50360
rect 53002 -50620 53480 -50558
rect 35690 -50733 41700 -50700
rect 25862 -50754 41700 -50733
rect 35900 -50800 41700 -50754
rect 53000 -50758 53480 -50620
rect 53510 -50568 53520 -50458
rect 53640 -50568 53800 -50458
rect 53510 -50688 53800 -50568
rect 53970 -50334 54040 -50318
rect 53970 -50372 53998 -50334
rect 54032 -50372 54040 -50334
rect 53970 -50568 54040 -50372
rect 54920 -50334 54990 -50318
rect 54920 -50372 54926 -50334
rect 54960 -50372 54990 -50334
rect 54079 -50400 54879 -50394
rect 54079 -50434 54091 -50400
rect 54867 -50434 54879 -50400
rect 54079 -50438 54879 -50434
rect 54079 -50440 54750 -50438
rect 54090 -50488 54750 -50440
rect 54740 -50518 54750 -50488
rect 54850 -50440 54879 -50438
rect 54850 -50508 54860 -50440
rect 54840 -50518 54860 -50508
rect 54750 -50528 54860 -50518
rect 54920 -50568 54990 -50372
rect 55430 -50418 55520 -50408
rect 55290 -50528 55390 -50518
rect 53970 -50598 55290 -50568
rect 55430 -50558 55520 -50488
rect 53970 -50608 55390 -50598
rect 54050 -50618 55380 -50608
rect 54050 -50628 54880 -50618
rect 54050 -50638 54091 -50628
rect 54079 -50662 54091 -50638
rect 54867 -50638 54880 -50628
rect 54867 -50662 54879 -50638
rect 54079 -50668 54879 -50662
rect 54920 -50678 54990 -50668
rect 53510 -50706 53630 -50688
rect 53510 -50738 53526 -50706
rect 53514 -50740 53526 -50738
rect 53614 -50738 53630 -50706
rect 53940 -50690 54038 -50678
rect 53940 -50698 53998 -50690
rect 53614 -50740 53626 -50738
rect 53514 -50746 53626 -50740
rect 35900 -51252 40800 -51200
rect 25860 -51271 40800 -51252
rect 25860 -51668 25882 -51271
rect 26996 -51668 27124 -51271
rect 28238 -51668 28366 -51271
rect 29480 -51668 29608 -51271
rect 30722 -51668 30850 -51271
rect 31964 -51668 32092 -51271
rect 33206 -51668 33334 -51271
rect 34448 -51668 34576 -51271
rect 35690 -51300 40800 -51271
rect 35690 -51668 36000 -51300
rect 25860 -51934 36000 -51668
rect 25860 -52331 25882 -51934
rect 26996 -52331 27124 -51934
rect 28238 -52331 28366 -51934
rect 29480 -52331 29608 -51934
rect 30722 -52331 30850 -51934
rect 31964 -52331 32092 -51934
rect 33206 -52331 33334 -51934
rect 34448 -52331 34576 -51934
rect 35690 -52300 36000 -51934
rect 40700 -52300 40800 -51300
rect 35690 -52331 40800 -52300
rect 25860 -52352 40800 -52331
rect 35900 -52400 40800 -52352
rect 53000 -52508 53050 -50758
rect 53250 -50768 53480 -50758
rect 53250 -52118 53330 -50768
rect 53400 -50778 53480 -50768
rect 53400 -50790 53504 -50778
rect 53400 -51566 53464 -50790
rect 53498 -51566 53504 -50790
rect 53400 -51578 53504 -51566
rect 53636 -50788 53682 -50778
rect 53636 -50790 53760 -50788
rect 53636 -51566 53642 -50790
rect 53676 -51566 53760 -50790
rect 53940 -50798 53950 -50698
rect 54032 -50728 54038 -50690
rect 54020 -50740 54038 -50728
rect 54020 -50798 54030 -50740
rect 54079 -50756 54879 -50750
rect 54079 -50790 54091 -50756
rect 54867 -50790 54879 -50756
rect 54920 -50778 54990 -50768
rect 55320 -50768 55380 -50618
rect 54079 -50796 54879 -50790
rect 53940 -50818 54030 -50798
rect 54090 -50828 54870 -50796
rect 55320 -50802 55334 -50768
rect 55368 -50802 55380 -50768
rect 55320 -50808 55380 -50802
rect 53840 -51128 53920 -51118
rect 53840 -51238 53860 -51128
rect 53840 -51248 53920 -51238
rect 53840 -51440 53900 -51248
rect 54320 -51328 54510 -50828
rect 55440 -50838 55520 -50558
rect 55410 -50840 55520 -50838
rect 55284 -50848 55330 -50840
rect 55230 -50852 55330 -50848
rect 55230 -50858 55290 -50852
rect 55324 -51028 55330 -50852
rect 55230 -51038 55330 -51028
rect 55284 -51040 55330 -51038
rect 55372 -50848 55520 -50840
rect 55372 -50852 55430 -50848
rect 55372 -51028 55378 -50852
rect 55412 -51018 55430 -50852
rect 55510 -51018 55520 -50848
rect 55412 -51028 55520 -51018
rect 55372 -51040 55418 -51028
rect 55580 -51128 55720 -49840
rect 72600 -49850 72820 -49670
rect 73040 -49850 73050 -49670
rect 79380 -49690 79710 -49660
rect 77960 -49770 78600 -49760
rect 77960 -49780 78170 -49770
rect 72600 -49860 73050 -49850
rect 77480 -49810 77590 -49800
rect 77480 -49900 77490 -49810
rect 77580 -49900 77590 -49810
rect 77960 -49820 77980 -49780
rect 78020 -49820 78170 -49780
rect 77480 -49910 77590 -49900
rect 77770 -49910 77780 -49850
rect 77840 -49910 77850 -49850
rect 77770 -49920 77850 -49910
rect 77960 -49900 78170 -49820
rect 77960 -49940 77980 -49900
rect 78020 -49940 78170 -49900
rect 58776 -50070 59306 -49950
rect 77400 -50000 77560 -49980
rect 58776 -50080 58966 -50070
rect 56146 -50180 57366 -50130
rect 55954 -50328 56046 -50316
rect 56146 -50328 56506 -50180
rect 55954 -50498 55960 -50328
rect 56040 -50498 56046 -50328
rect 55954 -50510 56046 -50498
rect 56120 -50358 56506 -50328
rect 56120 -50568 56190 -50358
rect 56390 -50430 56506 -50358
rect 57016 -50334 57366 -50180
rect 57586 -50230 58966 -50080
rect 59126 -50230 59306 -50070
rect 57586 -50250 59306 -50230
rect 59946 -50100 60386 -50000
rect 57586 -50280 58986 -50250
rect 59946 -50260 59956 -50100
rect 60166 -50260 60386 -50100
rect 72610 -50040 73050 -50030
rect 72610 -50220 72820 -50040
rect 73040 -50220 73050 -50040
rect 77400 -50080 77420 -50000
rect 72610 -50230 73050 -50220
rect 76900 -50100 77420 -50080
rect 57016 -50430 57368 -50334
rect 56390 -50470 57368 -50430
rect 56390 -50568 57126 -50470
rect 56120 -50574 57126 -50568
rect 56120 -50578 56750 -50574
rect 55880 -50618 55970 -50608
rect 55870 -50696 55880 -50650
rect 55970 -50696 55982 -50650
rect 55880 -50708 55970 -50698
rect 55000 -51138 55090 -51128
rect 55000 -51248 55090 -51238
rect 54710 -51328 54960 -51308
rect 53940 -51368 54960 -51328
rect 53940 -51372 54730 -51368
rect 53930 -51378 54730 -51372
rect 53930 -51412 53942 -51378
rect 54718 -51412 54730 -51378
rect 53930 -51418 54730 -51412
rect 53840 -51528 53858 -51440
rect 53892 -51528 53900 -51440
rect 53840 -51548 53900 -51528
rect 54762 -51438 54850 -51428
rect 54762 -51440 54770 -51438
rect 54762 -51528 54768 -51440
rect 54840 -51528 54850 -51438
rect 54762 -51540 54850 -51528
rect 54770 -51548 54850 -51540
rect 53636 -51578 53760 -51566
rect 53400 -51796 53480 -51578
rect 53514 -51616 53626 -51610
rect 53514 -51618 53526 -51616
rect 53510 -51650 53526 -51618
rect 53614 -51618 53626 -51616
rect 53614 -51650 53630 -51618
rect 53510 -51724 53630 -51650
rect 53510 -51758 53526 -51724
rect 53614 -51758 53630 -51724
rect 53680 -51638 53760 -51578
rect 53930 -51556 54730 -51550
rect 53930 -51590 53942 -51556
rect 54718 -51590 54730 -51556
rect 53930 -51596 54730 -51590
rect 53940 -51628 54720 -51596
rect 53920 -51638 54720 -51628
rect 53680 -51728 54720 -51638
rect 53514 -51764 53626 -51758
rect 53680 -51796 53760 -51728
rect 53920 -51738 54720 -51728
rect 53940 -51778 54720 -51738
rect 54900 -51768 54960 -51368
rect 55010 -51360 55090 -51248
rect 55540 -51138 55720 -51128
rect 55630 -51238 55720 -51138
rect 55130 -51274 55506 -51268
rect 55130 -51308 55142 -51274
rect 55494 -51308 55506 -51274
rect 55130 -51314 55506 -51308
rect 55010 -51394 55046 -51360
rect 55080 -51394 55090 -51360
rect 55010 -51408 55090 -51394
rect 55142 -51440 55494 -51314
rect 55540 -51360 55720 -51238
rect 55540 -51394 55556 -51360
rect 55590 -51394 55720 -51360
rect 55540 -51408 55720 -51394
rect 55780 -50740 55860 -50728
rect 55130 -51446 55506 -51440
rect 55130 -51480 55142 -51446
rect 55494 -51478 55506 -51446
rect 55494 -51480 55510 -51478
rect 55130 -51486 55510 -51480
rect 55140 -51498 55510 -51486
rect 55780 -51498 55820 -50740
rect 55140 -51516 55820 -51498
rect 55854 -51516 55860 -50740
rect 55140 -51528 55860 -51516
rect 55992 -50740 56038 -50728
rect 55992 -51516 55998 -50740
rect 56032 -50748 56038 -50740
rect 56120 -50748 56300 -50578
rect 57098 -50600 57126 -50574
rect 57356 -50600 57368 -50470
rect 57098 -50614 57368 -50600
rect 57096 -50645 57372 -50614
rect 57096 -50679 57125 -50645
rect 57159 -50679 57217 -50645
rect 57251 -50679 57309 -50645
rect 57343 -50679 57372 -50645
rect 57096 -50710 57372 -50679
rect 56032 -51106 56300 -50748
rect 56590 -50868 56660 -50858
rect 56660 -50934 57000 -50868
rect 57586 -50930 57706 -50280
rect 59946 -50290 60386 -50260
rect 76900 -50260 76920 -50100
rect 77060 -50260 77420 -50100
rect 76900 -50280 77420 -50260
rect 77400 -50290 77420 -50280
rect 77540 -50080 77560 -50000
rect 77960 -50000 78170 -49940
rect 77960 -50040 77980 -50000
rect 78020 -50040 78170 -50000
rect 78290 -50040 78530 -49770
rect 78590 -50040 78600 -49770
rect 77960 -50050 78600 -50040
rect 77540 -50115 78040 -50080
rect 77540 -50149 77607 -50115
rect 77641 -50149 77699 -50115
rect 77733 -50149 77791 -50115
rect 77825 -50149 77883 -50115
rect 77917 -50149 77975 -50115
rect 78009 -50149 78040 -50115
rect 77540 -50205 78040 -50149
rect 77540 -50239 77609 -50205
rect 77643 -50239 77701 -50205
rect 77735 -50239 77793 -50205
rect 77827 -50239 77885 -50205
rect 77919 -50239 77977 -50205
rect 78011 -50239 78040 -50205
rect 77540 -50280 78040 -50239
rect 77540 -50290 77560 -50280
rect 77400 -50310 77560 -50290
rect 77960 -50380 78310 -50370
rect 77960 -50420 77980 -50380
rect 78020 -50420 78060 -50380
rect 77460 -50450 77570 -50440
rect 57366 -50934 57706 -50930
rect 56660 -50938 57188 -50934
rect 56660 -50944 57190 -50938
rect 56660 -50994 57118 -50944
rect 57178 -50994 57190 -50944
rect 57314 -50940 57706 -50934
rect 57314 -50980 57326 -50940
rect 57366 -50980 57706 -50940
rect 57314 -50986 57706 -50980
rect 57366 -50990 57706 -50986
rect 58896 -50570 58986 -50550
rect 58896 -50630 58906 -50570
rect 58896 -50920 58926 -50630
rect 58966 -50920 58986 -50570
rect 59106 -50570 59516 -50560
rect 59106 -50630 59216 -50570
rect 59276 -50630 59326 -50570
rect 59386 -50630 59436 -50570
rect 59496 -50630 59516 -50570
rect 59106 -50647 59516 -50630
rect 59626 -50570 59706 -50530
rect 77460 -50540 77470 -50450
rect 77560 -50540 77570 -50450
rect 77770 -50480 77780 -50420
rect 77840 -50480 77850 -50420
rect 77770 -50490 77850 -50480
rect 77960 -50460 78060 -50420
rect 77460 -50550 77570 -50540
rect 77960 -50500 77980 -50460
rect 78020 -50500 78060 -50460
rect 59626 -50630 59636 -50570
rect 59626 -50640 59656 -50630
rect 59106 -50680 59125 -50647
rect 59113 -50681 59125 -50680
rect 59501 -50680 59516 -50647
rect 59501 -50681 59513 -50680
rect 59113 -50687 59513 -50681
rect 59546 -50690 59616 -50680
rect 59276 -50730 59356 -50720
rect 59276 -50749 59286 -50730
rect 59113 -50755 59286 -50749
rect 59346 -50749 59356 -50730
rect 59346 -50755 59513 -50749
rect 59113 -50789 59125 -50755
rect 59501 -50789 59513 -50755
rect 59606 -50750 59616 -50690
rect 59546 -50760 59616 -50750
rect 59113 -50790 59286 -50789
rect 59346 -50790 59513 -50789
rect 59016 -50800 59076 -50790
rect 59113 -50795 59513 -50790
rect 59276 -50800 59356 -50795
rect 59546 -50810 59616 -50800
rect 59016 -50870 59076 -50860
rect 59113 -50863 59513 -50857
rect 59113 -50897 59125 -50863
rect 59501 -50897 59513 -50863
rect 59606 -50870 59616 -50810
rect 59546 -50880 59616 -50870
rect 59113 -50900 59513 -50897
rect 59113 -50903 59516 -50900
rect 58896 -50930 58986 -50920
rect 58896 -50990 58906 -50930
rect 58966 -50990 58986 -50930
rect 58896 -50992 58986 -50990
rect 59116 -50920 59516 -50903
rect 59646 -50910 59656 -50640
rect 59116 -50980 59216 -50920
rect 59276 -50980 59336 -50920
rect 59396 -50980 59436 -50920
rect 59496 -50980 59516 -50920
rect 56660 -50998 57190 -50994
rect 56590 -51000 57190 -50998
rect 56590 -51004 57188 -51000
rect 56590 -51068 57000 -51004
rect 56032 -51118 56356 -51106
rect 56032 -51516 56280 -51118
rect 55992 -51528 56280 -51516
rect 55140 -51538 55200 -51528
rect 55450 -51558 55810 -51528
rect 55870 -51566 55982 -51560
rect 55870 -51600 55882 -51566
rect 55970 -51600 55982 -51566
rect 55870 -51606 55982 -51600
rect 55140 -51618 55200 -51608
rect 55024 -51648 55116 -51636
rect 55024 -51728 55030 -51648
rect 55110 -51728 55116 -51648
rect 55024 -51740 55116 -51728
rect 55734 -51648 55816 -51636
rect 55734 -51728 55740 -51648
rect 55810 -51728 55816 -51648
rect 55734 -51740 55816 -51728
rect 55880 -51638 55970 -51606
rect 55880 -51764 55970 -51728
rect 56060 -51748 56280 -51528
rect 56350 -51748 56356 -51118
rect 56480 -51188 56550 -51178
rect 56480 -51258 56550 -51248
rect 56590 -51287 56750 -51068
rect 58894 -51086 58988 -50992
rect 59116 -51000 59516 -50980
rect 59636 -50920 59656 -50910
rect 59696 -50920 59706 -50570
rect 77960 -50560 78060 -50500
rect 77960 -50600 77980 -50560
rect 78020 -50600 78060 -50560
rect 77960 -50640 78060 -50600
rect 77960 -50680 77980 -50640
rect 78020 -50680 78060 -50640
rect 78120 -50680 78310 -50380
rect 82790 -50530 91440 -50500
rect 77960 -50690 78310 -50680
rect 79380 -50680 79710 -50650
rect 77580 -50720 78040 -50718
rect 79380 -50720 79410 -50680
rect 59856 -50740 59976 -50730
rect 59856 -50830 59866 -50740
rect 59966 -50830 59976 -50740
rect 59856 -50840 59976 -50830
rect 60436 -50820 60446 -50720
rect 60526 -50820 60536 -50720
rect 60436 -50840 60536 -50820
rect 59636 -50930 59706 -50920
rect 59696 -50990 59706 -50930
rect 59636 -51010 59706 -50990
rect 59756 -50860 60536 -50840
rect 59756 -50900 59866 -50860
rect 60426 -50900 60536 -50860
rect 77570 -50749 79410 -50720
rect 77570 -50783 77609 -50749
rect 77643 -50783 77701 -50749
rect 77735 -50783 77793 -50749
rect 77827 -50783 77885 -50749
rect 77919 -50783 77977 -50749
rect 78011 -50750 79410 -50749
rect 78011 -50783 78940 -50750
rect 77570 -50821 78940 -50783
rect 77570 -50855 77607 -50821
rect 77641 -50855 77699 -50821
rect 77733 -50855 77791 -50821
rect 77825 -50855 77883 -50821
rect 77917 -50855 77975 -50821
rect 78009 -50855 78067 -50821
rect 78101 -50855 78159 -50821
rect 78193 -50855 78351 -50821
rect 78385 -50855 78443 -50821
rect 78477 -50855 78535 -50821
rect 78569 -50855 78627 -50821
rect 78661 -50855 78719 -50821
rect 78753 -50855 78811 -50821
rect 78845 -50855 78940 -50821
rect 77570 -50860 78940 -50855
rect 79050 -50860 79130 -50750
rect 79240 -50860 79410 -50750
rect 77570 -50870 79410 -50860
rect 77570 -50886 78222 -50870
rect 78320 -50880 79410 -50870
rect 78322 -50886 79410 -50880
rect 77570 -50890 78210 -50886
rect 78589 -50890 79410 -50886
rect 59756 -50910 60536 -50900
rect 59756 -50950 59826 -50910
rect 78238 -50920 78310 -50917
rect 59066 -51040 59176 -51030
rect 58896 -51150 58986 -51086
rect 59066 -51110 59076 -51040
rect 59166 -51110 59176 -51040
rect 59066 -51112 59103 -51110
rect 59137 -51112 59176 -51110
rect 59066 -51120 59176 -51112
rect 59756 -51140 59766 -50950
rect 59806 -51140 59826 -50950
rect 59956 -50968 60046 -50940
rect 59946 -50974 60046 -50968
rect 60126 -50968 60336 -50940
rect 60126 -50974 60346 -50968
rect 59856 -51010 59916 -51000
rect 59946 -51008 59958 -50974
rect 60334 -51008 60346 -50974
rect 59946 -51014 60346 -51008
rect 77460 -50970 77640 -50960
rect 60376 -51020 60446 -51010
rect 77460 -51040 77470 -50970
rect 77540 -50980 77640 -50970
rect 77540 -51030 77580 -50980
rect 77630 -51030 77640 -50980
rect 78230 -50980 78240 -50920
rect 78300 -50980 78310 -50920
rect 79380 -50920 79410 -50890
rect 79680 -50920 79710 -50680
rect 78830 -50960 79000 -50940
rect 79380 -50950 79710 -50920
rect 79980 -50950 80390 -50920
rect 78230 -50990 78300 -50980
rect 78830 -51010 78850 -50960
rect 77540 -51040 77640 -51030
rect 77460 -51050 77640 -51040
rect 78160 -51050 78230 -51030
rect 59856 -51090 59916 -51080
rect 59946 -51082 60346 -51076
rect 59946 -51116 59958 -51082
rect 60334 -51116 60346 -51082
rect 60376 -51090 60446 -51080
rect 77860 -51090 77920 -51080
rect 59946 -51122 59976 -51116
rect 57098 -51158 57368 -51154
rect 57096 -51164 57372 -51158
rect 57096 -51250 57098 -51164
rect 56424 -51288 56470 -51287
rect 56060 -51760 56356 -51748
rect 56410 -51299 56470 -51288
rect 53400 -51808 53504 -51796
rect 53400 -52118 53464 -51808
rect 53250 -52508 53464 -52118
rect 53000 -52584 53464 -52508
rect 53498 -52584 53504 -51808
rect 53000 -52588 53504 -52584
rect 53458 -52596 53504 -52588
rect 53636 -51808 53760 -51796
rect 53636 -52584 53642 -51808
rect 53676 -52584 53760 -51808
rect 53930 -51784 54730 -51778
rect 53930 -51818 53942 -51784
rect 54718 -51818 54730 -51784
rect 53930 -51824 54730 -51818
rect 53830 -51846 53900 -51828
rect 53830 -51934 53858 -51846
rect 53892 -51934 53900 -51846
rect 53830 -52128 53900 -51934
rect 54760 -51846 54850 -51828
rect 54760 -51934 54768 -51846
rect 54802 -51848 54850 -51846
rect 54900 -51838 55200 -51768
rect 55870 -51770 55982 -51764
rect 55870 -51804 55882 -51770
rect 55970 -51804 55982 -51770
rect 55450 -51838 55810 -51808
rect 55870 -51810 55982 -51804
rect 56060 -51838 56300 -51760
rect 54900 -51842 55820 -51838
rect 56000 -51842 56300 -51838
rect 54900 -51848 55860 -51842
rect 54840 -51928 54850 -51848
rect 54802 -51934 54850 -51928
rect 54760 -51948 54850 -51934
rect 55130 -51854 55860 -51848
rect 55130 -51878 55820 -51854
rect 55130 -51896 55510 -51878
rect 55130 -51930 55142 -51896
rect 55494 -51898 55510 -51896
rect 55494 -51930 55506 -51898
rect 55130 -51936 55506 -51930
rect 53930 -51962 54730 -51956
rect 53930 -51996 53942 -51962
rect 54718 -51996 54730 -51962
rect 55020 -51982 55090 -51968
rect 53930 -52002 54730 -51996
rect 53940 -52008 54730 -52002
rect 54920 -51998 54980 -51988
rect 53940 -52048 54920 -52008
rect 53830 -52138 53920 -52128
rect 53830 -52248 53850 -52138
rect 53830 -52258 53920 -52248
rect 54320 -52548 54510 -52048
rect 54710 -52068 54920 -52048
rect 54910 -52078 54980 -52068
rect 55020 -52016 55046 -51982
rect 55080 -52016 55090 -51982
rect 55020 -52128 55090 -52016
rect 55142 -52062 55494 -51936
rect 55540 -51982 55620 -51968
rect 55540 -52016 55556 -51982
rect 55590 -52016 55620 -51982
rect 55130 -52068 55506 -52062
rect 55130 -52102 55142 -52068
rect 55494 -52102 55506 -52068
rect 55130 -52108 55506 -52102
rect 55000 -52138 55090 -52128
rect 55000 -52248 55090 -52238
rect 55540 -52128 55620 -52016
rect 55540 -52138 55630 -52128
rect 55630 -52238 55680 -52148
rect 55540 -52248 55680 -52238
rect 55274 -52338 55320 -52336
rect 55220 -52348 55320 -52338
rect 55220 -52524 55280 -52518
rect 55314 -52524 55320 -52348
rect 55220 -52528 55320 -52524
rect 55274 -52536 55320 -52528
rect 55362 -52348 55408 -52336
rect 55362 -52524 55368 -52348
rect 55402 -52358 55510 -52348
rect 55402 -52524 55410 -52358
rect 55362 -52528 55410 -52524
rect 55500 -52528 55510 -52358
rect 55362 -52536 55510 -52528
rect 55390 -52538 55510 -52536
rect 53636 -52588 53760 -52584
rect 53636 -52596 53682 -52588
rect 53940 -52608 54020 -52568
rect 54080 -52582 54860 -52548
rect 55311 -52574 55371 -52568
rect 53514 -52634 53626 -52628
rect 53514 -52638 53526 -52634
rect 53510 -52668 53526 -52638
rect 53614 -52638 53626 -52634
rect 53614 -52668 53630 -52638
rect 53510 -52728 53630 -52668
rect 53940 -52688 53950 -52608
rect 54010 -52638 54020 -52608
rect 54069 -52588 54869 -52582
rect 54069 -52622 54081 -52588
rect 54857 -52622 54869 -52588
rect 54069 -52628 54869 -52622
rect 54910 -52598 54980 -52588
rect 54010 -52650 54028 -52638
rect 54022 -52688 54028 -52650
rect 53940 -52700 54028 -52688
rect 53940 -52708 54020 -52700
rect 54910 -52708 54980 -52698
rect 55311 -52608 55324 -52574
rect 55358 -52608 55371 -52574
rect 54070 -52710 54870 -52708
rect 35900 -52850 39900 -52800
rect 25860 -52869 39900 -52850
rect 54069 -52716 54870 -52710
rect 54069 -52738 54081 -52716
rect 54041 -52750 54081 -52738
rect 54857 -52718 54870 -52716
rect 54857 -52750 54880 -52718
rect 55311 -52748 55371 -52608
rect 54041 -52758 54880 -52750
rect 55240 -52758 55371 -52748
rect 54041 -52768 55240 -52758
rect 53510 -52858 53630 -52848
rect 53961 -52808 55240 -52768
rect 25860 -53266 25882 -52869
rect 26996 -53266 27124 -52869
rect 28238 -53266 28366 -52869
rect 29480 -53266 29608 -52869
rect 30722 -53266 30850 -52869
rect 31964 -53266 32092 -52869
rect 33206 -53266 33334 -52869
rect 34448 -53266 34576 -52869
rect 35690 -52900 39900 -52869
rect 35690 -53266 36000 -52900
rect 25860 -53536 36000 -53266
rect 25860 -53933 25884 -53536
rect 26998 -53933 27126 -53536
rect 28240 -53933 28368 -53536
rect 29482 -53933 29610 -53536
rect 30724 -53933 30852 -53536
rect 31966 -53933 32094 -53536
rect 33208 -53933 33336 -53536
rect 34450 -53933 34578 -53536
rect 35692 -53900 36000 -53536
rect 39800 -53900 39900 -52900
rect 53961 -53006 54031 -52808
rect 54730 -52868 54860 -52858
rect 54730 -52888 54740 -52868
rect 54080 -52938 54740 -52888
rect 54069 -52944 54740 -52938
rect 54850 -52938 54860 -52868
rect 54850 -52944 54869 -52938
rect 54069 -52978 54081 -52944
rect 54857 -52978 54869 -52944
rect 54069 -52984 54869 -52978
rect 54911 -52994 54981 -52808
rect 55370 -52808 55371 -52758
rect 55240 -52828 55370 -52818
rect 55410 -52848 55510 -52538
rect 55410 -52958 55510 -52938
rect 55570 -52868 55680 -52248
rect 55780 -52630 55820 -51878
rect 55854 -52630 55860 -51854
rect 55780 -52638 55860 -52630
rect 55814 -52642 55860 -52638
rect 55992 -51854 56300 -51842
rect 55992 -52630 55998 -51854
rect 56032 -52628 56300 -51854
rect 56410 -51898 56430 -51299
rect 56380 -52075 56430 -51898
rect 56464 -52075 56470 -51299
rect 56380 -52087 56470 -52075
rect 56552 -51299 56750 -51287
rect 56552 -52075 56558 -51299
rect 56592 -51438 56750 -51299
rect 57066 -51280 57098 -51250
rect 57368 -51250 57372 -51164
rect 58896 -51159 59076 -51150
rect 58896 -51160 59084 -51159
rect 59156 -51160 59202 -51159
rect 57368 -51280 57396 -51250
rect 57066 -51410 57086 -51280
rect 57376 -51410 57396 -51280
rect 56592 -52075 56610 -51438
rect 57066 -51440 57396 -51410
rect 56860 -51590 57060 -51578
rect 56860 -51618 57236 -51590
rect 56860 -51748 56900 -51618
rect 57020 -51748 57236 -51618
rect 56860 -51788 57236 -51748
rect 57036 -51790 57236 -51788
rect 58556 -51680 58756 -51660
rect 58556 -51840 58576 -51680
rect 58736 -51840 58756 -51680
rect 58556 -51860 58756 -51840
rect 56552 -52078 56610 -52075
rect 57036 -51940 57446 -51930
rect 56552 -52087 56598 -52078
rect 57036 -52080 57056 -51940
rect 57416 -52080 57446 -51940
rect 56380 -52358 56440 -52087
rect 57036 -52100 57098 -52080
rect 56480 -52128 56550 -52118
rect 56480 -52198 56550 -52188
rect 57096 -52214 57098 -52134
rect 57368 -52100 57446 -52080
rect 57368 -52214 57372 -52134
rect 57096 -52230 57372 -52214
rect 58896 -52290 58926 -51160
rect 58966 -51171 59086 -51160
rect 58966 -51547 59044 -51171
rect 59078 -51547 59086 -51171
rect 58966 -51570 59086 -51547
rect 59156 -51171 59256 -51160
rect 59756 -51170 59826 -51140
rect 59966 -51152 59976 -51122
rect 60316 -51122 60346 -51116
rect 61036 -51120 61466 -51110
rect 77190 -51120 77270 -51110
rect 60316 -51152 60326 -51122
rect 59966 -51160 60326 -51152
rect 59156 -51547 59162 -51171
rect 59196 -51240 59256 -51171
rect 59236 -51320 59256 -51240
rect 59196 -51440 59256 -51320
rect 59236 -51520 59256 -51440
rect 59196 -51547 59256 -51520
rect 59156 -51560 59256 -51547
rect 58966 -51880 59036 -51570
rect 59066 -51606 59176 -51600
rect 59066 -51610 59103 -51606
rect 59137 -51610 59176 -51606
rect 59066 -51680 59076 -51610
rect 59166 -51680 59176 -51610
rect 59066 -51690 59176 -51680
rect 59206 -51760 59256 -51560
rect 59376 -51190 59826 -51170
rect 59376 -51230 59476 -51190
rect 59656 -51230 59826 -51190
rect 59376 -51240 59826 -51230
rect 59376 -51290 59436 -51240
rect 59376 -51650 59386 -51290
rect 59426 -51650 59436 -51290
rect 59526 -51298 59576 -51270
rect 59526 -51332 59546 -51298
rect 59636 -51330 59706 -51270
rect 59580 -51332 59706 -51330
rect 59526 -51340 59706 -51332
rect 59476 -51382 59546 -51370
rect 59476 -51450 59502 -51382
rect 59476 -51558 59502 -51520
rect 59536 -51558 59546 -51382
rect 59476 -51570 59546 -51558
rect 59576 -51382 59636 -51370
rect 59576 -51390 59590 -51382
rect 59624 -51390 59636 -51382
rect 59576 -51570 59636 -51560
rect 59534 -51608 59592 -51602
rect 59534 -51610 59546 -51608
rect 59066 -51770 59176 -51760
rect 59066 -51840 59076 -51770
rect 59166 -51840 59176 -51770
rect 59066 -51842 59103 -51840
rect 59137 -51842 59176 -51840
rect 59066 -51850 59176 -51842
rect 59206 -51770 59266 -51760
rect 59206 -51850 59266 -51840
rect 59376 -51800 59436 -51650
rect 59516 -51642 59546 -51610
rect 59580 -51610 59592 -51608
rect 59666 -51610 59706 -51340
rect 59580 -51642 59706 -51610
rect 59516 -51680 59706 -51642
rect 59746 -51298 59936 -51270
rect 59746 -51332 59862 -51298
rect 59896 -51332 59936 -51298
rect 59746 -51340 59936 -51332
rect 61036 -51300 61206 -51120
rect 61346 -51300 61466 -51120
rect 75920 -51180 75940 -51120
rect 76050 -51180 77200 -51120
rect 77260 -51130 77830 -51120
rect 77260 -51170 77770 -51130
rect 77810 -51170 77830 -51130
rect 77260 -51180 77830 -51170
rect 77860 -51160 77920 -51150
rect 77190 -51190 77270 -51180
rect 77860 -51200 77870 -51160
rect 77910 -51200 77920 -51160
rect 61036 -51340 61466 -51300
rect 77390 -51250 77550 -51230
rect 77390 -51330 77410 -51250
rect 59746 -51600 59776 -51340
rect 60286 -51350 60476 -51340
rect 59806 -51382 59866 -51370
rect 59806 -51400 59818 -51382
rect 59852 -51400 59866 -51382
rect 59806 -51558 59818 -51540
rect 59852 -51558 59866 -51540
rect 59806 -51570 59866 -51558
rect 59900 -51380 60016 -51370
rect 59900 -51382 59916 -51380
rect 59900 -51558 59906 -51382
rect 59900 -51560 59916 -51558
rect 60006 -51560 60016 -51380
rect 60286 -51490 60306 -51350
rect 60456 -51490 60476 -51350
rect 76900 -51350 77410 -51330
rect 61176 -51400 61386 -51380
rect 60286 -51500 60476 -51490
rect 61026 -51420 61136 -51410
rect 59900 -51570 60016 -51560
rect 60076 -51557 60196 -51520
rect 60076 -51591 60127 -51557
rect 60161 -51591 60196 -51557
rect 59746 -51608 59926 -51600
rect 59746 -51610 59862 -51608
rect 59896 -51610 59926 -51608
rect 59746 -51680 59826 -51610
rect 59916 -51680 59926 -51610
rect 59746 -51690 59926 -51680
rect 60076 -51649 60196 -51591
rect 60336 -51560 60446 -51500
rect 60336 -51600 60366 -51560
rect 60406 -51600 60446 -51560
rect 60636 -51557 60816 -51520
rect 60636 -51591 60671 -51557
rect 60705 -51591 60747 -51557
rect 60781 -51591 60816 -51557
rect 60076 -51680 60127 -51649
rect 60161 -51680 60196 -51649
rect 59736 -51770 59936 -51760
rect 58966 -51901 59086 -51880
rect 58966 -52277 59044 -51901
rect 59078 -52277 59086 -51901
rect 58966 -52290 59086 -52277
rect 59156 -51890 59202 -51889
rect 59156 -51901 59236 -51890
rect 59156 -52277 59162 -51901
rect 59196 -51930 59236 -51901
rect 59226 -52010 59236 -51930
rect 59196 -52160 59236 -52010
rect 59226 -52240 59236 -52160
rect 59196 -52277 59236 -52240
rect 59376 -52170 59386 -51800
rect 59426 -52170 59436 -51800
rect 59516 -51811 59706 -51770
rect 59516 -51845 59545 -51811
rect 59579 -51845 59706 -51811
rect 59516 -51850 59706 -51845
rect 59533 -51851 59591 -51850
rect 59466 -51895 59546 -51880
rect 59586 -51883 59646 -51880
rect 59466 -51930 59501 -51895
rect 59466 -52071 59501 -52010
rect 59535 -52071 59546 -51895
rect 59466 -52080 59546 -52071
rect 59583 -51895 59646 -51883
rect 59583 -51910 59589 -51895
rect 59623 -51910 59646 -51895
rect 59583 -52050 59586 -51910
rect 59583 -52071 59589 -52050
rect 59623 -52071 59646 -52050
rect 59583 -52080 59646 -52071
rect 59495 -52083 59541 -52080
rect 59583 -52083 59629 -52080
rect 59533 -52120 59591 -52115
rect 59676 -52120 59706 -51850
rect 59376 -52210 59436 -52170
rect 59506 -52180 59516 -52120
rect 59596 -52180 59706 -52120
rect 59736 -51840 59826 -51770
rect 59926 -51840 59936 -51770
rect 59736 -51845 59861 -51840
rect 59895 -51845 59936 -51840
rect 59736 -51850 59936 -51845
rect 60076 -51840 60096 -51680
rect 60176 -51840 60196 -51680
rect 59736 -52120 59766 -51850
rect 59849 -51851 59907 -51850
rect 60076 -51867 60127 -51840
rect 60161 -51867 60196 -51840
rect 59796 -51883 59856 -51880
rect 59796 -51890 59857 -51883
rect 59856 -52070 59857 -51890
rect 59796 -52071 59817 -52070
rect 59851 -52071 59857 -52070
rect 59796 -52080 59857 -52071
rect 59811 -52083 59857 -52080
rect 59899 -51890 59945 -51883
rect 59899 -51895 59916 -51890
rect 59899 -52071 59905 -51895
rect 59899 -52080 59916 -52071
rect 60006 -52080 60016 -51890
rect 60076 -51925 60196 -51867
rect 60346 -51650 60426 -51600
rect 60346 -51690 60366 -51650
rect 60406 -51690 60426 -51650
rect 60346 -51740 60426 -51690
rect 60346 -51780 60366 -51740
rect 60406 -51780 60426 -51740
rect 60346 -51820 60426 -51780
rect 60346 -51860 60366 -51820
rect 60406 -51860 60426 -51820
rect 60346 -51870 60426 -51860
rect 60636 -51649 60816 -51591
rect 60636 -51683 60671 -51649
rect 60705 -51683 60747 -51649
rect 60781 -51683 60816 -51649
rect 60636 -51741 60816 -51683
rect 60636 -51775 60671 -51741
rect 60705 -51775 60747 -51741
rect 60781 -51775 60816 -51741
rect 60636 -51833 60816 -51775
rect 60636 -51867 60671 -51833
rect 60705 -51867 60747 -51833
rect 60781 -51867 60816 -51833
rect 60076 -51959 60127 -51925
rect 60161 -51959 60196 -51925
rect 60076 -51990 60196 -51959
rect 60276 -51910 60546 -51900
rect 60276 -51925 60476 -51910
rect 60276 -51959 60297 -51925
rect 60331 -51959 60369 -51925
rect 60405 -51959 60449 -51925
rect 60276 -51970 60476 -51959
rect 60536 -51970 60546 -51910
rect 60276 -51980 60546 -51970
rect 60636 -51925 60816 -51867
rect 61026 -51530 61036 -51420
rect 61126 -51530 61136 -51420
rect 61176 -51480 61196 -51400
rect 61366 -51480 61386 -51400
rect 61176 -51500 61386 -51480
rect 76900 -51490 76920 -51350
rect 77060 -51370 77410 -51350
rect 77530 -51330 77550 -51250
rect 77860 -51240 77920 -51200
rect 78160 -51220 78170 -51050
rect 78220 -51060 78230 -51050
rect 78220 -51080 78580 -51060
rect 78220 -51130 78470 -51080
rect 78560 -51130 78580 -51080
rect 78830 -51080 78860 -51010
rect 78220 -51140 78580 -51130
rect 78620 -51120 78710 -51110
rect 78220 -51220 78230 -51140
rect 78340 -51180 78410 -51170
rect 78620 -51180 78630 -51120
rect 78700 -51180 78710 -51120
rect 77860 -51280 77870 -51240
rect 77910 -51280 77920 -51240
rect 77860 -51300 77920 -51280
rect 77950 -51230 78030 -51220
rect 77950 -51290 77960 -51230
rect 78020 -51290 78030 -51230
rect 78160 -51240 78230 -51220
rect 78330 -51240 78340 -51180
rect 78410 -51240 78420 -51180
rect 78620 -51190 78710 -51180
rect 78830 -51130 78850 -51080
rect 78830 -51200 78860 -51130
rect 78830 -51250 78850 -51200
rect 78980 -51250 79000 -50960
rect 78830 -51270 79000 -51250
rect 77950 -51300 78030 -51290
rect 79980 -51330 80010 -50950
rect 80360 -51030 80390 -50950
rect 80360 -51230 80590 -51030
rect 82790 -51100 82820 -50530
rect 91410 -51100 91440 -50530
rect 82790 -51170 91440 -51100
rect 80360 -51330 80390 -51230
rect 77530 -51365 78880 -51330
rect 79980 -51360 80390 -51330
rect 82790 -51340 83450 -51170
rect 83620 -51340 85150 -51170
rect 85320 -51340 86530 -51170
rect 86700 -51340 87820 -51170
rect 87990 -51340 89340 -51170
rect 89510 -51340 90750 -51170
rect 90920 -51340 91440 -51170
rect 77530 -51370 77607 -51365
rect 77060 -51399 77607 -51370
rect 77641 -51399 77699 -51365
rect 77733 -51399 77791 -51365
rect 77825 -51399 77883 -51365
rect 77917 -51399 77975 -51365
rect 78009 -51399 78067 -51365
rect 78101 -51399 78159 -51365
rect 78193 -51399 78351 -51365
rect 78385 -51399 78443 -51365
rect 78477 -51399 78535 -51365
rect 78569 -51399 78627 -51365
rect 78661 -51399 78719 -51365
rect 78753 -51399 78811 -51365
rect 78845 -51399 78880 -51365
rect 77060 -51430 78880 -51399
rect 77060 -51490 77410 -51430
rect 61026 -51560 61136 -51530
rect 61026 -51600 61046 -51560
rect 61086 -51600 61136 -51560
rect 61026 -51650 61136 -51600
rect 61026 -51690 61046 -51650
rect 61086 -51690 61136 -51650
rect 61026 -51740 61136 -51690
rect 61026 -51780 61046 -51740
rect 61086 -51780 61136 -51740
rect 61026 -51820 61136 -51780
rect 61026 -51860 61046 -51820
rect 61086 -51860 61136 -51820
rect 61026 -51880 61136 -51860
rect 61256 -51557 61366 -51500
rect 76900 -51510 77410 -51490
rect 61256 -51591 61291 -51557
rect 61325 -51591 61366 -51557
rect 77390 -51550 77410 -51510
rect 77530 -51437 78880 -51430
rect 77530 -51471 77607 -51437
rect 77641 -51471 77699 -51437
rect 77733 -51471 77791 -51437
rect 77825 -51471 77883 -51437
rect 77917 -51471 77975 -51437
rect 78009 -51471 78067 -51437
rect 78101 -51471 78159 -51437
rect 78193 -51471 78880 -51437
rect 82790 -51381 91440 -51340
rect 82790 -51415 82867 -51381
rect 82901 -51415 82959 -51381
rect 82993 -51415 83051 -51381
rect 83085 -51415 83143 -51381
rect 83177 -51415 83235 -51381
rect 83269 -51415 83327 -51381
rect 83361 -51415 83419 -51381
rect 83453 -51415 83511 -51381
rect 83545 -51415 83603 -51381
rect 83637 -51415 83695 -51381
rect 83729 -51415 83787 -51381
rect 83821 -51415 83879 -51381
rect 83913 -51415 83971 -51381
rect 84005 -51415 84063 -51381
rect 84097 -51415 84155 -51381
rect 84189 -51415 84247 -51381
rect 84281 -51415 84339 -51381
rect 84373 -51415 84431 -51381
rect 84465 -51415 84523 -51381
rect 84557 -51415 84615 -51381
rect 84649 -51415 84707 -51381
rect 84741 -51415 84799 -51381
rect 84833 -51415 84891 -51381
rect 84925 -51415 84983 -51381
rect 85017 -51415 85075 -51381
rect 85109 -51415 85167 -51381
rect 85201 -51415 85259 -51381
rect 85293 -51415 85351 -51381
rect 85385 -51415 85443 -51381
rect 85477 -51415 85535 -51381
rect 85569 -51415 85627 -51381
rect 85661 -51415 85719 -51381
rect 85753 -51415 85811 -51381
rect 85845 -51415 85903 -51381
rect 85937 -51415 85995 -51381
rect 86029 -51415 86087 -51381
rect 86121 -51415 86179 -51381
rect 86213 -51415 86271 -51381
rect 86305 -51415 86363 -51381
rect 86397 -51415 86455 -51381
rect 86489 -51415 86547 -51381
rect 86581 -51415 86639 -51381
rect 86673 -51415 86731 -51381
rect 86765 -51415 86823 -51381
rect 86857 -51415 86915 -51381
rect 86949 -51415 87007 -51381
rect 87041 -51415 87099 -51381
rect 87133 -51415 87191 -51381
rect 87225 -51415 87283 -51381
rect 87317 -51415 87375 -51381
rect 87409 -51415 87467 -51381
rect 87501 -51415 87559 -51381
rect 87593 -51415 87651 -51381
rect 87685 -51415 87743 -51381
rect 87777 -51415 87835 -51381
rect 87869 -51415 87927 -51381
rect 87961 -51415 88019 -51381
rect 88053 -51415 88111 -51381
rect 88145 -51415 88203 -51381
rect 88237 -51415 88295 -51381
rect 88329 -51415 88387 -51381
rect 88421 -51415 88479 -51381
rect 88513 -51415 88571 -51381
rect 88605 -51415 88663 -51381
rect 88697 -51415 88755 -51381
rect 88789 -51415 88847 -51381
rect 88881 -51415 88939 -51381
rect 88973 -51415 89031 -51381
rect 89065 -51415 89123 -51381
rect 89157 -51415 89215 -51381
rect 89249 -51415 89307 -51381
rect 89341 -51415 89399 -51381
rect 89433 -51415 89491 -51381
rect 89525 -51415 89583 -51381
rect 89617 -51415 89675 -51381
rect 89709 -51415 89767 -51381
rect 89801 -51415 89859 -51381
rect 89893 -51415 89951 -51381
rect 89985 -51415 90043 -51381
rect 90077 -51415 90135 -51381
rect 90169 -51415 90227 -51381
rect 90261 -51415 90319 -51381
rect 90353 -51415 90411 -51381
rect 90445 -51415 90503 -51381
rect 90537 -51415 90595 -51381
rect 90629 -51415 90687 -51381
rect 90721 -51415 90779 -51381
rect 90813 -51415 90871 -51381
rect 90905 -51415 90963 -51381
rect 90997 -51415 91055 -51381
rect 91089 -51415 91147 -51381
rect 91181 -51415 91239 -51381
rect 91273 -51415 91331 -51381
rect 91365 -51415 91440 -51381
rect 82790 -51450 91440 -51415
rect 77530 -51510 78880 -51471
rect 77530 -51550 77550 -51510
rect 61256 -51649 61366 -51591
rect 77190 -51570 77270 -51560
rect 77390 -51570 77550 -51550
rect 77760 -51560 77820 -51540
rect 77190 -51630 77200 -51570
rect 77260 -51600 77270 -51570
rect 77760 -51600 77770 -51560
rect 77810 -51600 77820 -51560
rect 77260 -51630 77820 -51600
rect 77190 -51640 77820 -51630
rect 61256 -51650 61291 -51649
rect 61325 -51650 61366 -51649
rect 61256 -51860 61276 -51650
rect 61356 -51860 61366 -51650
rect 77760 -51650 77820 -51640
rect 77760 -51690 77770 -51650
rect 77810 -51690 77820 -51650
rect 77760 -51710 77820 -51690
rect 77850 -51710 77860 -51540
rect 77920 -51710 77930 -51540
rect 78170 -51550 78240 -51540
rect 78170 -51600 78200 -51550
rect 77850 -51720 77930 -51710
rect 77960 -51660 78030 -51650
rect 77960 -51720 77970 -51660
rect 77960 -51730 78030 -51720
rect 78170 -51690 78240 -51600
rect 78170 -51740 78200 -51690
rect 61256 -51867 61291 -51860
rect 61325 -51867 61366 -51860
rect 60636 -51959 60671 -51925
rect 60705 -51959 60747 -51925
rect 60781 -51959 60816 -51925
rect 60636 -52040 60816 -51959
rect 60966 -51924 61177 -51910
rect 60966 -51925 61129 -51924
rect 60966 -51959 60980 -51925
rect 61015 -51959 61053 -51925
rect 61088 -51958 61129 -51925
rect 61164 -51958 61177 -51924
rect 61088 -51959 61177 -51958
rect 60966 -51990 61177 -51959
rect 61256 -51925 61366 -51867
rect 77420 -51800 77510 -51790
rect 77420 -51870 77430 -51800
rect 77500 -51870 77510 -51800
rect 77420 -51880 77510 -51870
rect 78170 -51830 78240 -51740
rect 78170 -51880 78200 -51830
rect 78170 -51910 78240 -51880
rect 78300 -51910 78310 -51540
rect 86790 -51580 86880 -51570
rect 85310 -51600 85400 -51590
rect 82280 -51680 82950 -51670
rect 82280 -51790 82290 -51680
rect 82440 -51690 82950 -51680
rect 82440 -51780 82870 -51690
rect 82930 -51780 82950 -51690
rect 82440 -51790 82950 -51780
rect 82280 -51800 82950 -51790
rect 83020 -51680 83110 -51670
rect 83020 -51790 83030 -51680
rect 83100 -51790 83110 -51680
rect 83020 -51800 83110 -51790
rect 85310 -51790 85320 -51600
rect 85390 -51790 85400 -51600
rect 85580 -51660 86490 -51650
rect 85580 -51740 85590 -51660
rect 86480 -51740 86490 -51660
rect 85580 -51750 86490 -51740
rect 85310 -51800 85400 -51790
rect 86790 -51790 86800 -51580
rect 86870 -51790 86880 -51580
rect 88260 -51590 88350 -51580
rect 87030 -51660 87930 -51650
rect 87030 -51740 87040 -51660
rect 87920 -51740 87930 -51660
rect 87030 -51750 87930 -51740
rect 86790 -51800 86880 -51790
rect 88260 -51790 88270 -51590
rect 88340 -51790 88350 -51590
rect 89730 -51590 89820 -51580
rect 88500 -51670 89400 -51660
rect 88500 -51740 88510 -51670
rect 89390 -51740 89400 -51670
rect 88500 -51750 89400 -51740
rect 88260 -51800 88350 -51790
rect 89730 -51800 89740 -51590
rect 89810 -51800 89820 -51590
rect 91200 -51590 91290 -51580
rect 89970 -51669 90770 -51660
rect 89970 -51687 89982 -51669
rect 89970 -51689 89980 -51687
rect 89970 -51723 89978 -51689
rect 89970 -51741 89982 -51723
rect 90762 -51741 90770 -51669
rect 89970 -51750 90770 -51741
rect 89730 -51810 89820 -51800
rect 91200 -51800 91210 -51590
rect 91280 -51800 91290 -51590
rect 91200 -51810 91290 -51800
rect 92000 -51840 95800 -51000
rect 91750 -51870 95800 -51840
rect 78230 -51920 78310 -51910
rect 79380 -51900 79710 -51870
rect 61256 -51959 61291 -51925
rect 61325 -51959 61366 -51925
rect 79380 -51950 79410 -51900
rect 61256 -51990 61366 -51959
rect 77570 -51980 79410 -51950
rect 77570 -51981 78280 -51980
rect 60466 -52050 60546 -52040
rect 59899 -52083 59945 -52080
rect 60466 -52110 60476 -52050
rect 60536 -52110 60546 -52050
rect 59849 -52120 59907 -52115
rect 60466 -52120 60546 -52110
rect 60606 -52050 60826 -52040
rect 60606 -52110 60616 -52050
rect 60736 -52110 60756 -52050
rect 60816 -52110 60826 -52050
rect 60606 -52120 60826 -52110
rect 60886 -52050 60966 -52040
rect 60886 -52110 60896 -52050
rect 60956 -52110 60966 -52050
rect 60886 -52120 60966 -52110
rect 59736 -52121 59926 -52120
rect 59736 -52155 59861 -52121
rect 59895 -52155 59926 -52121
rect 59736 -52180 59926 -52155
rect 60636 -52170 60816 -52120
rect 59376 -52220 59826 -52210
rect 59376 -52260 59476 -52220
rect 59646 -52260 59826 -52220
rect 59376 -52270 59826 -52260
rect 59156 -52290 59236 -52277
rect 58896 -52300 59086 -52290
rect 56380 -52368 57000 -52358
rect 57356 -52364 57676 -52350
rect 56440 -52374 57000 -52368
rect 57314 -52370 57676 -52364
rect 56440 -52394 57178 -52374
rect 56440 -52444 57118 -52394
rect 57168 -52444 57178 -52394
rect 57314 -52410 57326 -52370
rect 57376 -52410 57676 -52370
rect 57314 -52416 57676 -52410
rect 57356 -52430 57676 -52416
rect 56440 -52454 57178 -52444
rect 56440 -52488 57000 -52454
rect 57112 -52456 57174 -52454
rect 56380 -52558 57000 -52488
rect 56032 -52630 56038 -52628
rect 55992 -52642 56038 -52630
rect 55880 -52674 55970 -52668
rect 55870 -52678 55982 -52674
rect 55870 -52720 55880 -52678
rect 55970 -52720 55982 -52678
rect 55880 -52768 55970 -52758
rect 56120 -52798 56300 -52628
rect 57096 -52709 57372 -52678
rect 57096 -52743 57125 -52709
rect 57159 -52743 57217 -52709
rect 57251 -52743 57309 -52709
rect 57343 -52720 57372 -52709
rect 57343 -52743 57376 -52720
rect 57096 -52780 57376 -52743
rect 57066 -52790 57376 -52780
rect 56426 -52798 57376 -52790
rect 56120 -52808 57376 -52798
rect 56014 -52858 56086 -52846
rect 55570 -52978 55830 -52868
rect 53961 -53044 53988 -53006
rect 54022 -53044 54031 -53006
rect 53961 -53058 54031 -53044
rect 54910 -53006 54981 -52994
rect 54910 -53044 54916 -53006
rect 54950 -53044 54981 -53006
rect 54910 -53056 54981 -53044
rect 54911 -53058 54981 -53056
rect 55220 -53018 55330 -53008
rect 54069 -53072 54869 -53066
rect 54069 -53106 54081 -53072
rect 54857 -53078 54869 -53072
rect 54857 -53106 54880 -53078
rect 54069 -53112 54880 -53106
rect 54090 -53188 54880 -53112
rect 55330 -53118 55380 -53018
rect 55330 -53128 55480 -53118
rect 55220 -53138 55480 -53128
rect 55280 -53152 55480 -53138
rect 55280 -53158 55488 -53152
rect 55280 -53178 55300 -53158
rect 54090 -53288 54150 -53188
rect 54840 -53288 54880 -53188
rect 55288 -53192 55300 -53178
rect 55476 -53192 55488 -53158
rect 55530 -53178 55610 -53168
rect 55288 -53198 55488 -53192
rect 55520 -53202 55530 -53190
rect 55520 -53236 55526 -53202
rect 55288 -53246 55488 -53240
rect 55288 -53280 55300 -53246
rect 55476 -53280 55488 -53246
rect 55520 -53248 55530 -53236
rect 55530 -53278 55610 -53268
rect 55288 -53286 55488 -53280
rect 54090 -53308 54140 -53288
rect 54100 -53548 54140 -53308
rect 54850 -53548 54880 -53288
rect 55300 -53328 55470 -53286
rect 55300 -53468 55320 -53328
rect 55470 -53414 55482 -53342
rect 55300 -53478 55470 -53468
rect 54100 -53588 54880 -53548
rect 55710 -53798 55830 -52978
rect 56014 -53008 56020 -52858
rect 56080 -53008 56086 -52858
rect 56014 -53020 56086 -53008
rect 56120 -53008 56170 -52808
rect 56390 -52860 57376 -52808
rect 56390 -52868 57156 -52860
rect 56390 -53008 56654 -52868
rect 56120 -53058 56654 -53008
rect 56306 -53086 56654 -53058
rect 56998 -53020 57156 -52868
rect 57316 -53020 57376 -52860
rect 56998 -53086 57376 -53020
rect 56306 -53500 57376 -53086
rect 57556 -53210 57676 -52430
rect 58896 -52460 58986 -52300
rect 59756 -52320 59826 -52270
rect 59066 -52336 59176 -52330
rect 59066 -52340 59103 -52336
rect 59137 -52340 59176 -52336
rect 59066 -52400 59076 -52340
rect 59166 -52400 59176 -52340
rect 59066 -52410 59176 -52400
rect 58896 -52830 58926 -52460
rect 58966 -52830 58986 -52530
rect 59116 -52460 59506 -52440
rect 59116 -52530 59146 -52460
rect 59226 -52530 59276 -52460
rect 59356 -52530 59396 -52460
rect 59476 -52530 59506 -52460
rect 59116 -52548 59506 -52530
rect 59646 -52460 59716 -52440
rect 59706 -52520 59716 -52460
rect 59646 -52530 59716 -52520
rect 59113 -52554 59513 -52548
rect 59113 -52588 59125 -52554
rect 59501 -52588 59513 -52554
rect 59113 -52594 59513 -52588
rect 59546 -52600 59616 -52590
rect 59246 -52656 59256 -52630
rect 59113 -52662 59256 -52656
rect 59366 -52656 59376 -52630
rect 59366 -52662 59513 -52656
rect 59016 -52700 59076 -52680
rect 59113 -52696 59125 -52662
rect 59501 -52696 59513 -52662
rect 59606 -52660 59616 -52600
rect 59546 -52670 59616 -52660
rect 59113 -52702 59513 -52696
rect 59016 -52790 59076 -52760
rect 59113 -52770 59513 -52764
rect 59113 -52804 59125 -52770
rect 59501 -52804 59513 -52770
rect 59113 -52810 59513 -52804
rect 58896 -52900 58906 -52830
rect 58896 -52920 58986 -52900
rect 59116 -52830 59516 -52810
rect 59116 -52900 59146 -52830
rect 59226 -52900 59276 -52830
rect 59356 -52900 59396 -52830
rect 59476 -52900 59516 -52830
rect 59116 -52920 59516 -52900
rect 59646 -52830 59656 -52530
rect 59706 -52830 59716 -52530
rect 59756 -52500 59766 -52320
rect 59806 -52500 59826 -52320
rect 59956 -52320 60336 -52310
rect 59956 -52334 59966 -52320
rect 59946 -52340 59966 -52334
rect 60326 -52334 60336 -52320
rect 60326 -52340 60346 -52334
rect 59856 -52380 59916 -52370
rect 59946 -52374 59958 -52340
rect 60334 -52374 60346 -52340
rect 61056 -52340 61176 -51990
rect 77570 -52015 77607 -51981
rect 77641 -52015 77699 -51981
rect 77733 -52015 77791 -51981
rect 77825 -52015 77883 -51981
rect 77917 -52015 77975 -51981
rect 78009 -52015 78067 -51981
rect 78101 -52015 78159 -51981
rect 78193 -52015 78280 -51981
rect 77570 -52053 78280 -52015
rect 77570 -52087 77607 -52053
rect 77641 -52087 77699 -52053
rect 77733 -52087 77791 -52053
rect 77825 -52087 77883 -52053
rect 77917 -52087 77975 -52053
rect 78009 -52087 78067 -52053
rect 78101 -52087 78159 -52053
rect 78193 -52087 78280 -52053
rect 77570 -52090 78280 -52087
rect 78390 -52090 78580 -51980
rect 78690 -52090 78880 -51980
rect 78990 -52090 79410 -51980
rect 77570 -52120 79410 -52090
rect 79380 -52140 79410 -52120
rect 79680 -52140 79710 -51900
rect 78160 -52170 78310 -52160
rect 79380 -52170 79710 -52140
rect 82790 -51925 91440 -51890
rect 82790 -51959 82867 -51925
rect 82901 -51959 82959 -51925
rect 82993 -51959 83051 -51925
rect 83085 -51959 83143 -51925
rect 83177 -51959 83235 -51925
rect 83269 -51959 83327 -51925
rect 83361 -51959 83419 -51925
rect 83453 -51959 83511 -51925
rect 83545 -51959 83603 -51925
rect 83637 -51959 83695 -51925
rect 83729 -51959 83787 -51925
rect 83821 -51959 83879 -51925
rect 83913 -51959 83971 -51925
rect 84005 -51959 84063 -51925
rect 84097 -51959 84155 -51925
rect 84189 -51959 84247 -51925
rect 84281 -51959 84339 -51925
rect 84373 -51959 84431 -51925
rect 84465 -51959 84523 -51925
rect 84557 -51959 84615 -51925
rect 84649 -51959 84707 -51925
rect 84741 -51959 84799 -51925
rect 84833 -51959 84891 -51925
rect 84925 -51959 84983 -51925
rect 85017 -51959 85075 -51925
rect 85109 -51959 85167 -51925
rect 85201 -51959 85259 -51925
rect 85293 -51959 85351 -51925
rect 85385 -51959 85443 -51925
rect 85477 -51959 85535 -51925
rect 85569 -51959 85627 -51925
rect 85661 -51959 85719 -51925
rect 85753 -51959 85811 -51925
rect 85845 -51959 85903 -51925
rect 85937 -51959 85995 -51925
rect 86029 -51959 86087 -51925
rect 86121 -51959 86179 -51925
rect 86213 -51959 86271 -51925
rect 86305 -51959 86363 -51925
rect 86397 -51959 86455 -51925
rect 86489 -51959 86547 -51925
rect 86581 -51959 86639 -51925
rect 86673 -51959 86731 -51925
rect 86765 -51959 86823 -51925
rect 86857 -51959 86915 -51925
rect 86949 -51959 87007 -51925
rect 87041 -51959 87099 -51925
rect 87133 -51959 87191 -51925
rect 87225 -51959 87283 -51925
rect 87317 -51959 87375 -51925
rect 87409 -51959 87467 -51925
rect 87501 -51959 87559 -51925
rect 87593 -51959 87651 -51925
rect 87685 -51959 87743 -51925
rect 87777 -51959 87835 -51925
rect 87869 -51959 87927 -51925
rect 87961 -51959 88019 -51925
rect 88053 -51959 88111 -51925
rect 88145 -51959 88203 -51925
rect 88237 -51959 88295 -51925
rect 88329 -51959 88387 -51925
rect 88421 -51959 88479 -51925
rect 88513 -51959 88571 -51925
rect 88605 -51959 88663 -51925
rect 88697 -51959 88755 -51925
rect 88789 -51959 88847 -51925
rect 88881 -51959 88939 -51925
rect 88973 -51959 89031 -51925
rect 89065 -51959 89123 -51925
rect 89157 -51959 89215 -51925
rect 89249 -51959 89307 -51925
rect 89341 -51959 89399 -51925
rect 89433 -51959 89491 -51925
rect 89525 -51959 89583 -51925
rect 89617 -51959 89675 -51925
rect 89709 -51959 89767 -51925
rect 89801 -51959 89859 -51925
rect 89893 -51959 89951 -51925
rect 89985 -51959 90043 -51925
rect 90077 -51959 90135 -51925
rect 90169 -51959 90227 -51925
rect 90261 -51959 90319 -51925
rect 90353 -51959 90411 -51925
rect 90445 -51959 90503 -51925
rect 90537 -51959 90595 -51925
rect 90629 -51959 90687 -51925
rect 90721 -51959 90779 -51925
rect 90813 -51959 90871 -51925
rect 90905 -51959 90963 -51925
rect 90997 -51959 91055 -51925
rect 91089 -51959 91147 -51925
rect 91181 -51959 91239 -51925
rect 91273 -51959 91331 -51925
rect 91365 -51959 91440 -51925
rect 82790 -52000 91440 -51959
rect 82790 -52170 83480 -52000
rect 83650 -52010 86530 -52000
rect 83650 -52170 85120 -52010
rect 75920 -52280 75940 -52190
rect 76050 -52210 77530 -52190
rect 76050 -52260 77470 -52210
rect 77510 -52260 77530 -52210
rect 76050 -52280 77530 -52260
rect 59946 -52380 59966 -52374
rect 60326 -52380 60346 -52374
rect 60376 -52380 60436 -52360
rect 59956 -52390 60336 -52380
rect 59856 -52460 59916 -52440
rect 59946 -52448 60346 -52442
rect 59756 -52540 59826 -52500
rect 59946 -52482 59958 -52448
rect 60334 -52482 60346 -52448
rect 60376 -52460 60436 -52440
rect 61126 -52440 61176 -52340
rect 75640 -52370 75660 -52310
rect 75760 -52340 77640 -52310
rect 75760 -52360 77920 -52340
rect 75760 -52370 77870 -52360
rect 77570 -52400 77870 -52370
rect 77910 -52400 77920 -52360
rect 61056 -52470 61176 -52440
rect 77380 -52420 77540 -52400
rect 77570 -52420 77920 -52400
rect 59946 -52488 60346 -52482
rect 59946 -52540 60336 -52488
rect 77380 -52540 77400 -52420
rect 77520 -52540 77540 -52420
rect 77860 -52450 77920 -52420
rect 77750 -52460 77830 -52450
rect 77750 -52520 77760 -52460
rect 77820 -52520 77830 -52460
rect 77750 -52530 77830 -52520
rect 77860 -52510 77870 -52450
rect 77910 -52510 77920 -52450
rect 77860 -52530 77920 -52510
rect 77960 -52390 78040 -52380
rect 77960 -52510 77970 -52390
rect 78030 -52510 78040 -52390
rect 77960 -52520 78040 -52510
rect 78160 -52510 78180 -52170
rect 78300 -52510 78310 -52170
rect 78160 -52520 78310 -52510
rect 82790 -52180 85120 -52170
rect 85290 -52170 86530 -52010
rect 86700 -52170 87910 -52000
rect 88080 -52010 91440 -52000
rect 88080 -52170 89450 -52010
rect 85290 -52180 89450 -52170
rect 89620 -52180 90730 -52010
rect 90900 -52180 91440 -52010
rect 82790 -52230 91440 -52180
rect 59756 -52560 60536 -52540
rect 59756 -52600 59866 -52560
rect 60426 -52600 60536 -52560
rect 59756 -52610 60536 -52600
rect 59796 -52720 59806 -52610
rect 59916 -52720 59926 -52610
rect 59796 -52730 59926 -52720
rect 60436 -52630 60536 -52610
rect 60436 -52750 60446 -52630
rect 60526 -52750 60536 -52630
rect 76900 -52560 77540 -52540
rect 76900 -52650 76920 -52560
rect 77060 -52597 78230 -52560
rect 77060 -52631 77607 -52597
rect 77641 -52631 77699 -52597
rect 77733 -52631 77791 -52597
rect 77825 -52631 77883 -52597
rect 77917 -52631 77975 -52597
rect 78009 -52631 78067 -52597
rect 78101 -52631 78159 -52597
rect 78193 -52631 78230 -52597
rect 77060 -52650 78230 -52631
rect 76900 -52670 78230 -52650
rect 60436 -52760 60536 -52750
rect 77380 -52790 77400 -52670
rect 77520 -52671 78230 -52670
rect 77520 -52705 77607 -52671
rect 77641 -52705 77699 -52671
rect 77733 -52705 77791 -52671
rect 77825 -52705 77883 -52671
rect 77917 -52705 77975 -52671
rect 78009 -52705 78067 -52671
rect 78101 -52705 78159 -52671
rect 78193 -52705 78230 -52671
rect 77520 -52740 78230 -52705
rect 77520 -52790 77540 -52740
rect 77380 -52810 77540 -52790
rect 77750 -52780 77830 -52770
rect 59646 -52840 59716 -52830
rect 59706 -52900 59716 -52840
rect 77750 -52840 77760 -52780
rect 77820 -52840 77830 -52780
rect 82790 -52800 82820 -52230
rect 91410 -52800 91440 -52230
rect 91750 -52250 91780 -51870
rect 92130 -52250 95800 -51870
rect 91750 -52280 95800 -52250
rect 82790 -52830 91440 -52800
rect 77750 -52850 77830 -52840
rect 77860 -52880 77920 -52870
rect 59646 -52920 59716 -52900
rect 75920 -52940 75940 -52880
rect 76050 -52890 77920 -52880
rect 76050 -52930 77870 -52890
rect 77910 -52930 77920 -52890
rect 76050 -52940 77920 -52930
rect 77860 -52950 77920 -52940
rect 77950 -52890 78030 -52880
rect 77950 -52960 77960 -52890
rect 78020 -52960 78030 -52890
rect 77950 -52970 78030 -52960
rect 77560 -52990 77640 -52970
rect 77560 -53010 77580 -52990
rect 75210 -53100 75230 -53010
rect 75330 -53080 77580 -53010
rect 77630 -53080 77640 -52990
rect 75330 -53100 77640 -53080
rect 78170 -52990 78760 -52980
rect 78170 -53120 78190 -52990
rect 78260 -53120 78640 -52990
rect 78170 -53130 78640 -53120
rect 78750 -53130 78760 -52990
rect 78170 -53140 78760 -53130
rect 79380 -53160 79710 -53130
rect 79380 -53180 79410 -53160
rect 58806 -53210 59356 -53180
rect 57556 -53220 59356 -53210
rect 57556 -53360 58986 -53220
rect 59126 -53360 59356 -53220
rect 59846 -53190 60256 -53180
rect 59846 -53300 59996 -53190
rect 60106 -53300 60256 -53190
rect 77570 -53215 79410 -53180
rect 77570 -53249 77607 -53215
rect 77641 -53249 77699 -53215
rect 77733 -53249 77791 -53215
rect 77825 -53249 77883 -53215
rect 77917 -53249 77975 -53215
rect 78009 -53249 78067 -53215
rect 78101 -53249 78159 -53215
rect 78193 -53220 79410 -53215
rect 78193 -53249 79120 -53220
rect 77570 -53291 79120 -53249
rect 57556 -53410 59356 -53360
rect 58806 -53490 59356 -53410
rect 55710 -53800 55910 -53798
rect 35692 -53933 39900 -53900
rect 25860 -53950 39900 -53933
rect 35900 -54000 39900 -53950
rect 55300 -53900 56200 -53800
rect 59600 -53900 60500 -53300
rect 77570 -53325 77607 -53291
rect 77641 -53325 77699 -53291
rect 77733 -53325 77791 -53291
rect 77825 -53325 77883 -53291
rect 77917 -53325 77975 -53291
rect 78009 -53325 78067 -53291
rect 78101 -53325 78159 -53291
rect 78193 -53325 78251 -53291
rect 78285 -53325 78343 -53291
rect 78377 -53325 78435 -53291
rect 78469 -53325 78527 -53291
rect 78561 -53325 78619 -53291
rect 78653 -53325 78711 -53291
rect 78745 -53325 78803 -53291
rect 78837 -53325 78895 -53291
rect 78929 -53325 78987 -53291
rect 79021 -53325 79120 -53291
rect 77570 -53330 79120 -53325
rect 79230 -53330 79410 -53220
rect 77570 -53356 79410 -53330
rect 77570 -53360 77720 -53356
rect 77880 -53360 79410 -53356
rect 77750 -53390 77850 -53385
rect 76480 -53460 76500 -53390
rect 76600 -53392 77850 -53390
rect 76600 -53432 77770 -53392
rect 77830 -53432 77850 -53392
rect 79380 -53400 79410 -53360
rect 79680 -53400 79710 -53160
rect 92000 -53200 95800 -52280
rect 76600 -53440 77850 -53432
rect 76600 -53460 77580 -53440
rect 77750 -53441 77850 -53440
rect 79000 -53410 79210 -53400
rect 78060 -53520 78150 -53510
rect 75210 -53610 75230 -53540
rect 75330 -53610 77880 -53540
rect 77800 -53630 77880 -53610
rect 77590 -53650 77720 -53640
rect 77380 -53660 77520 -53650
rect 76900 -53670 77520 -53660
rect 76900 -53680 77390 -53670
rect 76900 -53780 76920 -53680
rect 77060 -53780 77390 -53680
rect 76900 -53790 77390 -53780
rect 77510 -53790 77520 -53670
rect 77590 -53720 77600 -53650
rect 77710 -53720 77720 -53650
rect 77800 -53680 77820 -53630
rect 77860 -53680 77880 -53630
rect 78060 -53630 78070 -53520
rect 78140 -53630 78150 -53520
rect 78630 -53550 78750 -53540
rect 78060 -53640 78150 -53630
rect 78230 -53570 78310 -53560
rect 78230 -53630 78240 -53570
rect 78300 -53630 78310 -53570
rect 78230 -53640 78310 -53630
rect 78510 -53600 78590 -53580
rect 77800 -53690 77880 -53680
rect 78510 -53680 78530 -53600
rect 78570 -53680 78590 -53600
rect 78630 -53640 78640 -53550
rect 78740 -53640 78750 -53550
rect 78630 -53650 78750 -53640
rect 78800 -53590 78880 -53580
rect 78800 -53650 78810 -53590
rect 78870 -53650 78880 -53590
rect 78800 -53660 78880 -53650
rect 78510 -53710 78590 -53680
rect 77590 -53730 77720 -53720
rect 77970 -53720 78590 -53710
rect 77970 -53760 77990 -53720
rect 78030 -53760 78590 -53720
rect 79000 -53720 79020 -53410
rect 79070 -53420 79210 -53410
rect 79070 -53720 79080 -53420
rect 79190 -53720 79210 -53420
rect 79380 -53430 79710 -53400
rect 79000 -53740 79210 -53720
rect 79980 -53470 80390 -53440
rect 77970 -53770 78590 -53760
rect 76900 -53800 77520 -53790
rect 77380 -53835 79060 -53800
rect 77380 -53869 77607 -53835
rect 77641 -53869 77699 -53835
rect 77733 -53869 77791 -53835
rect 77825 -53869 77883 -53835
rect 77917 -53869 77975 -53835
rect 78009 -53869 78067 -53835
rect 78101 -53869 78159 -53835
rect 78193 -53869 78251 -53835
rect 78285 -53869 78343 -53835
rect 78377 -53869 78435 -53835
rect 78469 -53869 78527 -53835
rect 78561 -53869 78619 -53835
rect 78653 -53869 78711 -53835
rect 78745 -53869 78803 -53835
rect 78837 -53869 78895 -53835
rect 78929 -53869 78987 -53835
rect 79021 -53869 79060 -53835
rect 55300 -54300 55400 -53900
rect 56100 -54300 56200 -53900
rect 77380 -53920 79060 -53869
rect 79980 -53850 80010 -53470
rect 80360 -53570 80390 -53470
rect 80360 -53770 80590 -53570
rect 80360 -53850 80390 -53770
rect 79980 -53880 80390 -53850
rect 55300 -54400 56200 -54300
rect 35900 -54452 38900 -54400
rect 25862 -54471 38900 -54452
rect 25862 -54868 25884 -54471
rect 26998 -54868 27126 -54471
rect 28240 -54868 28368 -54471
rect 29482 -54868 29610 -54471
rect 30724 -54868 30852 -54471
rect 31966 -54868 32094 -54471
rect 33208 -54868 33336 -54471
rect 34450 -54868 34578 -54471
rect 35692 -54500 38900 -54471
rect 35692 -54868 36000 -54500
rect 25862 -55134 36000 -54868
rect 25862 -55531 25882 -55134
rect 26996 -55531 27124 -55134
rect 28238 -55531 28366 -55134
rect 29480 -55531 29608 -55134
rect 30722 -55531 30850 -55134
rect 31964 -55531 32092 -55134
rect 33206 -55531 33334 -55134
rect 34448 -55531 34576 -55134
rect 35690 -55500 36000 -55134
rect 38800 -55500 38900 -54500
rect 55380 -54880 55800 -54800
rect 55380 -55160 55460 -54880
rect 55720 -55160 55800 -54880
rect 55380 -55240 55800 -55160
rect 54090 -55338 54890 -55298
rect 54090 -55468 54150 -55338
rect 35690 -55531 38900 -55500
rect 53510 -55520 53800 -55518
rect 25862 -55552 38900 -55531
rect 35900 -55600 38900 -55552
rect 53460 -55540 53800 -55520
rect 53460 -55740 53480 -55540
rect 53780 -55740 53800 -55540
rect 54080 -55598 54150 -55468
rect 54860 -55578 54890 -55338
rect 54850 -55598 54890 -55578
rect 54080 -55666 54880 -55598
rect 54079 -55672 54880 -55666
rect 54079 -55706 54091 -55672
rect 54867 -55698 54880 -55672
rect 54867 -55706 54879 -55698
rect 54079 -55712 54879 -55706
rect 53460 -55760 53800 -55740
rect 53510 -55858 53800 -55760
rect 35900 -56050 37800 -56000
rect 53002 -56020 53480 -55958
rect 25860 -56069 37800 -56050
rect 25860 -56466 25882 -56069
rect 26996 -56466 27124 -56069
rect 28238 -56466 28366 -56069
rect 29480 -56466 29608 -56069
rect 30722 -56466 30850 -56069
rect 31964 -56466 32092 -56069
rect 33206 -56466 33334 -56069
rect 34448 -56466 34576 -56069
rect 35690 -56100 37800 -56069
rect 35690 -56466 36000 -56100
rect 25860 -56734 36000 -56466
rect 25860 -57131 25882 -56734
rect 26996 -57131 27124 -56734
rect 28238 -57131 28366 -56734
rect 29480 -57131 29608 -56734
rect 30722 -57131 30850 -56734
rect 31964 -57131 32092 -56734
rect 33206 -57131 33334 -56734
rect 34448 -57131 34576 -56734
rect 35690 -57100 36000 -56734
rect 37700 -57100 37800 -56100
rect 35690 -57131 37800 -57100
rect 25860 -57150 37800 -57131
rect 35900 -57200 37800 -57150
rect 53000 -56158 53480 -56020
rect 53510 -55968 53520 -55858
rect 53640 -55968 53800 -55858
rect 53510 -56088 53800 -55968
rect 53970 -55734 54040 -55718
rect 53970 -55772 53998 -55734
rect 54032 -55772 54040 -55734
rect 53970 -55968 54040 -55772
rect 54920 -55734 54990 -55718
rect 54920 -55772 54926 -55734
rect 54960 -55772 54990 -55734
rect 54079 -55800 54879 -55794
rect 54079 -55834 54091 -55800
rect 54867 -55834 54879 -55800
rect 54079 -55838 54879 -55834
rect 54079 -55840 54750 -55838
rect 54090 -55888 54750 -55840
rect 54740 -55918 54750 -55888
rect 54850 -55840 54879 -55838
rect 54850 -55908 54860 -55840
rect 54840 -55918 54860 -55908
rect 54750 -55928 54860 -55918
rect 54920 -55968 54990 -55772
rect 55430 -55818 55520 -55808
rect 55290 -55928 55390 -55918
rect 53970 -55998 55290 -55968
rect 55430 -55958 55520 -55888
rect 53970 -56008 55390 -55998
rect 54050 -56018 55380 -56008
rect 54050 -56028 54880 -56018
rect 54050 -56038 54091 -56028
rect 54079 -56062 54091 -56038
rect 54867 -56038 54880 -56028
rect 54867 -56062 54879 -56038
rect 54079 -56068 54879 -56062
rect 54920 -56078 54990 -56068
rect 53510 -56106 53630 -56088
rect 53510 -56138 53526 -56106
rect 53514 -56140 53526 -56138
rect 53614 -56138 53630 -56106
rect 53940 -56090 54038 -56078
rect 53940 -56098 53998 -56090
rect 53614 -56140 53626 -56138
rect 53514 -56146 53626 -56140
rect 25900 -57663 35740 -57580
rect 24380 -58020 25800 -57980
rect 25870 -57669 35740 -57663
rect 25870 -58066 25882 -57669
rect 26996 -58066 27124 -57669
rect 28238 -58066 28366 -57669
rect 29480 -58066 29608 -57669
rect 30722 -58066 30850 -57669
rect 31964 -58066 32092 -57669
rect 33206 -58066 33334 -57669
rect 34448 -58066 34576 -57669
rect 35690 -58066 35740 -57669
rect 53000 -57908 53050 -56158
rect 53250 -56168 53480 -56158
rect 53250 -57518 53330 -56168
rect 53400 -56178 53480 -56168
rect 53400 -56190 53504 -56178
rect 53400 -56966 53464 -56190
rect 53498 -56966 53504 -56190
rect 53400 -56978 53504 -56966
rect 53636 -56188 53682 -56178
rect 53636 -56190 53760 -56188
rect 53636 -56966 53642 -56190
rect 53676 -56966 53760 -56190
rect 53940 -56198 53950 -56098
rect 54032 -56128 54038 -56090
rect 54020 -56140 54038 -56128
rect 54020 -56198 54030 -56140
rect 54079 -56156 54879 -56150
rect 54079 -56190 54091 -56156
rect 54867 -56190 54879 -56156
rect 54920 -56178 54990 -56168
rect 55320 -56168 55380 -56018
rect 54079 -56196 54879 -56190
rect 53940 -56218 54030 -56198
rect 54090 -56228 54870 -56196
rect 55320 -56202 55334 -56168
rect 55368 -56202 55380 -56168
rect 55320 -56208 55380 -56202
rect 53840 -56528 53920 -56518
rect 53840 -56638 53860 -56528
rect 53840 -56648 53920 -56638
rect 53840 -56840 53900 -56648
rect 54320 -56728 54510 -56228
rect 55440 -56238 55520 -55958
rect 55410 -56240 55520 -56238
rect 55284 -56248 55330 -56240
rect 55230 -56252 55330 -56248
rect 55230 -56258 55290 -56252
rect 55324 -56428 55330 -56252
rect 55230 -56438 55330 -56428
rect 55284 -56440 55330 -56438
rect 55372 -56248 55520 -56240
rect 55372 -56252 55430 -56248
rect 55372 -56428 55378 -56252
rect 55412 -56418 55430 -56252
rect 55510 -56418 55520 -56248
rect 55412 -56428 55520 -56418
rect 55372 -56440 55418 -56428
rect 55580 -56528 55720 -55240
rect 58776 -55470 59306 -55350
rect 58776 -55480 58966 -55470
rect 56146 -55580 57366 -55530
rect 55954 -55728 56046 -55716
rect 56146 -55728 56506 -55580
rect 55954 -55898 55960 -55728
rect 56040 -55898 56046 -55728
rect 55954 -55910 56046 -55898
rect 56120 -55758 56506 -55728
rect 56120 -55968 56190 -55758
rect 56390 -55830 56506 -55758
rect 57016 -55734 57366 -55580
rect 57586 -55630 58966 -55480
rect 59126 -55630 59306 -55470
rect 57586 -55650 59306 -55630
rect 59946 -55500 60386 -55400
rect 57586 -55680 58986 -55650
rect 59946 -55660 59956 -55500
rect 60166 -55660 60386 -55500
rect 57016 -55830 57368 -55734
rect 56390 -55870 57368 -55830
rect 56390 -55968 57126 -55870
rect 56120 -55974 57126 -55968
rect 56120 -55978 56750 -55974
rect 55880 -56018 55970 -56008
rect 55870 -56096 55880 -56050
rect 55970 -56096 55982 -56050
rect 55880 -56108 55970 -56098
rect 55000 -56538 55090 -56528
rect 55000 -56648 55090 -56638
rect 54710 -56728 54960 -56708
rect 53940 -56768 54960 -56728
rect 53940 -56772 54730 -56768
rect 53930 -56778 54730 -56772
rect 53930 -56812 53942 -56778
rect 54718 -56812 54730 -56778
rect 53930 -56818 54730 -56812
rect 53840 -56928 53858 -56840
rect 53892 -56928 53900 -56840
rect 53840 -56948 53900 -56928
rect 54762 -56838 54850 -56828
rect 54762 -56840 54770 -56838
rect 54762 -56928 54768 -56840
rect 54840 -56928 54850 -56838
rect 54762 -56940 54850 -56928
rect 54770 -56948 54850 -56940
rect 53636 -56978 53760 -56966
rect 53400 -57196 53480 -56978
rect 53514 -57016 53626 -57010
rect 53514 -57018 53526 -57016
rect 53510 -57050 53526 -57018
rect 53614 -57018 53626 -57016
rect 53614 -57050 53630 -57018
rect 53510 -57124 53630 -57050
rect 53510 -57158 53526 -57124
rect 53614 -57158 53630 -57124
rect 53680 -57038 53760 -56978
rect 53930 -56956 54730 -56950
rect 53930 -56990 53942 -56956
rect 54718 -56990 54730 -56956
rect 53930 -56996 54730 -56990
rect 53940 -57028 54720 -56996
rect 53920 -57038 54720 -57028
rect 53680 -57128 54720 -57038
rect 53514 -57164 53626 -57158
rect 53680 -57196 53760 -57128
rect 53920 -57138 54720 -57128
rect 53940 -57178 54720 -57138
rect 54900 -57168 54960 -56768
rect 55010 -56760 55090 -56648
rect 55540 -56538 55720 -56528
rect 55630 -56638 55720 -56538
rect 55130 -56674 55506 -56668
rect 55130 -56708 55142 -56674
rect 55494 -56708 55506 -56674
rect 55130 -56714 55506 -56708
rect 55010 -56794 55046 -56760
rect 55080 -56794 55090 -56760
rect 55010 -56808 55090 -56794
rect 55142 -56840 55494 -56714
rect 55540 -56760 55720 -56638
rect 55540 -56794 55556 -56760
rect 55590 -56794 55720 -56760
rect 55540 -56808 55720 -56794
rect 55780 -56140 55860 -56128
rect 55130 -56846 55506 -56840
rect 55130 -56880 55142 -56846
rect 55494 -56878 55506 -56846
rect 55494 -56880 55510 -56878
rect 55130 -56886 55510 -56880
rect 55140 -56898 55510 -56886
rect 55780 -56898 55820 -56140
rect 55140 -56916 55820 -56898
rect 55854 -56916 55860 -56140
rect 55140 -56928 55860 -56916
rect 55992 -56140 56038 -56128
rect 55992 -56916 55998 -56140
rect 56032 -56148 56038 -56140
rect 56120 -56148 56300 -55978
rect 57098 -56000 57126 -55974
rect 57356 -56000 57368 -55870
rect 57098 -56014 57368 -56000
rect 57096 -56045 57372 -56014
rect 57096 -56079 57125 -56045
rect 57159 -56079 57217 -56045
rect 57251 -56079 57309 -56045
rect 57343 -56079 57372 -56045
rect 57096 -56110 57372 -56079
rect 56032 -56506 56300 -56148
rect 56590 -56268 56660 -56258
rect 56660 -56334 57000 -56268
rect 57586 -56330 57706 -55680
rect 59946 -55690 60386 -55660
rect 57366 -56334 57706 -56330
rect 56660 -56338 57188 -56334
rect 56660 -56344 57190 -56338
rect 56660 -56394 57118 -56344
rect 57178 -56394 57190 -56344
rect 57314 -56340 57706 -56334
rect 57314 -56380 57326 -56340
rect 57366 -56380 57706 -56340
rect 57314 -56386 57706 -56380
rect 57366 -56390 57706 -56386
rect 58896 -55970 58986 -55950
rect 58896 -56030 58906 -55970
rect 58896 -56320 58926 -56030
rect 58966 -56320 58986 -55970
rect 59106 -55970 59516 -55960
rect 59106 -56030 59216 -55970
rect 59276 -56030 59326 -55970
rect 59386 -56030 59436 -55970
rect 59496 -56030 59516 -55970
rect 59106 -56047 59516 -56030
rect 59626 -55970 59706 -55930
rect 59626 -56030 59636 -55970
rect 59626 -56040 59656 -56030
rect 59106 -56080 59125 -56047
rect 59113 -56081 59125 -56080
rect 59501 -56080 59516 -56047
rect 59501 -56081 59513 -56080
rect 59113 -56087 59513 -56081
rect 59546 -56090 59616 -56080
rect 59276 -56130 59356 -56120
rect 59276 -56149 59286 -56130
rect 59113 -56155 59286 -56149
rect 59346 -56149 59356 -56130
rect 59346 -56155 59513 -56149
rect 59113 -56189 59125 -56155
rect 59501 -56189 59513 -56155
rect 59606 -56150 59616 -56090
rect 59546 -56160 59616 -56150
rect 59113 -56190 59286 -56189
rect 59346 -56190 59513 -56189
rect 59016 -56200 59076 -56190
rect 59113 -56195 59513 -56190
rect 59276 -56200 59356 -56195
rect 59546 -56210 59616 -56200
rect 59016 -56270 59076 -56260
rect 59113 -56263 59513 -56257
rect 59113 -56297 59125 -56263
rect 59501 -56297 59513 -56263
rect 59606 -56270 59616 -56210
rect 59546 -56280 59616 -56270
rect 59113 -56300 59513 -56297
rect 59113 -56303 59516 -56300
rect 58896 -56330 58986 -56320
rect 58896 -56390 58906 -56330
rect 58966 -56390 58986 -56330
rect 58896 -56392 58986 -56390
rect 59116 -56320 59516 -56303
rect 59646 -56310 59656 -56040
rect 59116 -56380 59216 -56320
rect 59276 -56380 59336 -56320
rect 59396 -56380 59436 -56320
rect 59496 -56380 59516 -56320
rect 56660 -56398 57190 -56394
rect 56590 -56400 57190 -56398
rect 56590 -56404 57188 -56400
rect 56590 -56468 57000 -56404
rect 56032 -56518 56356 -56506
rect 56032 -56916 56280 -56518
rect 55992 -56928 56280 -56916
rect 55140 -56938 55200 -56928
rect 55450 -56958 55810 -56928
rect 55870 -56966 55982 -56960
rect 55870 -57000 55882 -56966
rect 55970 -57000 55982 -56966
rect 55870 -57006 55982 -57000
rect 55140 -57018 55200 -57008
rect 55024 -57048 55116 -57036
rect 55024 -57128 55030 -57048
rect 55110 -57128 55116 -57048
rect 55024 -57140 55116 -57128
rect 55734 -57048 55816 -57036
rect 55734 -57128 55740 -57048
rect 55810 -57128 55816 -57048
rect 55734 -57140 55816 -57128
rect 55880 -57038 55970 -57006
rect 55880 -57164 55970 -57128
rect 56060 -57148 56280 -56928
rect 56350 -57148 56356 -56518
rect 56480 -56588 56550 -56578
rect 56480 -56658 56550 -56648
rect 56590 -56687 56750 -56468
rect 58894 -56486 58988 -56392
rect 59116 -56400 59516 -56380
rect 59636 -56320 59656 -56310
rect 59696 -56320 59706 -55970
rect 59856 -56140 59976 -56130
rect 59856 -56230 59866 -56140
rect 59966 -56230 59976 -56140
rect 59856 -56240 59976 -56230
rect 60436 -56220 60446 -56120
rect 60526 -56220 60536 -56120
rect 60436 -56240 60536 -56220
rect 59636 -56330 59706 -56320
rect 59696 -56390 59706 -56330
rect 59636 -56410 59706 -56390
rect 59756 -56260 60536 -56240
rect 59756 -56300 59866 -56260
rect 60426 -56300 60536 -56260
rect 59756 -56310 60536 -56300
rect 59756 -56350 59826 -56310
rect 59066 -56440 59176 -56430
rect 58896 -56550 58986 -56486
rect 59066 -56510 59076 -56440
rect 59166 -56510 59176 -56440
rect 59066 -56512 59103 -56510
rect 59137 -56512 59176 -56510
rect 59066 -56520 59176 -56512
rect 59756 -56540 59766 -56350
rect 59806 -56540 59826 -56350
rect 59956 -56368 60046 -56340
rect 59946 -56374 60046 -56368
rect 60126 -56368 60336 -56340
rect 60126 -56374 60346 -56368
rect 59856 -56410 59916 -56400
rect 59946 -56408 59958 -56374
rect 60334 -56408 60346 -56374
rect 59946 -56414 60346 -56408
rect 60376 -56420 60446 -56410
rect 59856 -56490 59916 -56480
rect 59946 -56482 60346 -56476
rect 59946 -56516 59958 -56482
rect 60334 -56516 60346 -56482
rect 60376 -56490 60446 -56480
rect 59946 -56522 59976 -56516
rect 57098 -56558 57368 -56554
rect 57096 -56564 57372 -56558
rect 57096 -56650 57098 -56564
rect 56424 -56688 56470 -56687
rect 56060 -57160 56356 -57148
rect 56410 -56699 56470 -56688
rect 53400 -57208 53504 -57196
rect 53400 -57518 53464 -57208
rect 53250 -57908 53464 -57518
rect 53000 -57984 53464 -57908
rect 53498 -57984 53504 -57208
rect 53000 -57988 53504 -57984
rect 53458 -57996 53504 -57988
rect 53636 -57208 53760 -57196
rect 53636 -57984 53642 -57208
rect 53676 -57984 53760 -57208
rect 53930 -57184 54730 -57178
rect 53930 -57218 53942 -57184
rect 54718 -57218 54730 -57184
rect 53930 -57224 54730 -57218
rect 53830 -57246 53900 -57228
rect 53830 -57334 53858 -57246
rect 53892 -57334 53900 -57246
rect 53830 -57528 53900 -57334
rect 54760 -57246 54850 -57228
rect 54760 -57334 54768 -57246
rect 54802 -57248 54850 -57246
rect 54900 -57238 55200 -57168
rect 55870 -57170 55982 -57164
rect 55870 -57204 55882 -57170
rect 55970 -57204 55982 -57170
rect 55450 -57238 55810 -57208
rect 55870 -57210 55982 -57204
rect 56060 -57238 56300 -57160
rect 54900 -57242 55820 -57238
rect 56000 -57242 56300 -57238
rect 54900 -57248 55860 -57242
rect 54840 -57328 54850 -57248
rect 54802 -57334 54850 -57328
rect 54760 -57348 54850 -57334
rect 55130 -57254 55860 -57248
rect 55130 -57278 55820 -57254
rect 55130 -57296 55510 -57278
rect 55130 -57330 55142 -57296
rect 55494 -57298 55510 -57296
rect 55494 -57330 55506 -57298
rect 55130 -57336 55506 -57330
rect 53930 -57362 54730 -57356
rect 53930 -57396 53942 -57362
rect 54718 -57396 54730 -57362
rect 55020 -57382 55090 -57368
rect 53930 -57402 54730 -57396
rect 53940 -57408 54730 -57402
rect 54920 -57398 54980 -57388
rect 53940 -57448 54920 -57408
rect 53830 -57538 53920 -57528
rect 53830 -57648 53850 -57538
rect 53830 -57658 53920 -57648
rect 54320 -57948 54510 -57448
rect 54710 -57468 54920 -57448
rect 54910 -57478 54980 -57468
rect 55020 -57416 55046 -57382
rect 55080 -57416 55090 -57382
rect 55020 -57528 55090 -57416
rect 55142 -57462 55494 -57336
rect 55540 -57382 55620 -57368
rect 55540 -57416 55556 -57382
rect 55590 -57416 55620 -57382
rect 55130 -57468 55506 -57462
rect 55130 -57502 55142 -57468
rect 55494 -57502 55506 -57468
rect 55130 -57508 55506 -57502
rect 55000 -57538 55090 -57528
rect 55000 -57648 55090 -57638
rect 55540 -57528 55620 -57416
rect 55540 -57538 55630 -57528
rect 55630 -57638 55680 -57548
rect 55540 -57648 55680 -57638
rect 55274 -57738 55320 -57736
rect 55220 -57748 55320 -57738
rect 55220 -57924 55280 -57918
rect 55314 -57924 55320 -57748
rect 55220 -57928 55320 -57924
rect 55274 -57936 55320 -57928
rect 55362 -57748 55408 -57736
rect 55362 -57924 55368 -57748
rect 55402 -57758 55510 -57748
rect 55402 -57924 55410 -57758
rect 55362 -57928 55410 -57924
rect 55500 -57928 55510 -57758
rect 55362 -57936 55510 -57928
rect 55390 -57938 55510 -57936
rect 53636 -57988 53760 -57984
rect 53636 -57996 53682 -57988
rect 53940 -58008 54020 -57968
rect 54080 -57982 54860 -57948
rect 55311 -57974 55371 -57968
rect 53514 -58034 53626 -58028
rect 53514 -58038 53526 -58034
rect 25870 -58072 35740 -58066
rect 25900 -58200 35740 -58072
rect 53510 -58068 53526 -58038
rect 53614 -58038 53626 -58034
rect 53614 -58068 53630 -58038
rect 53510 -58128 53630 -58068
rect 53940 -58088 53950 -58008
rect 54010 -58038 54020 -58008
rect 54069 -57988 54869 -57982
rect 54069 -58022 54081 -57988
rect 54857 -58022 54869 -57988
rect 54069 -58028 54869 -58022
rect 54910 -57998 54980 -57988
rect 54010 -58050 54028 -58038
rect 54022 -58088 54028 -58050
rect 53940 -58100 54028 -58088
rect 53940 -58108 54020 -58100
rect 54910 -58108 54980 -58098
rect 55311 -58008 55324 -57974
rect 55358 -58008 55371 -57974
rect 54070 -58110 54870 -58108
rect 24400 -58800 36000 -58200
rect 54069 -58116 54870 -58110
rect 54069 -58138 54081 -58116
rect 54041 -58150 54081 -58138
rect 54857 -58118 54870 -58116
rect 54857 -58150 54880 -58118
rect 55311 -58148 55371 -58008
rect 54041 -58158 54880 -58150
rect 55240 -58158 55371 -58148
rect 54041 -58168 55240 -58158
rect 53510 -58258 53630 -58248
rect 53961 -58208 55240 -58168
rect 53961 -58406 54031 -58208
rect 54730 -58268 54860 -58258
rect 54730 -58288 54740 -58268
rect 54080 -58338 54740 -58288
rect 54069 -58344 54740 -58338
rect 54850 -58338 54860 -58268
rect 54850 -58344 54869 -58338
rect 54069 -58378 54081 -58344
rect 54857 -58378 54869 -58344
rect 54069 -58384 54869 -58378
rect 54911 -58394 54981 -58208
rect 55370 -58208 55371 -58158
rect 55240 -58228 55370 -58218
rect 55410 -58248 55510 -57938
rect 55410 -58358 55510 -58338
rect 55570 -58268 55680 -57648
rect 55780 -58030 55820 -57278
rect 55854 -58030 55860 -57254
rect 55780 -58038 55860 -58030
rect 55814 -58042 55860 -58038
rect 55992 -57254 56300 -57242
rect 55992 -58030 55998 -57254
rect 56032 -58028 56300 -57254
rect 56410 -57298 56430 -56699
rect 56380 -57475 56430 -57298
rect 56464 -57475 56470 -56699
rect 56380 -57487 56470 -57475
rect 56552 -56699 56750 -56687
rect 56552 -57475 56558 -56699
rect 56592 -56838 56750 -56699
rect 57066 -56680 57098 -56650
rect 57368 -56650 57372 -56564
rect 58896 -56559 59076 -56550
rect 58896 -56560 59084 -56559
rect 59156 -56560 59202 -56559
rect 57368 -56680 57396 -56650
rect 57066 -56810 57086 -56680
rect 57376 -56810 57396 -56680
rect 56592 -57475 56610 -56838
rect 57066 -56840 57396 -56810
rect 56860 -56990 57060 -56978
rect 56860 -57018 57236 -56990
rect 56860 -57148 56900 -57018
rect 57020 -57148 57236 -57018
rect 56860 -57188 57236 -57148
rect 57036 -57190 57236 -57188
rect 58556 -57080 58756 -57060
rect 58556 -57240 58576 -57080
rect 58736 -57240 58756 -57080
rect 58556 -57260 58756 -57240
rect 56552 -57478 56610 -57475
rect 57036 -57340 57446 -57330
rect 56552 -57487 56598 -57478
rect 57036 -57480 57056 -57340
rect 57416 -57480 57446 -57340
rect 56380 -57758 56440 -57487
rect 57036 -57500 57098 -57480
rect 56480 -57528 56550 -57518
rect 56480 -57598 56550 -57588
rect 57096 -57614 57098 -57534
rect 57368 -57500 57446 -57480
rect 57368 -57614 57372 -57534
rect 57096 -57630 57372 -57614
rect 58896 -57690 58926 -56560
rect 58966 -56571 59086 -56560
rect 58966 -56947 59044 -56571
rect 59078 -56947 59086 -56571
rect 58966 -56970 59086 -56947
rect 59156 -56571 59256 -56560
rect 59756 -56570 59826 -56540
rect 59966 -56552 59976 -56522
rect 60316 -56522 60346 -56516
rect 61036 -56520 61466 -56510
rect 60316 -56552 60326 -56522
rect 59966 -56560 60326 -56552
rect 59156 -56947 59162 -56571
rect 59196 -56640 59256 -56571
rect 59236 -56720 59256 -56640
rect 59196 -56840 59256 -56720
rect 59236 -56920 59256 -56840
rect 59196 -56947 59256 -56920
rect 59156 -56960 59256 -56947
rect 58966 -57280 59036 -56970
rect 59066 -57006 59176 -57000
rect 59066 -57010 59103 -57006
rect 59137 -57010 59176 -57006
rect 59066 -57080 59076 -57010
rect 59166 -57080 59176 -57010
rect 59066 -57090 59176 -57080
rect 59206 -57160 59256 -56960
rect 59376 -56590 59826 -56570
rect 59376 -56630 59476 -56590
rect 59656 -56630 59826 -56590
rect 59376 -56640 59826 -56630
rect 59376 -56690 59436 -56640
rect 59376 -57050 59386 -56690
rect 59426 -57050 59436 -56690
rect 59526 -56698 59576 -56670
rect 59526 -56732 59546 -56698
rect 59636 -56730 59706 -56670
rect 59580 -56732 59706 -56730
rect 59526 -56740 59706 -56732
rect 59476 -56782 59546 -56770
rect 59476 -56850 59502 -56782
rect 59476 -56958 59502 -56920
rect 59536 -56958 59546 -56782
rect 59476 -56970 59546 -56958
rect 59576 -56782 59636 -56770
rect 59576 -56790 59590 -56782
rect 59624 -56790 59636 -56782
rect 59576 -56970 59636 -56960
rect 59534 -57008 59592 -57002
rect 59534 -57010 59546 -57008
rect 59066 -57170 59176 -57160
rect 59066 -57240 59076 -57170
rect 59166 -57240 59176 -57170
rect 59066 -57242 59103 -57240
rect 59137 -57242 59176 -57240
rect 59066 -57250 59176 -57242
rect 59206 -57170 59266 -57160
rect 59206 -57250 59266 -57240
rect 59376 -57200 59436 -57050
rect 59516 -57042 59546 -57010
rect 59580 -57010 59592 -57008
rect 59666 -57010 59706 -56740
rect 59580 -57042 59706 -57010
rect 59516 -57080 59706 -57042
rect 59746 -56698 59936 -56670
rect 59746 -56732 59862 -56698
rect 59896 -56732 59936 -56698
rect 59746 -56740 59936 -56732
rect 61036 -56700 61206 -56520
rect 61346 -56700 61466 -56520
rect 61036 -56740 61466 -56700
rect 59746 -57000 59776 -56740
rect 60286 -56750 60476 -56740
rect 59806 -56782 59866 -56770
rect 59806 -56800 59818 -56782
rect 59852 -56800 59866 -56782
rect 59806 -56958 59818 -56940
rect 59852 -56958 59866 -56940
rect 59806 -56970 59866 -56958
rect 59900 -56780 60016 -56770
rect 59900 -56782 59916 -56780
rect 59900 -56958 59906 -56782
rect 59900 -56960 59916 -56958
rect 60006 -56960 60016 -56780
rect 60286 -56890 60306 -56750
rect 60456 -56890 60476 -56750
rect 61176 -56800 61386 -56780
rect 60286 -56900 60476 -56890
rect 61026 -56820 61136 -56810
rect 59900 -56970 60016 -56960
rect 60076 -56957 60196 -56920
rect 60076 -56991 60127 -56957
rect 60161 -56991 60196 -56957
rect 59746 -57008 59926 -57000
rect 59746 -57010 59862 -57008
rect 59896 -57010 59926 -57008
rect 59746 -57080 59826 -57010
rect 59916 -57080 59926 -57010
rect 59746 -57090 59926 -57080
rect 60076 -57049 60196 -56991
rect 60336 -56960 60446 -56900
rect 60336 -57000 60366 -56960
rect 60406 -57000 60446 -56960
rect 60636 -56957 60816 -56920
rect 60636 -56991 60671 -56957
rect 60705 -56991 60747 -56957
rect 60781 -56991 60816 -56957
rect 60076 -57080 60127 -57049
rect 60161 -57080 60196 -57049
rect 59736 -57170 59936 -57160
rect 58966 -57301 59086 -57280
rect 58966 -57677 59044 -57301
rect 59078 -57677 59086 -57301
rect 58966 -57690 59086 -57677
rect 59156 -57290 59202 -57289
rect 59156 -57301 59236 -57290
rect 59156 -57677 59162 -57301
rect 59196 -57330 59236 -57301
rect 59226 -57410 59236 -57330
rect 59196 -57560 59236 -57410
rect 59226 -57640 59236 -57560
rect 59196 -57677 59236 -57640
rect 59376 -57570 59386 -57200
rect 59426 -57570 59436 -57200
rect 59516 -57211 59706 -57170
rect 59516 -57245 59545 -57211
rect 59579 -57245 59706 -57211
rect 59516 -57250 59706 -57245
rect 59533 -57251 59591 -57250
rect 59466 -57295 59546 -57280
rect 59586 -57283 59646 -57280
rect 59466 -57330 59501 -57295
rect 59466 -57471 59501 -57410
rect 59535 -57471 59546 -57295
rect 59466 -57480 59546 -57471
rect 59583 -57295 59646 -57283
rect 59583 -57310 59589 -57295
rect 59623 -57310 59646 -57295
rect 59583 -57450 59586 -57310
rect 59583 -57471 59589 -57450
rect 59623 -57471 59646 -57450
rect 59583 -57480 59646 -57471
rect 59495 -57483 59541 -57480
rect 59583 -57483 59629 -57480
rect 59533 -57520 59591 -57515
rect 59676 -57520 59706 -57250
rect 59376 -57610 59436 -57570
rect 59506 -57580 59516 -57520
rect 59596 -57580 59706 -57520
rect 59736 -57240 59826 -57170
rect 59926 -57240 59936 -57170
rect 59736 -57245 59861 -57240
rect 59895 -57245 59936 -57240
rect 59736 -57250 59936 -57245
rect 60076 -57240 60096 -57080
rect 60176 -57240 60196 -57080
rect 59736 -57520 59766 -57250
rect 59849 -57251 59907 -57250
rect 60076 -57267 60127 -57240
rect 60161 -57267 60196 -57240
rect 59796 -57283 59856 -57280
rect 59796 -57290 59857 -57283
rect 59856 -57470 59857 -57290
rect 59796 -57471 59817 -57470
rect 59851 -57471 59857 -57470
rect 59796 -57480 59857 -57471
rect 59811 -57483 59857 -57480
rect 59899 -57290 59945 -57283
rect 59899 -57295 59916 -57290
rect 59899 -57471 59905 -57295
rect 59899 -57480 59916 -57471
rect 60006 -57480 60016 -57290
rect 60076 -57325 60196 -57267
rect 60346 -57050 60426 -57000
rect 60346 -57090 60366 -57050
rect 60406 -57090 60426 -57050
rect 60346 -57140 60426 -57090
rect 60346 -57180 60366 -57140
rect 60406 -57180 60426 -57140
rect 60346 -57220 60426 -57180
rect 60346 -57260 60366 -57220
rect 60406 -57260 60426 -57220
rect 60346 -57270 60426 -57260
rect 60636 -57049 60816 -56991
rect 60636 -57083 60671 -57049
rect 60705 -57083 60747 -57049
rect 60781 -57083 60816 -57049
rect 60636 -57141 60816 -57083
rect 60636 -57175 60671 -57141
rect 60705 -57175 60747 -57141
rect 60781 -57175 60816 -57141
rect 60636 -57233 60816 -57175
rect 60636 -57267 60671 -57233
rect 60705 -57267 60747 -57233
rect 60781 -57267 60816 -57233
rect 60076 -57359 60127 -57325
rect 60161 -57359 60196 -57325
rect 60076 -57390 60196 -57359
rect 60276 -57310 60546 -57300
rect 60276 -57325 60476 -57310
rect 60276 -57359 60297 -57325
rect 60331 -57359 60369 -57325
rect 60405 -57359 60449 -57325
rect 60276 -57370 60476 -57359
rect 60536 -57370 60546 -57310
rect 60276 -57380 60546 -57370
rect 60636 -57325 60816 -57267
rect 61026 -56930 61036 -56820
rect 61126 -56930 61136 -56820
rect 61176 -56880 61196 -56800
rect 61366 -56880 61386 -56800
rect 61176 -56900 61386 -56880
rect 61026 -56960 61136 -56930
rect 61026 -57000 61046 -56960
rect 61086 -57000 61136 -56960
rect 61026 -57050 61136 -57000
rect 61026 -57090 61046 -57050
rect 61086 -57090 61136 -57050
rect 61026 -57140 61136 -57090
rect 61026 -57180 61046 -57140
rect 61086 -57180 61136 -57140
rect 61026 -57220 61136 -57180
rect 61026 -57260 61046 -57220
rect 61086 -57260 61136 -57220
rect 61026 -57280 61136 -57260
rect 61256 -56957 61366 -56900
rect 61256 -56991 61291 -56957
rect 61325 -56991 61366 -56957
rect 61256 -57049 61366 -56991
rect 61256 -57050 61291 -57049
rect 61325 -57050 61366 -57049
rect 61256 -57260 61276 -57050
rect 61356 -57260 61366 -57050
rect 61256 -57267 61291 -57260
rect 61325 -57267 61366 -57260
rect 60636 -57359 60671 -57325
rect 60705 -57359 60747 -57325
rect 60781 -57359 60816 -57325
rect 60636 -57440 60816 -57359
rect 60966 -57324 61177 -57310
rect 60966 -57325 61129 -57324
rect 60966 -57359 60980 -57325
rect 61015 -57359 61053 -57325
rect 61088 -57358 61129 -57325
rect 61164 -57358 61177 -57324
rect 61088 -57359 61177 -57358
rect 60966 -57390 61177 -57359
rect 61256 -57325 61366 -57267
rect 61256 -57359 61291 -57325
rect 61325 -57359 61366 -57325
rect 61256 -57390 61366 -57359
rect 60466 -57450 60546 -57440
rect 59899 -57483 59945 -57480
rect 60466 -57510 60476 -57450
rect 60536 -57510 60546 -57450
rect 59849 -57520 59907 -57515
rect 60466 -57520 60546 -57510
rect 60606 -57450 60826 -57440
rect 60606 -57510 60616 -57450
rect 60736 -57510 60756 -57450
rect 60816 -57510 60826 -57450
rect 60606 -57520 60826 -57510
rect 60886 -57450 60966 -57440
rect 60886 -57510 60896 -57450
rect 60956 -57510 60966 -57450
rect 60886 -57520 60966 -57510
rect 59736 -57521 59926 -57520
rect 59736 -57555 59861 -57521
rect 59895 -57555 59926 -57521
rect 59736 -57580 59926 -57555
rect 60636 -57570 60816 -57520
rect 59376 -57620 59826 -57610
rect 59376 -57660 59476 -57620
rect 59646 -57660 59826 -57620
rect 59376 -57670 59826 -57660
rect 59156 -57690 59236 -57677
rect 58896 -57700 59086 -57690
rect 56380 -57768 57000 -57758
rect 57356 -57764 57676 -57750
rect 56440 -57774 57000 -57768
rect 57314 -57770 57676 -57764
rect 56440 -57794 57178 -57774
rect 56440 -57844 57118 -57794
rect 57168 -57844 57178 -57794
rect 57314 -57810 57326 -57770
rect 57376 -57810 57676 -57770
rect 57314 -57816 57676 -57810
rect 57356 -57830 57676 -57816
rect 56440 -57854 57178 -57844
rect 56440 -57888 57000 -57854
rect 57112 -57856 57174 -57854
rect 56380 -57958 57000 -57888
rect 56032 -58030 56038 -58028
rect 55992 -58042 56038 -58030
rect 55880 -58074 55970 -58068
rect 55870 -58078 55982 -58074
rect 55870 -58120 55880 -58078
rect 55970 -58120 55982 -58078
rect 55880 -58168 55970 -58158
rect 56120 -58198 56300 -58028
rect 57096 -58109 57372 -58078
rect 57096 -58143 57125 -58109
rect 57159 -58143 57217 -58109
rect 57251 -58143 57309 -58109
rect 57343 -58120 57372 -58109
rect 57343 -58143 57376 -58120
rect 57096 -58180 57376 -58143
rect 57066 -58190 57376 -58180
rect 56426 -58198 57376 -58190
rect 56120 -58208 57376 -58198
rect 56014 -58258 56086 -58246
rect 55570 -58378 55830 -58268
rect 53961 -58444 53988 -58406
rect 54022 -58444 54031 -58406
rect 53961 -58458 54031 -58444
rect 54910 -58406 54981 -58394
rect 54910 -58444 54916 -58406
rect 54950 -58444 54981 -58406
rect 54910 -58456 54981 -58444
rect 54911 -58458 54981 -58456
rect 55220 -58418 55330 -58408
rect 54069 -58472 54869 -58466
rect 54069 -58506 54081 -58472
rect 54857 -58478 54869 -58472
rect 54857 -58506 54880 -58478
rect 54069 -58512 54880 -58506
rect 54090 -58588 54880 -58512
rect 55330 -58518 55380 -58418
rect 55330 -58528 55480 -58518
rect 55220 -58538 55480 -58528
rect 55280 -58552 55480 -58538
rect 55280 -58558 55488 -58552
rect 55280 -58578 55300 -58558
rect 54090 -58688 54150 -58588
rect 54840 -58688 54880 -58588
rect 55288 -58592 55300 -58578
rect 55476 -58592 55488 -58558
rect 55530 -58578 55610 -58568
rect 55288 -58598 55488 -58592
rect 55520 -58602 55530 -58590
rect 55520 -58636 55526 -58602
rect 55288 -58646 55488 -58640
rect 55288 -58680 55300 -58646
rect 55476 -58680 55488 -58646
rect 55520 -58648 55530 -58636
rect 55530 -58678 55610 -58668
rect 55288 -58686 55488 -58680
rect 54090 -58708 54140 -58688
rect 14600 -60000 20200 -59400
rect 14600 -60800 15200 -60000
rect 10600 -64200 15200 -60800
rect 14600 -64800 15200 -64200
rect 19600 -64800 20200 -60000
rect 14600 -65400 20200 -64800
rect 24400 -64800 25000 -58800
rect 35400 -64800 36000 -58800
rect 54100 -58948 54140 -58708
rect 54850 -58948 54880 -58688
rect 55300 -58728 55470 -58686
rect 55300 -58868 55320 -58728
rect 55470 -58814 55482 -58742
rect 55300 -58878 55470 -58868
rect 54100 -58988 54880 -58948
rect 55710 -59198 55830 -58378
rect 56014 -58408 56020 -58258
rect 56080 -58408 56086 -58258
rect 56014 -58420 56086 -58408
rect 56120 -58408 56170 -58208
rect 56390 -58260 57376 -58208
rect 56390 -58268 57156 -58260
rect 56390 -58408 56654 -58268
rect 56120 -58458 56654 -58408
rect 56306 -58486 56654 -58458
rect 56998 -58420 57156 -58268
rect 57316 -58420 57376 -58260
rect 56998 -58486 57376 -58420
rect 56306 -58900 57376 -58486
rect 57556 -58610 57676 -57830
rect 58896 -57860 58986 -57700
rect 59756 -57720 59826 -57670
rect 59066 -57736 59176 -57730
rect 59066 -57740 59103 -57736
rect 59137 -57740 59176 -57736
rect 59066 -57800 59076 -57740
rect 59166 -57800 59176 -57740
rect 59066 -57810 59176 -57800
rect 58896 -58230 58926 -57860
rect 58966 -58230 58986 -57930
rect 59116 -57860 59506 -57840
rect 59116 -57930 59146 -57860
rect 59226 -57930 59276 -57860
rect 59356 -57930 59396 -57860
rect 59476 -57930 59506 -57860
rect 59116 -57948 59506 -57930
rect 59646 -57860 59716 -57840
rect 59706 -57920 59716 -57860
rect 59646 -57930 59716 -57920
rect 59113 -57954 59513 -57948
rect 59113 -57988 59125 -57954
rect 59501 -57988 59513 -57954
rect 59113 -57994 59513 -57988
rect 59546 -58000 59616 -57990
rect 59246 -58056 59256 -58030
rect 59113 -58062 59256 -58056
rect 59366 -58056 59376 -58030
rect 59366 -58062 59513 -58056
rect 59016 -58100 59076 -58080
rect 59113 -58096 59125 -58062
rect 59501 -58096 59513 -58062
rect 59606 -58060 59616 -58000
rect 59546 -58070 59616 -58060
rect 59113 -58102 59513 -58096
rect 59016 -58190 59076 -58160
rect 59113 -58170 59513 -58164
rect 59113 -58204 59125 -58170
rect 59501 -58204 59513 -58170
rect 59113 -58210 59513 -58204
rect 58896 -58300 58906 -58230
rect 58896 -58320 58986 -58300
rect 59116 -58230 59516 -58210
rect 59116 -58300 59146 -58230
rect 59226 -58300 59276 -58230
rect 59356 -58300 59396 -58230
rect 59476 -58300 59516 -58230
rect 59116 -58320 59516 -58300
rect 59646 -58230 59656 -57930
rect 59706 -58230 59716 -57930
rect 59756 -57900 59766 -57720
rect 59806 -57900 59826 -57720
rect 59956 -57720 60336 -57710
rect 59956 -57734 59966 -57720
rect 59946 -57740 59966 -57734
rect 60326 -57734 60336 -57720
rect 60326 -57740 60346 -57734
rect 59856 -57780 59916 -57770
rect 59946 -57774 59958 -57740
rect 60334 -57774 60346 -57740
rect 61056 -57740 61176 -57390
rect 59946 -57780 59966 -57774
rect 60326 -57780 60346 -57774
rect 60376 -57780 60436 -57760
rect 59956 -57790 60336 -57780
rect 59856 -57860 59916 -57840
rect 59946 -57848 60346 -57842
rect 59756 -57940 59826 -57900
rect 59946 -57882 59958 -57848
rect 60334 -57882 60346 -57848
rect 60376 -57860 60436 -57840
rect 61126 -57840 61176 -57740
rect 61056 -57870 61176 -57840
rect 59946 -57888 60346 -57882
rect 59946 -57940 60336 -57888
rect 59756 -57960 60536 -57940
rect 59756 -58000 59866 -57960
rect 60426 -58000 60536 -57960
rect 59756 -58010 60536 -58000
rect 59796 -58120 59806 -58010
rect 59916 -58120 59926 -58010
rect 59796 -58130 59926 -58120
rect 60436 -58030 60536 -58010
rect 60436 -58150 60446 -58030
rect 60526 -58150 60536 -58030
rect 60436 -58160 60536 -58150
rect 59646 -58240 59716 -58230
rect 59706 -58300 59716 -58240
rect 59646 -58320 59716 -58300
rect 58806 -58610 59356 -58580
rect 57556 -58620 59356 -58610
rect 57556 -58760 58986 -58620
rect 59126 -58760 59356 -58620
rect 59846 -58590 60256 -58580
rect 59846 -58700 59996 -58590
rect 60106 -58700 60256 -58590
rect 57556 -58810 59356 -58760
rect 58806 -58890 59356 -58810
rect 55710 -59200 55910 -59198
rect 55400 -59300 56200 -59200
rect 59600 -59300 60500 -58700
rect 55400 -59700 55500 -59300
rect 56100 -59700 56200 -59300
rect 55400 -59800 56200 -59700
rect 55380 -60280 55800 -60200
rect 55380 -60560 55460 -60280
rect 55720 -60560 55800 -60280
rect 55380 -60640 55800 -60560
rect 54090 -60738 54890 -60698
rect 54090 -60868 54150 -60738
rect 53510 -60920 53800 -60918
rect 53460 -60940 53800 -60920
rect 53460 -61140 53480 -60940
rect 53780 -61140 53800 -60940
rect 54080 -60998 54150 -60868
rect 54860 -60978 54890 -60738
rect 54850 -60998 54890 -60978
rect 54080 -61066 54880 -60998
rect 54079 -61072 54880 -61066
rect 54079 -61106 54091 -61072
rect 54867 -61098 54880 -61072
rect 54867 -61106 54879 -61098
rect 54079 -61112 54879 -61106
rect 53460 -61160 53800 -61140
rect 53510 -61258 53800 -61160
rect 53002 -61420 53480 -61358
rect 53000 -61558 53480 -61420
rect 53510 -61368 53520 -61258
rect 53640 -61368 53800 -61258
rect 53510 -61488 53800 -61368
rect 53970 -61134 54040 -61118
rect 53970 -61172 53998 -61134
rect 54032 -61172 54040 -61134
rect 53970 -61368 54040 -61172
rect 54920 -61134 54990 -61118
rect 54920 -61172 54926 -61134
rect 54960 -61172 54990 -61134
rect 54079 -61200 54879 -61194
rect 54079 -61234 54091 -61200
rect 54867 -61234 54879 -61200
rect 54079 -61238 54879 -61234
rect 54079 -61240 54750 -61238
rect 54090 -61288 54750 -61240
rect 54740 -61318 54750 -61288
rect 54850 -61240 54879 -61238
rect 54850 -61308 54860 -61240
rect 54840 -61318 54860 -61308
rect 54750 -61328 54860 -61318
rect 54920 -61368 54990 -61172
rect 55430 -61218 55520 -61208
rect 55290 -61328 55390 -61318
rect 53970 -61398 55290 -61368
rect 55430 -61358 55520 -61288
rect 53970 -61408 55390 -61398
rect 54050 -61418 55380 -61408
rect 54050 -61428 54880 -61418
rect 54050 -61438 54091 -61428
rect 54079 -61462 54091 -61438
rect 54867 -61438 54880 -61428
rect 54867 -61462 54879 -61438
rect 54079 -61468 54879 -61462
rect 54920 -61478 54990 -61468
rect 53510 -61506 53630 -61488
rect 53510 -61538 53526 -61506
rect 53514 -61540 53526 -61538
rect 53614 -61538 53630 -61506
rect 53940 -61490 54038 -61478
rect 53940 -61498 53998 -61490
rect 53614 -61540 53626 -61538
rect 53514 -61546 53626 -61540
rect 53000 -63308 53050 -61558
rect 53250 -61568 53480 -61558
rect 53250 -62918 53330 -61568
rect 53400 -61578 53480 -61568
rect 53400 -61590 53504 -61578
rect 53400 -62366 53464 -61590
rect 53498 -62366 53504 -61590
rect 53400 -62378 53504 -62366
rect 53636 -61588 53682 -61578
rect 53636 -61590 53760 -61588
rect 53636 -62366 53642 -61590
rect 53676 -62366 53760 -61590
rect 53940 -61598 53950 -61498
rect 54032 -61528 54038 -61490
rect 54020 -61540 54038 -61528
rect 54020 -61598 54030 -61540
rect 54079 -61556 54879 -61550
rect 54079 -61590 54091 -61556
rect 54867 -61590 54879 -61556
rect 54920 -61578 54990 -61568
rect 55320 -61568 55380 -61418
rect 54079 -61596 54879 -61590
rect 53940 -61618 54030 -61598
rect 54090 -61628 54870 -61596
rect 55320 -61602 55334 -61568
rect 55368 -61602 55380 -61568
rect 55320 -61608 55380 -61602
rect 53840 -61928 53920 -61918
rect 53840 -62038 53860 -61928
rect 53840 -62048 53920 -62038
rect 53840 -62240 53900 -62048
rect 54320 -62128 54510 -61628
rect 55440 -61638 55520 -61358
rect 55410 -61640 55520 -61638
rect 55284 -61648 55330 -61640
rect 55230 -61652 55330 -61648
rect 55230 -61658 55290 -61652
rect 55324 -61828 55330 -61652
rect 55230 -61838 55330 -61828
rect 55284 -61840 55330 -61838
rect 55372 -61648 55520 -61640
rect 55372 -61652 55430 -61648
rect 55372 -61828 55378 -61652
rect 55412 -61818 55430 -61652
rect 55510 -61818 55520 -61648
rect 55412 -61828 55520 -61818
rect 55372 -61840 55418 -61828
rect 55580 -61928 55720 -60640
rect 58776 -60870 59306 -60750
rect 58776 -60880 58966 -60870
rect 56146 -60980 57366 -60930
rect 55954 -61128 56046 -61116
rect 56146 -61128 56506 -60980
rect 55954 -61298 55960 -61128
rect 56040 -61298 56046 -61128
rect 55954 -61310 56046 -61298
rect 56120 -61158 56506 -61128
rect 56120 -61368 56190 -61158
rect 56390 -61230 56506 -61158
rect 57016 -61134 57366 -60980
rect 57586 -61030 58966 -60880
rect 59126 -61030 59306 -60870
rect 57586 -61050 59306 -61030
rect 59946 -60900 60386 -60800
rect 57586 -61080 58986 -61050
rect 59946 -61060 59956 -60900
rect 60166 -61060 60386 -60900
rect 57016 -61230 57368 -61134
rect 56390 -61270 57368 -61230
rect 56390 -61368 57126 -61270
rect 56120 -61374 57126 -61368
rect 56120 -61378 56750 -61374
rect 55880 -61418 55970 -61408
rect 55870 -61496 55880 -61450
rect 55970 -61496 55982 -61450
rect 55880 -61508 55970 -61498
rect 55000 -61938 55090 -61928
rect 55000 -62048 55090 -62038
rect 54710 -62128 54960 -62108
rect 53940 -62168 54960 -62128
rect 53940 -62172 54730 -62168
rect 53930 -62178 54730 -62172
rect 53930 -62212 53942 -62178
rect 54718 -62212 54730 -62178
rect 53930 -62218 54730 -62212
rect 53840 -62328 53858 -62240
rect 53892 -62328 53900 -62240
rect 53840 -62348 53900 -62328
rect 54762 -62238 54850 -62228
rect 54762 -62240 54770 -62238
rect 54762 -62328 54768 -62240
rect 54840 -62328 54850 -62238
rect 54762 -62340 54850 -62328
rect 54770 -62348 54850 -62340
rect 53636 -62378 53760 -62366
rect 53400 -62596 53480 -62378
rect 53514 -62416 53626 -62410
rect 53514 -62418 53526 -62416
rect 53510 -62450 53526 -62418
rect 53614 -62418 53626 -62416
rect 53614 -62450 53630 -62418
rect 53510 -62524 53630 -62450
rect 53510 -62558 53526 -62524
rect 53614 -62558 53630 -62524
rect 53680 -62438 53760 -62378
rect 53930 -62356 54730 -62350
rect 53930 -62390 53942 -62356
rect 54718 -62390 54730 -62356
rect 53930 -62396 54730 -62390
rect 53940 -62428 54720 -62396
rect 53920 -62438 54720 -62428
rect 53680 -62528 54720 -62438
rect 53514 -62564 53626 -62558
rect 53680 -62596 53760 -62528
rect 53920 -62538 54720 -62528
rect 53940 -62578 54720 -62538
rect 54900 -62568 54960 -62168
rect 55010 -62160 55090 -62048
rect 55540 -61938 55720 -61928
rect 55630 -62038 55720 -61938
rect 55130 -62074 55506 -62068
rect 55130 -62108 55142 -62074
rect 55494 -62108 55506 -62074
rect 55130 -62114 55506 -62108
rect 55010 -62194 55046 -62160
rect 55080 -62194 55090 -62160
rect 55010 -62208 55090 -62194
rect 55142 -62240 55494 -62114
rect 55540 -62160 55720 -62038
rect 55540 -62194 55556 -62160
rect 55590 -62194 55720 -62160
rect 55540 -62208 55720 -62194
rect 55780 -61540 55860 -61528
rect 55130 -62246 55506 -62240
rect 55130 -62280 55142 -62246
rect 55494 -62278 55506 -62246
rect 55494 -62280 55510 -62278
rect 55130 -62286 55510 -62280
rect 55140 -62298 55510 -62286
rect 55780 -62298 55820 -61540
rect 55140 -62316 55820 -62298
rect 55854 -62316 55860 -61540
rect 55140 -62328 55860 -62316
rect 55992 -61540 56038 -61528
rect 55992 -62316 55998 -61540
rect 56032 -61548 56038 -61540
rect 56120 -61548 56300 -61378
rect 57098 -61400 57126 -61374
rect 57356 -61400 57368 -61270
rect 57098 -61414 57368 -61400
rect 57096 -61445 57372 -61414
rect 57096 -61479 57125 -61445
rect 57159 -61479 57217 -61445
rect 57251 -61479 57309 -61445
rect 57343 -61479 57372 -61445
rect 57096 -61510 57372 -61479
rect 56032 -61906 56300 -61548
rect 56590 -61668 56660 -61658
rect 56660 -61734 57000 -61668
rect 57586 -61730 57706 -61080
rect 59946 -61090 60386 -61060
rect 57366 -61734 57706 -61730
rect 56660 -61738 57188 -61734
rect 56660 -61744 57190 -61738
rect 56660 -61794 57118 -61744
rect 57178 -61794 57190 -61744
rect 57314 -61740 57706 -61734
rect 57314 -61780 57326 -61740
rect 57366 -61780 57706 -61740
rect 57314 -61786 57706 -61780
rect 57366 -61790 57706 -61786
rect 58896 -61370 58986 -61350
rect 58896 -61430 58906 -61370
rect 58896 -61720 58926 -61430
rect 58966 -61720 58986 -61370
rect 59106 -61370 59516 -61360
rect 59106 -61430 59216 -61370
rect 59276 -61430 59326 -61370
rect 59386 -61430 59436 -61370
rect 59496 -61430 59516 -61370
rect 59106 -61447 59516 -61430
rect 59626 -61370 59706 -61330
rect 59626 -61430 59636 -61370
rect 59626 -61440 59656 -61430
rect 59106 -61480 59125 -61447
rect 59113 -61481 59125 -61480
rect 59501 -61480 59516 -61447
rect 59501 -61481 59513 -61480
rect 59113 -61487 59513 -61481
rect 59546 -61490 59616 -61480
rect 59276 -61530 59356 -61520
rect 59276 -61549 59286 -61530
rect 59113 -61555 59286 -61549
rect 59346 -61549 59356 -61530
rect 59346 -61555 59513 -61549
rect 59113 -61589 59125 -61555
rect 59501 -61589 59513 -61555
rect 59606 -61550 59616 -61490
rect 59546 -61560 59616 -61550
rect 59113 -61590 59286 -61589
rect 59346 -61590 59513 -61589
rect 59016 -61600 59076 -61590
rect 59113 -61595 59513 -61590
rect 59276 -61600 59356 -61595
rect 59546 -61610 59616 -61600
rect 59016 -61670 59076 -61660
rect 59113 -61663 59513 -61657
rect 59113 -61697 59125 -61663
rect 59501 -61697 59513 -61663
rect 59606 -61670 59616 -61610
rect 59546 -61680 59616 -61670
rect 59113 -61700 59513 -61697
rect 59113 -61703 59516 -61700
rect 58896 -61730 58986 -61720
rect 58896 -61790 58906 -61730
rect 58966 -61790 58986 -61730
rect 58896 -61792 58986 -61790
rect 59116 -61720 59516 -61703
rect 59646 -61710 59656 -61440
rect 59116 -61780 59216 -61720
rect 59276 -61780 59336 -61720
rect 59396 -61780 59436 -61720
rect 59496 -61780 59516 -61720
rect 56660 -61798 57190 -61794
rect 56590 -61800 57190 -61798
rect 56590 -61804 57188 -61800
rect 56590 -61868 57000 -61804
rect 56032 -61918 56356 -61906
rect 56032 -62316 56280 -61918
rect 55992 -62328 56280 -62316
rect 55140 -62338 55200 -62328
rect 55450 -62358 55810 -62328
rect 55870 -62366 55982 -62360
rect 55870 -62400 55882 -62366
rect 55970 -62400 55982 -62366
rect 55870 -62406 55982 -62400
rect 55140 -62418 55200 -62408
rect 55024 -62448 55116 -62436
rect 55024 -62528 55030 -62448
rect 55110 -62528 55116 -62448
rect 55024 -62540 55116 -62528
rect 55734 -62448 55816 -62436
rect 55734 -62528 55740 -62448
rect 55810 -62528 55816 -62448
rect 55734 -62540 55816 -62528
rect 55880 -62438 55970 -62406
rect 55880 -62564 55970 -62528
rect 56060 -62548 56280 -62328
rect 56350 -62548 56356 -61918
rect 56480 -61988 56550 -61978
rect 56480 -62058 56550 -62048
rect 56590 -62087 56750 -61868
rect 58894 -61886 58988 -61792
rect 59116 -61800 59516 -61780
rect 59636 -61720 59656 -61710
rect 59696 -61720 59706 -61370
rect 59856 -61540 59976 -61530
rect 59856 -61630 59866 -61540
rect 59966 -61630 59976 -61540
rect 59856 -61640 59976 -61630
rect 60436 -61620 60446 -61520
rect 60526 -61620 60536 -61520
rect 60436 -61640 60536 -61620
rect 59636 -61730 59706 -61720
rect 59696 -61790 59706 -61730
rect 59636 -61810 59706 -61790
rect 59756 -61660 60536 -61640
rect 59756 -61700 59866 -61660
rect 60426 -61700 60536 -61660
rect 59756 -61710 60536 -61700
rect 59756 -61750 59826 -61710
rect 59066 -61840 59176 -61830
rect 58896 -61950 58986 -61886
rect 59066 -61910 59076 -61840
rect 59166 -61910 59176 -61840
rect 59066 -61912 59103 -61910
rect 59137 -61912 59176 -61910
rect 59066 -61920 59176 -61912
rect 59756 -61940 59766 -61750
rect 59806 -61940 59826 -61750
rect 59956 -61768 60046 -61740
rect 59946 -61774 60046 -61768
rect 60126 -61768 60336 -61740
rect 60126 -61774 60346 -61768
rect 59856 -61810 59916 -61800
rect 59946 -61808 59958 -61774
rect 60334 -61808 60346 -61774
rect 59946 -61814 60346 -61808
rect 60376 -61820 60446 -61810
rect 59856 -61890 59916 -61880
rect 59946 -61882 60346 -61876
rect 59946 -61916 59958 -61882
rect 60334 -61916 60346 -61882
rect 60376 -61890 60446 -61880
rect 59946 -61922 59976 -61916
rect 57098 -61958 57368 -61954
rect 57096 -61964 57372 -61958
rect 57096 -62050 57098 -61964
rect 56424 -62088 56470 -62087
rect 56060 -62560 56356 -62548
rect 56410 -62099 56470 -62088
rect 53400 -62608 53504 -62596
rect 53400 -62918 53464 -62608
rect 53250 -63308 53464 -62918
rect 53000 -63384 53464 -63308
rect 53498 -63384 53504 -62608
rect 53000 -63388 53504 -63384
rect 53458 -63396 53504 -63388
rect 53636 -62608 53760 -62596
rect 53636 -63384 53642 -62608
rect 53676 -63384 53760 -62608
rect 53930 -62584 54730 -62578
rect 53930 -62618 53942 -62584
rect 54718 -62618 54730 -62584
rect 53930 -62624 54730 -62618
rect 53830 -62646 53900 -62628
rect 53830 -62734 53858 -62646
rect 53892 -62734 53900 -62646
rect 53830 -62928 53900 -62734
rect 54760 -62646 54850 -62628
rect 54760 -62734 54768 -62646
rect 54802 -62648 54850 -62646
rect 54900 -62638 55200 -62568
rect 55870 -62570 55982 -62564
rect 55870 -62604 55882 -62570
rect 55970 -62604 55982 -62570
rect 55450 -62638 55810 -62608
rect 55870 -62610 55982 -62604
rect 56060 -62638 56300 -62560
rect 54900 -62642 55820 -62638
rect 56000 -62642 56300 -62638
rect 54900 -62648 55860 -62642
rect 54840 -62728 54850 -62648
rect 54802 -62734 54850 -62728
rect 54760 -62748 54850 -62734
rect 55130 -62654 55860 -62648
rect 55130 -62678 55820 -62654
rect 55130 -62696 55510 -62678
rect 55130 -62730 55142 -62696
rect 55494 -62698 55510 -62696
rect 55494 -62730 55506 -62698
rect 55130 -62736 55506 -62730
rect 53930 -62762 54730 -62756
rect 53930 -62796 53942 -62762
rect 54718 -62796 54730 -62762
rect 55020 -62782 55090 -62768
rect 53930 -62802 54730 -62796
rect 53940 -62808 54730 -62802
rect 54920 -62798 54980 -62788
rect 53940 -62848 54920 -62808
rect 53830 -62938 53920 -62928
rect 53830 -63048 53850 -62938
rect 53830 -63058 53920 -63048
rect 54320 -63348 54510 -62848
rect 54710 -62868 54920 -62848
rect 54910 -62878 54980 -62868
rect 55020 -62816 55046 -62782
rect 55080 -62816 55090 -62782
rect 55020 -62928 55090 -62816
rect 55142 -62862 55494 -62736
rect 55540 -62782 55620 -62768
rect 55540 -62816 55556 -62782
rect 55590 -62816 55620 -62782
rect 55130 -62868 55506 -62862
rect 55130 -62902 55142 -62868
rect 55494 -62902 55506 -62868
rect 55130 -62908 55506 -62902
rect 55000 -62938 55090 -62928
rect 55000 -63048 55090 -63038
rect 55540 -62928 55620 -62816
rect 55540 -62938 55630 -62928
rect 55630 -63038 55680 -62948
rect 55540 -63048 55680 -63038
rect 55274 -63138 55320 -63136
rect 55220 -63148 55320 -63138
rect 55220 -63324 55280 -63318
rect 55314 -63324 55320 -63148
rect 55220 -63328 55320 -63324
rect 55274 -63336 55320 -63328
rect 55362 -63148 55408 -63136
rect 55362 -63324 55368 -63148
rect 55402 -63158 55510 -63148
rect 55402 -63324 55410 -63158
rect 55362 -63328 55410 -63324
rect 55500 -63328 55510 -63158
rect 55362 -63336 55510 -63328
rect 55390 -63338 55510 -63336
rect 53636 -63388 53760 -63384
rect 53636 -63396 53682 -63388
rect 53940 -63408 54020 -63368
rect 54080 -63382 54860 -63348
rect 55311 -63374 55371 -63368
rect 53514 -63434 53626 -63428
rect 53514 -63438 53526 -63434
rect 53510 -63468 53526 -63438
rect 53614 -63438 53626 -63434
rect 53614 -63468 53630 -63438
rect 53510 -63528 53630 -63468
rect 53940 -63488 53950 -63408
rect 54010 -63438 54020 -63408
rect 54069 -63388 54869 -63382
rect 54069 -63422 54081 -63388
rect 54857 -63422 54869 -63388
rect 54069 -63428 54869 -63422
rect 54910 -63398 54980 -63388
rect 54010 -63450 54028 -63438
rect 54022 -63488 54028 -63450
rect 53940 -63500 54028 -63488
rect 53940 -63508 54020 -63500
rect 54910 -63508 54980 -63498
rect 55311 -63408 55324 -63374
rect 55358 -63408 55371 -63374
rect 54070 -63510 54870 -63508
rect 54069 -63516 54870 -63510
rect 54069 -63538 54081 -63516
rect 54041 -63550 54081 -63538
rect 54857 -63518 54870 -63516
rect 54857 -63550 54880 -63518
rect 55311 -63548 55371 -63408
rect 54041 -63558 54880 -63550
rect 55240 -63558 55371 -63548
rect 54041 -63568 55240 -63558
rect 53510 -63658 53630 -63648
rect 53961 -63608 55240 -63568
rect 53961 -63806 54031 -63608
rect 54730 -63668 54860 -63658
rect 54730 -63688 54740 -63668
rect 54080 -63738 54740 -63688
rect 54069 -63744 54740 -63738
rect 54850 -63738 54860 -63668
rect 54850 -63744 54869 -63738
rect 54069 -63778 54081 -63744
rect 54857 -63778 54869 -63744
rect 54069 -63784 54869 -63778
rect 54911 -63794 54981 -63608
rect 55370 -63608 55371 -63558
rect 55240 -63628 55370 -63618
rect 55410 -63648 55510 -63338
rect 55410 -63758 55510 -63738
rect 55570 -63668 55680 -63048
rect 55780 -63430 55820 -62678
rect 55854 -63430 55860 -62654
rect 55780 -63438 55860 -63430
rect 55814 -63442 55860 -63438
rect 55992 -62654 56300 -62642
rect 55992 -63430 55998 -62654
rect 56032 -63428 56300 -62654
rect 56410 -62698 56430 -62099
rect 56380 -62875 56430 -62698
rect 56464 -62875 56470 -62099
rect 56380 -62887 56470 -62875
rect 56552 -62099 56750 -62087
rect 56552 -62875 56558 -62099
rect 56592 -62238 56750 -62099
rect 57066 -62080 57098 -62050
rect 57368 -62050 57372 -61964
rect 58896 -61959 59076 -61950
rect 58896 -61960 59084 -61959
rect 59156 -61960 59202 -61959
rect 57368 -62080 57396 -62050
rect 57066 -62210 57086 -62080
rect 57376 -62210 57396 -62080
rect 56592 -62875 56610 -62238
rect 57066 -62240 57396 -62210
rect 56860 -62390 57060 -62378
rect 56860 -62418 57236 -62390
rect 56860 -62548 56900 -62418
rect 57020 -62548 57236 -62418
rect 56860 -62588 57236 -62548
rect 57036 -62590 57236 -62588
rect 58556 -62480 58756 -62460
rect 58556 -62640 58576 -62480
rect 58736 -62640 58756 -62480
rect 58556 -62660 58756 -62640
rect 56552 -62878 56610 -62875
rect 57036 -62740 57446 -62730
rect 56552 -62887 56598 -62878
rect 57036 -62880 57056 -62740
rect 57416 -62880 57446 -62740
rect 56380 -63158 56440 -62887
rect 57036 -62900 57098 -62880
rect 56480 -62928 56550 -62918
rect 56480 -62998 56550 -62988
rect 57096 -63014 57098 -62934
rect 57368 -62900 57446 -62880
rect 57368 -63014 57372 -62934
rect 57096 -63030 57372 -63014
rect 58896 -63090 58926 -61960
rect 58966 -61971 59086 -61960
rect 58966 -62347 59044 -61971
rect 59078 -62347 59086 -61971
rect 58966 -62370 59086 -62347
rect 59156 -61971 59256 -61960
rect 59756 -61970 59826 -61940
rect 59966 -61952 59976 -61922
rect 60316 -61922 60346 -61916
rect 61036 -61920 61466 -61910
rect 60316 -61952 60326 -61922
rect 59966 -61960 60326 -61952
rect 59156 -62347 59162 -61971
rect 59196 -62040 59256 -61971
rect 59236 -62120 59256 -62040
rect 59196 -62240 59256 -62120
rect 59236 -62320 59256 -62240
rect 59196 -62347 59256 -62320
rect 59156 -62360 59256 -62347
rect 58966 -62680 59036 -62370
rect 59066 -62406 59176 -62400
rect 59066 -62410 59103 -62406
rect 59137 -62410 59176 -62406
rect 59066 -62480 59076 -62410
rect 59166 -62480 59176 -62410
rect 59066 -62490 59176 -62480
rect 59206 -62560 59256 -62360
rect 59376 -61990 59826 -61970
rect 59376 -62030 59476 -61990
rect 59656 -62030 59826 -61990
rect 59376 -62040 59826 -62030
rect 59376 -62090 59436 -62040
rect 59376 -62450 59386 -62090
rect 59426 -62450 59436 -62090
rect 59526 -62098 59576 -62070
rect 59526 -62132 59546 -62098
rect 59636 -62130 59706 -62070
rect 59580 -62132 59706 -62130
rect 59526 -62140 59706 -62132
rect 59476 -62182 59546 -62170
rect 59476 -62250 59502 -62182
rect 59476 -62358 59502 -62320
rect 59536 -62358 59546 -62182
rect 59476 -62370 59546 -62358
rect 59576 -62182 59636 -62170
rect 59576 -62190 59590 -62182
rect 59624 -62190 59636 -62182
rect 59576 -62370 59636 -62360
rect 59534 -62408 59592 -62402
rect 59534 -62410 59546 -62408
rect 59066 -62570 59176 -62560
rect 59066 -62640 59076 -62570
rect 59166 -62640 59176 -62570
rect 59066 -62642 59103 -62640
rect 59137 -62642 59176 -62640
rect 59066 -62650 59176 -62642
rect 59206 -62570 59266 -62560
rect 59206 -62650 59266 -62640
rect 59376 -62600 59436 -62450
rect 59516 -62442 59546 -62410
rect 59580 -62410 59592 -62408
rect 59666 -62410 59706 -62140
rect 59580 -62442 59706 -62410
rect 59516 -62480 59706 -62442
rect 59746 -62098 59936 -62070
rect 59746 -62132 59862 -62098
rect 59896 -62132 59936 -62098
rect 59746 -62140 59936 -62132
rect 61036 -62100 61206 -61920
rect 61346 -62100 61466 -61920
rect 61036 -62140 61466 -62100
rect 59746 -62400 59776 -62140
rect 60286 -62150 60476 -62140
rect 59806 -62182 59866 -62170
rect 59806 -62200 59818 -62182
rect 59852 -62200 59866 -62182
rect 59806 -62358 59818 -62340
rect 59852 -62358 59866 -62340
rect 59806 -62370 59866 -62358
rect 59900 -62180 60016 -62170
rect 59900 -62182 59916 -62180
rect 59900 -62358 59906 -62182
rect 59900 -62360 59916 -62358
rect 60006 -62360 60016 -62180
rect 60286 -62290 60306 -62150
rect 60456 -62290 60476 -62150
rect 61176 -62200 61386 -62180
rect 60286 -62300 60476 -62290
rect 61026 -62220 61136 -62210
rect 59900 -62370 60016 -62360
rect 60076 -62357 60196 -62320
rect 60076 -62391 60127 -62357
rect 60161 -62391 60196 -62357
rect 59746 -62408 59926 -62400
rect 59746 -62410 59862 -62408
rect 59896 -62410 59926 -62408
rect 59746 -62480 59826 -62410
rect 59916 -62480 59926 -62410
rect 59746 -62490 59926 -62480
rect 60076 -62449 60196 -62391
rect 60336 -62360 60446 -62300
rect 60336 -62400 60366 -62360
rect 60406 -62400 60446 -62360
rect 60636 -62357 60816 -62320
rect 60636 -62391 60671 -62357
rect 60705 -62391 60747 -62357
rect 60781 -62391 60816 -62357
rect 60076 -62480 60127 -62449
rect 60161 -62480 60196 -62449
rect 59736 -62570 59936 -62560
rect 58966 -62701 59086 -62680
rect 58966 -63077 59044 -62701
rect 59078 -63077 59086 -62701
rect 58966 -63090 59086 -63077
rect 59156 -62690 59202 -62689
rect 59156 -62701 59236 -62690
rect 59156 -63077 59162 -62701
rect 59196 -62730 59236 -62701
rect 59226 -62810 59236 -62730
rect 59196 -62960 59236 -62810
rect 59226 -63040 59236 -62960
rect 59196 -63077 59236 -63040
rect 59376 -62970 59386 -62600
rect 59426 -62970 59436 -62600
rect 59516 -62611 59706 -62570
rect 59516 -62645 59545 -62611
rect 59579 -62645 59706 -62611
rect 59516 -62650 59706 -62645
rect 59533 -62651 59591 -62650
rect 59466 -62695 59546 -62680
rect 59586 -62683 59646 -62680
rect 59466 -62730 59501 -62695
rect 59466 -62871 59501 -62810
rect 59535 -62871 59546 -62695
rect 59466 -62880 59546 -62871
rect 59583 -62695 59646 -62683
rect 59583 -62710 59589 -62695
rect 59623 -62710 59646 -62695
rect 59583 -62850 59586 -62710
rect 59583 -62871 59589 -62850
rect 59623 -62871 59646 -62850
rect 59583 -62880 59646 -62871
rect 59495 -62883 59541 -62880
rect 59583 -62883 59629 -62880
rect 59533 -62920 59591 -62915
rect 59676 -62920 59706 -62650
rect 59376 -63010 59436 -62970
rect 59506 -62980 59516 -62920
rect 59596 -62980 59706 -62920
rect 59736 -62640 59826 -62570
rect 59926 -62640 59936 -62570
rect 59736 -62645 59861 -62640
rect 59895 -62645 59936 -62640
rect 59736 -62650 59936 -62645
rect 60076 -62640 60096 -62480
rect 60176 -62640 60196 -62480
rect 59736 -62920 59766 -62650
rect 59849 -62651 59907 -62650
rect 60076 -62667 60127 -62640
rect 60161 -62667 60196 -62640
rect 59796 -62683 59856 -62680
rect 59796 -62690 59857 -62683
rect 59856 -62870 59857 -62690
rect 59796 -62871 59817 -62870
rect 59851 -62871 59857 -62870
rect 59796 -62880 59857 -62871
rect 59811 -62883 59857 -62880
rect 59899 -62690 59945 -62683
rect 59899 -62695 59916 -62690
rect 59899 -62871 59905 -62695
rect 59899 -62880 59916 -62871
rect 60006 -62880 60016 -62690
rect 60076 -62725 60196 -62667
rect 60346 -62450 60426 -62400
rect 60346 -62490 60366 -62450
rect 60406 -62490 60426 -62450
rect 60346 -62540 60426 -62490
rect 60346 -62580 60366 -62540
rect 60406 -62580 60426 -62540
rect 60346 -62620 60426 -62580
rect 60346 -62660 60366 -62620
rect 60406 -62660 60426 -62620
rect 60346 -62670 60426 -62660
rect 60636 -62449 60816 -62391
rect 60636 -62483 60671 -62449
rect 60705 -62483 60747 -62449
rect 60781 -62483 60816 -62449
rect 60636 -62541 60816 -62483
rect 60636 -62575 60671 -62541
rect 60705 -62575 60747 -62541
rect 60781 -62575 60816 -62541
rect 60636 -62633 60816 -62575
rect 60636 -62667 60671 -62633
rect 60705 -62667 60747 -62633
rect 60781 -62667 60816 -62633
rect 60076 -62759 60127 -62725
rect 60161 -62759 60196 -62725
rect 60076 -62790 60196 -62759
rect 60276 -62710 60546 -62700
rect 60276 -62725 60476 -62710
rect 60276 -62759 60297 -62725
rect 60331 -62759 60369 -62725
rect 60405 -62759 60449 -62725
rect 60276 -62770 60476 -62759
rect 60536 -62770 60546 -62710
rect 60276 -62780 60546 -62770
rect 60636 -62725 60816 -62667
rect 61026 -62330 61036 -62220
rect 61126 -62330 61136 -62220
rect 61176 -62280 61196 -62200
rect 61366 -62280 61386 -62200
rect 61176 -62300 61386 -62280
rect 61026 -62360 61136 -62330
rect 61026 -62400 61046 -62360
rect 61086 -62400 61136 -62360
rect 61026 -62450 61136 -62400
rect 61026 -62490 61046 -62450
rect 61086 -62490 61136 -62450
rect 61026 -62540 61136 -62490
rect 61026 -62580 61046 -62540
rect 61086 -62580 61136 -62540
rect 61026 -62620 61136 -62580
rect 61026 -62660 61046 -62620
rect 61086 -62660 61136 -62620
rect 61026 -62680 61136 -62660
rect 61256 -62357 61366 -62300
rect 61256 -62391 61291 -62357
rect 61325 -62391 61366 -62357
rect 61256 -62449 61366 -62391
rect 61256 -62450 61291 -62449
rect 61325 -62450 61366 -62449
rect 61256 -62660 61276 -62450
rect 61356 -62660 61366 -62450
rect 61256 -62667 61291 -62660
rect 61325 -62667 61366 -62660
rect 60636 -62759 60671 -62725
rect 60705 -62759 60747 -62725
rect 60781 -62759 60816 -62725
rect 60636 -62840 60816 -62759
rect 60966 -62724 61177 -62710
rect 60966 -62725 61129 -62724
rect 60966 -62759 60980 -62725
rect 61015 -62759 61053 -62725
rect 61088 -62758 61129 -62725
rect 61164 -62758 61177 -62724
rect 61088 -62759 61177 -62758
rect 60966 -62790 61177 -62759
rect 61256 -62725 61366 -62667
rect 61256 -62759 61291 -62725
rect 61325 -62759 61366 -62725
rect 61256 -62790 61366 -62759
rect 60466 -62850 60546 -62840
rect 59899 -62883 59945 -62880
rect 60466 -62910 60476 -62850
rect 60536 -62910 60546 -62850
rect 59849 -62920 59907 -62915
rect 60466 -62920 60546 -62910
rect 60606 -62850 60826 -62840
rect 60606 -62910 60616 -62850
rect 60736 -62910 60756 -62850
rect 60816 -62910 60826 -62850
rect 60606 -62920 60826 -62910
rect 60886 -62850 60966 -62840
rect 60886 -62910 60896 -62850
rect 60956 -62910 60966 -62850
rect 60886 -62920 60966 -62910
rect 59736 -62921 59926 -62920
rect 59736 -62955 59861 -62921
rect 59895 -62955 59926 -62921
rect 59736 -62980 59926 -62955
rect 60636 -62970 60816 -62920
rect 59376 -63020 59826 -63010
rect 59376 -63060 59476 -63020
rect 59646 -63060 59826 -63020
rect 59376 -63070 59826 -63060
rect 59156 -63090 59236 -63077
rect 58896 -63100 59086 -63090
rect 56380 -63168 57000 -63158
rect 57356 -63164 57676 -63150
rect 56440 -63174 57000 -63168
rect 57314 -63170 57676 -63164
rect 56440 -63194 57178 -63174
rect 56440 -63244 57118 -63194
rect 57168 -63244 57178 -63194
rect 57314 -63210 57326 -63170
rect 57376 -63210 57676 -63170
rect 57314 -63216 57676 -63210
rect 57356 -63230 57676 -63216
rect 56440 -63254 57178 -63244
rect 56440 -63288 57000 -63254
rect 57112 -63256 57174 -63254
rect 56380 -63358 57000 -63288
rect 56032 -63430 56038 -63428
rect 55992 -63442 56038 -63430
rect 55880 -63474 55970 -63468
rect 55870 -63478 55982 -63474
rect 55870 -63520 55880 -63478
rect 55970 -63520 55982 -63478
rect 55880 -63568 55970 -63558
rect 56120 -63598 56300 -63428
rect 57096 -63509 57372 -63478
rect 57096 -63543 57125 -63509
rect 57159 -63543 57217 -63509
rect 57251 -63543 57309 -63509
rect 57343 -63520 57372 -63509
rect 57343 -63543 57376 -63520
rect 57096 -63580 57376 -63543
rect 57066 -63590 57376 -63580
rect 56426 -63598 57376 -63590
rect 56120 -63608 57376 -63598
rect 56014 -63658 56086 -63646
rect 55570 -63778 55830 -63668
rect 53961 -63844 53988 -63806
rect 54022 -63844 54031 -63806
rect 53961 -63858 54031 -63844
rect 54910 -63806 54981 -63794
rect 54910 -63844 54916 -63806
rect 54950 -63844 54981 -63806
rect 54910 -63856 54981 -63844
rect 54911 -63858 54981 -63856
rect 55220 -63818 55330 -63808
rect 54069 -63872 54869 -63866
rect 54069 -63906 54081 -63872
rect 54857 -63878 54869 -63872
rect 54857 -63906 54880 -63878
rect 54069 -63912 54880 -63906
rect 54090 -63988 54880 -63912
rect 55330 -63918 55380 -63818
rect 55330 -63928 55480 -63918
rect 55220 -63938 55480 -63928
rect 55280 -63952 55480 -63938
rect 55280 -63958 55488 -63952
rect 55280 -63978 55300 -63958
rect 54090 -64088 54150 -63988
rect 54840 -64088 54880 -63988
rect 55288 -63992 55300 -63978
rect 55476 -63992 55488 -63958
rect 55530 -63978 55610 -63968
rect 55288 -63998 55488 -63992
rect 55520 -64002 55530 -63990
rect 55520 -64036 55526 -64002
rect 55288 -64046 55488 -64040
rect 55288 -64080 55300 -64046
rect 55476 -64080 55488 -64046
rect 55520 -64048 55530 -64036
rect 55530 -64078 55610 -64068
rect 55288 -64086 55488 -64080
rect 54090 -64108 54140 -64088
rect 54100 -64348 54140 -64108
rect 54850 -64348 54880 -64088
rect 55300 -64128 55470 -64086
rect 55300 -64268 55320 -64128
rect 55470 -64214 55482 -64142
rect 55300 -64278 55470 -64268
rect 54100 -64388 54880 -64348
rect 55710 -64598 55830 -63778
rect 56014 -63808 56020 -63658
rect 56080 -63808 56086 -63658
rect 56014 -63820 56086 -63808
rect 56120 -63808 56170 -63608
rect 56390 -63660 57376 -63608
rect 56390 -63668 57156 -63660
rect 56390 -63808 56654 -63668
rect 56120 -63858 56654 -63808
rect 56306 -63886 56654 -63858
rect 56998 -63820 57156 -63668
rect 57316 -63820 57376 -63660
rect 56998 -63886 57376 -63820
rect 56306 -64300 57376 -63886
rect 57556 -64010 57676 -63230
rect 58896 -63260 58986 -63100
rect 59756 -63120 59826 -63070
rect 59066 -63136 59176 -63130
rect 59066 -63140 59103 -63136
rect 59137 -63140 59176 -63136
rect 59066 -63200 59076 -63140
rect 59166 -63200 59176 -63140
rect 59066 -63210 59176 -63200
rect 58896 -63630 58926 -63260
rect 58966 -63630 58986 -63330
rect 59116 -63260 59506 -63240
rect 59116 -63330 59146 -63260
rect 59226 -63330 59276 -63260
rect 59356 -63330 59396 -63260
rect 59476 -63330 59506 -63260
rect 59116 -63348 59506 -63330
rect 59646 -63260 59716 -63240
rect 59706 -63320 59716 -63260
rect 59646 -63330 59716 -63320
rect 59113 -63354 59513 -63348
rect 59113 -63388 59125 -63354
rect 59501 -63388 59513 -63354
rect 59113 -63394 59513 -63388
rect 59546 -63400 59616 -63390
rect 59246 -63456 59256 -63430
rect 59113 -63462 59256 -63456
rect 59366 -63456 59376 -63430
rect 59366 -63462 59513 -63456
rect 59016 -63500 59076 -63480
rect 59113 -63496 59125 -63462
rect 59501 -63496 59513 -63462
rect 59606 -63460 59616 -63400
rect 59546 -63470 59616 -63460
rect 59113 -63502 59513 -63496
rect 59016 -63590 59076 -63560
rect 59113 -63570 59513 -63564
rect 59113 -63604 59125 -63570
rect 59501 -63604 59513 -63570
rect 59113 -63610 59513 -63604
rect 58896 -63700 58906 -63630
rect 58896 -63720 58986 -63700
rect 59116 -63630 59516 -63610
rect 59116 -63700 59146 -63630
rect 59226 -63700 59276 -63630
rect 59356 -63700 59396 -63630
rect 59476 -63700 59516 -63630
rect 59116 -63720 59516 -63700
rect 59646 -63630 59656 -63330
rect 59706 -63630 59716 -63330
rect 59756 -63300 59766 -63120
rect 59806 -63300 59826 -63120
rect 59956 -63120 60336 -63110
rect 59956 -63134 59966 -63120
rect 59946 -63140 59966 -63134
rect 60326 -63134 60336 -63120
rect 60326 -63140 60346 -63134
rect 59856 -63180 59916 -63170
rect 59946 -63174 59958 -63140
rect 60334 -63174 60346 -63140
rect 61056 -63140 61176 -62790
rect 59946 -63180 59966 -63174
rect 60326 -63180 60346 -63174
rect 60376 -63180 60436 -63160
rect 59956 -63190 60336 -63180
rect 59856 -63260 59916 -63240
rect 59946 -63248 60346 -63242
rect 59756 -63340 59826 -63300
rect 59946 -63282 59958 -63248
rect 60334 -63282 60346 -63248
rect 60376 -63260 60436 -63240
rect 61126 -63240 61176 -63140
rect 61056 -63270 61176 -63240
rect 59946 -63288 60346 -63282
rect 59946 -63340 60336 -63288
rect 59756 -63360 60536 -63340
rect 59756 -63400 59866 -63360
rect 60426 -63400 60536 -63360
rect 59756 -63410 60536 -63400
rect 59796 -63520 59806 -63410
rect 59916 -63520 59926 -63410
rect 59796 -63530 59926 -63520
rect 60436 -63430 60536 -63410
rect 60436 -63550 60446 -63430
rect 60526 -63550 60536 -63430
rect 60436 -63560 60536 -63550
rect 59646 -63640 59716 -63630
rect 59706 -63700 59716 -63640
rect 59646 -63720 59716 -63700
rect 58806 -64010 59356 -63980
rect 57556 -64020 59356 -64010
rect 57556 -64160 58986 -64020
rect 59126 -64160 59356 -64020
rect 59846 -63990 60256 -63980
rect 59846 -64100 59996 -63990
rect 60106 -64100 60256 -63990
rect 57556 -64210 59356 -64160
rect 58806 -64290 59356 -64210
rect 55710 -64600 55910 -64598
rect 24400 -65400 36000 -64800
rect 55400 -64700 56200 -64600
rect 59600 -64700 60500 -64100
rect 55400 -65100 55500 -64700
rect 56100 -65100 56200 -64700
rect 55400 -65200 56200 -65100
rect 55360 -65680 55800 -65600
rect 55360 -65960 55440 -65680
rect 55720 -65960 55800 -65680
rect 55360 -66040 55800 -65960
rect 54090 -66138 54890 -66098
rect 54090 -66268 54150 -66138
rect 53510 -66320 53800 -66318
rect 53460 -66340 53800 -66320
rect 53460 -66540 53480 -66340
rect 53780 -66540 53800 -66340
rect 54080 -66398 54150 -66268
rect 54860 -66378 54890 -66138
rect 54850 -66398 54890 -66378
rect 54080 -66466 54880 -66398
rect 54079 -66472 54880 -66466
rect 54079 -66506 54091 -66472
rect 54867 -66498 54880 -66472
rect 54867 -66506 54879 -66498
rect 54079 -66512 54879 -66506
rect 53460 -66560 53800 -66540
rect 53510 -66658 53800 -66560
rect 53002 -66820 53480 -66758
rect 53000 -66958 53480 -66820
rect 53510 -66768 53520 -66658
rect 53640 -66768 53800 -66658
rect 53510 -66888 53800 -66768
rect 53970 -66534 54040 -66518
rect 53970 -66572 53998 -66534
rect 54032 -66572 54040 -66534
rect 53970 -66768 54040 -66572
rect 54920 -66534 54990 -66518
rect 54920 -66572 54926 -66534
rect 54960 -66572 54990 -66534
rect 54079 -66600 54879 -66594
rect 54079 -66634 54091 -66600
rect 54867 -66634 54879 -66600
rect 54079 -66638 54879 -66634
rect 54079 -66640 54750 -66638
rect 54090 -66688 54750 -66640
rect 54740 -66718 54750 -66688
rect 54850 -66640 54879 -66638
rect 54850 -66708 54860 -66640
rect 54840 -66718 54860 -66708
rect 54750 -66728 54860 -66718
rect 54920 -66768 54990 -66572
rect 55430 -66618 55520 -66608
rect 55290 -66728 55390 -66718
rect 53970 -66798 55290 -66768
rect 55430 -66758 55520 -66688
rect 53970 -66808 55390 -66798
rect 54050 -66818 55380 -66808
rect 54050 -66828 54880 -66818
rect 54050 -66838 54091 -66828
rect 54079 -66862 54091 -66838
rect 54867 -66838 54880 -66828
rect 54867 -66862 54879 -66838
rect 54079 -66868 54879 -66862
rect 54920 -66878 54990 -66868
rect 53510 -66906 53630 -66888
rect 53510 -66938 53526 -66906
rect 53514 -66940 53526 -66938
rect 53614 -66938 53630 -66906
rect 53940 -66890 54038 -66878
rect 53940 -66898 53998 -66890
rect 53614 -66940 53626 -66938
rect 53514 -66946 53626 -66940
rect 53000 -68708 53050 -66958
rect 53250 -66968 53480 -66958
rect 53250 -68318 53330 -66968
rect 53400 -66978 53480 -66968
rect 53400 -66990 53504 -66978
rect 53400 -67766 53464 -66990
rect 53498 -67766 53504 -66990
rect 53400 -67778 53504 -67766
rect 53636 -66988 53682 -66978
rect 53636 -66990 53760 -66988
rect 53636 -67766 53642 -66990
rect 53676 -67766 53760 -66990
rect 53940 -66998 53950 -66898
rect 54032 -66928 54038 -66890
rect 54020 -66940 54038 -66928
rect 54020 -66998 54030 -66940
rect 54079 -66956 54879 -66950
rect 54079 -66990 54091 -66956
rect 54867 -66990 54879 -66956
rect 54920 -66978 54990 -66968
rect 55320 -66968 55380 -66818
rect 54079 -66996 54879 -66990
rect 53940 -67018 54030 -66998
rect 54090 -67028 54870 -66996
rect 55320 -67002 55334 -66968
rect 55368 -67002 55380 -66968
rect 55320 -67008 55380 -67002
rect 53840 -67328 53920 -67318
rect 53840 -67438 53860 -67328
rect 53840 -67448 53920 -67438
rect 53840 -67640 53900 -67448
rect 54320 -67528 54510 -67028
rect 55440 -67038 55520 -66758
rect 55410 -67040 55520 -67038
rect 55284 -67048 55330 -67040
rect 55230 -67052 55330 -67048
rect 55230 -67058 55290 -67052
rect 55324 -67228 55330 -67052
rect 55230 -67238 55330 -67228
rect 55284 -67240 55330 -67238
rect 55372 -67048 55520 -67040
rect 55372 -67052 55430 -67048
rect 55372 -67228 55378 -67052
rect 55412 -67218 55430 -67052
rect 55510 -67218 55520 -67048
rect 55412 -67228 55520 -67218
rect 55372 -67240 55418 -67228
rect 55580 -67328 55720 -66040
rect 58776 -66270 59306 -66150
rect 58776 -66280 58966 -66270
rect 56146 -66380 57366 -66330
rect 55954 -66528 56046 -66516
rect 56146 -66528 56506 -66380
rect 55954 -66698 55960 -66528
rect 56040 -66698 56046 -66528
rect 55954 -66710 56046 -66698
rect 56120 -66558 56506 -66528
rect 56120 -66768 56190 -66558
rect 56390 -66630 56506 -66558
rect 57016 -66534 57366 -66380
rect 57586 -66430 58966 -66280
rect 59126 -66430 59306 -66270
rect 57586 -66450 59306 -66430
rect 59946 -66300 60386 -66200
rect 57586 -66480 58986 -66450
rect 59946 -66460 59956 -66300
rect 60166 -66460 60386 -66300
rect 57016 -66630 57368 -66534
rect 56390 -66670 57368 -66630
rect 56390 -66768 57126 -66670
rect 56120 -66774 57126 -66768
rect 56120 -66778 56750 -66774
rect 55880 -66818 55970 -66808
rect 55870 -66896 55880 -66850
rect 55970 -66896 55982 -66850
rect 55880 -66908 55970 -66898
rect 55000 -67338 55090 -67328
rect 55000 -67448 55090 -67438
rect 54710 -67528 54960 -67508
rect 53940 -67568 54960 -67528
rect 53940 -67572 54730 -67568
rect 53930 -67578 54730 -67572
rect 53930 -67612 53942 -67578
rect 54718 -67612 54730 -67578
rect 53930 -67618 54730 -67612
rect 53840 -67728 53858 -67640
rect 53892 -67728 53900 -67640
rect 53840 -67748 53900 -67728
rect 54762 -67638 54850 -67628
rect 54762 -67640 54770 -67638
rect 54762 -67728 54768 -67640
rect 54840 -67728 54850 -67638
rect 54762 -67740 54850 -67728
rect 54770 -67748 54850 -67740
rect 53636 -67778 53760 -67766
rect 53400 -67996 53480 -67778
rect 53514 -67816 53626 -67810
rect 53514 -67818 53526 -67816
rect 53510 -67850 53526 -67818
rect 53614 -67818 53626 -67816
rect 53614 -67850 53630 -67818
rect 53510 -67924 53630 -67850
rect 53510 -67958 53526 -67924
rect 53614 -67958 53630 -67924
rect 53680 -67838 53760 -67778
rect 53930 -67756 54730 -67750
rect 53930 -67790 53942 -67756
rect 54718 -67790 54730 -67756
rect 53930 -67796 54730 -67790
rect 53940 -67828 54720 -67796
rect 53920 -67838 54720 -67828
rect 53680 -67928 54720 -67838
rect 53514 -67964 53626 -67958
rect 53680 -67996 53760 -67928
rect 53920 -67938 54720 -67928
rect 53940 -67978 54720 -67938
rect 54900 -67968 54960 -67568
rect 55010 -67560 55090 -67448
rect 55540 -67338 55720 -67328
rect 55630 -67438 55720 -67338
rect 55130 -67474 55506 -67468
rect 55130 -67508 55142 -67474
rect 55494 -67508 55506 -67474
rect 55130 -67514 55506 -67508
rect 55010 -67594 55046 -67560
rect 55080 -67594 55090 -67560
rect 55010 -67608 55090 -67594
rect 55142 -67640 55494 -67514
rect 55540 -67560 55720 -67438
rect 55540 -67594 55556 -67560
rect 55590 -67594 55720 -67560
rect 55540 -67608 55720 -67594
rect 55780 -66940 55860 -66928
rect 55130 -67646 55506 -67640
rect 55130 -67680 55142 -67646
rect 55494 -67678 55506 -67646
rect 55494 -67680 55510 -67678
rect 55130 -67686 55510 -67680
rect 55140 -67698 55510 -67686
rect 55780 -67698 55820 -66940
rect 55140 -67716 55820 -67698
rect 55854 -67716 55860 -66940
rect 55140 -67728 55860 -67716
rect 55992 -66940 56038 -66928
rect 55992 -67716 55998 -66940
rect 56032 -66948 56038 -66940
rect 56120 -66948 56300 -66778
rect 57098 -66800 57126 -66774
rect 57356 -66800 57368 -66670
rect 57098 -66814 57368 -66800
rect 57096 -66845 57372 -66814
rect 57096 -66879 57125 -66845
rect 57159 -66879 57217 -66845
rect 57251 -66879 57309 -66845
rect 57343 -66879 57372 -66845
rect 57096 -66910 57372 -66879
rect 56032 -67306 56300 -66948
rect 56590 -67068 56660 -67058
rect 56660 -67134 57000 -67068
rect 57586 -67130 57706 -66480
rect 59946 -66490 60386 -66460
rect 57366 -67134 57706 -67130
rect 56660 -67138 57188 -67134
rect 56660 -67144 57190 -67138
rect 56660 -67194 57118 -67144
rect 57178 -67194 57190 -67144
rect 57314 -67140 57706 -67134
rect 57314 -67180 57326 -67140
rect 57366 -67180 57706 -67140
rect 57314 -67186 57706 -67180
rect 57366 -67190 57706 -67186
rect 58896 -66770 58986 -66750
rect 58896 -66830 58906 -66770
rect 58896 -67120 58926 -66830
rect 58966 -67120 58986 -66770
rect 59106 -66770 59516 -66760
rect 59106 -66830 59216 -66770
rect 59276 -66830 59326 -66770
rect 59386 -66830 59436 -66770
rect 59496 -66830 59516 -66770
rect 59106 -66847 59516 -66830
rect 59626 -66770 59706 -66730
rect 59626 -66830 59636 -66770
rect 59626 -66840 59656 -66830
rect 59106 -66880 59125 -66847
rect 59113 -66881 59125 -66880
rect 59501 -66880 59516 -66847
rect 59501 -66881 59513 -66880
rect 59113 -66887 59513 -66881
rect 59546 -66890 59616 -66880
rect 59276 -66930 59356 -66920
rect 59276 -66949 59286 -66930
rect 59113 -66955 59286 -66949
rect 59346 -66949 59356 -66930
rect 59346 -66955 59513 -66949
rect 59113 -66989 59125 -66955
rect 59501 -66989 59513 -66955
rect 59606 -66950 59616 -66890
rect 59546 -66960 59616 -66950
rect 59113 -66990 59286 -66989
rect 59346 -66990 59513 -66989
rect 59016 -67000 59076 -66990
rect 59113 -66995 59513 -66990
rect 59276 -67000 59356 -66995
rect 59546 -67010 59616 -67000
rect 59016 -67070 59076 -67060
rect 59113 -67063 59513 -67057
rect 59113 -67097 59125 -67063
rect 59501 -67097 59513 -67063
rect 59606 -67070 59616 -67010
rect 59546 -67080 59616 -67070
rect 59113 -67100 59513 -67097
rect 59113 -67103 59516 -67100
rect 58896 -67130 58986 -67120
rect 58896 -67190 58906 -67130
rect 58966 -67190 58986 -67130
rect 58896 -67192 58986 -67190
rect 59116 -67120 59516 -67103
rect 59646 -67110 59656 -66840
rect 59116 -67180 59216 -67120
rect 59276 -67180 59336 -67120
rect 59396 -67180 59436 -67120
rect 59496 -67180 59516 -67120
rect 56660 -67198 57190 -67194
rect 56590 -67200 57190 -67198
rect 56590 -67204 57188 -67200
rect 56590 -67268 57000 -67204
rect 56032 -67318 56356 -67306
rect 56032 -67716 56280 -67318
rect 55992 -67728 56280 -67716
rect 55140 -67738 55200 -67728
rect 55450 -67758 55810 -67728
rect 55870 -67766 55982 -67760
rect 55870 -67800 55882 -67766
rect 55970 -67800 55982 -67766
rect 55870 -67806 55982 -67800
rect 55140 -67818 55200 -67808
rect 55024 -67848 55116 -67836
rect 55024 -67928 55030 -67848
rect 55110 -67928 55116 -67848
rect 55024 -67940 55116 -67928
rect 55734 -67848 55816 -67836
rect 55734 -67928 55740 -67848
rect 55810 -67928 55816 -67848
rect 55734 -67940 55816 -67928
rect 55880 -67838 55970 -67806
rect 55880 -67964 55970 -67928
rect 56060 -67948 56280 -67728
rect 56350 -67948 56356 -67318
rect 56480 -67388 56550 -67378
rect 56480 -67458 56550 -67448
rect 56590 -67487 56750 -67268
rect 58894 -67286 58988 -67192
rect 59116 -67200 59516 -67180
rect 59636 -67120 59656 -67110
rect 59696 -67120 59706 -66770
rect 59856 -66940 59976 -66930
rect 59856 -67030 59866 -66940
rect 59966 -67030 59976 -66940
rect 59856 -67040 59976 -67030
rect 60436 -67020 60446 -66920
rect 60526 -67020 60536 -66920
rect 60436 -67040 60536 -67020
rect 59636 -67130 59706 -67120
rect 59696 -67190 59706 -67130
rect 59636 -67210 59706 -67190
rect 59756 -67060 60536 -67040
rect 59756 -67100 59866 -67060
rect 60426 -67100 60536 -67060
rect 59756 -67110 60536 -67100
rect 59756 -67150 59826 -67110
rect 59066 -67240 59176 -67230
rect 58896 -67350 58986 -67286
rect 59066 -67310 59076 -67240
rect 59166 -67310 59176 -67240
rect 59066 -67312 59103 -67310
rect 59137 -67312 59176 -67310
rect 59066 -67320 59176 -67312
rect 59756 -67340 59766 -67150
rect 59806 -67340 59826 -67150
rect 59956 -67168 60046 -67140
rect 59946 -67174 60046 -67168
rect 60126 -67168 60336 -67140
rect 60126 -67174 60346 -67168
rect 59856 -67210 59916 -67200
rect 59946 -67208 59958 -67174
rect 60334 -67208 60346 -67174
rect 59946 -67214 60346 -67208
rect 60376 -67220 60446 -67210
rect 59856 -67290 59916 -67280
rect 59946 -67282 60346 -67276
rect 59946 -67316 59958 -67282
rect 60334 -67316 60346 -67282
rect 60376 -67290 60446 -67280
rect 59946 -67322 59976 -67316
rect 57098 -67358 57368 -67354
rect 57096 -67364 57372 -67358
rect 57096 -67450 57098 -67364
rect 56424 -67488 56470 -67487
rect 56060 -67960 56356 -67948
rect 56410 -67499 56470 -67488
rect 53400 -68008 53504 -67996
rect 53400 -68318 53464 -68008
rect 53250 -68708 53464 -68318
rect 53000 -68784 53464 -68708
rect 53498 -68784 53504 -68008
rect 53000 -68788 53504 -68784
rect 53458 -68796 53504 -68788
rect 53636 -68008 53760 -67996
rect 53636 -68784 53642 -68008
rect 53676 -68784 53760 -68008
rect 53930 -67984 54730 -67978
rect 53930 -68018 53942 -67984
rect 54718 -68018 54730 -67984
rect 53930 -68024 54730 -68018
rect 53830 -68046 53900 -68028
rect 53830 -68134 53858 -68046
rect 53892 -68134 53900 -68046
rect 53830 -68328 53900 -68134
rect 54760 -68046 54850 -68028
rect 54760 -68134 54768 -68046
rect 54802 -68048 54850 -68046
rect 54900 -68038 55200 -67968
rect 55870 -67970 55982 -67964
rect 55870 -68004 55882 -67970
rect 55970 -68004 55982 -67970
rect 55450 -68038 55810 -68008
rect 55870 -68010 55982 -68004
rect 56060 -68038 56300 -67960
rect 54900 -68042 55820 -68038
rect 56000 -68042 56300 -68038
rect 54900 -68048 55860 -68042
rect 54840 -68128 54850 -68048
rect 54802 -68134 54850 -68128
rect 54760 -68148 54850 -68134
rect 55130 -68054 55860 -68048
rect 55130 -68078 55820 -68054
rect 55130 -68096 55510 -68078
rect 55130 -68130 55142 -68096
rect 55494 -68098 55510 -68096
rect 55494 -68130 55506 -68098
rect 55130 -68136 55506 -68130
rect 53930 -68162 54730 -68156
rect 53930 -68196 53942 -68162
rect 54718 -68196 54730 -68162
rect 55020 -68182 55090 -68168
rect 53930 -68202 54730 -68196
rect 53940 -68208 54730 -68202
rect 54920 -68198 54980 -68188
rect 53940 -68248 54920 -68208
rect 53830 -68338 53920 -68328
rect 53830 -68448 53850 -68338
rect 53830 -68458 53920 -68448
rect 54320 -68748 54510 -68248
rect 54710 -68268 54920 -68248
rect 54910 -68278 54980 -68268
rect 55020 -68216 55046 -68182
rect 55080 -68216 55090 -68182
rect 55020 -68328 55090 -68216
rect 55142 -68262 55494 -68136
rect 55540 -68182 55620 -68168
rect 55540 -68216 55556 -68182
rect 55590 -68216 55620 -68182
rect 55130 -68268 55506 -68262
rect 55130 -68302 55142 -68268
rect 55494 -68302 55506 -68268
rect 55130 -68308 55506 -68302
rect 55000 -68338 55090 -68328
rect 55000 -68448 55090 -68438
rect 55540 -68328 55620 -68216
rect 55540 -68338 55630 -68328
rect 55630 -68438 55680 -68348
rect 55540 -68448 55680 -68438
rect 55274 -68538 55320 -68536
rect 55220 -68548 55320 -68538
rect 55220 -68724 55280 -68718
rect 55314 -68724 55320 -68548
rect 55220 -68728 55320 -68724
rect 55274 -68736 55320 -68728
rect 55362 -68548 55408 -68536
rect 55362 -68724 55368 -68548
rect 55402 -68558 55510 -68548
rect 55402 -68724 55410 -68558
rect 55362 -68728 55410 -68724
rect 55500 -68728 55510 -68558
rect 55362 -68736 55510 -68728
rect 55390 -68738 55510 -68736
rect 53636 -68788 53760 -68784
rect 53636 -68796 53682 -68788
rect 53940 -68808 54020 -68768
rect 54080 -68782 54860 -68748
rect 55311 -68774 55371 -68768
rect 53514 -68834 53626 -68828
rect 53514 -68838 53526 -68834
rect 53510 -68868 53526 -68838
rect 53614 -68838 53626 -68834
rect 53614 -68868 53630 -68838
rect 53510 -68928 53630 -68868
rect 53940 -68888 53950 -68808
rect 54010 -68838 54020 -68808
rect 54069 -68788 54869 -68782
rect 54069 -68822 54081 -68788
rect 54857 -68822 54869 -68788
rect 54069 -68828 54869 -68822
rect 54910 -68798 54980 -68788
rect 54010 -68850 54028 -68838
rect 54022 -68888 54028 -68850
rect 53940 -68900 54028 -68888
rect 53940 -68908 54020 -68900
rect 54910 -68908 54980 -68898
rect 55311 -68808 55324 -68774
rect 55358 -68808 55371 -68774
rect 54070 -68910 54870 -68908
rect 54069 -68916 54870 -68910
rect 54069 -68938 54081 -68916
rect 54041 -68950 54081 -68938
rect 54857 -68918 54870 -68916
rect 54857 -68950 54880 -68918
rect 55311 -68948 55371 -68808
rect 54041 -68958 54880 -68950
rect 55240 -68958 55371 -68948
rect 54041 -68968 55240 -68958
rect 53510 -69058 53630 -69048
rect 53961 -69008 55240 -68968
rect 53961 -69206 54031 -69008
rect 54730 -69068 54860 -69058
rect 54730 -69088 54740 -69068
rect 54080 -69138 54740 -69088
rect 54069 -69144 54740 -69138
rect 54850 -69138 54860 -69068
rect 54850 -69144 54869 -69138
rect 54069 -69178 54081 -69144
rect 54857 -69178 54869 -69144
rect 54069 -69184 54869 -69178
rect 54911 -69194 54981 -69008
rect 55370 -69008 55371 -68958
rect 55240 -69028 55370 -69018
rect 55410 -69048 55510 -68738
rect 55410 -69158 55510 -69138
rect 55570 -69068 55680 -68448
rect 55780 -68830 55820 -68078
rect 55854 -68830 55860 -68054
rect 55780 -68838 55860 -68830
rect 55814 -68842 55860 -68838
rect 55992 -68054 56300 -68042
rect 55992 -68830 55998 -68054
rect 56032 -68828 56300 -68054
rect 56410 -68098 56430 -67499
rect 56380 -68275 56430 -68098
rect 56464 -68275 56470 -67499
rect 56380 -68287 56470 -68275
rect 56552 -67499 56750 -67487
rect 56552 -68275 56558 -67499
rect 56592 -67638 56750 -67499
rect 57066 -67480 57098 -67450
rect 57368 -67450 57372 -67364
rect 58896 -67359 59076 -67350
rect 58896 -67360 59084 -67359
rect 59156 -67360 59202 -67359
rect 57368 -67480 57396 -67450
rect 57066 -67610 57086 -67480
rect 57376 -67610 57396 -67480
rect 56592 -68275 56610 -67638
rect 57066 -67640 57396 -67610
rect 56860 -67790 57060 -67778
rect 56860 -67818 57236 -67790
rect 56860 -67948 56900 -67818
rect 57020 -67948 57236 -67818
rect 56860 -67988 57236 -67948
rect 57036 -67990 57236 -67988
rect 58556 -67880 58756 -67860
rect 58556 -68040 58576 -67880
rect 58736 -68040 58756 -67880
rect 58556 -68060 58756 -68040
rect 56552 -68278 56610 -68275
rect 57036 -68140 57446 -68130
rect 56552 -68287 56598 -68278
rect 57036 -68280 57056 -68140
rect 57416 -68280 57446 -68140
rect 56380 -68558 56440 -68287
rect 57036 -68300 57098 -68280
rect 56480 -68328 56550 -68318
rect 56480 -68398 56550 -68388
rect 57096 -68414 57098 -68334
rect 57368 -68300 57446 -68280
rect 57368 -68414 57372 -68334
rect 57096 -68430 57372 -68414
rect 58896 -68490 58926 -67360
rect 58966 -67371 59086 -67360
rect 58966 -67747 59044 -67371
rect 59078 -67747 59086 -67371
rect 58966 -67770 59086 -67747
rect 59156 -67371 59256 -67360
rect 59756 -67370 59826 -67340
rect 59966 -67352 59976 -67322
rect 60316 -67322 60346 -67316
rect 61036 -67320 61466 -67310
rect 60316 -67352 60326 -67322
rect 59966 -67360 60326 -67352
rect 59156 -67747 59162 -67371
rect 59196 -67440 59256 -67371
rect 59236 -67520 59256 -67440
rect 59196 -67640 59256 -67520
rect 59236 -67720 59256 -67640
rect 59196 -67747 59256 -67720
rect 59156 -67760 59256 -67747
rect 58966 -68080 59036 -67770
rect 59066 -67806 59176 -67800
rect 59066 -67810 59103 -67806
rect 59137 -67810 59176 -67806
rect 59066 -67880 59076 -67810
rect 59166 -67880 59176 -67810
rect 59066 -67890 59176 -67880
rect 59206 -67960 59256 -67760
rect 59376 -67390 59826 -67370
rect 59376 -67430 59476 -67390
rect 59656 -67430 59826 -67390
rect 59376 -67440 59826 -67430
rect 59376 -67490 59436 -67440
rect 59376 -67850 59386 -67490
rect 59426 -67850 59436 -67490
rect 59526 -67498 59576 -67470
rect 59526 -67532 59546 -67498
rect 59636 -67530 59706 -67470
rect 59580 -67532 59706 -67530
rect 59526 -67540 59706 -67532
rect 59476 -67582 59546 -67570
rect 59476 -67650 59502 -67582
rect 59476 -67758 59502 -67720
rect 59536 -67758 59546 -67582
rect 59476 -67770 59546 -67758
rect 59576 -67582 59636 -67570
rect 59576 -67590 59590 -67582
rect 59624 -67590 59636 -67582
rect 59576 -67770 59636 -67760
rect 59534 -67808 59592 -67802
rect 59534 -67810 59546 -67808
rect 59066 -67970 59176 -67960
rect 59066 -68040 59076 -67970
rect 59166 -68040 59176 -67970
rect 59066 -68042 59103 -68040
rect 59137 -68042 59176 -68040
rect 59066 -68050 59176 -68042
rect 59206 -67970 59266 -67960
rect 59206 -68050 59266 -68040
rect 59376 -68000 59436 -67850
rect 59516 -67842 59546 -67810
rect 59580 -67810 59592 -67808
rect 59666 -67810 59706 -67540
rect 59580 -67842 59706 -67810
rect 59516 -67880 59706 -67842
rect 59746 -67498 59936 -67470
rect 59746 -67532 59862 -67498
rect 59896 -67532 59936 -67498
rect 59746 -67540 59936 -67532
rect 61036 -67500 61206 -67320
rect 61346 -67500 61466 -67320
rect 61036 -67540 61466 -67500
rect 59746 -67800 59776 -67540
rect 60286 -67550 60476 -67540
rect 59806 -67582 59866 -67570
rect 59806 -67600 59818 -67582
rect 59852 -67600 59866 -67582
rect 59806 -67758 59818 -67740
rect 59852 -67758 59866 -67740
rect 59806 -67770 59866 -67758
rect 59900 -67580 60016 -67570
rect 59900 -67582 59916 -67580
rect 59900 -67758 59906 -67582
rect 59900 -67760 59916 -67758
rect 60006 -67760 60016 -67580
rect 60286 -67690 60306 -67550
rect 60456 -67690 60476 -67550
rect 61176 -67600 61386 -67580
rect 60286 -67700 60476 -67690
rect 61026 -67620 61136 -67610
rect 59900 -67770 60016 -67760
rect 60076 -67757 60196 -67720
rect 60076 -67791 60127 -67757
rect 60161 -67791 60196 -67757
rect 59746 -67808 59926 -67800
rect 59746 -67810 59862 -67808
rect 59896 -67810 59926 -67808
rect 59746 -67880 59826 -67810
rect 59916 -67880 59926 -67810
rect 59746 -67890 59926 -67880
rect 60076 -67849 60196 -67791
rect 60336 -67760 60446 -67700
rect 60336 -67800 60366 -67760
rect 60406 -67800 60446 -67760
rect 60636 -67757 60816 -67720
rect 60636 -67791 60671 -67757
rect 60705 -67791 60747 -67757
rect 60781 -67791 60816 -67757
rect 60076 -67880 60127 -67849
rect 60161 -67880 60196 -67849
rect 59736 -67970 59936 -67960
rect 58966 -68101 59086 -68080
rect 58966 -68477 59044 -68101
rect 59078 -68477 59086 -68101
rect 58966 -68490 59086 -68477
rect 59156 -68090 59202 -68089
rect 59156 -68101 59236 -68090
rect 59156 -68477 59162 -68101
rect 59196 -68130 59236 -68101
rect 59226 -68210 59236 -68130
rect 59196 -68360 59236 -68210
rect 59226 -68440 59236 -68360
rect 59196 -68477 59236 -68440
rect 59376 -68370 59386 -68000
rect 59426 -68370 59436 -68000
rect 59516 -68011 59706 -67970
rect 59516 -68045 59545 -68011
rect 59579 -68045 59706 -68011
rect 59516 -68050 59706 -68045
rect 59533 -68051 59591 -68050
rect 59466 -68095 59546 -68080
rect 59586 -68083 59646 -68080
rect 59466 -68130 59501 -68095
rect 59466 -68271 59501 -68210
rect 59535 -68271 59546 -68095
rect 59466 -68280 59546 -68271
rect 59583 -68095 59646 -68083
rect 59583 -68110 59589 -68095
rect 59623 -68110 59646 -68095
rect 59583 -68250 59586 -68110
rect 59583 -68271 59589 -68250
rect 59623 -68271 59646 -68250
rect 59583 -68280 59646 -68271
rect 59495 -68283 59541 -68280
rect 59583 -68283 59629 -68280
rect 59533 -68320 59591 -68315
rect 59676 -68320 59706 -68050
rect 59376 -68410 59436 -68370
rect 59506 -68380 59516 -68320
rect 59596 -68380 59706 -68320
rect 59736 -68040 59826 -67970
rect 59926 -68040 59936 -67970
rect 59736 -68045 59861 -68040
rect 59895 -68045 59936 -68040
rect 59736 -68050 59936 -68045
rect 60076 -68040 60096 -67880
rect 60176 -68040 60196 -67880
rect 59736 -68320 59766 -68050
rect 59849 -68051 59907 -68050
rect 60076 -68067 60127 -68040
rect 60161 -68067 60196 -68040
rect 59796 -68083 59856 -68080
rect 59796 -68090 59857 -68083
rect 59856 -68270 59857 -68090
rect 59796 -68271 59817 -68270
rect 59851 -68271 59857 -68270
rect 59796 -68280 59857 -68271
rect 59811 -68283 59857 -68280
rect 59899 -68090 59945 -68083
rect 59899 -68095 59916 -68090
rect 59899 -68271 59905 -68095
rect 59899 -68280 59916 -68271
rect 60006 -68280 60016 -68090
rect 60076 -68125 60196 -68067
rect 60346 -67850 60426 -67800
rect 60346 -67890 60366 -67850
rect 60406 -67890 60426 -67850
rect 60346 -67940 60426 -67890
rect 60346 -67980 60366 -67940
rect 60406 -67980 60426 -67940
rect 60346 -68020 60426 -67980
rect 60346 -68060 60366 -68020
rect 60406 -68060 60426 -68020
rect 60346 -68070 60426 -68060
rect 60636 -67849 60816 -67791
rect 60636 -67883 60671 -67849
rect 60705 -67883 60747 -67849
rect 60781 -67883 60816 -67849
rect 60636 -67941 60816 -67883
rect 60636 -67975 60671 -67941
rect 60705 -67975 60747 -67941
rect 60781 -67975 60816 -67941
rect 60636 -68033 60816 -67975
rect 60636 -68067 60671 -68033
rect 60705 -68067 60747 -68033
rect 60781 -68067 60816 -68033
rect 60076 -68159 60127 -68125
rect 60161 -68159 60196 -68125
rect 60076 -68190 60196 -68159
rect 60276 -68110 60546 -68100
rect 60276 -68125 60476 -68110
rect 60276 -68159 60297 -68125
rect 60331 -68159 60369 -68125
rect 60405 -68159 60449 -68125
rect 60276 -68170 60476 -68159
rect 60536 -68170 60546 -68110
rect 60276 -68180 60546 -68170
rect 60636 -68125 60816 -68067
rect 61026 -67730 61036 -67620
rect 61126 -67730 61136 -67620
rect 61176 -67680 61196 -67600
rect 61366 -67680 61386 -67600
rect 61176 -67700 61386 -67680
rect 61026 -67760 61136 -67730
rect 61026 -67800 61046 -67760
rect 61086 -67800 61136 -67760
rect 61026 -67850 61136 -67800
rect 61026 -67890 61046 -67850
rect 61086 -67890 61136 -67850
rect 61026 -67940 61136 -67890
rect 61026 -67980 61046 -67940
rect 61086 -67980 61136 -67940
rect 61026 -68020 61136 -67980
rect 61026 -68060 61046 -68020
rect 61086 -68060 61136 -68020
rect 61026 -68080 61136 -68060
rect 61256 -67757 61366 -67700
rect 61256 -67791 61291 -67757
rect 61325 -67791 61366 -67757
rect 61256 -67849 61366 -67791
rect 61256 -67850 61291 -67849
rect 61325 -67850 61366 -67849
rect 61256 -68060 61276 -67850
rect 61356 -68060 61366 -67850
rect 61256 -68067 61291 -68060
rect 61325 -68067 61366 -68060
rect 60636 -68159 60671 -68125
rect 60705 -68159 60747 -68125
rect 60781 -68159 60816 -68125
rect 60636 -68240 60816 -68159
rect 60966 -68124 61177 -68110
rect 60966 -68125 61129 -68124
rect 60966 -68159 60980 -68125
rect 61015 -68159 61053 -68125
rect 61088 -68158 61129 -68125
rect 61164 -68158 61177 -68124
rect 61088 -68159 61177 -68158
rect 60966 -68190 61177 -68159
rect 61256 -68125 61366 -68067
rect 61256 -68159 61291 -68125
rect 61325 -68159 61366 -68125
rect 61256 -68190 61366 -68159
rect 60466 -68250 60546 -68240
rect 59899 -68283 59945 -68280
rect 60466 -68310 60476 -68250
rect 60536 -68310 60546 -68250
rect 59849 -68320 59907 -68315
rect 60466 -68320 60546 -68310
rect 60606 -68250 60826 -68240
rect 60606 -68310 60616 -68250
rect 60736 -68310 60756 -68250
rect 60816 -68310 60826 -68250
rect 60606 -68320 60826 -68310
rect 60886 -68250 60966 -68240
rect 60886 -68310 60896 -68250
rect 60956 -68310 60966 -68250
rect 60886 -68320 60966 -68310
rect 59736 -68321 59926 -68320
rect 59736 -68355 59861 -68321
rect 59895 -68355 59926 -68321
rect 59736 -68380 59926 -68355
rect 60636 -68370 60816 -68320
rect 59376 -68420 59826 -68410
rect 59376 -68460 59476 -68420
rect 59646 -68460 59826 -68420
rect 59376 -68470 59826 -68460
rect 59156 -68490 59236 -68477
rect 58896 -68500 59086 -68490
rect 56380 -68568 57000 -68558
rect 57356 -68564 57676 -68550
rect 56440 -68574 57000 -68568
rect 57314 -68570 57676 -68564
rect 56440 -68594 57178 -68574
rect 56440 -68644 57118 -68594
rect 57168 -68644 57178 -68594
rect 57314 -68610 57326 -68570
rect 57376 -68610 57676 -68570
rect 57314 -68616 57676 -68610
rect 57356 -68630 57676 -68616
rect 56440 -68654 57178 -68644
rect 56440 -68688 57000 -68654
rect 57112 -68656 57174 -68654
rect 56380 -68758 57000 -68688
rect 56032 -68830 56038 -68828
rect 55992 -68842 56038 -68830
rect 55880 -68874 55970 -68868
rect 55870 -68878 55982 -68874
rect 55870 -68920 55880 -68878
rect 55970 -68920 55982 -68878
rect 55880 -68968 55970 -68958
rect 56120 -68998 56300 -68828
rect 57096 -68909 57372 -68878
rect 57096 -68943 57125 -68909
rect 57159 -68943 57217 -68909
rect 57251 -68943 57309 -68909
rect 57343 -68920 57372 -68909
rect 57343 -68943 57376 -68920
rect 57096 -68980 57376 -68943
rect 57066 -68990 57376 -68980
rect 56426 -68998 57376 -68990
rect 56120 -69008 57376 -68998
rect 56014 -69058 56086 -69046
rect 55570 -69178 55830 -69068
rect 53961 -69244 53988 -69206
rect 54022 -69244 54031 -69206
rect 53961 -69258 54031 -69244
rect 54910 -69206 54981 -69194
rect 54910 -69244 54916 -69206
rect 54950 -69244 54981 -69206
rect 54910 -69256 54981 -69244
rect 54911 -69258 54981 -69256
rect 55220 -69218 55330 -69208
rect 54069 -69272 54869 -69266
rect 54069 -69306 54081 -69272
rect 54857 -69278 54869 -69272
rect 54857 -69306 54880 -69278
rect 54069 -69312 54880 -69306
rect 54090 -69388 54880 -69312
rect 55330 -69318 55380 -69218
rect 55330 -69328 55480 -69318
rect 55220 -69338 55480 -69328
rect 55280 -69352 55480 -69338
rect 55280 -69358 55488 -69352
rect 55280 -69378 55300 -69358
rect 54090 -69488 54150 -69388
rect 54840 -69488 54880 -69388
rect 55288 -69392 55300 -69378
rect 55476 -69392 55488 -69358
rect 55530 -69378 55610 -69368
rect 55288 -69398 55488 -69392
rect 55520 -69402 55530 -69390
rect 55520 -69436 55526 -69402
rect 55288 -69446 55488 -69440
rect 55288 -69480 55300 -69446
rect 55476 -69480 55488 -69446
rect 55520 -69448 55530 -69436
rect 55530 -69478 55610 -69468
rect 55288 -69486 55488 -69480
rect 54090 -69508 54140 -69488
rect 54100 -69748 54140 -69508
rect 54850 -69748 54880 -69488
rect 55300 -69528 55470 -69486
rect 55300 -69668 55320 -69528
rect 55470 -69614 55482 -69542
rect 55300 -69678 55470 -69668
rect 54100 -69788 54880 -69748
rect 55710 -69998 55830 -69178
rect 56014 -69208 56020 -69058
rect 56080 -69208 56086 -69058
rect 56014 -69220 56086 -69208
rect 56120 -69208 56170 -69008
rect 56390 -69060 57376 -69008
rect 56390 -69068 57156 -69060
rect 56390 -69208 56654 -69068
rect 56120 -69258 56654 -69208
rect 56306 -69286 56654 -69258
rect 56998 -69220 57156 -69068
rect 57316 -69220 57376 -69060
rect 56998 -69286 57376 -69220
rect 56306 -69700 57376 -69286
rect 57556 -69410 57676 -68630
rect 58896 -68660 58986 -68500
rect 59756 -68520 59826 -68470
rect 59066 -68536 59176 -68530
rect 59066 -68540 59103 -68536
rect 59137 -68540 59176 -68536
rect 59066 -68600 59076 -68540
rect 59166 -68600 59176 -68540
rect 59066 -68610 59176 -68600
rect 58896 -69030 58926 -68660
rect 58966 -69030 58986 -68730
rect 59116 -68660 59506 -68640
rect 59116 -68730 59146 -68660
rect 59226 -68730 59276 -68660
rect 59356 -68730 59396 -68660
rect 59476 -68730 59506 -68660
rect 59116 -68748 59506 -68730
rect 59646 -68660 59716 -68640
rect 59706 -68720 59716 -68660
rect 59646 -68730 59716 -68720
rect 59113 -68754 59513 -68748
rect 59113 -68788 59125 -68754
rect 59501 -68788 59513 -68754
rect 59113 -68794 59513 -68788
rect 59546 -68800 59616 -68790
rect 59246 -68856 59256 -68830
rect 59113 -68862 59256 -68856
rect 59366 -68856 59376 -68830
rect 59366 -68862 59513 -68856
rect 59016 -68900 59076 -68880
rect 59113 -68896 59125 -68862
rect 59501 -68896 59513 -68862
rect 59606 -68860 59616 -68800
rect 59546 -68870 59616 -68860
rect 59113 -68902 59513 -68896
rect 59016 -68990 59076 -68960
rect 59113 -68970 59513 -68964
rect 59113 -69004 59125 -68970
rect 59501 -69004 59513 -68970
rect 59113 -69010 59513 -69004
rect 58896 -69100 58906 -69030
rect 58896 -69120 58986 -69100
rect 59116 -69030 59516 -69010
rect 59116 -69100 59146 -69030
rect 59226 -69100 59276 -69030
rect 59356 -69100 59396 -69030
rect 59476 -69100 59516 -69030
rect 59116 -69120 59516 -69100
rect 59646 -69030 59656 -68730
rect 59706 -69030 59716 -68730
rect 59756 -68700 59766 -68520
rect 59806 -68700 59826 -68520
rect 59956 -68520 60336 -68510
rect 59956 -68534 59966 -68520
rect 59946 -68540 59966 -68534
rect 60326 -68534 60336 -68520
rect 60326 -68540 60346 -68534
rect 59856 -68580 59916 -68570
rect 59946 -68574 59958 -68540
rect 60334 -68574 60346 -68540
rect 61056 -68540 61176 -68190
rect 59946 -68580 59966 -68574
rect 60326 -68580 60346 -68574
rect 60376 -68580 60436 -68560
rect 59956 -68590 60336 -68580
rect 59856 -68660 59916 -68640
rect 59946 -68648 60346 -68642
rect 59756 -68740 59826 -68700
rect 59946 -68682 59958 -68648
rect 60334 -68682 60346 -68648
rect 60376 -68660 60436 -68640
rect 61126 -68640 61176 -68540
rect 61056 -68670 61176 -68640
rect 59946 -68688 60346 -68682
rect 59946 -68740 60336 -68688
rect 59756 -68760 60536 -68740
rect 59756 -68800 59866 -68760
rect 60426 -68800 60536 -68760
rect 59756 -68810 60536 -68800
rect 59796 -68920 59806 -68810
rect 59916 -68920 59926 -68810
rect 59796 -68930 59926 -68920
rect 60436 -68830 60536 -68810
rect 60436 -68950 60446 -68830
rect 60526 -68950 60536 -68830
rect 60436 -68960 60536 -68950
rect 59646 -69040 59716 -69030
rect 59706 -69100 59716 -69040
rect 59646 -69120 59716 -69100
rect 58806 -69410 59356 -69380
rect 57556 -69420 59356 -69410
rect 57556 -69560 58986 -69420
rect 59126 -69560 59356 -69420
rect 59846 -69390 60256 -69380
rect 59846 -69500 59996 -69390
rect 60106 -69500 60256 -69390
rect 57556 -69610 59356 -69560
rect 58806 -69690 59356 -69610
rect 55710 -70000 55910 -69998
rect 55400 -70100 56200 -70000
rect 59600 -70100 60500 -69500
rect 55400 -70500 55500 -70100
rect 56100 -70500 56200 -70100
rect 55400 -70600 56200 -70500
rect 55380 -71080 55800 -71000
rect 55380 -71360 55460 -71080
rect 55720 -71360 55800 -71080
rect 55380 -71440 55800 -71360
rect 54090 -71538 54890 -71498
rect 54090 -71668 54150 -71538
rect 53510 -71720 53800 -71718
rect 53460 -71740 53800 -71720
rect 53460 -71940 53480 -71740
rect 53780 -71940 53800 -71740
rect 54080 -71798 54150 -71668
rect 54860 -71778 54890 -71538
rect 54850 -71798 54890 -71778
rect 54080 -71866 54880 -71798
rect 54079 -71872 54880 -71866
rect 54079 -71906 54091 -71872
rect 54867 -71898 54880 -71872
rect 54867 -71906 54879 -71898
rect 54079 -71912 54879 -71906
rect 53460 -71960 53800 -71940
rect 53510 -72058 53800 -71960
rect 53002 -72220 53480 -72158
rect 53000 -72358 53480 -72220
rect 53510 -72168 53520 -72058
rect 53640 -72168 53800 -72058
rect 53510 -72288 53800 -72168
rect 53970 -71934 54040 -71918
rect 53970 -71972 53998 -71934
rect 54032 -71972 54040 -71934
rect 53970 -72168 54040 -71972
rect 54920 -71934 54990 -71918
rect 54920 -71972 54926 -71934
rect 54960 -71972 54990 -71934
rect 54079 -72000 54879 -71994
rect 54079 -72034 54091 -72000
rect 54867 -72034 54879 -72000
rect 54079 -72038 54879 -72034
rect 54079 -72040 54750 -72038
rect 54090 -72088 54750 -72040
rect 54740 -72118 54750 -72088
rect 54850 -72040 54879 -72038
rect 54850 -72108 54860 -72040
rect 54840 -72118 54860 -72108
rect 54750 -72128 54860 -72118
rect 54920 -72168 54990 -71972
rect 55430 -72018 55520 -72008
rect 55290 -72128 55390 -72118
rect 53970 -72198 55290 -72168
rect 55430 -72158 55520 -72088
rect 53970 -72208 55390 -72198
rect 54050 -72218 55380 -72208
rect 54050 -72228 54880 -72218
rect 54050 -72238 54091 -72228
rect 54079 -72262 54091 -72238
rect 54867 -72238 54880 -72228
rect 54867 -72262 54879 -72238
rect 54079 -72268 54879 -72262
rect 54920 -72278 54990 -72268
rect 53510 -72306 53630 -72288
rect 53510 -72338 53526 -72306
rect 53514 -72340 53526 -72338
rect 53614 -72338 53630 -72306
rect 53940 -72290 54038 -72278
rect 53940 -72298 53998 -72290
rect 53614 -72340 53626 -72338
rect 53514 -72346 53626 -72340
rect 53000 -74108 53050 -72358
rect 53250 -72368 53480 -72358
rect 53250 -73718 53330 -72368
rect 53400 -72378 53480 -72368
rect 53400 -72390 53504 -72378
rect 53400 -73166 53464 -72390
rect 53498 -73166 53504 -72390
rect 53400 -73178 53504 -73166
rect 53636 -72388 53682 -72378
rect 53636 -72390 53760 -72388
rect 53636 -73166 53642 -72390
rect 53676 -73166 53760 -72390
rect 53940 -72398 53950 -72298
rect 54032 -72328 54038 -72290
rect 54020 -72340 54038 -72328
rect 54020 -72398 54030 -72340
rect 54079 -72356 54879 -72350
rect 54079 -72390 54091 -72356
rect 54867 -72390 54879 -72356
rect 54920 -72378 54990 -72368
rect 55320 -72368 55380 -72218
rect 54079 -72396 54879 -72390
rect 53940 -72418 54030 -72398
rect 54090 -72428 54870 -72396
rect 55320 -72402 55334 -72368
rect 55368 -72402 55380 -72368
rect 55320 -72408 55380 -72402
rect 53840 -72728 53920 -72718
rect 53840 -72838 53860 -72728
rect 53840 -72848 53920 -72838
rect 53840 -73040 53900 -72848
rect 54320 -72928 54510 -72428
rect 55440 -72438 55520 -72158
rect 55410 -72440 55520 -72438
rect 55284 -72448 55330 -72440
rect 55230 -72452 55330 -72448
rect 55230 -72458 55290 -72452
rect 55324 -72628 55330 -72452
rect 55230 -72638 55330 -72628
rect 55284 -72640 55330 -72638
rect 55372 -72448 55520 -72440
rect 55372 -72452 55430 -72448
rect 55372 -72628 55378 -72452
rect 55412 -72618 55430 -72452
rect 55510 -72618 55520 -72448
rect 55412 -72628 55520 -72618
rect 55372 -72640 55418 -72628
rect 55580 -72728 55720 -71440
rect 58776 -71670 59306 -71550
rect 58776 -71680 58966 -71670
rect 56146 -71780 57366 -71730
rect 55954 -71928 56046 -71916
rect 56146 -71928 56506 -71780
rect 55954 -72098 55960 -71928
rect 56040 -72098 56046 -71928
rect 55954 -72110 56046 -72098
rect 56120 -71958 56506 -71928
rect 56120 -72168 56190 -71958
rect 56390 -72030 56506 -71958
rect 57016 -71934 57366 -71780
rect 57586 -71830 58966 -71680
rect 59126 -71830 59306 -71670
rect 57586 -71850 59306 -71830
rect 59946 -71700 60386 -71600
rect 57586 -71880 58986 -71850
rect 59946 -71860 59956 -71700
rect 60166 -71860 60386 -71700
rect 57016 -72030 57368 -71934
rect 56390 -72070 57368 -72030
rect 56390 -72168 57126 -72070
rect 56120 -72174 57126 -72168
rect 56120 -72178 56750 -72174
rect 55880 -72218 55970 -72208
rect 55870 -72296 55880 -72250
rect 55970 -72296 55982 -72250
rect 55880 -72308 55970 -72298
rect 55000 -72738 55090 -72728
rect 55000 -72848 55090 -72838
rect 54710 -72928 54960 -72908
rect 53940 -72968 54960 -72928
rect 53940 -72972 54730 -72968
rect 53930 -72978 54730 -72972
rect 53930 -73012 53942 -72978
rect 54718 -73012 54730 -72978
rect 53930 -73018 54730 -73012
rect 53840 -73128 53858 -73040
rect 53892 -73128 53900 -73040
rect 53840 -73148 53900 -73128
rect 54762 -73038 54850 -73028
rect 54762 -73040 54770 -73038
rect 54762 -73128 54768 -73040
rect 54840 -73128 54850 -73038
rect 54762 -73140 54850 -73128
rect 54770 -73148 54850 -73140
rect 53636 -73178 53760 -73166
rect 53400 -73396 53480 -73178
rect 53514 -73216 53626 -73210
rect 53514 -73218 53526 -73216
rect 53510 -73250 53526 -73218
rect 53614 -73218 53626 -73216
rect 53614 -73250 53630 -73218
rect 53510 -73324 53630 -73250
rect 53510 -73358 53526 -73324
rect 53614 -73358 53630 -73324
rect 53680 -73238 53760 -73178
rect 53930 -73156 54730 -73150
rect 53930 -73190 53942 -73156
rect 54718 -73190 54730 -73156
rect 53930 -73196 54730 -73190
rect 53940 -73228 54720 -73196
rect 53920 -73238 54720 -73228
rect 53680 -73328 54720 -73238
rect 53514 -73364 53626 -73358
rect 53680 -73396 53760 -73328
rect 53920 -73338 54720 -73328
rect 53940 -73378 54720 -73338
rect 54900 -73368 54960 -72968
rect 55010 -72960 55090 -72848
rect 55540 -72738 55720 -72728
rect 55630 -72838 55720 -72738
rect 55130 -72874 55506 -72868
rect 55130 -72908 55142 -72874
rect 55494 -72908 55506 -72874
rect 55130 -72914 55506 -72908
rect 55010 -72994 55046 -72960
rect 55080 -72994 55090 -72960
rect 55010 -73008 55090 -72994
rect 55142 -73040 55494 -72914
rect 55540 -72960 55720 -72838
rect 55540 -72994 55556 -72960
rect 55590 -72994 55720 -72960
rect 55540 -73008 55720 -72994
rect 55780 -72340 55860 -72328
rect 55130 -73046 55506 -73040
rect 55130 -73080 55142 -73046
rect 55494 -73078 55506 -73046
rect 55494 -73080 55510 -73078
rect 55130 -73086 55510 -73080
rect 55140 -73098 55510 -73086
rect 55780 -73098 55820 -72340
rect 55140 -73116 55820 -73098
rect 55854 -73116 55860 -72340
rect 55140 -73128 55860 -73116
rect 55992 -72340 56038 -72328
rect 55992 -73116 55998 -72340
rect 56032 -72348 56038 -72340
rect 56120 -72348 56300 -72178
rect 57098 -72200 57126 -72174
rect 57356 -72200 57368 -72070
rect 57098 -72214 57368 -72200
rect 57096 -72245 57372 -72214
rect 57096 -72279 57125 -72245
rect 57159 -72279 57217 -72245
rect 57251 -72279 57309 -72245
rect 57343 -72279 57372 -72245
rect 57096 -72310 57372 -72279
rect 56032 -72706 56300 -72348
rect 56590 -72468 56660 -72458
rect 56660 -72534 57000 -72468
rect 57586 -72530 57706 -71880
rect 59946 -71890 60386 -71860
rect 57366 -72534 57706 -72530
rect 56660 -72538 57188 -72534
rect 56660 -72544 57190 -72538
rect 56660 -72594 57118 -72544
rect 57178 -72594 57190 -72544
rect 57314 -72540 57706 -72534
rect 57314 -72580 57326 -72540
rect 57366 -72580 57706 -72540
rect 57314 -72586 57706 -72580
rect 57366 -72590 57706 -72586
rect 58896 -72170 58986 -72150
rect 58896 -72230 58906 -72170
rect 58896 -72520 58926 -72230
rect 58966 -72520 58986 -72170
rect 59106 -72170 59516 -72160
rect 59106 -72230 59216 -72170
rect 59276 -72230 59326 -72170
rect 59386 -72230 59436 -72170
rect 59496 -72230 59516 -72170
rect 59106 -72247 59516 -72230
rect 59626 -72170 59706 -72130
rect 59626 -72230 59636 -72170
rect 59626 -72240 59656 -72230
rect 59106 -72280 59125 -72247
rect 59113 -72281 59125 -72280
rect 59501 -72280 59516 -72247
rect 59501 -72281 59513 -72280
rect 59113 -72287 59513 -72281
rect 59546 -72290 59616 -72280
rect 59276 -72330 59356 -72320
rect 59276 -72349 59286 -72330
rect 59113 -72355 59286 -72349
rect 59346 -72349 59356 -72330
rect 59346 -72355 59513 -72349
rect 59113 -72389 59125 -72355
rect 59501 -72389 59513 -72355
rect 59606 -72350 59616 -72290
rect 59546 -72360 59616 -72350
rect 59113 -72390 59286 -72389
rect 59346 -72390 59513 -72389
rect 59016 -72400 59076 -72390
rect 59113 -72395 59513 -72390
rect 59276 -72400 59356 -72395
rect 59546 -72410 59616 -72400
rect 59016 -72470 59076 -72460
rect 59113 -72463 59513 -72457
rect 59113 -72497 59125 -72463
rect 59501 -72497 59513 -72463
rect 59606 -72470 59616 -72410
rect 59546 -72480 59616 -72470
rect 59113 -72500 59513 -72497
rect 59113 -72503 59516 -72500
rect 58896 -72530 58986 -72520
rect 58896 -72590 58906 -72530
rect 58966 -72590 58986 -72530
rect 58896 -72592 58986 -72590
rect 59116 -72520 59516 -72503
rect 59646 -72510 59656 -72240
rect 59116 -72580 59216 -72520
rect 59276 -72580 59336 -72520
rect 59396 -72580 59436 -72520
rect 59496 -72580 59516 -72520
rect 56660 -72598 57190 -72594
rect 56590 -72600 57190 -72598
rect 56590 -72604 57188 -72600
rect 56590 -72668 57000 -72604
rect 56032 -72718 56356 -72706
rect 56032 -73116 56280 -72718
rect 55992 -73128 56280 -73116
rect 55140 -73138 55200 -73128
rect 55450 -73158 55810 -73128
rect 55870 -73166 55982 -73160
rect 55870 -73200 55882 -73166
rect 55970 -73200 55982 -73166
rect 55870 -73206 55982 -73200
rect 55140 -73218 55200 -73208
rect 55024 -73248 55116 -73236
rect 55024 -73328 55030 -73248
rect 55110 -73328 55116 -73248
rect 55024 -73340 55116 -73328
rect 55734 -73248 55816 -73236
rect 55734 -73328 55740 -73248
rect 55810 -73328 55816 -73248
rect 55734 -73340 55816 -73328
rect 55880 -73238 55970 -73206
rect 55880 -73364 55970 -73328
rect 56060 -73348 56280 -73128
rect 56350 -73348 56356 -72718
rect 56480 -72788 56550 -72778
rect 56480 -72858 56550 -72848
rect 56590 -72887 56750 -72668
rect 58894 -72686 58988 -72592
rect 59116 -72600 59516 -72580
rect 59636 -72520 59656 -72510
rect 59696 -72520 59706 -72170
rect 59856 -72340 59976 -72330
rect 59856 -72430 59866 -72340
rect 59966 -72430 59976 -72340
rect 59856 -72440 59976 -72430
rect 60436 -72420 60446 -72320
rect 60526 -72420 60536 -72320
rect 60436 -72440 60536 -72420
rect 59636 -72530 59706 -72520
rect 59696 -72590 59706 -72530
rect 59636 -72610 59706 -72590
rect 59756 -72460 60536 -72440
rect 59756 -72500 59866 -72460
rect 60426 -72500 60536 -72460
rect 59756 -72510 60536 -72500
rect 59756 -72550 59826 -72510
rect 59066 -72640 59176 -72630
rect 58896 -72750 58986 -72686
rect 59066 -72710 59076 -72640
rect 59166 -72710 59176 -72640
rect 59066 -72712 59103 -72710
rect 59137 -72712 59176 -72710
rect 59066 -72720 59176 -72712
rect 59756 -72740 59766 -72550
rect 59806 -72740 59826 -72550
rect 59956 -72568 60046 -72540
rect 59946 -72574 60046 -72568
rect 60126 -72568 60336 -72540
rect 60126 -72574 60346 -72568
rect 59856 -72610 59916 -72600
rect 59946 -72608 59958 -72574
rect 60334 -72608 60346 -72574
rect 59946 -72614 60346 -72608
rect 60376 -72620 60446 -72610
rect 59856 -72690 59916 -72680
rect 59946 -72682 60346 -72676
rect 59946 -72716 59958 -72682
rect 60334 -72716 60346 -72682
rect 60376 -72690 60446 -72680
rect 59946 -72722 59976 -72716
rect 57098 -72758 57368 -72754
rect 57096 -72764 57372 -72758
rect 57096 -72850 57098 -72764
rect 56424 -72888 56470 -72887
rect 56060 -73360 56356 -73348
rect 56410 -72899 56470 -72888
rect 53400 -73408 53504 -73396
rect 53400 -73718 53464 -73408
rect 53250 -74108 53464 -73718
rect 53000 -74184 53464 -74108
rect 53498 -74184 53504 -73408
rect 53000 -74188 53504 -74184
rect 53458 -74196 53504 -74188
rect 53636 -73408 53760 -73396
rect 53636 -74184 53642 -73408
rect 53676 -74184 53760 -73408
rect 53930 -73384 54730 -73378
rect 53930 -73418 53942 -73384
rect 54718 -73418 54730 -73384
rect 53930 -73424 54730 -73418
rect 53830 -73446 53900 -73428
rect 53830 -73534 53858 -73446
rect 53892 -73534 53900 -73446
rect 53830 -73728 53900 -73534
rect 54760 -73446 54850 -73428
rect 54760 -73534 54768 -73446
rect 54802 -73448 54850 -73446
rect 54900 -73438 55200 -73368
rect 55870 -73370 55982 -73364
rect 55870 -73404 55882 -73370
rect 55970 -73404 55982 -73370
rect 55450 -73438 55810 -73408
rect 55870 -73410 55982 -73404
rect 56060 -73438 56300 -73360
rect 54900 -73442 55820 -73438
rect 56000 -73442 56300 -73438
rect 54900 -73448 55860 -73442
rect 54840 -73528 54850 -73448
rect 54802 -73534 54850 -73528
rect 54760 -73548 54850 -73534
rect 55130 -73454 55860 -73448
rect 55130 -73478 55820 -73454
rect 55130 -73496 55510 -73478
rect 55130 -73530 55142 -73496
rect 55494 -73498 55510 -73496
rect 55494 -73530 55506 -73498
rect 55130 -73536 55506 -73530
rect 53930 -73562 54730 -73556
rect 53930 -73596 53942 -73562
rect 54718 -73596 54730 -73562
rect 55020 -73582 55090 -73568
rect 53930 -73602 54730 -73596
rect 53940 -73608 54730 -73602
rect 54920 -73598 54980 -73588
rect 53940 -73648 54920 -73608
rect 53830 -73738 53920 -73728
rect 53830 -73848 53850 -73738
rect 53830 -73858 53920 -73848
rect 54320 -74148 54510 -73648
rect 54710 -73668 54920 -73648
rect 54910 -73678 54980 -73668
rect 55020 -73616 55046 -73582
rect 55080 -73616 55090 -73582
rect 55020 -73728 55090 -73616
rect 55142 -73662 55494 -73536
rect 55540 -73582 55620 -73568
rect 55540 -73616 55556 -73582
rect 55590 -73616 55620 -73582
rect 55130 -73668 55506 -73662
rect 55130 -73702 55142 -73668
rect 55494 -73702 55506 -73668
rect 55130 -73708 55506 -73702
rect 55000 -73738 55090 -73728
rect 55000 -73848 55090 -73838
rect 55540 -73728 55620 -73616
rect 55540 -73738 55630 -73728
rect 55630 -73838 55680 -73748
rect 55540 -73848 55680 -73838
rect 55274 -73938 55320 -73936
rect 55220 -73948 55320 -73938
rect 55220 -74124 55280 -74118
rect 55314 -74124 55320 -73948
rect 55220 -74128 55320 -74124
rect 55274 -74136 55320 -74128
rect 55362 -73948 55408 -73936
rect 55362 -74124 55368 -73948
rect 55402 -73958 55510 -73948
rect 55402 -74124 55410 -73958
rect 55362 -74128 55410 -74124
rect 55500 -74128 55510 -73958
rect 55362 -74136 55510 -74128
rect 55390 -74138 55510 -74136
rect 53636 -74188 53760 -74184
rect 53636 -74196 53682 -74188
rect 53940 -74208 54020 -74168
rect 54080 -74182 54860 -74148
rect 55311 -74174 55371 -74168
rect 53514 -74234 53626 -74228
rect 53514 -74238 53526 -74234
rect 53510 -74268 53526 -74238
rect 53614 -74238 53626 -74234
rect 53614 -74268 53630 -74238
rect 53510 -74328 53630 -74268
rect 53940 -74288 53950 -74208
rect 54010 -74238 54020 -74208
rect 54069 -74188 54869 -74182
rect 54069 -74222 54081 -74188
rect 54857 -74222 54869 -74188
rect 54069 -74228 54869 -74222
rect 54910 -74198 54980 -74188
rect 54010 -74250 54028 -74238
rect 54022 -74288 54028 -74250
rect 53940 -74300 54028 -74288
rect 53940 -74308 54020 -74300
rect 54910 -74308 54980 -74298
rect 55311 -74208 55324 -74174
rect 55358 -74208 55371 -74174
rect 54070 -74310 54870 -74308
rect 54069 -74316 54870 -74310
rect 54069 -74338 54081 -74316
rect 54041 -74350 54081 -74338
rect 54857 -74318 54870 -74316
rect 54857 -74350 54880 -74318
rect 55311 -74348 55371 -74208
rect 54041 -74358 54880 -74350
rect 55240 -74358 55371 -74348
rect 54041 -74368 55240 -74358
rect 53510 -74458 53630 -74448
rect 53961 -74408 55240 -74368
rect 53961 -74606 54031 -74408
rect 54730 -74468 54860 -74458
rect 54730 -74488 54740 -74468
rect 54080 -74538 54740 -74488
rect 54069 -74544 54740 -74538
rect 54850 -74538 54860 -74468
rect 54850 -74544 54869 -74538
rect 54069 -74578 54081 -74544
rect 54857 -74578 54869 -74544
rect 54069 -74584 54869 -74578
rect 54911 -74594 54981 -74408
rect 55370 -74408 55371 -74358
rect 55240 -74428 55370 -74418
rect 55410 -74448 55510 -74138
rect 55410 -74558 55510 -74538
rect 55570 -74468 55680 -73848
rect 55780 -74230 55820 -73478
rect 55854 -74230 55860 -73454
rect 55780 -74238 55860 -74230
rect 55814 -74242 55860 -74238
rect 55992 -73454 56300 -73442
rect 55992 -74230 55998 -73454
rect 56032 -74228 56300 -73454
rect 56410 -73498 56430 -72899
rect 56380 -73675 56430 -73498
rect 56464 -73675 56470 -72899
rect 56380 -73687 56470 -73675
rect 56552 -72899 56750 -72887
rect 56552 -73675 56558 -72899
rect 56592 -73038 56750 -72899
rect 57066 -72880 57098 -72850
rect 57368 -72850 57372 -72764
rect 58896 -72759 59076 -72750
rect 58896 -72760 59084 -72759
rect 59156 -72760 59202 -72759
rect 57368 -72880 57396 -72850
rect 57066 -73010 57086 -72880
rect 57376 -73010 57396 -72880
rect 56592 -73675 56610 -73038
rect 57066 -73040 57396 -73010
rect 56860 -73190 57060 -73178
rect 56860 -73218 57236 -73190
rect 56860 -73348 56900 -73218
rect 57020 -73348 57236 -73218
rect 56860 -73388 57236 -73348
rect 57036 -73390 57236 -73388
rect 58556 -73280 58756 -73260
rect 58556 -73440 58576 -73280
rect 58736 -73440 58756 -73280
rect 58556 -73460 58756 -73440
rect 56552 -73678 56610 -73675
rect 57036 -73540 57446 -73530
rect 56552 -73687 56598 -73678
rect 57036 -73680 57056 -73540
rect 57416 -73680 57446 -73540
rect 56380 -73958 56440 -73687
rect 57036 -73700 57098 -73680
rect 56480 -73728 56550 -73718
rect 56480 -73798 56550 -73788
rect 57096 -73814 57098 -73734
rect 57368 -73700 57446 -73680
rect 57368 -73814 57372 -73734
rect 57096 -73830 57372 -73814
rect 58896 -73890 58926 -72760
rect 58966 -72771 59086 -72760
rect 58966 -73147 59044 -72771
rect 59078 -73147 59086 -72771
rect 58966 -73170 59086 -73147
rect 59156 -72771 59256 -72760
rect 59756 -72770 59826 -72740
rect 59966 -72752 59976 -72722
rect 60316 -72722 60346 -72716
rect 61036 -72720 61466 -72710
rect 60316 -72752 60326 -72722
rect 59966 -72760 60326 -72752
rect 59156 -73147 59162 -72771
rect 59196 -72840 59256 -72771
rect 59236 -72920 59256 -72840
rect 59196 -73040 59256 -72920
rect 59236 -73120 59256 -73040
rect 59196 -73147 59256 -73120
rect 59156 -73160 59256 -73147
rect 58966 -73480 59036 -73170
rect 59066 -73206 59176 -73200
rect 59066 -73210 59103 -73206
rect 59137 -73210 59176 -73206
rect 59066 -73280 59076 -73210
rect 59166 -73280 59176 -73210
rect 59066 -73290 59176 -73280
rect 59206 -73360 59256 -73160
rect 59376 -72790 59826 -72770
rect 59376 -72830 59476 -72790
rect 59656 -72830 59826 -72790
rect 59376 -72840 59826 -72830
rect 59376 -72890 59436 -72840
rect 59376 -73250 59386 -72890
rect 59426 -73250 59436 -72890
rect 59526 -72898 59576 -72870
rect 59526 -72932 59546 -72898
rect 59636 -72930 59706 -72870
rect 59580 -72932 59706 -72930
rect 59526 -72940 59706 -72932
rect 59476 -72982 59546 -72970
rect 59476 -73050 59502 -72982
rect 59476 -73158 59502 -73120
rect 59536 -73158 59546 -72982
rect 59476 -73170 59546 -73158
rect 59576 -72982 59636 -72970
rect 59576 -72990 59590 -72982
rect 59624 -72990 59636 -72982
rect 59576 -73170 59636 -73160
rect 59534 -73208 59592 -73202
rect 59534 -73210 59546 -73208
rect 59066 -73370 59176 -73360
rect 59066 -73440 59076 -73370
rect 59166 -73440 59176 -73370
rect 59066 -73442 59103 -73440
rect 59137 -73442 59176 -73440
rect 59066 -73450 59176 -73442
rect 59206 -73370 59266 -73360
rect 59206 -73450 59266 -73440
rect 59376 -73400 59436 -73250
rect 59516 -73242 59546 -73210
rect 59580 -73210 59592 -73208
rect 59666 -73210 59706 -72940
rect 59580 -73242 59706 -73210
rect 59516 -73280 59706 -73242
rect 59746 -72898 59936 -72870
rect 59746 -72932 59862 -72898
rect 59896 -72932 59936 -72898
rect 59746 -72940 59936 -72932
rect 61036 -72900 61206 -72720
rect 61346 -72900 61466 -72720
rect 61036 -72940 61466 -72900
rect 59746 -73200 59776 -72940
rect 60286 -72950 60476 -72940
rect 59806 -72982 59866 -72970
rect 59806 -73000 59818 -72982
rect 59852 -73000 59866 -72982
rect 59806 -73158 59818 -73140
rect 59852 -73158 59866 -73140
rect 59806 -73170 59866 -73158
rect 59900 -72980 60016 -72970
rect 59900 -72982 59916 -72980
rect 59900 -73158 59906 -72982
rect 59900 -73160 59916 -73158
rect 60006 -73160 60016 -72980
rect 60286 -73090 60306 -72950
rect 60456 -73090 60476 -72950
rect 61176 -73000 61386 -72980
rect 60286 -73100 60476 -73090
rect 61026 -73020 61136 -73010
rect 59900 -73170 60016 -73160
rect 60076 -73157 60196 -73120
rect 60076 -73191 60127 -73157
rect 60161 -73191 60196 -73157
rect 59746 -73208 59926 -73200
rect 59746 -73210 59862 -73208
rect 59896 -73210 59926 -73208
rect 59746 -73280 59826 -73210
rect 59916 -73280 59926 -73210
rect 59746 -73290 59926 -73280
rect 60076 -73249 60196 -73191
rect 60336 -73160 60446 -73100
rect 60336 -73200 60366 -73160
rect 60406 -73200 60446 -73160
rect 60636 -73157 60816 -73120
rect 60636 -73191 60671 -73157
rect 60705 -73191 60747 -73157
rect 60781 -73191 60816 -73157
rect 60076 -73280 60127 -73249
rect 60161 -73280 60196 -73249
rect 59736 -73370 59936 -73360
rect 58966 -73501 59086 -73480
rect 58966 -73877 59044 -73501
rect 59078 -73877 59086 -73501
rect 58966 -73890 59086 -73877
rect 59156 -73490 59202 -73489
rect 59156 -73501 59236 -73490
rect 59156 -73877 59162 -73501
rect 59196 -73530 59236 -73501
rect 59226 -73610 59236 -73530
rect 59196 -73760 59236 -73610
rect 59226 -73840 59236 -73760
rect 59196 -73877 59236 -73840
rect 59376 -73770 59386 -73400
rect 59426 -73770 59436 -73400
rect 59516 -73411 59706 -73370
rect 59516 -73445 59545 -73411
rect 59579 -73445 59706 -73411
rect 59516 -73450 59706 -73445
rect 59533 -73451 59591 -73450
rect 59466 -73495 59546 -73480
rect 59586 -73483 59646 -73480
rect 59466 -73530 59501 -73495
rect 59466 -73671 59501 -73610
rect 59535 -73671 59546 -73495
rect 59466 -73680 59546 -73671
rect 59583 -73495 59646 -73483
rect 59583 -73510 59589 -73495
rect 59623 -73510 59646 -73495
rect 59583 -73650 59586 -73510
rect 59583 -73671 59589 -73650
rect 59623 -73671 59646 -73650
rect 59583 -73680 59646 -73671
rect 59495 -73683 59541 -73680
rect 59583 -73683 59629 -73680
rect 59533 -73720 59591 -73715
rect 59676 -73720 59706 -73450
rect 59376 -73810 59436 -73770
rect 59506 -73780 59516 -73720
rect 59596 -73780 59706 -73720
rect 59736 -73440 59826 -73370
rect 59926 -73440 59936 -73370
rect 59736 -73445 59861 -73440
rect 59895 -73445 59936 -73440
rect 59736 -73450 59936 -73445
rect 60076 -73440 60096 -73280
rect 60176 -73440 60196 -73280
rect 59736 -73720 59766 -73450
rect 59849 -73451 59907 -73450
rect 60076 -73467 60127 -73440
rect 60161 -73467 60196 -73440
rect 59796 -73483 59856 -73480
rect 59796 -73490 59857 -73483
rect 59856 -73670 59857 -73490
rect 59796 -73671 59817 -73670
rect 59851 -73671 59857 -73670
rect 59796 -73680 59857 -73671
rect 59811 -73683 59857 -73680
rect 59899 -73490 59945 -73483
rect 59899 -73495 59916 -73490
rect 59899 -73671 59905 -73495
rect 59899 -73680 59916 -73671
rect 60006 -73680 60016 -73490
rect 60076 -73525 60196 -73467
rect 60346 -73250 60426 -73200
rect 60346 -73290 60366 -73250
rect 60406 -73290 60426 -73250
rect 60346 -73340 60426 -73290
rect 60346 -73380 60366 -73340
rect 60406 -73380 60426 -73340
rect 60346 -73420 60426 -73380
rect 60346 -73460 60366 -73420
rect 60406 -73460 60426 -73420
rect 60346 -73470 60426 -73460
rect 60636 -73249 60816 -73191
rect 60636 -73283 60671 -73249
rect 60705 -73283 60747 -73249
rect 60781 -73283 60816 -73249
rect 60636 -73341 60816 -73283
rect 60636 -73375 60671 -73341
rect 60705 -73375 60747 -73341
rect 60781 -73375 60816 -73341
rect 60636 -73433 60816 -73375
rect 60636 -73467 60671 -73433
rect 60705 -73467 60747 -73433
rect 60781 -73467 60816 -73433
rect 60076 -73559 60127 -73525
rect 60161 -73559 60196 -73525
rect 60076 -73590 60196 -73559
rect 60276 -73510 60546 -73500
rect 60276 -73525 60476 -73510
rect 60276 -73559 60297 -73525
rect 60331 -73559 60369 -73525
rect 60405 -73559 60449 -73525
rect 60276 -73570 60476 -73559
rect 60536 -73570 60546 -73510
rect 60276 -73580 60546 -73570
rect 60636 -73525 60816 -73467
rect 61026 -73130 61036 -73020
rect 61126 -73130 61136 -73020
rect 61176 -73080 61196 -73000
rect 61366 -73080 61386 -73000
rect 61176 -73100 61386 -73080
rect 61026 -73160 61136 -73130
rect 61026 -73200 61046 -73160
rect 61086 -73200 61136 -73160
rect 61026 -73250 61136 -73200
rect 61026 -73290 61046 -73250
rect 61086 -73290 61136 -73250
rect 61026 -73340 61136 -73290
rect 61026 -73380 61046 -73340
rect 61086 -73380 61136 -73340
rect 61026 -73420 61136 -73380
rect 61026 -73460 61046 -73420
rect 61086 -73460 61136 -73420
rect 61026 -73480 61136 -73460
rect 61256 -73157 61366 -73100
rect 61256 -73191 61291 -73157
rect 61325 -73191 61366 -73157
rect 61256 -73249 61366 -73191
rect 61256 -73250 61291 -73249
rect 61325 -73250 61366 -73249
rect 61256 -73460 61276 -73250
rect 61356 -73460 61366 -73250
rect 61256 -73467 61291 -73460
rect 61325 -73467 61366 -73460
rect 60636 -73559 60671 -73525
rect 60705 -73559 60747 -73525
rect 60781 -73559 60816 -73525
rect 60636 -73640 60816 -73559
rect 60966 -73524 61177 -73510
rect 60966 -73525 61129 -73524
rect 60966 -73559 60980 -73525
rect 61015 -73559 61053 -73525
rect 61088 -73558 61129 -73525
rect 61164 -73558 61177 -73524
rect 61088 -73559 61177 -73558
rect 60966 -73590 61177 -73559
rect 61256 -73525 61366 -73467
rect 61256 -73559 61291 -73525
rect 61325 -73559 61366 -73525
rect 61256 -73590 61366 -73559
rect 60466 -73650 60546 -73640
rect 59899 -73683 59945 -73680
rect 60466 -73710 60476 -73650
rect 60536 -73710 60546 -73650
rect 59849 -73720 59907 -73715
rect 60466 -73720 60546 -73710
rect 60606 -73650 60826 -73640
rect 60606 -73710 60616 -73650
rect 60736 -73710 60756 -73650
rect 60816 -73710 60826 -73650
rect 60606 -73720 60826 -73710
rect 60886 -73650 60966 -73640
rect 60886 -73710 60896 -73650
rect 60956 -73710 60966 -73650
rect 60886 -73720 60966 -73710
rect 59736 -73721 59926 -73720
rect 59736 -73755 59861 -73721
rect 59895 -73755 59926 -73721
rect 59736 -73780 59926 -73755
rect 60636 -73770 60816 -73720
rect 59376 -73820 59826 -73810
rect 59376 -73860 59476 -73820
rect 59646 -73860 59826 -73820
rect 59376 -73870 59826 -73860
rect 59156 -73890 59236 -73877
rect 58896 -73900 59086 -73890
rect 56380 -73968 57000 -73958
rect 57356 -73964 57676 -73950
rect 56440 -73974 57000 -73968
rect 57314 -73970 57676 -73964
rect 56440 -73994 57178 -73974
rect 56440 -74044 57118 -73994
rect 57168 -74044 57178 -73994
rect 57314 -74010 57326 -73970
rect 57376 -74010 57676 -73970
rect 57314 -74016 57676 -74010
rect 57356 -74030 57676 -74016
rect 56440 -74054 57178 -74044
rect 56440 -74088 57000 -74054
rect 57112 -74056 57174 -74054
rect 56380 -74158 57000 -74088
rect 56032 -74230 56038 -74228
rect 55992 -74242 56038 -74230
rect 55880 -74274 55970 -74268
rect 55870 -74278 55982 -74274
rect 55870 -74320 55880 -74278
rect 55970 -74320 55982 -74278
rect 55880 -74368 55970 -74358
rect 56120 -74398 56300 -74228
rect 57096 -74309 57372 -74278
rect 57096 -74343 57125 -74309
rect 57159 -74343 57217 -74309
rect 57251 -74343 57309 -74309
rect 57343 -74320 57372 -74309
rect 57343 -74343 57376 -74320
rect 57096 -74380 57376 -74343
rect 57066 -74390 57376 -74380
rect 56426 -74398 57376 -74390
rect 56120 -74408 57376 -74398
rect 56014 -74458 56086 -74446
rect 55570 -74578 55830 -74468
rect 53961 -74644 53988 -74606
rect 54022 -74644 54031 -74606
rect 53961 -74658 54031 -74644
rect 54910 -74606 54981 -74594
rect 54910 -74644 54916 -74606
rect 54950 -74644 54981 -74606
rect 54910 -74656 54981 -74644
rect 54911 -74658 54981 -74656
rect 55220 -74618 55330 -74608
rect 54069 -74672 54869 -74666
rect 54069 -74706 54081 -74672
rect 54857 -74678 54869 -74672
rect 54857 -74706 54880 -74678
rect 54069 -74712 54880 -74706
rect 54090 -74788 54880 -74712
rect 55330 -74718 55380 -74618
rect 55330 -74728 55480 -74718
rect 55220 -74738 55480 -74728
rect 55280 -74752 55480 -74738
rect 55280 -74758 55488 -74752
rect 55280 -74778 55300 -74758
rect 54090 -74888 54150 -74788
rect 54840 -74888 54880 -74788
rect 55288 -74792 55300 -74778
rect 55476 -74792 55488 -74758
rect 55530 -74778 55610 -74768
rect 55288 -74798 55488 -74792
rect 55520 -74802 55530 -74790
rect 55520 -74836 55526 -74802
rect 55288 -74846 55488 -74840
rect 55288 -74880 55300 -74846
rect 55476 -74880 55488 -74846
rect 55520 -74848 55530 -74836
rect 55530 -74878 55610 -74868
rect 55288 -74886 55488 -74880
rect 54090 -74908 54140 -74888
rect 54100 -75148 54140 -74908
rect 54850 -75148 54880 -74888
rect 55300 -74928 55470 -74886
rect 55300 -75068 55320 -74928
rect 55470 -75014 55482 -74942
rect 55300 -75078 55470 -75068
rect 54100 -75188 54880 -75148
rect 55710 -75398 55830 -74578
rect 56014 -74608 56020 -74458
rect 56080 -74608 56086 -74458
rect 56014 -74620 56086 -74608
rect 56120 -74608 56170 -74408
rect 56390 -74460 57376 -74408
rect 56390 -74468 57156 -74460
rect 56390 -74608 56654 -74468
rect 56120 -74658 56654 -74608
rect 56306 -74686 56654 -74658
rect 56998 -74620 57156 -74468
rect 57316 -74620 57376 -74460
rect 56998 -74686 57376 -74620
rect 56306 -75100 57376 -74686
rect 57556 -74810 57676 -74030
rect 58896 -74060 58986 -73900
rect 59756 -73920 59826 -73870
rect 59066 -73936 59176 -73930
rect 59066 -73940 59103 -73936
rect 59137 -73940 59176 -73936
rect 59066 -74000 59076 -73940
rect 59166 -74000 59176 -73940
rect 59066 -74010 59176 -74000
rect 58896 -74430 58926 -74060
rect 58966 -74430 58986 -74130
rect 59116 -74060 59506 -74040
rect 59116 -74130 59146 -74060
rect 59226 -74130 59276 -74060
rect 59356 -74130 59396 -74060
rect 59476 -74130 59506 -74060
rect 59116 -74148 59506 -74130
rect 59646 -74060 59716 -74040
rect 59706 -74120 59716 -74060
rect 59646 -74130 59716 -74120
rect 59113 -74154 59513 -74148
rect 59113 -74188 59125 -74154
rect 59501 -74188 59513 -74154
rect 59113 -74194 59513 -74188
rect 59546 -74200 59616 -74190
rect 59246 -74256 59256 -74230
rect 59113 -74262 59256 -74256
rect 59366 -74256 59376 -74230
rect 59366 -74262 59513 -74256
rect 59016 -74300 59076 -74280
rect 59113 -74296 59125 -74262
rect 59501 -74296 59513 -74262
rect 59606 -74260 59616 -74200
rect 59546 -74270 59616 -74260
rect 59113 -74302 59513 -74296
rect 59016 -74390 59076 -74360
rect 59113 -74370 59513 -74364
rect 59113 -74404 59125 -74370
rect 59501 -74404 59513 -74370
rect 59113 -74410 59513 -74404
rect 58896 -74500 58906 -74430
rect 58896 -74520 58986 -74500
rect 59116 -74430 59516 -74410
rect 59116 -74500 59146 -74430
rect 59226 -74500 59276 -74430
rect 59356 -74500 59396 -74430
rect 59476 -74500 59516 -74430
rect 59116 -74520 59516 -74500
rect 59646 -74430 59656 -74130
rect 59706 -74430 59716 -74130
rect 59756 -74100 59766 -73920
rect 59806 -74100 59826 -73920
rect 59956 -73920 60336 -73910
rect 59956 -73934 59966 -73920
rect 59946 -73940 59966 -73934
rect 60326 -73934 60336 -73920
rect 60326 -73940 60346 -73934
rect 59856 -73980 59916 -73970
rect 59946 -73974 59958 -73940
rect 60334 -73974 60346 -73940
rect 61056 -73940 61176 -73590
rect 59946 -73980 59966 -73974
rect 60326 -73980 60346 -73974
rect 60376 -73980 60436 -73960
rect 59956 -73990 60336 -73980
rect 59856 -74060 59916 -74040
rect 59946 -74048 60346 -74042
rect 59756 -74140 59826 -74100
rect 59946 -74082 59958 -74048
rect 60334 -74082 60346 -74048
rect 60376 -74060 60436 -74040
rect 61126 -74040 61176 -73940
rect 61056 -74070 61176 -74040
rect 59946 -74088 60346 -74082
rect 59946 -74140 60336 -74088
rect 59756 -74160 60536 -74140
rect 59756 -74200 59866 -74160
rect 60426 -74200 60536 -74160
rect 59756 -74210 60536 -74200
rect 59796 -74320 59806 -74210
rect 59916 -74320 59926 -74210
rect 59796 -74330 59926 -74320
rect 60436 -74230 60536 -74210
rect 60436 -74350 60446 -74230
rect 60526 -74350 60536 -74230
rect 60436 -74360 60536 -74350
rect 59646 -74440 59716 -74430
rect 59706 -74500 59716 -74440
rect 59646 -74520 59716 -74500
rect 58806 -74810 59356 -74780
rect 57556 -74820 59356 -74810
rect 57556 -74960 58986 -74820
rect 59126 -74960 59356 -74820
rect 59846 -74790 60256 -74780
rect 59846 -74900 59996 -74790
rect 60106 -74900 60256 -74790
rect 57556 -75010 59356 -74960
rect 58806 -75090 59356 -75010
rect 55710 -75400 55910 -75398
rect 55400 -75500 56200 -75400
rect 59600 -75500 60500 -74900
rect 55400 -75900 55500 -75500
rect 56100 -75900 56200 -75500
rect 55400 -76000 56200 -75900
rect 55320 -76480 55800 -76400
rect 55320 -76760 55400 -76480
rect 55720 -76760 55800 -76480
rect 55320 -76840 55800 -76760
rect 54090 -76938 54890 -76898
rect 54090 -77068 54150 -76938
rect 53510 -77120 53800 -77118
rect 53460 -77140 53800 -77120
rect 53460 -77340 53480 -77140
rect 53780 -77340 53800 -77140
rect 54080 -77198 54150 -77068
rect 54860 -77178 54890 -76938
rect 54850 -77198 54890 -77178
rect 54080 -77266 54880 -77198
rect 54079 -77272 54880 -77266
rect 54079 -77306 54091 -77272
rect 54867 -77298 54880 -77272
rect 54867 -77306 54879 -77298
rect 54079 -77312 54879 -77306
rect 53460 -77360 53800 -77340
rect 53510 -77458 53800 -77360
rect 53002 -77620 53480 -77558
rect 53000 -77758 53480 -77620
rect 53510 -77568 53520 -77458
rect 53640 -77568 53800 -77458
rect 53510 -77688 53800 -77568
rect 53970 -77334 54040 -77318
rect 53970 -77372 53998 -77334
rect 54032 -77372 54040 -77334
rect 53970 -77568 54040 -77372
rect 54920 -77334 54990 -77318
rect 54920 -77372 54926 -77334
rect 54960 -77372 54990 -77334
rect 54079 -77400 54879 -77394
rect 54079 -77434 54091 -77400
rect 54867 -77434 54879 -77400
rect 54079 -77438 54879 -77434
rect 54079 -77440 54750 -77438
rect 54090 -77488 54750 -77440
rect 54740 -77518 54750 -77488
rect 54850 -77440 54879 -77438
rect 54850 -77508 54860 -77440
rect 54840 -77518 54860 -77508
rect 54750 -77528 54860 -77518
rect 54920 -77568 54990 -77372
rect 55430 -77418 55520 -77408
rect 55290 -77528 55390 -77518
rect 53970 -77598 55290 -77568
rect 55430 -77558 55520 -77488
rect 53970 -77608 55390 -77598
rect 54050 -77618 55380 -77608
rect 54050 -77628 54880 -77618
rect 54050 -77638 54091 -77628
rect 54079 -77662 54091 -77638
rect 54867 -77638 54880 -77628
rect 54867 -77662 54879 -77638
rect 54079 -77668 54879 -77662
rect 54920 -77678 54990 -77668
rect 53510 -77706 53630 -77688
rect 53510 -77738 53526 -77706
rect 53514 -77740 53526 -77738
rect 53614 -77738 53630 -77706
rect 53940 -77690 54038 -77678
rect 53940 -77698 53998 -77690
rect 53614 -77740 53626 -77738
rect 53514 -77746 53626 -77740
rect 53000 -79508 53050 -77758
rect 53250 -77768 53480 -77758
rect 53250 -79118 53330 -77768
rect 53400 -77778 53480 -77768
rect 53400 -77790 53504 -77778
rect 53400 -78566 53464 -77790
rect 53498 -78566 53504 -77790
rect 53400 -78578 53504 -78566
rect 53636 -77788 53682 -77778
rect 53636 -77790 53760 -77788
rect 53636 -78566 53642 -77790
rect 53676 -78566 53760 -77790
rect 53940 -77798 53950 -77698
rect 54032 -77728 54038 -77690
rect 54020 -77740 54038 -77728
rect 54020 -77798 54030 -77740
rect 54079 -77756 54879 -77750
rect 54079 -77790 54091 -77756
rect 54867 -77790 54879 -77756
rect 54920 -77778 54990 -77768
rect 55320 -77768 55380 -77618
rect 54079 -77796 54879 -77790
rect 53940 -77818 54030 -77798
rect 54090 -77828 54870 -77796
rect 55320 -77802 55334 -77768
rect 55368 -77802 55380 -77768
rect 55320 -77808 55380 -77802
rect 53840 -78128 53920 -78118
rect 53840 -78238 53860 -78128
rect 53840 -78248 53920 -78238
rect 53840 -78440 53900 -78248
rect 54320 -78328 54510 -77828
rect 55440 -77838 55520 -77558
rect 55410 -77840 55520 -77838
rect 55284 -77848 55330 -77840
rect 55230 -77852 55330 -77848
rect 55230 -77858 55290 -77852
rect 55324 -78028 55330 -77852
rect 55230 -78038 55330 -78028
rect 55284 -78040 55330 -78038
rect 55372 -77848 55520 -77840
rect 55372 -77852 55430 -77848
rect 55372 -78028 55378 -77852
rect 55412 -78018 55430 -77852
rect 55510 -78018 55520 -77848
rect 55412 -78028 55520 -78018
rect 55372 -78040 55418 -78028
rect 55580 -78128 55720 -76840
rect 58776 -77070 59306 -76950
rect 58776 -77080 58966 -77070
rect 56146 -77180 57366 -77130
rect 55954 -77328 56046 -77316
rect 56146 -77328 56506 -77180
rect 55954 -77498 55960 -77328
rect 56040 -77498 56046 -77328
rect 55954 -77510 56046 -77498
rect 56120 -77358 56506 -77328
rect 56120 -77568 56190 -77358
rect 56390 -77430 56506 -77358
rect 57016 -77334 57366 -77180
rect 57586 -77230 58966 -77080
rect 59126 -77230 59306 -77070
rect 57586 -77250 59306 -77230
rect 59946 -77100 60386 -77000
rect 57586 -77280 58986 -77250
rect 59946 -77260 59956 -77100
rect 60166 -77260 60386 -77100
rect 57016 -77430 57368 -77334
rect 56390 -77470 57368 -77430
rect 56390 -77568 57126 -77470
rect 56120 -77574 57126 -77568
rect 56120 -77578 56750 -77574
rect 55880 -77618 55970 -77608
rect 55870 -77696 55880 -77650
rect 55970 -77696 55982 -77650
rect 55880 -77708 55970 -77698
rect 55000 -78138 55090 -78128
rect 55000 -78248 55090 -78238
rect 54710 -78328 54960 -78308
rect 53940 -78368 54960 -78328
rect 53940 -78372 54730 -78368
rect 53930 -78378 54730 -78372
rect 53930 -78412 53942 -78378
rect 54718 -78412 54730 -78378
rect 53930 -78418 54730 -78412
rect 53840 -78528 53858 -78440
rect 53892 -78528 53900 -78440
rect 53840 -78548 53900 -78528
rect 54762 -78438 54850 -78428
rect 54762 -78440 54770 -78438
rect 54762 -78528 54768 -78440
rect 54840 -78528 54850 -78438
rect 54762 -78540 54850 -78528
rect 54770 -78548 54850 -78540
rect 53636 -78578 53760 -78566
rect 53400 -78796 53480 -78578
rect 53514 -78616 53626 -78610
rect 53514 -78618 53526 -78616
rect 53510 -78650 53526 -78618
rect 53614 -78618 53626 -78616
rect 53614 -78650 53630 -78618
rect 53510 -78724 53630 -78650
rect 53510 -78758 53526 -78724
rect 53614 -78758 53630 -78724
rect 53680 -78638 53760 -78578
rect 53930 -78556 54730 -78550
rect 53930 -78590 53942 -78556
rect 54718 -78590 54730 -78556
rect 53930 -78596 54730 -78590
rect 53940 -78628 54720 -78596
rect 53920 -78638 54720 -78628
rect 53680 -78728 54720 -78638
rect 53514 -78764 53626 -78758
rect 53680 -78796 53760 -78728
rect 53920 -78738 54720 -78728
rect 53940 -78778 54720 -78738
rect 54900 -78768 54960 -78368
rect 55010 -78360 55090 -78248
rect 55540 -78138 55720 -78128
rect 55630 -78238 55720 -78138
rect 55130 -78274 55506 -78268
rect 55130 -78308 55142 -78274
rect 55494 -78308 55506 -78274
rect 55130 -78314 55506 -78308
rect 55010 -78394 55046 -78360
rect 55080 -78394 55090 -78360
rect 55010 -78408 55090 -78394
rect 55142 -78440 55494 -78314
rect 55540 -78360 55720 -78238
rect 55540 -78394 55556 -78360
rect 55590 -78394 55720 -78360
rect 55540 -78408 55720 -78394
rect 55780 -77740 55860 -77728
rect 55130 -78446 55506 -78440
rect 55130 -78480 55142 -78446
rect 55494 -78478 55506 -78446
rect 55494 -78480 55510 -78478
rect 55130 -78486 55510 -78480
rect 55140 -78498 55510 -78486
rect 55780 -78498 55820 -77740
rect 55140 -78516 55820 -78498
rect 55854 -78516 55860 -77740
rect 55140 -78528 55860 -78516
rect 55992 -77740 56038 -77728
rect 55992 -78516 55998 -77740
rect 56032 -77748 56038 -77740
rect 56120 -77748 56300 -77578
rect 57098 -77600 57126 -77574
rect 57356 -77600 57368 -77470
rect 56032 -78106 56300 -77748
rect 56580 -77868 57066 -77610
rect 57098 -77614 57368 -77600
rect 57096 -77645 57372 -77614
rect 57096 -77679 57125 -77645
rect 57159 -77679 57217 -77645
rect 57251 -77679 57309 -77645
rect 57343 -77679 57372 -77645
rect 57096 -77710 57372 -77679
rect 56580 -77892 56590 -77868
rect 56660 -77892 57066 -77868
rect 56660 -77934 57000 -77892
rect 57586 -77930 57706 -77280
rect 59946 -77290 60386 -77260
rect 57366 -77934 57706 -77930
rect 56660 -77938 57188 -77934
rect 56660 -77944 57190 -77938
rect 56660 -77994 57118 -77944
rect 57178 -77994 57190 -77944
rect 57314 -77940 57706 -77934
rect 57314 -77980 57326 -77940
rect 57366 -77980 57706 -77940
rect 57314 -77986 57706 -77980
rect 57366 -77990 57706 -77986
rect 58896 -77570 58986 -77550
rect 58896 -77630 58906 -77570
rect 58896 -77920 58926 -77630
rect 58966 -77920 58986 -77570
rect 59106 -77570 59516 -77560
rect 59106 -77630 59216 -77570
rect 59276 -77630 59326 -77570
rect 59386 -77630 59436 -77570
rect 59496 -77630 59516 -77570
rect 59106 -77647 59516 -77630
rect 59626 -77570 59706 -77530
rect 59626 -77630 59636 -77570
rect 59626 -77640 59656 -77630
rect 59106 -77680 59125 -77647
rect 59113 -77681 59125 -77680
rect 59501 -77680 59516 -77647
rect 59501 -77681 59513 -77680
rect 59113 -77687 59513 -77681
rect 59546 -77690 59616 -77680
rect 59276 -77730 59356 -77720
rect 59276 -77749 59286 -77730
rect 59113 -77755 59286 -77749
rect 59346 -77749 59356 -77730
rect 59346 -77755 59513 -77749
rect 59113 -77789 59125 -77755
rect 59501 -77789 59513 -77755
rect 59606 -77750 59616 -77690
rect 59546 -77760 59616 -77750
rect 59113 -77790 59286 -77789
rect 59346 -77790 59513 -77789
rect 59016 -77800 59076 -77790
rect 59113 -77795 59513 -77790
rect 59276 -77800 59356 -77795
rect 59546 -77810 59616 -77800
rect 59016 -77870 59076 -77860
rect 59113 -77863 59513 -77857
rect 59113 -77897 59125 -77863
rect 59501 -77897 59513 -77863
rect 59606 -77870 59616 -77810
rect 59546 -77880 59616 -77870
rect 59113 -77900 59513 -77897
rect 59113 -77903 59516 -77900
rect 58896 -77930 58986 -77920
rect 58896 -77990 58906 -77930
rect 58966 -77990 58986 -77930
rect 58896 -77992 58986 -77990
rect 59116 -77920 59516 -77903
rect 59646 -77910 59656 -77640
rect 59116 -77980 59216 -77920
rect 59276 -77980 59336 -77920
rect 59396 -77980 59436 -77920
rect 59496 -77980 59516 -77920
rect 56660 -77998 57190 -77994
rect 56590 -78000 57190 -77998
rect 56590 -78004 57188 -78000
rect 56590 -78068 57000 -78004
rect 56032 -78118 56356 -78106
rect 56032 -78516 56280 -78118
rect 55992 -78528 56280 -78516
rect 55140 -78538 55200 -78528
rect 55450 -78558 55810 -78528
rect 55870 -78566 55982 -78560
rect 55870 -78600 55882 -78566
rect 55970 -78600 55982 -78566
rect 55870 -78606 55982 -78600
rect 55140 -78618 55200 -78608
rect 55024 -78648 55116 -78636
rect 55024 -78728 55030 -78648
rect 55110 -78728 55116 -78648
rect 55024 -78740 55116 -78728
rect 55734 -78648 55816 -78636
rect 55734 -78728 55740 -78648
rect 55810 -78728 55816 -78648
rect 55734 -78740 55816 -78728
rect 55880 -78638 55970 -78606
rect 55880 -78764 55970 -78728
rect 56060 -78748 56280 -78528
rect 56350 -78748 56356 -78118
rect 56480 -78188 56550 -78178
rect 56480 -78258 56550 -78248
rect 56590 -78287 56750 -78068
rect 58894 -78086 58988 -77992
rect 59116 -78000 59516 -77980
rect 59636 -77920 59656 -77910
rect 59696 -77920 59706 -77570
rect 59856 -77740 59976 -77730
rect 59856 -77830 59866 -77740
rect 59966 -77830 59976 -77740
rect 59856 -77840 59976 -77830
rect 60436 -77820 60446 -77720
rect 60526 -77820 60536 -77720
rect 60436 -77840 60536 -77820
rect 59636 -77930 59706 -77920
rect 59696 -77990 59706 -77930
rect 59636 -78010 59706 -77990
rect 59756 -77860 60536 -77840
rect 59756 -77900 59866 -77860
rect 60426 -77900 60536 -77860
rect 59756 -77910 60536 -77900
rect 59756 -77950 59826 -77910
rect 59066 -78040 59176 -78030
rect 58896 -78150 58986 -78086
rect 59066 -78110 59076 -78040
rect 59166 -78110 59176 -78040
rect 59066 -78112 59103 -78110
rect 59137 -78112 59176 -78110
rect 59066 -78120 59176 -78112
rect 59756 -78140 59766 -77950
rect 59806 -78140 59826 -77950
rect 59956 -77968 60046 -77940
rect 59946 -77974 60046 -77968
rect 60126 -77968 60336 -77940
rect 60126 -77974 60346 -77968
rect 59856 -78010 59916 -78000
rect 59946 -78008 59958 -77974
rect 60334 -78008 60346 -77974
rect 59946 -78014 60346 -78008
rect 60376 -78020 60446 -78010
rect 59856 -78090 59916 -78080
rect 59946 -78082 60346 -78076
rect 59946 -78116 59958 -78082
rect 60334 -78116 60346 -78082
rect 60376 -78090 60446 -78080
rect 59946 -78122 59976 -78116
rect 57098 -78158 57368 -78154
rect 57096 -78164 57372 -78158
rect 57096 -78250 57098 -78164
rect 56424 -78288 56470 -78287
rect 56060 -78760 56356 -78748
rect 56410 -78299 56470 -78288
rect 53400 -78808 53504 -78796
rect 53400 -79118 53464 -78808
rect 53250 -79508 53464 -79118
rect 53000 -79584 53464 -79508
rect 53498 -79584 53504 -78808
rect 53000 -79588 53504 -79584
rect 53458 -79596 53504 -79588
rect 53636 -78808 53760 -78796
rect 53636 -79584 53642 -78808
rect 53676 -79584 53760 -78808
rect 53930 -78784 54730 -78778
rect 53930 -78818 53942 -78784
rect 54718 -78818 54730 -78784
rect 53930 -78824 54730 -78818
rect 53830 -78846 53900 -78828
rect 53830 -78934 53858 -78846
rect 53892 -78934 53900 -78846
rect 53830 -79128 53900 -78934
rect 54760 -78846 54850 -78828
rect 54760 -78934 54768 -78846
rect 54802 -78848 54850 -78846
rect 54900 -78838 55200 -78768
rect 55870 -78770 55982 -78764
rect 55870 -78804 55882 -78770
rect 55970 -78804 55982 -78770
rect 55450 -78838 55810 -78808
rect 55870 -78810 55982 -78804
rect 56060 -78838 56300 -78760
rect 54900 -78842 55820 -78838
rect 56000 -78842 56300 -78838
rect 54900 -78848 55860 -78842
rect 54840 -78928 54850 -78848
rect 54802 -78934 54850 -78928
rect 54760 -78948 54850 -78934
rect 55130 -78854 55860 -78848
rect 55130 -78878 55820 -78854
rect 55130 -78896 55510 -78878
rect 55130 -78930 55142 -78896
rect 55494 -78898 55510 -78896
rect 55494 -78930 55506 -78898
rect 55130 -78936 55506 -78930
rect 53930 -78962 54730 -78956
rect 53930 -78996 53942 -78962
rect 54718 -78996 54730 -78962
rect 55020 -78982 55090 -78968
rect 53930 -79002 54730 -78996
rect 53940 -79008 54730 -79002
rect 54920 -78998 54980 -78988
rect 53940 -79048 54920 -79008
rect 53830 -79138 53920 -79128
rect 53830 -79248 53850 -79138
rect 53830 -79258 53920 -79248
rect 54320 -79548 54510 -79048
rect 54710 -79068 54920 -79048
rect 54910 -79078 54980 -79068
rect 55020 -79016 55046 -78982
rect 55080 -79016 55090 -78982
rect 55020 -79128 55090 -79016
rect 55142 -79062 55494 -78936
rect 55540 -78982 55620 -78968
rect 55540 -79016 55556 -78982
rect 55590 -79016 55620 -78982
rect 55130 -79068 55506 -79062
rect 55130 -79102 55142 -79068
rect 55494 -79102 55506 -79068
rect 55130 -79108 55506 -79102
rect 55000 -79138 55090 -79128
rect 55000 -79248 55090 -79238
rect 55540 -79128 55620 -79016
rect 55540 -79138 55630 -79128
rect 55630 -79238 55680 -79148
rect 55540 -79248 55680 -79238
rect 55274 -79338 55320 -79336
rect 55220 -79348 55320 -79338
rect 55220 -79524 55280 -79518
rect 55314 -79524 55320 -79348
rect 55220 -79528 55320 -79524
rect 55274 -79536 55320 -79528
rect 55362 -79348 55408 -79336
rect 55362 -79524 55368 -79348
rect 55402 -79358 55510 -79348
rect 55402 -79524 55410 -79358
rect 55362 -79528 55410 -79524
rect 55500 -79528 55510 -79358
rect 55362 -79536 55510 -79528
rect 55390 -79538 55510 -79536
rect 53636 -79588 53760 -79584
rect 53636 -79596 53682 -79588
rect 53940 -79608 54020 -79568
rect 54080 -79582 54860 -79548
rect 55311 -79574 55371 -79568
rect 53514 -79634 53626 -79628
rect 53514 -79638 53526 -79634
rect 53510 -79668 53526 -79638
rect 53614 -79638 53626 -79634
rect 53614 -79668 53630 -79638
rect 53510 -79728 53630 -79668
rect 53940 -79688 53950 -79608
rect 54010 -79638 54020 -79608
rect 54069 -79588 54869 -79582
rect 54069 -79622 54081 -79588
rect 54857 -79622 54869 -79588
rect 54069 -79628 54869 -79622
rect 54910 -79598 54980 -79588
rect 54010 -79650 54028 -79638
rect 54022 -79688 54028 -79650
rect 53940 -79700 54028 -79688
rect 53940 -79708 54020 -79700
rect 54910 -79708 54980 -79698
rect 55311 -79608 55324 -79574
rect 55358 -79608 55371 -79574
rect 54070 -79710 54870 -79708
rect 54069 -79716 54870 -79710
rect 54069 -79738 54081 -79716
rect 54041 -79750 54081 -79738
rect 54857 -79718 54870 -79716
rect 54857 -79750 54880 -79718
rect 55311 -79748 55371 -79608
rect 54041 -79758 54880 -79750
rect 55240 -79758 55371 -79748
rect 54041 -79768 55240 -79758
rect 53510 -79858 53630 -79848
rect 53961 -79808 55240 -79768
rect 53961 -80006 54031 -79808
rect 54730 -79868 54860 -79858
rect 54730 -79888 54740 -79868
rect 54080 -79938 54740 -79888
rect 54069 -79944 54740 -79938
rect 54850 -79938 54860 -79868
rect 54850 -79944 54869 -79938
rect 54069 -79978 54081 -79944
rect 54857 -79978 54869 -79944
rect 54069 -79984 54869 -79978
rect 54911 -79994 54981 -79808
rect 55370 -79808 55371 -79758
rect 55240 -79828 55370 -79818
rect 55410 -79848 55510 -79538
rect 55410 -79958 55510 -79938
rect 55570 -79868 55680 -79248
rect 55780 -79630 55820 -78878
rect 55854 -79630 55860 -78854
rect 55780 -79638 55860 -79630
rect 55814 -79642 55860 -79638
rect 55992 -78854 56300 -78842
rect 55992 -79630 55998 -78854
rect 56032 -79628 56300 -78854
rect 56410 -78898 56430 -78299
rect 56380 -79075 56430 -78898
rect 56464 -79075 56470 -78299
rect 56380 -79087 56470 -79075
rect 56552 -78299 56750 -78287
rect 56552 -79075 56558 -78299
rect 56592 -78438 56750 -78299
rect 57066 -78280 57098 -78250
rect 57368 -78250 57372 -78164
rect 58896 -78159 59076 -78150
rect 58896 -78160 59084 -78159
rect 59156 -78160 59202 -78159
rect 57368 -78280 57396 -78250
rect 57066 -78410 57086 -78280
rect 57376 -78410 57396 -78280
rect 56592 -79075 56610 -78438
rect 57066 -78440 57396 -78410
rect 56860 -78590 57060 -78578
rect 56860 -78618 57236 -78590
rect 56860 -78748 56900 -78618
rect 57020 -78748 57236 -78618
rect 56860 -78788 57236 -78748
rect 57036 -78790 57236 -78788
rect 58556 -78680 58756 -78660
rect 58556 -78840 58576 -78680
rect 58736 -78840 58756 -78680
rect 58556 -78860 58756 -78840
rect 56552 -79078 56610 -79075
rect 57036 -78940 57446 -78930
rect 56552 -79087 56598 -79078
rect 57036 -79080 57056 -78940
rect 57416 -79080 57446 -78940
rect 56380 -79358 56440 -79087
rect 57036 -79100 57098 -79080
rect 56480 -79128 56550 -79118
rect 56480 -79198 56550 -79188
rect 57096 -79214 57098 -79134
rect 57368 -79100 57446 -79080
rect 57368 -79214 57372 -79134
rect 57096 -79230 57372 -79214
rect 58896 -79290 58926 -78160
rect 58966 -78171 59086 -78160
rect 58966 -78547 59044 -78171
rect 59078 -78547 59086 -78171
rect 58966 -78570 59086 -78547
rect 59156 -78171 59256 -78160
rect 59756 -78170 59826 -78140
rect 59966 -78152 59976 -78122
rect 60316 -78122 60346 -78116
rect 61036 -78120 61466 -78110
rect 60316 -78152 60326 -78122
rect 59966 -78160 60326 -78152
rect 59156 -78547 59162 -78171
rect 59196 -78240 59256 -78171
rect 59236 -78320 59256 -78240
rect 59196 -78440 59256 -78320
rect 59236 -78520 59256 -78440
rect 59196 -78547 59256 -78520
rect 59156 -78560 59256 -78547
rect 58966 -78880 59036 -78570
rect 59066 -78606 59176 -78600
rect 59066 -78610 59103 -78606
rect 59137 -78610 59176 -78606
rect 59066 -78680 59076 -78610
rect 59166 -78680 59176 -78610
rect 59066 -78690 59176 -78680
rect 59206 -78760 59256 -78560
rect 59376 -78190 59826 -78170
rect 59376 -78230 59476 -78190
rect 59656 -78230 59826 -78190
rect 59376 -78240 59826 -78230
rect 59376 -78290 59436 -78240
rect 59376 -78650 59386 -78290
rect 59426 -78650 59436 -78290
rect 59526 -78298 59576 -78270
rect 59526 -78332 59546 -78298
rect 59636 -78330 59706 -78270
rect 59580 -78332 59706 -78330
rect 59526 -78340 59706 -78332
rect 59476 -78382 59546 -78370
rect 59476 -78450 59502 -78382
rect 59476 -78558 59502 -78520
rect 59536 -78558 59546 -78382
rect 59476 -78570 59546 -78558
rect 59576 -78382 59636 -78370
rect 59576 -78390 59590 -78382
rect 59624 -78390 59636 -78382
rect 59576 -78570 59636 -78560
rect 59534 -78608 59592 -78602
rect 59534 -78610 59546 -78608
rect 59066 -78770 59176 -78760
rect 59066 -78840 59076 -78770
rect 59166 -78840 59176 -78770
rect 59066 -78842 59103 -78840
rect 59137 -78842 59176 -78840
rect 59066 -78850 59176 -78842
rect 59206 -78770 59266 -78760
rect 59206 -78850 59266 -78840
rect 59376 -78800 59436 -78650
rect 59516 -78642 59546 -78610
rect 59580 -78610 59592 -78608
rect 59666 -78610 59706 -78340
rect 59580 -78642 59706 -78610
rect 59516 -78680 59706 -78642
rect 59746 -78298 59936 -78270
rect 59746 -78332 59862 -78298
rect 59896 -78332 59936 -78298
rect 59746 -78340 59936 -78332
rect 61036 -78300 61206 -78120
rect 61346 -78300 61466 -78120
rect 61036 -78340 61466 -78300
rect 59746 -78600 59776 -78340
rect 60286 -78350 60476 -78340
rect 59806 -78382 59866 -78370
rect 59806 -78400 59818 -78382
rect 59852 -78400 59866 -78382
rect 59806 -78558 59818 -78540
rect 59852 -78558 59866 -78540
rect 59806 -78570 59866 -78558
rect 59900 -78380 60016 -78370
rect 59900 -78382 59916 -78380
rect 59900 -78558 59906 -78382
rect 59900 -78560 59916 -78558
rect 60006 -78560 60016 -78380
rect 60286 -78490 60306 -78350
rect 60456 -78490 60476 -78350
rect 61176 -78400 61386 -78380
rect 60286 -78500 60476 -78490
rect 61026 -78420 61136 -78410
rect 59900 -78570 60016 -78560
rect 60076 -78557 60196 -78520
rect 60076 -78591 60127 -78557
rect 60161 -78591 60196 -78557
rect 59746 -78608 59926 -78600
rect 59746 -78610 59862 -78608
rect 59896 -78610 59926 -78608
rect 59746 -78680 59826 -78610
rect 59916 -78680 59926 -78610
rect 59746 -78690 59926 -78680
rect 60076 -78649 60196 -78591
rect 60336 -78560 60446 -78500
rect 60336 -78600 60366 -78560
rect 60406 -78600 60446 -78560
rect 60636 -78557 60816 -78520
rect 60636 -78591 60671 -78557
rect 60705 -78591 60747 -78557
rect 60781 -78591 60816 -78557
rect 60076 -78680 60127 -78649
rect 60161 -78680 60196 -78649
rect 59736 -78770 59936 -78760
rect 58966 -78901 59086 -78880
rect 58966 -79277 59044 -78901
rect 59078 -79277 59086 -78901
rect 58966 -79290 59086 -79277
rect 59156 -78890 59202 -78889
rect 59156 -78901 59236 -78890
rect 59156 -79277 59162 -78901
rect 59196 -78930 59236 -78901
rect 59226 -79010 59236 -78930
rect 59196 -79160 59236 -79010
rect 59226 -79240 59236 -79160
rect 59196 -79277 59236 -79240
rect 59376 -79170 59386 -78800
rect 59426 -79170 59436 -78800
rect 59516 -78811 59706 -78770
rect 59516 -78845 59545 -78811
rect 59579 -78845 59706 -78811
rect 59516 -78850 59706 -78845
rect 59533 -78851 59591 -78850
rect 59466 -78895 59546 -78880
rect 59586 -78883 59646 -78880
rect 59466 -78930 59501 -78895
rect 59466 -79071 59501 -79010
rect 59535 -79071 59546 -78895
rect 59466 -79080 59546 -79071
rect 59583 -78895 59646 -78883
rect 59583 -78910 59589 -78895
rect 59623 -78910 59646 -78895
rect 59583 -79050 59586 -78910
rect 59583 -79071 59589 -79050
rect 59623 -79071 59646 -79050
rect 59583 -79080 59646 -79071
rect 59495 -79083 59541 -79080
rect 59583 -79083 59629 -79080
rect 59533 -79120 59591 -79115
rect 59676 -79120 59706 -78850
rect 59376 -79210 59436 -79170
rect 59506 -79180 59516 -79120
rect 59596 -79180 59706 -79120
rect 59736 -78840 59826 -78770
rect 59926 -78840 59936 -78770
rect 59736 -78845 59861 -78840
rect 59895 -78845 59936 -78840
rect 59736 -78850 59936 -78845
rect 60076 -78840 60096 -78680
rect 60176 -78840 60196 -78680
rect 59736 -79120 59766 -78850
rect 59849 -78851 59907 -78850
rect 60076 -78867 60127 -78840
rect 60161 -78867 60196 -78840
rect 59796 -78883 59856 -78880
rect 59796 -78890 59857 -78883
rect 59856 -79070 59857 -78890
rect 59796 -79071 59817 -79070
rect 59851 -79071 59857 -79070
rect 59796 -79080 59857 -79071
rect 59811 -79083 59857 -79080
rect 59899 -78890 59945 -78883
rect 59899 -78895 59916 -78890
rect 59899 -79071 59905 -78895
rect 59899 -79080 59916 -79071
rect 60006 -79080 60016 -78890
rect 60076 -78925 60196 -78867
rect 60346 -78650 60426 -78600
rect 60346 -78690 60366 -78650
rect 60406 -78690 60426 -78650
rect 60346 -78740 60426 -78690
rect 60346 -78780 60366 -78740
rect 60406 -78780 60426 -78740
rect 60346 -78820 60426 -78780
rect 60346 -78860 60366 -78820
rect 60406 -78860 60426 -78820
rect 60346 -78870 60426 -78860
rect 60636 -78649 60816 -78591
rect 60636 -78683 60671 -78649
rect 60705 -78683 60747 -78649
rect 60781 -78683 60816 -78649
rect 60636 -78741 60816 -78683
rect 60636 -78775 60671 -78741
rect 60705 -78775 60747 -78741
rect 60781 -78775 60816 -78741
rect 60636 -78833 60816 -78775
rect 60636 -78867 60671 -78833
rect 60705 -78867 60747 -78833
rect 60781 -78867 60816 -78833
rect 60076 -78959 60127 -78925
rect 60161 -78959 60196 -78925
rect 60076 -78990 60196 -78959
rect 60276 -78910 60546 -78900
rect 60276 -78925 60476 -78910
rect 60276 -78959 60297 -78925
rect 60331 -78959 60369 -78925
rect 60405 -78959 60449 -78925
rect 60276 -78970 60476 -78959
rect 60536 -78970 60546 -78910
rect 60276 -78980 60546 -78970
rect 60636 -78925 60816 -78867
rect 61026 -78530 61036 -78420
rect 61126 -78530 61136 -78420
rect 61176 -78480 61196 -78400
rect 61366 -78480 61386 -78400
rect 61176 -78500 61386 -78480
rect 61026 -78560 61136 -78530
rect 61026 -78600 61046 -78560
rect 61086 -78600 61136 -78560
rect 61026 -78650 61136 -78600
rect 61026 -78690 61046 -78650
rect 61086 -78690 61136 -78650
rect 61026 -78740 61136 -78690
rect 61026 -78780 61046 -78740
rect 61086 -78780 61136 -78740
rect 61026 -78820 61136 -78780
rect 61026 -78860 61046 -78820
rect 61086 -78860 61136 -78820
rect 61026 -78880 61136 -78860
rect 61256 -78557 61366 -78500
rect 61256 -78591 61291 -78557
rect 61325 -78591 61366 -78557
rect 61256 -78649 61366 -78591
rect 61256 -78650 61291 -78649
rect 61325 -78650 61366 -78649
rect 61256 -78860 61276 -78650
rect 61356 -78860 61366 -78650
rect 61256 -78867 61291 -78860
rect 61325 -78867 61366 -78860
rect 60636 -78959 60671 -78925
rect 60705 -78959 60747 -78925
rect 60781 -78959 60816 -78925
rect 60636 -79040 60816 -78959
rect 60966 -78924 61177 -78910
rect 60966 -78925 61129 -78924
rect 60966 -78959 60980 -78925
rect 61015 -78959 61053 -78925
rect 61088 -78958 61129 -78925
rect 61164 -78958 61177 -78924
rect 61088 -78959 61177 -78958
rect 60966 -78990 61177 -78959
rect 61256 -78925 61366 -78867
rect 61256 -78959 61291 -78925
rect 61325 -78959 61366 -78925
rect 61256 -78990 61366 -78959
rect 60466 -79050 60546 -79040
rect 59899 -79083 59945 -79080
rect 60466 -79110 60476 -79050
rect 60536 -79110 60546 -79050
rect 59849 -79120 59907 -79115
rect 60466 -79120 60546 -79110
rect 60606 -79050 60826 -79040
rect 60606 -79110 60616 -79050
rect 60736 -79110 60756 -79050
rect 60816 -79110 60826 -79050
rect 60606 -79120 60826 -79110
rect 60886 -79050 60966 -79040
rect 60886 -79110 60896 -79050
rect 60956 -79110 60966 -79050
rect 60886 -79120 60966 -79110
rect 59736 -79121 59926 -79120
rect 59736 -79155 59861 -79121
rect 59895 -79155 59926 -79121
rect 59736 -79180 59926 -79155
rect 60636 -79170 60816 -79120
rect 59376 -79220 59826 -79210
rect 59376 -79260 59476 -79220
rect 59646 -79260 59826 -79220
rect 59376 -79270 59826 -79260
rect 59156 -79290 59236 -79277
rect 58896 -79300 59086 -79290
rect 56380 -79368 57000 -79358
rect 57356 -79364 57676 -79350
rect 56440 -79374 57000 -79368
rect 57314 -79370 57676 -79364
rect 56440 -79394 57178 -79374
rect 56440 -79444 57118 -79394
rect 57168 -79444 57178 -79394
rect 57314 -79410 57326 -79370
rect 57376 -79410 57676 -79370
rect 57314 -79416 57676 -79410
rect 57356 -79430 57676 -79416
rect 56440 -79454 57178 -79444
rect 56440 -79488 57000 -79454
rect 57112 -79456 57174 -79454
rect 56380 -79558 57000 -79488
rect 56032 -79630 56038 -79628
rect 55992 -79642 56038 -79630
rect 55880 -79674 55970 -79668
rect 55870 -79678 55982 -79674
rect 55870 -79720 55880 -79678
rect 55970 -79720 55982 -79678
rect 55880 -79768 55970 -79758
rect 56120 -79798 56300 -79628
rect 56362 -79722 57006 -79558
rect 57096 -79709 57372 -79678
rect 57096 -79743 57125 -79709
rect 57159 -79743 57217 -79709
rect 57251 -79743 57309 -79709
rect 57343 -79720 57372 -79709
rect 57343 -79743 57376 -79720
rect 57096 -79780 57376 -79743
rect 57066 -79790 57376 -79780
rect 56426 -79798 57376 -79790
rect 56120 -79808 57376 -79798
rect 56014 -79858 56086 -79846
rect 55570 -79978 55830 -79868
rect 53961 -80044 53988 -80006
rect 54022 -80044 54031 -80006
rect 53961 -80058 54031 -80044
rect 54910 -80006 54981 -79994
rect 54910 -80044 54916 -80006
rect 54950 -80044 54981 -80006
rect 54910 -80056 54981 -80044
rect 54911 -80058 54981 -80056
rect 55220 -80018 55330 -80008
rect 54069 -80072 54869 -80066
rect 54069 -80106 54081 -80072
rect 54857 -80078 54869 -80072
rect 54857 -80106 54880 -80078
rect 54069 -80112 54880 -80106
rect 54090 -80188 54880 -80112
rect 55330 -80118 55380 -80018
rect 55330 -80128 55480 -80118
rect 55220 -80138 55480 -80128
rect 55280 -80152 55480 -80138
rect 55280 -80158 55488 -80152
rect 55280 -80178 55300 -80158
rect 54090 -80288 54150 -80188
rect 54840 -80288 54880 -80188
rect 55288 -80192 55300 -80178
rect 55476 -80192 55488 -80158
rect 55530 -80178 55610 -80168
rect 55288 -80198 55488 -80192
rect 55520 -80202 55530 -80190
rect 55520 -80236 55526 -80202
rect 55288 -80246 55488 -80240
rect 55288 -80280 55300 -80246
rect 55476 -80280 55488 -80246
rect 55520 -80248 55530 -80236
rect 55530 -80278 55610 -80268
rect 55288 -80286 55488 -80280
rect 54090 -80308 54140 -80288
rect 54100 -80548 54140 -80308
rect 54850 -80548 54880 -80288
rect 55300 -80328 55470 -80286
rect 55300 -80468 55320 -80328
rect 55470 -80414 55482 -80342
rect 55300 -80478 55470 -80468
rect 54100 -80588 54880 -80548
rect 55710 -80798 55830 -79978
rect 56014 -80008 56020 -79858
rect 56080 -80008 56086 -79858
rect 56014 -80020 56086 -80008
rect 56120 -80008 56170 -79808
rect 56390 -79860 57376 -79808
rect 56390 -79868 57156 -79860
rect 56390 -80008 56654 -79868
rect 56120 -80058 56654 -80008
rect 56306 -80086 56654 -80058
rect 56998 -80020 57156 -79868
rect 57316 -80020 57376 -79860
rect 56998 -80086 57376 -80020
rect 56306 -80500 57376 -80086
rect 57556 -80210 57676 -79430
rect 58896 -79460 58986 -79300
rect 59756 -79320 59826 -79270
rect 59066 -79336 59176 -79330
rect 59066 -79340 59103 -79336
rect 59137 -79340 59176 -79336
rect 59066 -79400 59076 -79340
rect 59166 -79400 59176 -79340
rect 59066 -79410 59176 -79400
rect 58896 -79830 58926 -79460
rect 58966 -79830 58986 -79530
rect 59116 -79460 59506 -79440
rect 59116 -79530 59146 -79460
rect 59226 -79530 59276 -79460
rect 59356 -79530 59396 -79460
rect 59476 -79530 59506 -79460
rect 59116 -79548 59506 -79530
rect 59646 -79460 59716 -79440
rect 59706 -79520 59716 -79460
rect 59646 -79530 59716 -79520
rect 59113 -79554 59513 -79548
rect 59113 -79588 59125 -79554
rect 59501 -79588 59513 -79554
rect 59113 -79594 59513 -79588
rect 59546 -79600 59616 -79590
rect 59246 -79656 59256 -79630
rect 59113 -79662 59256 -79656
rect 59366 -79656 59376 -79630
rect 59366 -79662 59513 -79656
rect 59016 -79700 59076 -79680
rect 59113 -79696 59125 -79662
rect 59501 -79696 59513 -79662
rect 59606 -79660 59616 -79600
rect 59546 -79670 59616 -79660
rect 59113 -79702 59513 -79696
rect 59016 -79790 59076 -79760
rect 59113 -79770 59513 -79764
rect 59113 -79804 59125 -79770
rect 59501 -79804 59513 -79770
rect 59113 -79810 59513 -79804
rect 58896 -79900 58906 -79830
rect 58896 -79920 58986 -79900
rect 59116 -79830 59516 -79810
rect 59116 -79900 59146 -79830
rect 59226 -79900 59276 -79830
rect 59356 -79900 59396 -79830
rect 59476 -79900 59516 -79830
rect 59116 -79920 59516 -79900
rect 59646 -79830 59656 -79530
rect 59706 -79830 59716 -79530
rect 59756 -79500 59766 -79320
rect 59806 -79500 59826 -79320
rect 59956 -79320 60336 -79310
rect 59956 -79334 59966 -79320
rect 59946 -79340 59966 -79334
rect 60326 -79334 60336 -79320
rect 60326 -79340 60346 -79334
rect 59856 -79380 59916 -79370
rect 59946 -79374 59958 -79340
rect 60334 -79374 60346 -79340
rect 61056 -79340 61176 -78990
rect 59946 -79380 59966 -79374
rect 60326 -79380 60346 -79374
rect 60376 -79380 60436 -79360
rect 59956 -79390 60336 -79380
rect 59856 -79460 59916 -79440
rect 59946 -79448 60346 -79442
rect 59756 -79540 59826 -79500
rect 59946 -79482 59958 -79448
rect 60334 -79482 60346 -79448
rect 60376 -79460 60436 -79440
rect 61126 -79440 61176 -79340
rect 61056 -79470 61176 -79440
rect 59946 -79488 60346 -79482
rect 59946 -79540 60336 -79488
rect 59756 -79560 60536 -79540
rect 59756 -79600 59866 -79560
rect 60426 -79600 60536 -79560
rect 59756 -79610 60536 -79600
rect 59796 -79720 59806 -79610
rect 59916 -79720 59926 -79610
rect 59796 -79730 59926 -79720
rect 60436 -79630 60536 -79610
rect 60436 -79750 60446 -79630
rect 60526 -79750 60536 -79630
rect 60436 -79760 60536 -79750
rect 59646 -79840 59716 -79830
rect 59706 -79900 59716 -79840
rect 59646 -79920 59716 -79900
rect 58806 -80210 59356 -80180
rect 57556 -80220 59356 -80210
rect 57556 -80360 58986 -80220
rect 59126 -80360 59356 -80220
rect 59846 -80190 60256 -80180
rect 59846 -80300 59996 -80190
rect 60106 -80300 60256 -80190
rect 57556 -80410 59356 -80360
rect 58806 -80490 59356 -80410
rect 55710 -80800 55910 -80798
rect 55400 -80900 56300 -80800
rect 59600 -80900 60500 -80300
rect 55400 -81300 55500 -80900
rect 56200 -81300 56300 -80900
rect 55400 -81400 56300 -81300
rect 55360 -81880 55800 -81800
rect 55360 -82160 55440 -81880
rect 55720 -82160 55800 -81880
rect 55360 -82240 55800 -82160
rect 54090 -82338 54890 -82298
rect 54090 -82468 54150 -82338
rect 53510 -82520 53800 -82518
rect 53460 -82540 53800 -82520
rect 53460 -82740 53480 -82540
rect 53780 -82740 53800 -82540
rect 54080 -82598 54150 -82468
rect 54860 -82578 54890 -82338
rect 54850 -82598 54890 -82578
rect 54080 -82666 54880 -82598
rect 54079 -82672 54880 -82666
rect 54079 -82706 54091 -82672
rect 54867 -82698 54880 -82672
rect 54867 -82706 54879 -82698
rect 54079 -82712 54879 -82706
rect 53460 -82760 53800 -82740
rect 53510 -82858 53800 -82760
rect 53002 -83020 53480 -82958
rect 53000 -83158 53480 -83020
rect 53510 -82968 53520 -82858
rect 53640 -82968 53800 -82858
rect 53510 -83088 53800 -82968
rect 53970 -82734 54040 -82718
rect 53970 -82772 53998 -82734
rect 54032 -82772 54040 -82734
rect 53970 -82968 54040 -82772
rect 54920 -82734 54990 -82718
rect 54920 -82772 54926 -82734
rect 54960 -82772 54990 -82734
rect 54079 -82800 54879 -82794
rect 54079 -82834 54091 -82800
rect 54867 -82834 54879 -82800
rect 54079 -82838 54879 -82834
rect 54079 -82840 54750 -82838
rect 54090 -82888 54750 -82840
rect 54740 -82918 54750 -82888
rect 54850 -82840 54879 -82838
rect 54850 -82908 54860 -82840
rect 54840 -82918 54860 -82908
rect 54750 -82928 54860 -82918
rect 54920 -82968 54990 -82772
rect 55430 -82818 55520 -82808
rect 55290 -82928 55390 -82918
rect 53970 -82998 55290 -82968
rect 55430 -82958 55520 -82888
rect 53970 -83008 55390 -82998
rect 54050 -83018 55380 -83008
rect 54050 -83028 54880 -83018
rect 54050 -83038 54091 -83028
rect 54079 -83062 54091 -83038
rect 54867 -83038 54880 -83028
rect 54867 -83062 54879 -83038
rect 54079 -83068 54879 -83062
rect 54920 -83078 54990 -83068
rect 53510 -83106 53630 -83088
rect 53510 -83138 53526 -83106
rect 53514 -83140 53526 -83138
rect 53614 -83138 53630 -83106
rect 53940 -83090 54038 -83078
rect 53940 -83098 53998 -83090
rect 53614 -83140 53626 -83138
rect 53514 -83146 53626 -83140
rect 53000 -84908 53050 -83158
rect 53250 -83168 53480 -83158
rect 53250 -84518 53330 -83168
rect 53400 -83178 53480 -83168
rect 53400 -83190 53504 -83178
rect 53400 -83966 53464 -83190
rect 53498 -83966 53504 -83190
rect 53400 -83978 53504 -83966
rect 53636 -83188 53682 -83178
rect 53636 -83190 53760 -83188
rect 53636 -83966 53642 -83190
rect 53676 -83966 53760 -83190
rect 53940 -83198 53950 -83098
rect 54032 -83128 54038 -83090
rect 54020 -83140 54038 -83128
rect 54020 -83198 54030 -83140
rect 54079 -83156 54879 -83150
rect 54079 -83190 54091 -83156
rect 54867 -83190 54879 -83156
rect 54920 -83178 54990 -83168
rect 55320 -83168 55380 -83018
rect 54079 -83196 54879 -83190
rect 53940 -83218 54030 -83198
rect 54090 -83228 54870 -83196
rect 55320 -83202 55334 -83168
rect 55368 -83202 55380 -83168
rect 55320 -83208 55380 -83202
rect 53840 -83528 53920 -83518
rect 53840 -83638 53860 -83528
rect 53840 -83648 53920 -83638
rect 53840 -83840 53900 -83648
rect 54320 -83728 54510 -83228
rect 55440 -83238 55520 -82958
rect 55410 -83240 55520 -83238
rect 55284 -83248 55330 -83240
rect 55230 -83252 55330 -83248
rect 55230 -83258 55290 -83252
rect 55324 -83428 55330 -83252
rect 55230 -83438 55330 -83428
rect 55284 -83440 55330 -83438
rect 55372 -83248 55520 -83240
rect 55372 -83252 55430 -83248
rect 55372 -83428 55378 -83252
rect 55412 -83418 55430 -83252
rect 55510 -83418 55520 -83248
rect 55412 -83428 55520 -83418
rect 55372 -83440 55418 -83428
rect 55580 -83528 55720 -82240
rect 58776 -82470 59306 -82350
rect 58776 -82480 58966 -82470
rect 56146 -82580 57366 -82530
rect 55954 -82728 56046 -82716
rect 56146 -82728 56506 -82580
rect 55954 -82898 55960 -82728
rect 56040 -82898 56046 -82728
rect 55954 -82910 56046 -82898
rect 56120 -82758 56506 -82728
rect 56120 -82968 56190 -82758
rect 56390 -82830 56506 -82758
rect 57016 -82734 57366 -82580
rect 57586 -82630 58966 -82480
rect 59126 -82630 59306 -82470
rect 57586 -82650 59306 -82630
rect 59946 -82500 60386 -82400
rect 57586 -82680 58986 -82650
rect 59946 -82660 59956 -82500
rect 60166 -82660 60386 -82500
rect 57016 -82830 57368 -82734
rect 56390 -82870 57368 -82830
rect 56390 -82968 57126 -82870
rect 56120 -82974 57126 -82968
rect 56120 -82978 56750 -82974
rect 55880 -83018 55970 -83008
rect 55870 -83096 55880 -83050
rect 55970 -83096 55982 -83050
rect 55880 -83108 55970 -83098
rect 55000 -83538 55090 -83528
rect 55000 -83648 55090 -83638
rect 54710 -83728 54960 -83708
rect 53940 -83768 54960 -83728
rect 53940 -83772 54730 -83768
rect 53930 -83778 54730 -83772
rect 53930 -83812 53942 -83778
rect 54718 -83812 54730 -83778
rect 53930 -83818 54730 -83812
rect 53840 -83928 53858 -83840
rect 53892 -83928 53900 -83840
rect 53840 -83948 53900 -83928
rect 54762 -83838 54850 -83828
rect 54762 -83840 54770 -83838
rect 54762 -83928 54768 -83840
rect 54840 -83928 54850 -83838
rect 54762 -83940 54850 -83928
rect 54770 -83948 54850 -83940
rect 53636 -83978 53760 -83966
rect 53400 -84196 53480 -83978
rect 53514 -84016 53626 -84010
rect 53514 -84018 53526 -84016
rect 53510 -84050 53526 -84018
rect 53614 -84018 53626 -84016
rect 53614 -84050 53630 -84018
rect 53510 -84124 53630 -84050
rect 53510 -84158 53526 -84124
rect 53614 -84158 53630 -84124
rect 53680 -84038 53760 -83978
rect 53930 -83956 54730 -83950
rect 53930 -83990 53942 -83956
rect 54718 -83990 54730 -83956
rect 53930 -83996 54730 -83990
rect 53940 -84028 54720 -83996
rect 53920 -84038 54720 -84028
rect 53680 -84128 54720 -84038
rect 53514 -84164 53626 -84158
rect 53680 -84196 53760 -84128
rect 53920 -84138 54720 -84128
rect 53940 -84178 54720 -84138
rect 54900 -84168 54960 -83768
rect 55010 -83760 55090 -83648
rect 55540 -83538 55720 -83528
rect 55630 -83638 55720 -83538
rect 55130 -83674 55506 -83668
rect 55130 -83708 55142 -83674
rect 55494 -83708 55506 -83674
rect 55130 -83714 55506 -83708
rect 55010 -83794 55046 -83760
rect 55080 -83794 55090 -83760
rect 55010 -83808 55090 -83794
rect 55142 -83840 55494 -83714
rect 55540 -83760 55720 -83638
rect 55540 -83794 55556 -83760
rect 55590 -83794 55720 -83760
rect 55540 -83808 55720 -83794
rect 55780 -83140 55860 -83128
rect 55130 -83846 55506 -83840
rect 55130 -83880 55142 -83846
rect 55494 -83878 55506 -83846
rect 55494 -83880 55510 -83878
rect 55130 -83886 55510 -83880
rect 55140 -83898 55510 -83886
rect 55780 -83898 55820 -83140
rect 55140 -83916 55820 -83898
rect 55854 -83916 55860 -83140
rect 55140 -83928 55860 -83916
rect 55992 -83140 56038 -83128
rect 55992 -83916 55998 -83140
rect 56032 -83148 56038 -83140
rect 56120 -83148 56300 -82978
rect 57098 -83000 57126 -82974
rect 57356 -83000 57368 -82870
rect 57098 -83014 57368 -83000
rect 56592 -83034 57024 -83024
rect 56032 -83506 56300 -83148
rect 56584 -83258 57024 -83034
rect 57096 -83045 57372 -83014
rect 57096 -83079 57125 -83045
rect 57159 -83079 57217 -83045
rect 57251 -83079 57309 -83045
rect 57343 -83079 57372 -83045
rect 57096 -83110 57372 -83079
rect 56584 -83268 57016 -83258
rect 56660 -83334 57000 -83268
rect 57586 -83330 57706 -82680
rect 59946 -82690 60386 -82660
rect 57366 -83334 57706 -83330
rect 56660 -83338 57188 -83334
rect 56660 -83344 57190 -83338
rect 56660 -83394 57118 -83344
rect 57178 -83394 57190 -83344
rect 57314 -83340 57706 -83334
rect 57314 -83380 57326 -83340
rect 57366 -83380 57706 -83340
rect 57314 -83386 57706 -83380
rect 57366 -83390 57706 -83386
rect 58896 -82970 58986 -82950
rect 58896 -83030 58906 -82970
rect 58896 -83320 58926 -83030
rect 58966 -83320 58986 -82970
rect 59106 -82970 59516 -82960
rect 59106 -83030 59216 -82970
rect 59276 -83030 59326 -82970
rect 59386 -83030 59436 -82970
rect 59496 -83030 59516 -82970
rect 59106 -83047 59516 -83030
rect 59626 -82970 59706 -82930
rect 59626 -83030 59636 -82970
rect 59626 -83040 59656 -83030
rect 59106 -83080 59125 -83047
rect 59113 -83081 59125 -83080
rect 59501 -83080 59516 -83047
rect 59501 -83081 59513 -83080
rect 59113 -83087 59513 -83081
rect 59546 -83090 59616 -83080
rect 59276 -83130 59356 -83120
rect 59276 -83149 59286 -83130
rect 59113 -83155 59286 -83149
rect 59346 -83149 59356 -83130
rect 59346 -83155 59513 -83149
rect 59113 -83189 59125 -83155
rect 59501 -83189 59513 -83155
rect 59606 -83150 59616 -83090
rect 59546 -83160 59616 -83150
rect 59113 -83190 59286 -83189
rect 59346 -83190 59513 -83189
rect 59016 -83200 59076 -83190
rect 59113 -83195 59513 -83190
rect 59276 -83200 59356 -83195
rect 59546 -83210 59616 -83200
rect 59016 -83270 59076 -83260
rect 59113 -83263 59513 -83257
rect 59113 -83297 59125 -83263
rect 59501 -83297 59513 -83263
rect 59606 -83270 59616 -83210
rect 59546 -83280 59616 -83270
rect 59113 -83300 59513 -83297
rect 59113 -83303 59516 -83300
rect 58896 -83330 58986 -83320
rect 58896 -83390 58906 -83330
rect 58966 -83390 58986 -83330
rect 58896 -83392 58986 -83390
rect 59116 -83320 59516 -83303
rect 59646 -83310 59656 -83040
rect 59116 -83380 59216 -83320
rect 59276 -83380 59336 -83320
rect 59396 -83380 59436 -83320
rect 59496 -83380 59516 -83320
rect 56660 -83398 57190 -83394
rect 56590 -83400 57190 -83398
rect 56590 -83404 57188 -83400
rect 56590 -83468 57000 -83404
rect 56032 -83518 56356 -83506
rect 56032 -83916 56280 -83518
rect 55992 -83928 56280 -83916
rect 55140 -83938 55200 -83928
rect 55450 -83958 55810 -83928
rect 55870 -83966 55982 -83960
rect 55870 -84000 55882 -83966
rect 55970 -84000 55982 -83966
rect 55870 -84006 55982 -84000
rect 55140 -84018 55200 -84008
rect 55024 -84048 55116 -84036
rect 55024 -84128 55030 -84048
rect 55110 -84128 55116 -84048
rect 55024 -84140 55116 -84128
rect 55734 -84048 55816 -84036
rect 55734 -84128 55740 -84048
rect 55810 -84128 55816 -84048
rect 55734 -84140 55816 -84128
rect 55880 -84038 55970 -84006
rect 55880 -84164 55970 -84128
rect 56060 -84148 56280 -83928
rect 56350 -84148 56356 -83518
rect 56480 -83588 56550 -83578
rect 56480 -83658 56550 -83648
rect 56590 -83687 56750 -83468
rect 58894 -83486 58988 -83392
rect 59116 -83400 59516 -83380
rect 59636 -83320 59656 -83310
rect 59696 -83320 59706 -82970
rect 59856 -83140 59976 -83130
rect 59856 -83230 59866 -83140
rect 59966 -83230 59976 -83140
rect 59856 -83240 59976 -83230
rect 60436 -83220 60446 -83120
rect 60526 -83220 60536 -83120
rect 60436 -83240 60536 -83220
rect 59636 -83330 59706 -83320
rect 59696 -83390 59706 -83330
rect 59636 -83410 59706 -83390
rect 59756 -83260 60536 -83240
rect 59756 -83300 59866 -83260
rect 60426 -83300 60536 -83260
rect 59756 -83310 60536 -83300
rect 59756 -83350 59826 -83310
rect 59066 -83440 59176 -83430
rect 58896 -83550 58986 -83486
rect 59066 -83510 59076 -83440
rect 59166 -83510 59176 -83440
rect 59066 -83512 59103 -83510
rect 59137 -83512 59176 -83510
rect 59066 -83520 59176 -83512
rect 59756 -83540 59766 -83350
rect 59806 -83540 59826 -83350
rect 59956 -83368 60046 -83340
rect 59946 -83374 60046 -83368
rect 60126 -83368 60336 -83340
rect 60126 -83374 60346 -83368
rect 59856 -83410 59916 -83400
rect 59946 -83408 59958 -83374
rect 60334 -83408 60346 -83374
rect 59946 -83414 60346 -83408
rect 60376 -83420 60446 -83410
rect 59856 -83490 59916 -83480
rect 59946 -83482 60346 -83476
rect 59946 -83516 59958 -83482
rect 60334 -83516 60346 -83482
rect 60376 -83490 60446 -83480
rect 59946 -83522 59976 -83516
rect 57098 -83558 57368 -83554
rect 57096 -83564 57372 -83558
rect 57096 -83650 57098 -83564
rect 56424 -83688 56470 -83687
rect 56060 -84160 56356 -84148
rect 56410 -83699 56470 -83688
rect 53400 -84208 53504 -84196
rect 53400 -84518 53464 -84208
rect 53250 -84908 53464 -84518
rect 53000 -84984 53464 -84908
rect 53498 -84984 53504 -84208
rect 53000 -84988 53504 -84984
rect 53458 -84996 53504 -84988
rect 53636 -84208 53760 -84196
rect 53636 -84984 53642 -84208
rect 53676 -84984 53760 -84208
rect 53930 -84184 54730 -84178
rect 53930 -84218 53942 -84184
rect 54718 -84218 54730 -84184
rect 53930 -84224 54730 -84218
rect 53830 -84246 53900 -84228
rect 53830 -84334 53858 -84246
rect 53892 -84334 53900 -84246
rect 53830 -84528 53900 -84334
rect 54760 -84246 54850 -84228
rect 54760 -84334 54768 -84246
rect 54802 -84248 54850 -84246
rect 54900 -84238 55200 -84168
rect 55870 -84170 55982 -84164
rect 55870 -84204 55882 -84170
rect 55970 -84204 55982 -84170
rect 55450 -84238 55810 -84208
rect 55870 -84210 55982 -84204
rect 56060 -84238 56300 -84160
rect 54900 -84242 55820 -84238
rect 56000 -84242 56300 -84238
rect 54900 -84248 55860 -84242
rect 54840 -84328 54850 -84248
rect 54802 -84334 54850 -84328
rect 54760 -84348 54850 -84334
rect 55130 -84254 55860 -84248
rect 55130 -84278 55820 -84254
rect 55130 -84296 55510 -84278
rect 55130 -84330 55142 -84296
rect 55494 -84298 55510 -84296
rect 55494 -84330 55506 -84298
rect 55130 -84336 55506 -84330
rect 53930 -84362 54730 -84356
rect 53930 -84396 53942 -84362
rect 54718 -84396 54730 -84362
rect 55020 -84382 55090 -84368
rect 53930 -84402 54730 -84396
rect 53940 -84408 54730 -84402
rect 54920 -84398 54980 -84388
rect 53940 -84448 54920 -84408
rect 53830 -84538 53920 -84528
rect 53830 -84648 53850 -84538
rect 53830 -84658 53920 -84648
rect 54320 -84948 54510 -84448
rect 54710 -84468 54920 -84448
rect 54910 -84478 54980 -84468
rect 55020 -84416 55046 -84382
rect 55080 -84416 55090 -84382
rect 55020 -84528 55090 -84416
rect 55142 -84462 55494 -84336
rect 55540 -84382 55620 -84368
rect 55540 -84416 55556 -84382
rect 55590 -84416 55620 -84382
rect 55130 -84468 55506 -84462
rect 55130 -84502 55142 -84468
rect 55494 -84502 55506 -84468
rect 55130 -84508 55506 -84502
rect 55000 -84538 55090 -84528
rect 55000 -84648 55090 -84638
rect 55540 -84528 55620 -84416
rect 55540 -84538 55630 -84528
rect 55630 -84638 55680 -84548
rect 55540 -84648 55680 -84638
rect 55274 -84738 55320 -84736
rect 55220 -84748 55320 -84738
rect 55220 -84924 55280 -84918
rect 55314 -84924 55320 -84748
rect 55220 -84928 55320 -84924
rect 55274 -84936 55320 -84928
rect 55362 -84748 55408 -84736
rect 55362 -84924 55368 -84748
rect 55402 -84758 55510 -84748
rect 55402 -84924 55410 -84758
rect 55362 -84928 55410 -84924
rect 55500 -84928 55510 -84758
rect 55362 -84936 55510 -84928
rect 55390 -84938 55510 -84936
rect 53636 -84988 53760 -84984
rect 53636 -84996 53682 -84988
rect 53940 -85008 54020 -84968
rect 54080 -84982 54860 -84948
rect 55311 -84974 55371 -84968
rect 53514 -85034 53626 -85028
rect 53514 -85038 53526 -85034
rect 53510 -85068 53526 -85038
rect 53614 -85038 53626 -85034
rect 53614 -85068 53630 -85038
rect 53510 -85128 53630 -85068
rect 53940 -85088 53950 -85008
rect 54010 -85038 54020 -85008
rect 54069 -84988 54869 -84982
rect 54069 -85022 54081 -84988
rect 54857 -85022 54869 -84988
rect 54069 -85028 54869 -85022
rect 54910 -84998 54980 -84988
rect 54010 -85050 54028 -85038
rect 54022 -85088 54028 -85050
rect 53940 -85100 54028 -85088
rect 53940 -85108 54020 -85100
rect 54910 -85108 54980 -85098
rect 55311 -85008 55324 -84974
rect 55358 -85008 55371 -84974
rect 54070 -85110 54870 -85108
rect 54069 -85116 54870 -85110
rect 54069 -85138 54081 -85116
rect 54041 -85150 54081 -85138
rect 54857 -85118 54870 -85116
rect 54857 -85150 54880 -85118
rect 55311 -85148 55371 -85008
rect 54041 -85158 54880 -85150
rect 55240 -85158 55371 -85148
rect 54041 -85168 55240 -85158
rect 53510 -85258 53630 -85248
rect 53961 -85208 55240 -85168
rect 53961 -85406 54031 -85208
rect 54730 -85268 54860 -85258
rect 54730 -85288 54740 -85268
rect 54080 -85338 54740 -85288
rect 54069 -85344 54740 -85338
rect 54850 -85338 54860 -85268
rect 54850 -85344 54869 -85338
rect 54069 -85378 54081 -85344
rect 54857 -85378 54869 -85344
rect 54069 -85384 54869 -85378
rect 54911 -85394 54981 -85208
rect 55370 -85208 55371 -85158
rect 55240 -85228 55370 -85218
rect 55410 -85248 55510 -84938
rect 55410 -85358 55510 -85338
rect 55570 -85268 55680 -84648
rect 55780 -85030 55820 -84278
rect 55854 -85030 55860 -84254
rect 55780 -85038 55860 -85030
rect 55814 -85042 55860 -85038
rect 55992 -84254 56300 -84242
rect 55992 -85030 55998 -84254
rect 56032 -85028 56300 -84254
rect 56410 -84298 56430 -83699
rect 56380 -84475 56430 -84298
rect 56464 -84475 56470 -83699
rect 56380 -84487 56470 -84475
rect 56552 -83699 56750 -83687
rect 56552 -84475 56558 -83699
rect 56592 -83838 56750 -83699
rect 57066 -83680 57098 -83650
rect 57368 -83650 57372 -83564
rect 58896 -83559 59076 -83550
rect 58896 -83560 59084 -83559
rect 59156 -83560 59202 -83559
rect 57368 -83680 57396 -83650
rect 57066 -83810 57086 -83680
rect 57376 -83810 57396 -83680
rect 56592 -84475 56610 -83838
rect 57066 -83840 57396 -83810
rect 56860 -83990 57060 -83978
rect 56860 -84018 57236 -83990
rect 56860 -84148 56900 -84018
rect 57020 -84148 57236 -84018
rect 56860 -84188 57236 -84148
rect 57036 -84190 57236 -84188
rect 58556 -84080 58756 -84060
rect 58556 -84240 58576 -84080
rect 58736 -84240 58756 -84080
rect 58556 -84260 58756 -84240
rect 56552 -84478 56610 -84475
rect 57036 -84340 57446 -84330
rect 56552 -84487 56598 -84478
rect 57036 -84480 57056 -84340
rect 57416 -84480 57446 -84340
rect 56380 -84758 56440 -84487
rect 57036 -84500 57098 -84480
rect 56480 -84528 56550 -84518
rect 56480 -84598 56550 -84588
rect 57096 -84614 57098 -84534
rect 57368 -84500 57446 -84480
rect 57368 -84614 57372 -84534
rect 57096 -84630 57372 -84614
rect 58896 -84690 58926 -83560
rect 58966 -83571 59086 -83560
rect 58966 -83947 59044 -83571
rect 59078 -83947 59086 -83571
rect 58966 -83970 59086 -83947
rect 59156 -83571 59256 -83560
rect 59756 -83570 59826 -83540
rect 59966 -83552 59976 -83522
rect 60316 -83522 60346 -83516
rect 61036 -83520 61466 -83510
rect 60316 -83552 60326 -83522
rect 59966 -83560 60326 -83552
rect 59156 -83947 59162 -83571
rect 59196 -83640 59256 -83571
rect 59236 -83720 59256 -83640
rect 59196 -83840 59256 -83720
rect 59236 -83920 59256 -83840
rect 59196 -83947 59256 -83920
rect 59156 -83960 59256 -83947
rect 58966 -84280 59036 -83970
rect 59066 -84006 59176 -84000
rect 59066 -84010 59103 -84006
rect 59137 -84010 59176 -84006
rect 59066 -84080 59076 -84010
rect 59166 -84080 59176 -84010
rect 59066 -84090 59176 -84080
rect 59206 -84160 59256 -83960
rect 59376 -83590 59826 -83570
rect 59376 -83630 59476 -83590
rect 59656 -83630 59826 -83590
rect 59376 -83640 59826 -83630
rect 59376 -83690 59436 -83640
rect 59376 -84050 59386 -83690
rect 59426 -84050 59436 -83690
rect 59526 -83698 59576 -83670
rect 59526 -83732 59546 -83698
rect 59636 -83730 59706 -83670
rect 59580 -83732 59706 -83730
rect 59526 -83740 59706 -83732
rect 59476 -83782 59546 -83770
rect 59476 -83850 59502 -83782
rect 59476 -83958 59502 -83920
rect 59536 -83958 59546 -83782
rect 59476 -83970 59546 -83958
rect 59576 -83782 59636 -83770
rect 59576 -83790 59590 -83782
rect 59624 -83790 59636 -83782
rect 59576 -83970 59636 -83960
rect 59534 -84008 59592 -84002
rect 59534 -84010 59546 -84008
rect 59066 -84170 59176 -84160
rect 59066 -84240 59076 -84170
rect 59166 -84240 59176 -84170
rect 59066 -84242 59103 -84240
rect 59137 -84242 59176 -84240
rect 59066 -84250 59176 -84242
rect 59206 -84170 59266 -84160
rect 59206 -84250 59266 -84240
rect 59376 -84200 59436 -84050
rect 59516 -84042 59546 -84010
rect 59580 -84010 59592 -84008
rect 59666 -84010 59706 -83740
rect 59580 -84042 59706 -84010
rect 59516 -84080 59706 -84042
rect 59746 -83698 59936 -83670
rect 59746 -83732 59862 -83698
rect 59896 -83732 59936 -83698
rect 59746 -83740 59936 -83732
rect 61036 -83700 61206 -83520
rect 61346 -83700 61466 -83520
rect 61036 -83740 61466 -83700
rect 59746 -84000 59776 -83740
rect 60286 -83750 60476 -83740
rect 59806 -83782 59866 -83770
rect 59806 -83800 59818 -83782
rect 59852 -83800 59866 -83782
rect 59806 -83958 59818 -83940
rect 59852 -83958 59866 -83940
rect 59806 -83970 59866 -83958
rect 59900 -83780 60016 -83770
rect 59900 -83782 59916 -83780
rect 59900 -83958 59906 -83782
rect 59900 -83960 59916 -83958
rect 60006 -83960 60016 -83780
rect 60286 -83890 60306 -83750
rect 60456 -83890 60476 -83750
rect 61176 -83800 61386 -83780
rect 60286 -83900 60476 -83890
rect 61026 -83820 61136 -83810
rect 59900 -83970 60016 -83960
rect 60076 -83957 60196 -83920
rect 60076 -83991 60127 -83957
rect 60161 -83991 60196 -83957
rect 59746 -84008 59926 -84000
rect 59746 -84010 59862 -84008
rect 59896 -84010 59926 -84008
rect 59746 -84080 59826 -84010
rect 59916 -84080 59926 -84010
rect 59746 -84090 59926 -84080
rect 60076 -84049 60196 -83991
rect 60336 -83960 60446 -83900
rect 60336 -84000 60366 -83960
rect 60406 -84000 60446 -83960
rect 60636 -83957 60816 -83920
rect 60636 -83991 60671 -83957
rect 60705 -83991 60747 -83957
rect 60781 -83991 60816 -83957
rect 60076 -84080 60127 -84049
rect 60161 -84080 60196 -84049
rect 59736 -84170 59936 -84160
rect 58966 -84301 59086 -84280
rect 58966 -84677 59044 -84301
rect 59078 -84677 59086 -84301
rect 58966 -84690 59086 -84677
rect 59156 -84290 59202 -84289
rect 59156 -84301 59236 -84290
rect 59156 -84677 59162 -84301
rect 59196 -84330 59236 -84301
rect 59226 -84410 59236 -84330
rect 59196 -84560 59236 -84410
rect 59226 -84640 59236 -84560
rect 59196 -84677 59236 -84640
rect 59376 -84570 59386 -84200
rect 59426 -84570 59436 -84200
rect 59516 -84211 59706 -84170
rect 59516 -84245 59545 -84211
rect 59579 -84245 59706 -84211
rect 59516 -84250 59706 -84245
rect 59533 -84251 59591 -84250
rect 59466 -84295 59546 -84280
rect 59586 -84283 59646 -84280
rect 59466 -84330 59501 -84295
rect 59466 -84471 59501 -84410
rect 59535 -84471 59546 -84295
rect 59466 -84480 59546 -84471
rect 59583 -84295 59646 -84283
rect 59583 -84310 59589 -84295
rect 59623 -84310 59646 -84295
rect 59583 -84450 59586 -84310
rect 59583 -84471 59589 -84450
rect 59623 -84471 59646 -84450
rect 59583 -84480 59646 -84471
rect 59495 -84483 59541 -84480
rect 59583 -84483 59629 -84480
rect 59533 -84520 59591 -84515
rect 59676 -84520 59706 -84250
rect 59376 -84610 59436 -84570
rect 59506 -84580 59516 -84520
rect 59596 -84580 59706 -84520
rect 59736 -84240 59826 -84170
rect 59926 -84240 59936 -84170
rect 59736 -84245 59861 -84240
rect 59895 -84245 59936 -84240
rect 59736 -84250 59936 -84245
rect 60076 -84240 60096 -84080
rect 60176 -84240 60196 -84080
rect 59736 -84520 59766 -84250
rect 59849 -84251 59907 -84250
rect 60076 -84267 60127 -84240
rect 60161 -84267 60196 -84240
rect 59796 -84283 59856 -84280
rect 59796 -84290 59857 -84283
rect 59856 -84470 59857 -84290
rect 59796 -84471 59817 -84470
rect 59851 -84471 59857 -84470
rect 59796 -84480 59857 -84471
rect 59811 -84483 59857 -84480
rect 59899 -84290 59945 -84283
rect 59899 -84295 59916 -84290
rect 59899 -84471 59905 -84295
rect 59899 -84480 59916 -84471
rect 60006 -84480 60016 -84290
rect 60076 -84325 60196 -84267
rect 60346 -84050 60426 -84000
rect 60346 -84090 60366 -84050
rect 60406 -84090 60426 -84050
rect 60346 -84140 60426 -84090
rect 60346 -84180 60366 -84140
rect 60406 -84180 60426 -84140
rect 60346 -84220 60426 -84180
rect 60346 -84260 60366 -84220
rect 60406 -84260 60426 -84220
rect 60346 -84270 60426 -84260
rect 60636 -84049 60816 -83991
rect 60636 -84083 60671 -84049
rect 60705 -84083 60747 -84049
rect 60781 -84083 60816 -84049
rect 60636 -84141 60816 -84083
rect 60636 -84175 60671 -84141
rect 60705 -84175 60747 -84141
rect 60781 -84175 60816 -84141
rect 60636 -84233 60816 -84175
rect 60636 -84267 60671 -84233
rect 60705 -84267 60747 -84233
rect 60781 -84267 60816 -84233
rect 60076 -84359 60127 -84325
rect 60161 -84359 60196 -84325
rect 60076 -84390 60196 -84359
rect 60276 -84310 60546 -84300
rect 60276 -84325 60476 -84310
rect 60276 -84359 60297 -84325
rect 60331 -84359 60369 -84325
rect 60405 -84359 60449 -84325
rect 60276 -84370 60476 -84359
rect 60536 -84370 60546 -84310
rect 60276 -84380 60546 -84370
rect 60636 -84325 60816 -84267
rect 61026 -83930 61036 -83820
rect 61126 -83930 61136 -83820
rect 61176 -83880 61196 -83800
rect 61366 -83880 61386 -83800
rect 61176 -83900 61386 -83880
rect 61026 -83960 61136 -83930
rect 61026 -84000 61046 -83960
rect 61086 -84000 61136 -83960
rect 61026 -84050 61136 -84000
rect 61026 -84090 61046 -84050
rect 61086 -84090 61136 -84050
rect 61026 -84140 61136 -84090
rect 61026 -84180 61046 -84140
rect 61086 -84180 61136 -84140
rect 61026 -84220 61136 -84180
rect 61026 -84260 61046 -84220
rect 61086 -84260 61136 -84220
rect 61026 -84280 61136 -84260
rect 61256 -83957 61366 -83900
rect 61256 -83991 61291 -83957
rect 61325 -83991 61366 -83957
rect 61256 -84049 61366 -83991
rect 61256 -84050 61291 -84049
rect 61325 -84050 61366 -84049
rect 61256 -84260 61276 -84050
rect 61356 -84260 61366 -84050
rect 61256 -84267 61291 -84260
rect 61325 -84267 61366 -84260
rect 60636 -84359 60671 -84325
rect 60705 -84359 60747 -84325
rect 60781 -84359 60816 -84325
rect 60636 -84440 60816 -84359
rect 60966 -84324 61177 -84310
rect 60966 -84325 61129 -84324
rect 60966 -84359 60980 -84325
rect 61015 -84359 61053 -84325
rect 61088 -84358 61129 -84325
rect 61164 -84358 61177 -84324
rect 61088 -84359 61177 -84358
rect 60966 -84390 61177 -84359
rect 61256 -84325 61366 -84267
rect 61256 -84359 61291 -84325
rect 61325 -84359 61366 -84325
rect 61256 -84390 61366 -84359
rect 60466 -84450 60546 -84440
rect 59899 -84483 59945 -84480
rect 60466 -84510 60476 -84450
rect 60536 -84510 60546 -84450
rect 59849 -84520 59907 -84515
rect 60466 -84520 60546 -84510
rect 60606 -84450 60826 -84440
rect 60606 -84510 60616 -84450
rect 60736 -84510 60756 -84450
rect 60816 -84510 60826 -84450
rect 60606 -84520 60826 -84510
rect 60886 -84450 60966 -84440
rect 60886 -84510 60896 -84450
rect 60956 -84510 60966 -84450
rect 60886 -84520 60966 -84510
rect 59736 -84521 59926 -84520
rect 59736 -84555 59861 -84521
rect 59895 -84555 59926 -84521
rect 59736 -84580 59926 -84555
rect 60636 -84570 60816 -84520
rect 59376 -84620 59826 -84610
rect 59376 -84660 59476 -84620
rect 59646 -84660 59826 -84620
rect 59376 -84670 59826 -84660
rect 59156 -84690 59236 -84677
rect 58896 -84700 59086 -84690
rect 56380 -84768 57000 -84758
rect 57356 -84764 57676 -84750
rect 56440 -84774 57000 -84768
rect 57314 -84770 57676 -84764
rect 56440 -84794 57178 -84774
rect 56440 -84844 57118 -84794
rect 57168 -84844 57178 -84794
rect 57314 -84810 57326 -84770
rect 57376 -84810 57676 -84770
rect 57314 -84816 57676 -84810
rect 57356 -84830 57676 -84816
rect 56440 -84854 57178 -84844
rect 56440 -84888 57000 -84854
rect 57112 -84856 57174 -84854
rect 56380 -84958 57000 -84888
rect 56032 -85030 56038 -85028
rect 55992 -85042 56038 -85030
rect 55880 -85074 55970 -85068
rect 55870 -85078 55982 -85074
rect 55870 -85120 55880 -85078
rect 55970 -85120 55982 -85078
rect 55880 -85168 55970 -85158
rect 56120 -85198 56300 -85028
rect 56374 -85082 57010 -84958
rect 57096 -85109 57372 -85078
rect 57096 -85143 57125 -85109
rect 57159 -85143 57217 -85109
rect 57251 -85143 57309 -85109
rect 57343 -85120 57372 -85109
rect 57343 -85143 57376 -85120
rect 57096 -85180 57376 -85143
rect 57066 -85190 57376 -85180
rect 56426 -85198 57376 -85190
rect 56120 -85208 57376 -85198
rect 56014 -85258 56086 -85246
rect 55570 -85378 55830 -85268
rect 53961 -85444 53988 -85406
rect 54022 -85444 54031 -85406
rect 53961 -85458 54031 -85444
rect 54910 -85406 54981 -85394
rect 54910 -85444 54916 -85406
rect 54950 -85444 54981 -85406
rect 54910 -85456 54981 -85444
rect 54911 -85458 54981 -85456
rect 55220 -85418 55330 -85408
rect 54069 -85472 54869 -85466
rect 54069 -85506 54081 -85472
rect 54857 -85478 54869 -85472
rect 54857 -85506 54880 -85478
rect 54069 -85512 54880 -85506
rect 54090 -85588 54880 -85512
rect 55330 -85518 55380 -85418
rect 55330 -85528 55480 -85518
rect 55220 -85538 55480 -85528
rect 55280 -85552 55480 -85538
rect 55280 -85558 55488 -85552
rect 55280 -85578 55300 -85558
rect 54090 -85688 54150 -85588
rect 54840 -85688 54880 -85588
rect 55288 -85592 55300 -85578
rect 55476 -85592 55488 -85558
rect 55530 -85578 55610 -85568
rect 55288 -85598 55488 -85592
rect 55520 -85602 55530 -85590
rect 55520 -85636 55526 -85602
rect 55288 -85646 55488 -85640
rect 55288 -85680 55300 -85646
rect 55476 -85680 55488 -85646
rect 55520 -85648 55530 -85636
rect 55530 -85678 55610 -85668
rect 55288 -85686 55488 -85680
rect 54090 -85708 54140 -85688
rect 54100 -85948 54140 -85708
rect 54850 -85948 54880 -85688
rect 55300 -85728 55470 -85686
rect 55300 -85868 55320 -85728
rect 55470 -85814 55482 -85742
rect 55300 -85878 55470 -85868
rect 54100 -85988 54880 -85948
rect 55710 -86198 55830 -85378
rect 56014 -85408 56020 -85258
rect 56080 -85408 56086 -85258
rect 56014 -85420 56086 -85408
rect 56120 -85408 56170 -85208
rect 56390 -85260 57376 -85208
rect 56390 -85268 57156 -85260
rect 56390 -85408 56654 -85268
rect 56120 -85458 56654 -85408
rect 56306 -85486 56654 -85458
rect 56998 -85420 57156 -85268
rect 57316 -85420 57376 -85260
rect 56998 -85486 57376 -85420
rect 56306 -85900 57376 -85486
rect 57556 -85610 57676 -84830
rect 58896 -84860 58986 -84700
rect 59756 -84720 59826 -84670
rect 59066 -84736 59176 -84730
rect 59066 -84740 59103 -84736
rect 59137 -84740 59176 -84736
rect 59066 -84800 59076 -84740
rect 59166 -84800 59176 -84740
rect 59066 -84810 59176 -84800
rect 58896 -85230 58926 -84860
rect 58966 -85230 58986 -84930
rect 59116 -84860 59506 -84840
rect 59116 -84930 59146 -84860
rect 59226 -84930 59276 -84860
rect 59356 -84930 59396 -84860
rect 59476 -84930 59506 -84860
rect 59116 -84948 59506 -84930
rect 59646 -84860 59716 -84840
rect 59706 -84920 59716 -84860
rect 59646 -84930 59716 -84920
rect 59113 -84954 59513 -84948
rect 59113 -84988 59125 -84954
rect 59501 -84988 59513 -84954
rect 59113 -84994 59513 -84988
rect 59546 -85000 59616 -84990
rect 59246 -85056 59256 -85030
rect 59113 -85062 59256 -85056
rect 59366 -85056 59376 -85030
rect 59366 -85062 59513 -85056
rect 59016 -85100 59076 -85080
rect 59113 -85096 59125 -85062
rect 59501 -85096 59513 -85062
rect 59606 -85060 59616 -85000
rect 59546 -85070 59616 -85060
rect 59113 -85102 59513 -85096
rect 59016 -85190 59076 -85160
rect 59113 -85170 59513 -85164
rect 59113 -85204 59125 -85170
rect 59501 -85204 59513 -85170
rect 59113 -85210 59513 -85204
rect 58896 -85300 58906 -85230
rect 58896 -85320 58986 -85300
rect 59116 -85230 59516 -85210
rect 59116 -85300 59146 -85230
rect 59226 -85300 59276 -85230
rect 59356 -85300 59396 -85230
rect 59476 -85300 59516 -85230
rect 59116 -85320 59516 -85300
rect 59646 -85230 59656 -84930
rect 59706 -85230 59716 -84930
rect 59756 -84900 59766 -84720
rect 59806 -84900 59826 -84720
rect 59956 -84720 60336 -84710
rect 59956 -84734 59966 -84720
rect 59946 -84740 59966 -84734
rect 60326 -84734 60336 -84720
rect 60326 -84740 60346 -84734
rect 59856 -84780 59916 -84770
rect 59946 -84774 59958 -84740
rect 60334 -84774 60346 -84740
rect 61056 -84740 61176 -84390
rect 59946 -84780 59966 -84774
rect 60326 -84780 60346 -84774
rect 60376 -84780 60436 -84760
rect 59956 -84790 60336 -84780
rect 59856 -84860 59916 -84840
rect 59946 -84848 60346 -84842
rect 59756 -84940 59826 -84900
rect 59946 -84882 59958 -84848
rect 60334 -84882 60346 -84848
rect 60376 -84860 60436 -84840
rect 61126 -84840 61176 -84740
rect 61056 -84870 61176 -84840
rect 59946 -84888 60346 -84882
rect 59946 -84940 60336 -84888
rect 59756 -84960 60536 -84940
rect 59756 -85000 59866 -84960
rect 60426 -85000 60536 -84960
rect 59756 -85010 60536 -85000
rect 59796 -85120 59806 -85010
rect 59916 -85120 59926 -85010
rect 59796 -85130 59926 -85120
rect 60436 -85030 60536 -85010
rect 60436 -85150 60446 -85030
rect 60526 -85150 60536 -85030
rect 60436 -85160 60536 -85150
rect 59646 -85240 59716 -85230
rect 59706 -85300 59716 -85240
rect 59646 -85320 59716 -85300
rect 58806 -85610 59356 -85580
rect 57556 -85620 59356 -85610
rect 57556 -85760 58986 -85620
rect 59126 -85760 59356 -85620
rect 59846 -85590 60256 -85580
rect 59846 -85700 59996 -85590
rect 60106 -85700 60256 -85590
rect 57556 -85810 59356 -85760
rect 58806 -85890 59356 -85810
rect 55710 -86200 55910 -86198
rect 55400 -86300 56200 -86200
rect 59600 -86300 60500 -85700
rect 55400 -86600 55500 -86300
rect 56100 -86600 56200 -86300
rect 55400 -86700 56200 -86600
<< via1 >>
rect 38000 1400 41400 2800
rect 37900 -3600 41500 -400
rect 43000 1000 46400 2400
rect 43000 -1400 46400 0
rect 50900 -20 53100 820
rect 56880 -40 59080 1020
rect 55400 -1000 55700 -600
rect 53400 -1600 53700 -1400
rect 54150 -1508 54860 -1338
rect 54150 -1578 54850 -1508
rect 54850 -1578 54860 -1508
rect 53520 -1968 53640 -1858
rect 54750 -1908 54850 -1838
rect 54750 -1918 54840 -1908
rect 55430 -1888 55520 -1818
rect 55290 -1998 55390 -1928
rect 53050 -3908 53250 -2158
rect 53950 -2128 53998 -2098
rect 53998 -2128 54020 -2098
rect 53950 -2198 54020 -2128
rect 54920 -2090 54990 -2078
rect 54920 -2128 54926 -2090
rect 54926 -2128 54960 -2090
rect 54960 -2128 54990 -2090
rect 54920 -2168 54990 -2128
rect 53860 -2638 53920 -2528
rect 55230 -2428 55290 -2258
rect 55290 -2428 55320 -2258
rect 55430 -2418 55510 -2248
rect 55960 -1888 56040 -1738
rect 56190 -1968 56390 -1758
rect 56506 -1830 57016 -1580
rect 58966 -1630 59126 -1470
rect 59956 -1660 60166 -1500
rect 55880 -2056 55970 -2018
rect 55880 -2090 55882 -2056
rect 55882 -2090 55970 -2056
rect 55880 -2098 55970 -2090
rect 55000 -2638 55090 -2538
rect 54770 -2840 54840 -2838
rect 54770 -2928 54802 -2840
rect 54802 -2928 54840 -2840
rect 55540 -2638 55630 -2538
rect 56590 -2398 56660 -2268
rect 58906 -2020 58966 -1970
rect 58906 -2030 58926 -2020
rect 58926 -2030 58966 -2020
rect 59216 -2030 59276 -1970
rect 59326 -2030 59386 -1970
rect 59436 -2030 59496 -1970
rect 59636 -2030 59696 -1970
rect 59546 -2101 59606 -2090
rect 59286 -2155 59346 -2130
rect 59546 -2135 59560 -2101
rect 59560 -2135 59594 -2101
rect 59594 -2135 59606 -2101
rect 59286 -2189 59346 -2155
rect 59546 -2150 59606 -2135
rect 59286 -2190 59346 -2189
rect 59016 -2209 59076 -2200
rect 59016 -2243 59032 -2209
rect 59032 -2243 59066 -2209
rect 59066 -2243 59076 -2209
rect 59016 -2260 59076 -2243
rect 59546 -2270 59606 -2210
rect 58906 -2390 58966 -2330
rect 59216 -2380 59276 -2320
rect 59336 -2380 59396 -2320
rect 59436 -2380 59496 -2320
rect 55140 -3008 55200 -2938
rect 55030 -3128 55110 -3048
rect 55740 -3128 55810 -3048
rect 55880 -3128 55970 -3038
rect 56480 -2606 56550 -2588
rect 56480 -2640 56492 -2606
rect 56492 -2640 56530 -2606
rect 56530 -2640 56550 -2606
rect 56480 -2648 56550 -2640
rect 59866 -2230 59966 -2140
rect 60446 -2220 60526 -2120
rect 59636 -2390 59696 -2330
rect 59076 -2478 59166 -2440
rect 59076 -2510 59103 -2478
rect 59103 -2510 59137 -2478
rect 59137 -2510 59166 -2478
rect 60046 -2374 60126 -2340
rect 59856 -2428 59916 -2410
rect 60046 -2400 60126 -2374
rect 59856 -2462 59874 -2428
rect 59874 -2462 59908 -2428
rect 59908 -2462 59916 -2428
rect 59856 -2480 59916 -2462
rect 60376 -2428 60446 -2420
rect 60376 -2462 60384 -2428
rect 60384 -2462 60418 -2428
rect 60418 -2462 60446 -2428
rect 59976 -2516 60316 -2500
rect 60376 -2480 60446 -2462
rect 57098 -2589 57368 -2564
rect 57098 -2623 57125 -2589
rect 57125 -2623 57159 -2589
rect 57159 -2623 57217 -2589
rect 57217 -2623 57251 -2589
rect 57251 -2623 57309 -2589
rect 57309 -2623 57343 -2589
rect 57343 -2623 57368 -2589
rect 54770 -3328 54802 -3248
rect 54802 -3328 54840 -3248
rect 53850 -3648 53920 -3538
rect 54920 -3468 54980 -3398
rect 55000 -3638 55090 -3538
rect 55540 -3638 55630 -3538
rect 55220 -3918 55280 -3748
rect 55280 -3918 55310 -3748
rect 55410 -3928 55500 -3758
rect 53950 -4050 54010 -4008
rect 53950 -4088 53988 -4050
rect 53988 -4088 54010 -4050
rect 54910 -4050 54980 -3998
rect 54910 -4088 54916 -4050
rect 54916 -4088 54950 -4050
rect 54950 -4088 54980 -4050
rect 54910 -4098 54980 -4088
rect 53510 -4248 53630 -4128
rect 54740 -4344 54850 -4268
rect 54740 -4358 54850 -4344
rect 55240 -4218 55370 -4158
rect 55410 -4338 55510 -4248
rect 57098 -2680 57368 -2623
rect 57098 -2704 57368 -2680
rect 56900 -3148 57020 -3018
rect 58576 -3240 58736 -3080
rect 57098 -3480 57368 -3474
rect 56480 -3534 56550 -3528
rect 56480 -3568 56492 -3534
rect 56492 -3568 56530 -3534
rect 56530 -3568 56550 -3534
rect 56480 -3588 56550 -3568
rect 57098 -3565 57368 -3480
rect 57098 -3599 57125 -3565
rect 57125 -3599 57159 -3565
rect 57159 -3599 57217 -3565
rect 57217 -3599 57251 -3565
rect 57251 -3599 57309 -3565
rect 57309 -3599 57343 -3565
rect 57343 -3599 57368 -3565
rect 57098 -3614 57368 -3599
rect 59976 -2552 60316 -2516
rect 59176 -2720 59196 -2640
rect 59196 -2720 59236 -2640
rect 59176 -2920 59196 -2840
rect 59196 -2920 59236 -2840
rect 59076 -3040 59103 -3010
rect 59103 -3040 59137 -3010
rect 59137 -3040 59166 -3010
rect 59076 -3080 59166 -3040
rect 59576 -2698 59636 -2670
rect 59576 -2730 59580 -2698
rect 59580 -2730 59636 -2698
rect 59476 -2920 59502 -2850
rect 59502 -2920 59536 -2850
rect 59576 -2958 59590 -2790
rect 59590 -2958 59624 -2790
rect 59624 -2958 59636 -2790
rect 59576 -2960 59636 -2958
rect 59076 -3208 59166 -3170
rect 59076 -3240 59103 -3208
rect 59103 -3240 59137 -3208
rect 59137 -3240 59166 -3208
rect 59206 -3240 59266 -3170
rect 61206 -2700 61346 -2520
rect 59806 -2940 59818 -2800
rect 59818 -2940 59852 -2800
rect 59852 -2940 59866 -2800
rect 59916 -2782 60006 -2780
rect 59916 -2958 59940 -2782
rect 59940 -2958 60006 -2782
rect 59916 -2960 60006 -2958
rect 60306 -2890 60456 -2750
rect 59826 -3042 59862 -3010
rect 59862 -3042 59896 -3010
rect 59896 -3042 59916 -3010
rect 59826 -3080 59916 -3042
rect 59166 -3410 59196 -3330
rect 59196 -3410 59226 -3330
rect 59166 -3640 59196 -3560
rect 59196 -3640 59226 -3560
rect 59466 -3410 59501 -3330
rect 59501 -3410 59526 -3330
rect 59586 -3450 59589 -3310
rect 59589 -3450 59623 -3310
rect 59623 -3450 59646 -3310
rect 59516 -3521 59596 -3520
rect 59516 -3555 59545 -3521
rect 59545 -3555 59579 -3521
rect 59579 -3555 59596 -3521
rect 59516 -3580 59596 -3555
rect 59826 -3211 59926 -3170
rect 59826 -3240 59861 -3211
rect 59861 -3240 59895 -3211
rect 59895 -3240 59926 -3211
rect 60096 -3083 60127 -3080
rect 60127 -3083 60161 -3080
rect 60161 -3083 60176 -3080
rect 60096 -3141 60176 -3083
rect 60096 -3175 60127 -3141
rect 60127 -3175 60161 -3141
rect 60161 -3175 60176 -3141
rect 60096 -3233 60176 -3175
rect 60096 -3240 60127 -3233
rect 60127 -3240 60161 -3233
rect 60161 -3240 60176 -3233
rect 59796 -3295 59856 -3290
rect 59796 -3470 59817 -3295
rect 59817 -3470 59851 -3295
rect 59851 -3470 59856 -3295
rect 59916 -3295 60006 -3290
rect 59916 -3471 59939 -3295
rect 59939 -3471 60006 -3295
rect 59916 -3480 60006 -3471
rect 60476 -3325 60536 -3310
rect 60476 -3359 60484 -3325
rect 60484 -3359 60536 -3325
rect 60476 -3370 60536 -3359
rect 61036 -2930 61126 -2820
rect 61276 -3083 61291 -3050
rect 61291 -3083 61325 -3050
rect 61325 -3083 61356 -3050
rect 61276 -3141 61356 -3083
rect 61276 -3175 61291 -3141
rect 61291 -3175 61325 -3141
rect 61325 -3175 61356 -3141
rect 61276 -3233 61356 -3175
rect 61276 -3260 61291 -3233
rect 61291 -3260 61325 -3233
rect 61325 -3260 61356 -3233
rect 60476 -3460 60536 -3450
rect 60476 -3500 60486 -3460
rect 60486 -3500 60526 -3460
rect 60526 -3500 60536 -3460
rect 60476 -3510 60536 -3500
rect 60616 -3460 60736 -3450
rect 60616 -3500 60626 -3460
rect 60626 -3500 60666 -3460
rect 60666 -3500 60736 -3460
rect 60616 -3510 60736 -3500
rect 60756 -3460 60816 -3450
rect 60756 -3500 60766 -3460
rect 60766 -3500 60806 -3460
rect 60806 -3500 60816 -3460
rect 60756 -3510 60816 -3500
rect 60896 -3460 60956 -3450
rect 60896 -3500 60906 -3460
rect 60906 -3500 60946 -3460
rect 60946 -3500 60956 -3460
rect 60896 -3510 60956 -3500
rect 56380 -3888 56440 -3768
rect 55880 -4080 55970 -4078
rect 55880 -4114 55882 -4080
rect 55882 -4114 55970 -4080
rect 55880 -4158 55970 -4114
rect 55220 -4528 55330 -4418
rect 55530 -4602 55610 -4578
rect 55530 -4636 55560 -4602
rect 55560 -4636 55610 -4602
rect 55530 -4668 55610 -4636
rect 54140 -4708 54150 -4688
rect 54150 -4708 54840 -4688
rect 54840 -4708 54850 -4688
rect 54140 -4948 54850 -4708
rect 55320 -4748 55470 -4728
rect 55320 -4808 55470 -4748
rect 55320 -4868 55470 -4808
rect 56020 -4408 56080 -4258
rect 56170 -4408 56390 -4208
rect 56654 -4486 56998 -4268
rect 59076 -3770 59103 -3740
rect 59103 -3770 59137 -3740
rect 59137 -3770 59166 -3740
rect 59076 -3800 59166 -3770
rect 58926 -3910 58986 -3860
rect 58926 -3930 58966 -3910
rect 58966 -3930 58986 -3910
rect 59146 -3930 59226 -3860
rect 59276 -3930 59356 -3860
rect 59396 -3930 59476 -3860
rect 59646 -3920 59706 -3860
rect 59546 -4008 59606 -4000
rect 59256 -4062 59366 -4030
rect 59546 -4042 59560 -4008
rect 59560 -4042 59594 -4008
rect 59594 -4042 59606 -4008
rect 59016 -4116 59076 -4100
rect 59256 -4090 59366 -4062
rect 59546 -4060 59606 -4042
rect 59016 -4150 59032 -4116
rect 59032 -4150 59066 -4116
rect 59066 -4150 59076 -4116
rect 59016 -4160 59076 -4150
rect 58906 -4300 58926 -4230
rect 58926 -4300 58966 -4230
rect 58966 -4300 58986 -4230
rect 59146 -4300 59226 -4230
rect 59276 -4300 59356 -4230
rect 59396 -4300 59476 -4230
rect 59966 -3740 60326 -3720
rect 59966 -3774 60326 -3740
rect 59966 -3780 60326 -3774
rect 59856 -3794 59916 -3780
rect 59856 -3828 59874 -3794
rect 59874 -3828 59908 -3794
rect 59908 -3828 59916 -3794
rect 59856 -3840 59916 -3828
rect 60376 -3794 60436 -3780
rect 60376 -3828 60384 -3794
rect 60384 -3828 60418 -3794
rect 60418 -3828 60436 -3794
rect 60376 -3840 60436 -3828
rect 61056 -3840 61126 -3740
rect 59806 -4120 59916 -4010
rect 60446 -4150 60526 -4030
rect 59646 -4300 59706 -4240
rect 58986 -4760 59126 -4620
rect 59996 -4700 60106 -4590
rect 59700 -5200 60400 -4900
rect 55600 -5600 55900 -5300
rect 55400 -6500 55700 -6200
rect 21000 -7400 22000 -6600
rect 53520 -7120 53780 -6860
rect 54150 -6908 54860 -6738
rect 54150 -6978 54850 -6908
rect 54850 -6978 54860 -6908
rect 21390 -7612 21620 -7482
rect 53520 -7368 53640 -7258
rect 54750 -7308 54850 -7238
rect 54750 -7318 54840 -7308
rect 55430 -7288 55520 -7218
rect 55290 -7398 55390 -7328
rect 20804 -11629 20846 -7875
rect 20846 -11629 20878 -7875
rect 21186 -11479 21206 -7969
rect 21206 -11479 21256 -7969
rect 21256 -11479 21276 -7969
rect 21726 -11479 21756 -7969
rect 21756 -11479 21816 -7969
rect 22070 -11632 22076 -7872
rect 22076 -11632 22110 -7872
rect 22110 -11632 22140 -7872
rect 53050 -9308 53250 -7558
rect 53950 -7528 53998 -7498
rect 53998 -7528 54020 -7498
rect 53950 -7598 54020 -7528
rect 54920 -7490 54990 -7478
rect 54920 -7528 54926 -7490
rect 54926 -7528 54960 -7490
rect 54960 -7528 54990 -7490
rect 54920 -7568 54990 -7528
rect 53860 -8038 53920 -7928
rect 55230 -7828 55290 -7658
rect 55290 -7828 55320 -7658
rect 55430 -7818 55510 -7648
rect 55960 -7288 56040 -7138
rect 56190 -7368 56390 -7158
rect 56506 -7230 57016 -6980
rect 58966 -7030 59126 -6870
rect 59956 -7060 60166 -6900
rect 55880 -7456 55970 -7418
rect 55880 -7490 55882 -7456
rect 55882 -7490 55970 -7456
rect 55880 -7498 55970 -7490
rect 55000 -8038 55090 -7938
rect 54770 -8240 54840 -8238
rect 54770 -8328 54802 -8240
rect 54802 -8328 54840 -8240
rect 55540 -8038 55630 -7938
rect 56590 -7798 56660 -7668
rect 58906 -7420 58966 -7370
rect 58906 -7430 58926 -7420
rect 58926 -7430 58966 -7420
rect 59216 -7430 59276 -7370
rect 59326 -7430 59386 -7370
rect 59436 -7430 59496 -7370
rect 59636 -7430 59696 -7370
rect 59546 -7501 59606 -7490
rect 59286 -7555 59346 -7530
rect 59546 -7535 59560 -7501
rect 59560 -7535 59594 -7501
rect 59594 -7535 59606 -7501
rect 59286 -7589 59346 -7555
rect 59546 -7550 59606 -7535
rect 59286 -7590 59346 -7589
rect 59016 -7609 59076 -7600
rect 59016 -7643 59032 -7609
rect 59032 -7643 59066 -7609
rect 59066 -7643 59076 -7609
rect 59016 -7660 59076 -7643
rect 59546 -7670 59606 -7610
rect 58906 -7790 58966 -7730
rect 59216 -7780 59276 -7720
rect 59336 -7780 59396 -7720
rect 59436 -7780 59496 -7720
rect 55140 -8408 55200 -8338
rect 55030 -8528 55110 -8448
rect 55740 -8528 55810 -8448
rect 55880 -8528 55970 -8438
rect 56480 -8006 56550 -7988
rect 56480 -8040 56492 -8006
rect 56492 -8040 56530 -8006
rect 56530 -8040 56550 -8006
rect 56480 -8048 56550 -8040
rect 59866 -7630 59966 -7540
rect 60446 -7620 60526 -7520
rect 59636 -7790 59696 -7730
rect 59076 -7878 59166 -7840
rect 59076 -7910 59103 -7878
rect 59103 -7910 59137 -7878
rect 59137 -7910 59166 -7878
rect 60046 -7774 60126 -7740
rect 59856 -7828 59916 -7810
rect 60046 -7800 60126 -7774
rect 59856 -7862 59874 -7828
rect 59874 -7862 59908 -7828
rect 59908 -7862 59916 -7828
rect 59856 -7880 59916 -7862
rect 60376 -7828 60446 -7820
rect 60376 -7862 60384 -7828
rect 60384 -7862 60418 -7828
rect 60418 -7862 60446 -7828
rect 59976 -7916 60316 -7900
rect 60376 -7880 60446 -7862
rect 57098 -7989 57368 -7964
rect 57098 -8023 57125 -7989
rect 57125 -8023 57159 -7989
rect 57159 -8023 57217 -7989
rect 57217 -8023 57251 -7989
rect 57251 -8023 57309 -7989
rect 57309 -8023 57343 -7989
rect 57343 -8023 57368 -7989
rect 54770 -8728 54802 -8648
rect 54802 -8728 54840 -8648
rect 53850 -9048 53920 -8938
rect 54920 -8868 54980 -8798
rect 55000 -9038 55090 -8938
rect 55540 -9038 55630 -8938
rect 55220 -9318 55280 -9148
rect 55280 -9318 55310 -9148
rect 55410 -9328 55500 -9158
rect 53950 -9450 54010 -9408
rect 53950 -9488 53988 -9450
rect 53988 -9488 54010 -9450
rect 54910 -9450 54980 -9398
rect 54910 -9488 54916 -9450
rect 54916 -9488 54950 -9450
rect 54950 -9488 54980 -9450
rect 54910 -9498 54980 -9488
rect 53510 -9648 53630 -9528
rect 54740 -9744 54850 -9668
rect 54740 -9758 54850 -9744
rect 55240 -9618 55370 -9558
rect 55410 -9738 55510 -9648
rect 57098 -8080 57368 -8023
rect 57098 -8104 57368 -8080
rect 56900 -8548 57020 -8418
rect 58576 -8640 58736 -8480
rect 57098 -8880 57368 -8874
rect 56480 -8934 56550 -8928
rect 56480 -8968 56492 -8934
rect 56492 -8968 56530 -8934
rect 56530 -8968 56550 -8934
rect 56480 -8988 56550 -8968
rect 57098 -8965 57368 -8880
rect 57098 -8999 57125 -8965
rect 57125 -8999 57159 -8965
rect 57159 -8999 57217 -8965
rect 57217 -8999 57251 -8965
rect 57251 -8999 57309 -8965
rect 57309 -8999 57343 -8965
rect 57343 -8999 57368 -8965
rect 57098 -9014 57368 -8999
rect 59976 -7952 60316 -7916
rect 59176 -8120 59196 -8040
rect 59196 -8120 59236 -8040
rect 59176 -8320 59196 -8240
rect 59196 -8320 59236 -8240
rect 59076 -8440 59103 -8410
rect 59103 -8440 59137 -8410
rect 59137 -8440 59166 -8410
rect 59076 -8480 59166 -8440
rect 59576 -8098 59636 -8070
rect 59576 -8130 59580 -8098
rect 59580 -8130 59636 -8098
rect 59476 -8320 59502 -8250
rect 59502 -8320 59536 -8250
rect 59576 -8358 59590 -8190
rect 59590 -8358 59624 -8190
rect 59624 -8358 59636 -8190
rect 59576 -8360 59636 -8358
rect 59076 -8608 59166 -8570
rect 59076 -8640 59103 -8608
rect 59103 -8640 59137 -8608
rect 59137 -8640 59166 -8608
rect 59206 -8640 59266 -8570
rect 61206 -8100 61346 -7920
rect 59806 -8340 59818 -8200
rect 59818 -8340 59852 -8200
rect 59852 -8340 59866 -8200
rect 59916 -8182 60006 -8180
rect 59916 -8358 59940 -8182
rect 59940 -8358 60006 -8182
rect 59916 -8360 60006 -8358
rect 60306 -8290 60456 -8150
rect 59826 -8442 59862 -8410
rect 59862 -8442 59896 -8410
rect 59896 -8442 59916 -8410
rect 59826 -8480 59916 -8442
rect 59166 -8810 59196 -8730
rect 59196 -8810 59226 -8730
rect 59166 -9040 59196 -8960
rect 59196 -9040 59226 -8960
rect 59466 -8810 59501 -8730
rect 59501 -8810 59526 -8730
rect 59586 -8850 59589 -8710
rect 59589 -8850 59623 -8710
rect 59623 -8850 59646 -8710
rect 59516 -8921 59596 -8920
rect 59516 -8955 59545 -8921
rect 59545 -8955 59579 -8921
rect 59579 -8955 59596 -8921
rect 59516 -8980 59596 -8955
rect 59826 -8611 59926 -8570
rect 59826 -8640 59861 -8611
rect 59861 -8640 59895 -8611
rect 59895 -8640 59926 -8611
rect 60096 -8483 60127 -8480
rect 60127 -8483 60161 -8480
rect 60161 -8483 60176 -8480
rect 60096 -8541 60176 -8483
rect 60096 -8575 60127 -8541
rect 60127 -8575 60161 -8541
rect 60161 -8575 60176 -8541
rect 60096 -8633 60176 -8575
rect 60096 -8640 60127 -8633
rect 60127 -8640 60161 -8633
rect 60161 -8640 60176 -8633
rect 59796 -8695 59856 -8690
rect 59796 -8870 59817 -8695
rect 59817 -8870 59851 -8695
rect 59851 -8870 59856 -8695
rect 59916 -8695 60006 -8690
rect 59916 -8871 59939 -8695
rect 59939 -8871 60006 -8695
rect 59916 -8880 60006 -8871
rect 60476 -8725 60536 -8710
rect 60476 -8759 60484 -8725
rect 60484 -8759 60536 -8725
rect 60476 -8770 60536 -8759
rect 61036 -8330 61126 -8220
rect 61276 -8483 61291 -8450
rect 61291 -8483 61325 -8450
rect 61325 -8483 61356 -8450
rect 61276 -8541 61356 -8483
rect 61276 -8575 61291 -8541
rect 61291 -8575 61325 -8541
rect 61325 -8575 61356 -8541
rect 61276 -8633 61356 -8575
rect 61276 -8660 61291 -8633
rect 61291 -8660 61325 -8633
rect 61325 -8660 61356 -8633
rect 60476 -8860 60536 -8850
rect 60476 -8900 60486 -8860
rect 60486 -8900 60526 -8860
rect 60526 -8900 60536 -8860
rect 60476 -8910 60536 -8900
rect 60616 -8860 60736 -8850
rect 60616 -8900 60626 -8860
rect 60626 -8900 60666 -8860
rect 60666 -8900 60736 -8860
rect 60616 -8910 60736 -8900
rect 60756 -8860 60816 -8850
rect 60756 -8900 60766 -8860
rect 60766 -8900 60806 -8860
rect 60806 -8900 60816 -8860
rect 60756 -8910 60816 -8900
rect 60896 -8860 60956 -8850
rect 60896 -8900 60906 -8860
rect 60906 -8900 60946 -8860
rect 60946 -8900 60956 -8860
rect 60896 -8910 60956 -8900
rect 56380 -9288 56440 -9168
rect 55880 -9480 55970 -9478
rect 55880 -9514 55882 -9480
rect 55882 -9514 55970 -9480
rect 55880 -9558 55970 -9514
rect 55220 -9928 55330 -9818
rect 55530 -10002 55610 -9978
rect 55530 -10036 55560 -10002
rect 55560 -10036 55610 -10002
rect 55530 -10068 55610 -10036
rect 54140 -10108 54150 -10088
rect 54150 -10108 54840 -10088
rect 54840 -10108 54850 -10088
rect 54140 -10348 54850 -10108
rect 55320 -10148 55470 -10128
rect 55320 -10208 55470 -10148
rect 55320 -10268 55470 -10208
rect 56020 -9808 56080 -9658
rect 56170 -9808 56390 -9608
rect 56654 -9886 56998 -9668
rect 59076 -9170 59103 -9140
rect 59103 -9170 59137 -9140
rect 59137 -9170 59166 -9140
rect 59076 -9200 59166 -9170
rect 58926 -9310 58986 -9260
rect 58926 -9330 58966 -9310
rect 58966 -9330 58986 -9310
rect 59146 -9330 59226 -9260
rect 59276 -9330 59356 -9260
rect 59396 -9330 59476 -9260
rect 59646 -9320 59706 -9260
rect 59546 -9408 59606 -9400
rect 59256 -9462 59366 -9430
rect 59546 -9442 59560 -9408
rect 59560 -9442 59594 -9408
rect 59594 -9442 59606 -9408
rect 59016 -9516 59076 -9500
rect 59256 -9490 59366 -9462
rect 59546 -9460 59606 -9442
rect 59016 -9550 59032 -9516
rect 59032 -9550 59066 -9516
rect 59066 -9550 59076 -9516
rect 59016 -9560 59076 -9550
rect 58906 -9700 58926 -9630
rect 58926 -9700 58966 -9630
rect 58966 -9700 58986 -9630
rect 59146 -9700 59226 -9630
rect 59276 -9700 59356 -9630
rect 59396 -9700 59476 -9630
rect 59966 -9140 60326 -9120
rect 59966 -9174 60326 -9140
rect 59966 -9180 60326 -9174
rect 59856 -9194 59916 -9180
rect 59856 -9228 59874 -9194
rect 59874 -9228 59908 -9194
rect 59908 -9228 59916 -9194
rect 59856 -9240 59916 -9228
rect 60376 -9194 60436 -9180
rect 60376 -9228 60384 -9194
rect 60384 -9228 60418 -9194
rect 60418 -9228 60436 -9194
rect 60376 -9240 60436 -9228
rect 61056 -9240 61126 -9140
rect 59806 -9520 59916 -9410
rect 60446 -9550 60526 -9430
rect 59646 -9700 59706 -9640
rect 58986 -10160 59126 -10020
rect 59996 -10100 60106 -9990
rect 24730 -11632 25190 -11432
rect 21070 -11703 21910 -11702
rect 21070 -11737 21076 -11703
rect 21076 -11737 21394 -11703
rect 21394 -11737 21562 -11703
rect 21562 -11737 21880 -11703
rect 21880 -11737 21910 -11703
rect 21070 -11772 21910 -11737
rect 20260 -12052 20280 -12022
rect 20280 -12052 20340 -12022
rect 20260 -12082 20340 -12052
rect 16527 -13105 16553 -12329
rect 16553 -13105 16586 -12329
rect 16527 -13106 16586 -13105
rect 16730 -13105 16731 -12330
rect 16731 -13105 16765 -12330
rect 16765 -13105 16789 -12330
rect 16730 -13107 16789 -13105
rect 16933 -13105 16959 -12329
rect 16959 -13105 16992 -12329
rect 16933 -13106 16992 -13105
rect 17136 -13105 17137 -12330
rect 17137 -13105 17171 -12330
rect 17171 -13105 17195 -12330
rect 17136 -13107 17195 -13105
rect 17339 -13105 17365 -12329
rect 17365 -13105 17398 -12329
rect 17339 -13106 17398 -13105
rect 17542 -13105 17543 -12330
rect 17543 -13105 17577 -12330
rect 17577 -13105 17601 -12330
rect 17542 -13107 17601 -13105
rect 17745 -13105 17771 -12329
rect 17771 -13105 17804 -12329
rect 17745 -13106 17804 -13105
rect 17948 -13105 17949 -12330
rect 17949 -13105 17983 -12330
rect 17983 -13105 18007 -12330
rect 17948 -13107 18007 -13105
rect 18151 -13105 18177 -12329
rect 18177 -13105 18210 -12329
rect 18151 -13106 18210 -13105
rect 18354 -13105 18355 -12330
rect 18355 -13105 18389 -12330
rect 18389 -13105 18413 -12330
rect 18354 -13107 18413 -13105
rect 18557 -13105 18583 -12329
rect 18583 -13105 18616 -12329
rect 18557 -13106 18616 -13105
rect 18760 -13105 18761 -12330
rect 18761 -13105 18795 -12330
rect 18795 -13105 18819 -12330
rect 18760 -13107 18819 -13105
rect 18963 -13105 18989 -12329
rect 18989 -13105 19022 -12329
rect 18963 -13106 19022 -13105
rect 19166 -13105 19167 -12330
rect 19167 -13105 19201 -12330
rect 19201 -13105 19225 -12330
rect 19166 -13107 19225 -13105
rect 19369 -13105 19395 -12329
rect 19395 -13105 19428 -12329
rect 19369 -13106 19428 -13105
rect 19572 -13105 19573 -12330
rect 19573 -13105 19607 -12330
rect 19607 -13105 19631 -12330
rect 19572 -13107 19631 -13105
rect 19775 -13105 19801 -12329
rect 19801 -13105 19834 -12329
rect 19775 -13106 19834 -13105
rect 19978 -13105 19979 -12330
rect 19979 -13105 20013 -12330
rect 20013 -13105 20037 -12330
rect 19978 -13107 20037 -13105
rect 20181 -13105 20207 -12329
rect 20207 -13105 20240 -12329
rect 20181 -13106 20240 -13105
rect 20384 -13105 20385 -12330
rect 20385 -13105 20419 -12330
rect 20419 -13105 20443 -12330
rect 20384 -13107 20443 -13105
rect 20580 -13042 20613 -12352
rect 20613 -13042 20640 -12352
rect 20801 -13041 20825 -12351
rect 20825 -13041 20861 -12351
rect 20993 -13105 21019 -12329
rect 21019 -13105 21052 -12329
rect 20993 -13106 21052 -13105
rect 21196 -13105 21197 -12330
rect 21197 -13105 21231 -12330
rect 21231 -13105 21255 -12330
rect 21196 -13107 21255 -13105
rect 21399 -13105 21425 -12329
rect 21425 -13105 21458 -12329
rect 21399 -13106 21458 -13105
rect 21602 -13105 21603 -12330
rect 21603 -13105 21637 -12330
rect 21637 -13105 21661 -12330
rect 21602 -13107 21661 -13105
rect 21805 -13105 21831 -12329
rect 21831 -13105 21864 -12329
rect 21805 -13106 21864 -13105
rect 22008 -13105 22009 -12330
rect 22009 -13105 22043 -12330
rect 22043 -13105 22067 -12330
rect 22008 -13107 22067 -13105
rect 22211 -13105 22237 -12329
rect 22237 -13105 22270 -12329
rect 22211 -13106 22270 -13105
rect 22414 -13105 22415 -12330
rect 22415 -13105 22449 -12330
rect 22449 -13105 22473 -12330
rect 22414 -13107 22473 -13105
rect 22617 -13105 22643 -12329
rect 22643 -13105 22676 -12329
rect 22617 -13106 22676 -13105
rect 22820 -13105 22821 -12330
rect 22821 -13105 22855 -12330
rect 22855 -13105 22879 -12330
rect 22820 -13107 22879 -13105
rect 23023 -13105 23049 -12329
rect 23049 -13105 23082 -12329
rect 23023 -13106 23082 -13105
rect 23226 -13105 23227 -12330
rect 23227 -13105 23261 -12330
rect 23261 -13105 23285 -12330
rect 23226 -13107 23285 -13105
rect 23429 -13105 23455 -12329
rect 23455 -13105 23488 -12329
rect 23429 -13106 23488 -13105
rect 23632 -13105 23633 -12330
rect 23633 -13105 23667 -12330
rect 23667 -13105 23691 -12330
rect 23632 -13107 23691 -13105
rect 23835 -13105 23861 -12329
rect 23861 -13105 23894 -12329
rect 23835 -13106 23894 -13105
rect 24038 -13105 24039 -12330
rect 24039 -13105 24073 -12330
rect 24073 -13105 24097 -12330
rect 24038 -13107 24097 -13105
rect 24241 -13105 24267 -12329
rect 24267 -13105 24300 -12329
rect 24241 -13106 24300 -13105
rect 24444 -13105 24445 -12330
rect 24445 -13105 24479 -12330
rect 24479 -13105 24503 -12330
rect 24444 -13107 24503 -13105
rect 24647 -13105 24673 -12329
rect 24673 -13105 24706 -12329
rect 24647 -13106 24706 -13105
rect 24850 -13105 24851 -12330
rect 24851 -13105 24885 -12330
rect 24885 -13105 24909 -12330
rect 24850 -13107 24909 -13105
rect 25090 -12245 25210 -12222
rect 25090 -12279 25141 -12245
rect 25141 -12279 25210 -12245
rect 25090 -12292 25210 -12279
rect 27200 -13000 34400 -10600
rect 55500 -11100 56000 -10700
rect 59700 -10700 60400 -10300
rect 55380 -11980 55740 -11660
rect 53480 -12540 53780 -12340
rect 54150 -12308 54860 -12138
rect 54150 -12378 54850 -12308
rect 54850 -12378 54860 -12308
rect 20570 -13314 20670 -13312
rect 20570 -13362 20670 -13314
rect 20570 -13392 20670 -13362
rect 16580 -14642 16584 -13532
rect 16584 -14642 16981 -13532
rect 16981 -14642 16990 -13532
rect 53520 -12768 53640 -12658
rect 54750 -12708 54850 -12638
rect 54750 -12718 54840 -12708
rect 55430 -12688 55520 -12618
rect 55290 -12798 55390 -12728
rect 53050 -14708 53250 -12958
rect 53950 -12928 53998 -12898
rect 53998 -12928 54020 -12898
rect 53950 -12998 54020 -12928
rect 54920 -12890 54990 -12878
rect 54920 -12928 54926 -12890
rect 54926 -12928 54960 -12890
rect 54960 -12928 54990 -12890
rect 54920 -12968 54990 -12928
rect 53860 -13438 53920 -13328
rect 55230 -13228 55290 -13058
rect 55290 -13228 55320 -13058
rect 55430 -13218 55510 -13048
rect 55960 -12688 56040 -12538
rect 56190 -12768 56390 -12558
rect 56506 -12630 57016 -12380
rect 58966 -12430 59126 -12270
rect 59956 -12460 60166 -12300
rect 55880 -12856 55970 -12818
rect 55880 -12890 55882 -12856
rect 55882 -12890 55970 -12856
rect 55880 -12898 55970 -12890
rect 55000 -13438 55090 -13338
rect 54770 -13640 54840 -13638
rect 54770 -13728 54802 -13640
rect 54802 -13728 54840 -13640
rect 55540 -13438 55630 -13338
rect 56590 -13198 56660 -13068
rect 58906 -12820 58966 -12770
rect 58906 -12830 58926 -12820
rect 58926 -12830 58966 -12820
rect 59216 -12830 59276 -12770
rect 59326 -12830 59386 -12770
rect 59436 -12830 59496 -12770
rect 59636 -12830 59696 -12770
rect 59546 -12901 59606 -12890
rect 59286 -12955 59346 -12930
rect 59546 -12935 59560 -12901
rect 59560 -12935 59594 -12901
rect 59594 -12935 59606 -12901
rect 59286 -12989 59346 -12955
rect 59546 -12950 59606 -12935
rect 59286 -12990 59346 -12989
rect 59016 -13009 59076 -13000
rect 59016 -13043 59032 -13009
rect 59032 -13043 59066 -13009
rect 59066 -13043 59076 -13009
rect 59016 -13060 59076 -13043
rect 59546 -13070 59606 -13010
rect 58906 -13190 58966 -13130
rect 59216 -13180 59276 -13120
rect 59336 -13180 59396 -13120
rect 59436 -13180 59496 -13120
rect 55140 -13808 55200 -13738
rect 55030 -13928 55110 -13848
rect 55740 -13928 55810 -13848
rect 55880 -13928 55970 -13838
rect 56480 -13406 56550 -13388
rect 56480 -13440 56492 -13406
rect 56492 -13440 56530 -13406
rect 56530 -13440 56550 -13406
rect 56480 -13448 56550 -13440
rect 59866 -13030 59966 -12940
rect 60446 -13020 60526 -12920
rect 59636 -13190 59696 -13130
rect 59076 -13278 59166 -13240
rect 59076 -13310 59103 -13278
rect 59103 -13310 59137 -13278
rect 59137 -13310 59166 -13278
rect 60046 -13174 60126 -13140
rect 59856 -13228 59916 -13210
rect 60046 -13200 60126 -13174
rect 59856 -13262 59874 -13228
rect 59874 -13262 59908 -13228
rect 59908 -13262 59916 -13228
rect 59856 -13280 59916 -13262
rect 60376 -13228 60446 -13220
rect 60376 -13262 60384 -13228
rect 60384 -13262 60418 -13228
rect 60418 -13262 60446 -13228
rect 59976 -13316 60316 -13300
rect 60376 -13280 60446 -13262
rect 57098 -13389 57368 -13364
rect 57098 -13423 57125 -13389
rect 57125 -13423 57159 -13389
rect 57159 -13423 57217 -13389
rect 57217 -13423 57251 -13389
rect 57251 -13423 57309 -13389
rect 57309 -13423 57343 -13389
rect 57343 -13423 57368 -13389
rect 54770 -14128 54802 -14048
rect 54802 -14128 54840 -14048
rect 53850 -14448 53920 -14338
rect 54920 -14268 54980 -14198
rect 55000 -14438 55090 -14338
rect 55540 -14438 55630 -14338
rect 55220 -14718 55280 -14548
rect 55280 -14718 55310 -14548
rect 55410 -14728 55500 -14558
rect 16580 -16018 16584 -14912
rect 16584 -16018 16981 -14912
rect 16981 -16018 16990 -14912
rect 16580 -16022 16990 -16018
rect 53950 -14850 54010 -14808
rect 53950 -14888 53988 -14850
rect 53988 -14888 54010 -14850
rect 54910 -14850 54980 -14798
rect 54910 -14888 54916 -14850
rect 54916 -14888 54950 -14850
rect 54950 -14888 54980 -14850
rect 54910 -14898 54980 -14888
rect 53510 -15048 53630 -14928
rect 54740 -15144 54850 -15068
rect 54740 -15158 54850 -15144
rect 55240 -15018 55370 -14958
rect 55410 -15138 55510 -15048
rect 57098 -13480 57368 -13423
rect 57098 -13504 57368 -13480
rect 56900 -13948 57020 -13818
rect 58576 -14040 58736 -13880
rect 57098 -14280 57368 -14274
rect 56480 -14334 56550 -14328
rect 56480 -14368 56492 -14334
rect 56492 -14368 56530 -14334
rect 56530 -14368 56550 -14334
rect 56480 -14388 56550 -14368
rect 57098 -14365 57368 -14280
rect 57098 -14399 57125 -14365
rect 57125 -14399 57159 -14365
rect 57159 -14399 57217 -14365
rect 57217 -14399 57251 -14365
rect 57251 -14399 57309 -14365
rect 57309 -14399 57343 -14365
rect 57343 -14399 57368 -14365
rect 57098 -14414 57368 -14399
rect 59976 -13352 60316 -13316
rect 59176 -13520 59196 -13440
rect 59196 -13520 59236 -13440
rect 59176 -13720 59196 -13640
rect 59196 -13720 59236 -13640
rect 59076 -13840 59103 -13810
rect 59103 -13840 59137 -13810
rect 59137 -13840 59166 -13810
rect 59076 -13880 59166 -13840
rect 59576 -13498 59636 -13470
rect 59576 -13530 59580 -13498
rect 59580 -13530 59636 -13498
rect 59476 -13720 59502 -13650
rect 59502 -13720 59536 -13650
rect 59576 -13758 59590 -13590
rect 59590 -13758 59624 -13590
rect 59624 -13758 59636 -13590
rect 59576 -13760 59636 -13758
rect 59076 -14008 59166 -13970
rect 59076 -14040 59103 -14008
rect 59103 -14040 59137 -14008
rect 59137 -14040 59166 -14008
rect 59206 -14040 59266 -13970
rect 61206 -13500 61346 -13320
rect 59806 -13740 59818 -13600
rect 59818 -13740 59852 -13600
rect 59852 -13740 59866 -13600
rect 59916 -13582 60006 -13580
rect 59916 -13758 59940 -13582
rect 59940 -13758 60006 -13582
rect 59916 -13760 60006 -13758
rect 60306 -13690 60456 -13550
rect 59826 -13842 59862 -13810
rect 59862 -13842 59896 -13810
rect 59896 -13842 59916 -13810
rect 59826 -13880 59916 -13842
rect 59166 -14210 59196 -14130
rect 59196 -14210 59226 -14130
rect 59166 -14440 59196 -14360
rect 59196 -14440 59226 -14360
rect 59466 -14210 59501 -14130
rect 59501 -14210 59526 -14130
rect 59586 -14250 59589 -14110
rect 59589 -14250 59623 -14110
rect 59623 -14250 59646 -14110
rect 59516 -14321 59596 -14320
rect 59516 -14355 59545 -14321
rect 59545 -14355 59579 -14321
rect 59579 -14355 59596 -14321
rect 59516 -14380 59596 -14355
rect 59826 -14011 59926 -13970
rect 59826 -14040 59861 -14011
rect 59861 -14040 59895 -14011
rect 59895 -14040 59926 -14011
rect 60096 -13883 60127 -13880
rect 60127 -13883 60161 -13880
rect 60161 -13883 60176 -13880
rect 60096 -13941 60176 -13883
rect 60096 -13975 60127 -13941
rect 60127 -13975 60161 -13941
rect 60161 -13975 60176 -13941
rect 60096 -14033 60176 -13975
rect 60096 -14040 60127 -14033
rect 60127 -14040 60161 -14033
rect 60161 -14040 60176 -14033
rect 59796 -14095 59856 -14090
rect 59796 -14270 59817 -14095
rect 59817 -14270 59851 -14095
rect 59851 -14270 59856 -14095
rect 59916 -14095 60006 -14090
rect 59916 -14271 59939 -14095
rect 59939 -14271 60006 -14095
rect 59916 -14280 60006 -14271
rect 60476 -14125 60536 -14110
rect 60476 -14159 60484 -14125
rect 60484 -14159 60536 -14125
rect 60476 -14170 60536 -14159
rect 61036 -13730 61126 -13620
rect 61276 -13883 61291 -13850
rect 61291 -13883 61325 -13850
rect 61325 -13883 61356 -13850
rect 61276 -13941 61356 -13883
rect 61276 -13975 61291 -13941
rect 61291 -13975 61325 -13941
rect 61325 -13975 61356 -13941
rect 61276 -14033 61356 -13975
rect 61276 -14060 61291 -14033
rect 61291 -14060 61325 -14033
rect 61325 -14060 61356 -14033
rect 60476 -14260 60536 -14250
rect 60476 -14300 60486 -14260
rect 60486 -14300 60526 -14260
rect 60526 -14300 60536 -14260
rect 60476 -14310 60536 -14300
rect 60616 -14260 60736 -14250
rect 60616 -14300 60626 -14260
rect 60626 -14300 60666 -14260
rect 60666 -14300 60736 -14260
rect 60616 -14310 60736 -14300
rect 60756 -14260 60816 -14250
rect 60756 -14300 60766 -14260
rect 60766 -14300 60806 -14260
rect 60806 -14300 60816 -14260
rect 60756 -14310 60816 -14300
rect 60896 -14260 60956 -14250
rect 60896 -14300 60906 -14260
rect 60906 -14300 60946 -14260
rect 60946 -14300 60956 -14260
rect 60896 -14310 60956 -14300
rect 56380 -14688 56440 -14568
rect 55880 -14880 55970 -14878
rect 55880 -14914 55882 -14880
rect 55882 -14914 55970 -14880
rect 55880 -14958 55970 -14914
rect 55220 -15328 55330 -15218
rect 55530 -15402 55610 -15378
rect 55530 -15436 55560 -15402
rect 55560 -15436 55610 -15402
rect 55530 -15468 55610 -15436
rect 54140 -15508 54150 -15488
rect 54150 -15508 54840 -15488
rect 54840 -15508 54850 -15488
rect 54140 -15748 54850 -15508
rect 55320 -15548 55470 -15528
rect 55320 -15608 55470 -15548
rect 55320 -15668 55470 -15608
rect 56020 -15208 56080 -15058
rect 56170 -15208 56390 -15008
rect 56654 -15286 56998 -15068
rect 59076 -14570 59103 -14540
rect 59103 -14570 59137 -14540
rect 59137 -14570 59166 -14540
rect 59076 -14600 59166 -14570
rect 58926 -14710 58986 -14660
rect 58926 -14730 58966 -14710
rect 58966 -14730 58986 -14710
rect 59146 -14730 59226 -14660
rect 59276 -14730 59356 -14660
rect 59396 -14730 59476 -14660
rect 59646 -14720 59706 -14660
rect 59546 -14808 59606 -14800
rect 59256 -14862 59366 -14830
rect 59546 -14842 59560 -14808
rect 59560 -14842 59594 -14808
rect 59594 -14842 59606 -14808
rect 59016 -14916 59076 -14900
rect 59256 -14890 59366 -14862
rect 59546 -14860 59606 -14842
rect 59016 -14950 59032 -14916
rect 59032 -14950 59066 -14916
rect 59066 -14950 59076 -14916
rect 59016 -14960 59076 -14950
rect 58906 -15100 58926 -15030
rect 58926 -15100 58966 -15030
rect 58966 -15100 58986 -15030
rect 59146 -15100 59226 -15030
rect 59276 -15100 59356 -15030
rect 59396 -15100 59476 -15030
rect 59966 -14540 60326 -14520
rect 59966 -14574 60326 -14540
rect 59966 -14580 60326 -14574
rect 59856 -14594 59916 -14580
rect 59856 -14628 59874 -14594
rect 59874 -14628 59908 -14594
rect 59908 -14628 59916 -14594
rect 59856 -14640 59916 -14628
rect 60376 -14594 60436 -14580
rect 60376 -14628 60384 -14594
rect 60384 -14628 60418 -14594
rect 60418 -14628 60436 -14594
rect 60376 -14640 60436 -14628
rect 61056 -14640 61126 -14540
rect 59806 -14920 59916 -14810
rect 60446 -14950 60526 -14830
rect 59646 -15100 59706 -15040
rect 58986 -15560 59126 -15420
rect 59996 -15500 60106 -15390
rect 59800 -15900 60300 -15600
rect 55500 -16500 56000 -16100
rect 55400 -17400 55700 -17100
rect 53500 -17940 53780 -17740
rect 54150 -17708 54860 -17538
rect 54150 -17778 54850 -17708
rect 54850 -17778 54860 -17708
rect 53520 -18168 53640 -18058
rect 54750 -18108 54850 -18038
rect 54750 -18118 54840 -18108
rect 55430 -18088 55520 -18018
rect 55290 -18198 55390 -18128
rect 53050 -20108 53250 -18358
rect 53950 -18328 53998 -18298
rect 53998 -18328 54020 -18298
rect 53950 -18398 54020 -18328
rect 54920 -18290 54990 -18278
rect 54920 -18328 54926 -18290
rect 54926 -18328 54960 -18290
rect 54960 -18328 54990 -18290
rect 54920 -18368 54990 -18328
rect 53860 -18838 53920 -18728
rect 55230 -18628 55290 -18458
rect 55290 -18628 55320 -18458
rect 55430 -18618 55510 -18448
rect 55960 -18088 56040 -17938
rect 56190 -18168 56390 -17958
rect 56506 -18030 57016 -17780
rect 58966 -17830 59126 -17670
rect 59956 -17860 60166 -17700
rect 55880 -18256 55970 -18218
rect 55880 -18290 55882 -18256
rect 55882 -18290 55970 -18256
rect 55880 -18298 55970 -18290
rect 55000 -18838 55090 -18738
rect 54770 -19040 54840 -19038
rect 54770 -19128 54802 -19040
rect 54802 -19128 54840 -19040
rect 55540 -18838 55630 -18738
rect 56590 -18598 56660 -18468
rect 58906 -18220 58966 -18170
rect 58906 -18230 58926 -18220
rect 58926 -18230 58966 -18220
rect 59216 -18230 59276 -18170
rect 59326 -18230 59386 -18170
rect 59436 -18230 59496 -18170
rect 59636 -18230 59696 -18170
rect 59546 -18301 59606 -18290
rect 59286 -18355 59346 -18330
rect 59546 -18335 59560 -18301
rect 59560 -18335 59594 -18301
rect 59594 -18335 59606 -18301
rect 59286 -18389 59346 -18355
rect 59546 -18350 59606 -18335
rect 59286 -18390 59346 -18389
rect 59016 -18409 59076 -18400
rect 59016 -18443 59032 -18409
rect 59032 -18443 59066 -18409
rect 59066 -18443 59076 -18409
rect 59016 -18460 59076 -18443
rect 59546 -18470 59606 -18410
rect 58906 -18590 58966 -18530
rect 59216 -18580 59276 -18520
rect 59336 -18580 59396 -18520
rect 59436 -18580 59496 -18520
rect 55140 -19208 55200 -19138
rect 55030 -19328 55110 -19248
rect 55740 -19328 55810 -19248
rect 55880 -19328 55970 -19238
rect 56480 -18806 56550 -18788
rect 56480 -18840 56492 -18806
rect 56492 -18840 56530 -18806
rect 56530 -18840 56550 -18806
rect 56480 -18848 56550 -18840
rect 59866 -18430 59966 -18340
rect 60446 -18420 60526 -18320
rect 59636 -18590 59696 -18530
rect 59076 -18678 59166 -18640
rect 59076 -18710 59103 -18678
rect 59103 -18710 59137 -18678
rect 59137 -18710 59166 -18678
rect 60046 -18574 60126 -18540
rect 59856 -18628 59916 -18610
rect 60046 -18600 60126 -18574
rect 59856 -18662 59874 -18628
rect 59874 -18662 59908 -18628
rect 59908 -18662 59916 -18628
rect 59856 -18680 59916 -18662
rect 60376 -18628 60446 -18620
rect 60376 -18662 60384 -18628
rect 60384 -18662 60418 -18628
rect 60418 -18662 60446 -18628
rect 59976 -18716 60316 -18700
rect 60376 -18680 60446 -18662
rect 57098 -18789 57368 -18764
rect 57098 -18823 57125 -18789
rect 57125 -18823 57159 -18789
rect 57159 -18823 57217 -18789
rect 57217 -18823 57251 -18789
rect 57251 -18823 57309 -18789
rect 57309 -18823 57343 -18789
rect 57343 -18823 57368 -18789
rect 54770 -19528 54802 -19448
rect 54802 -19528 54840 -19448
rect 53850 -19848 53920 -19738
rect 54920 -19668 54980 -19598
rect 55000 -19838 55090 -19738
rect 55540 -19838 55630 -19738
rect 55220 -20118 55280 -19948
rect 55280 -20118 55310 -19948
rect 55410 -20128 55500 -19958
rect 53950 -20250 54010 -20208
rect 53950 -20288 53988 -20250
rect 53988 -20288 54010 -20250
rect 54910 -20250 54980 -20198
rect 54910 -20288 54916 -20250
rect 54916 -20288 54950 -20250
rect 54950 -20288 54980 -20250
rect 54910 -20298 54980 -20288
rect 53510 -20448 53630 -20328
rect 54740 -20544 54850 -20468
rect 54740 -20558 54850 -20544
rect 55240 -20418 55370 -20358
rect 55410 -20538 55510 -20448
rect 57098 -18880 57368 -18823
rect 57098 -18904 57368 -18880
rect 56900 -19348 57020 -19218
rect 58576 -19440 58736 -19280
rect 57098 -19680 57368 -19674
rect 56480 -19734 56550 -19728
rect 56480 -19768 56492 -19734
rect 56492 -19768 56530 -19734
rect 56530 -19768 56550 -19734
rect 56480 -19788 56550 -19768
rect 57098 -19765 57368 -19680
rect 57098 -19799 57125 -19765
rect 57125 -19799 57159 -19765
rect 57159 -19799 57217 -19765
rect 57217 -19799 57251 -19765
rect 57251 -19799 57309 -19765
rect 57309 -19799 57343 -19765
rect 57343 -19799 57368 -19765
rect 57098 -19814 57368 -19799
rect 59976 -18752 60316 -18716
rect 59176 -18920 59196 -18840
rect 59196 -18920 59236 -18840
rect 59176 -19120 59196 -19040
rect 59196 -19120 59236 -19040
rect 59076 -19240 59103 -19210
rect 59103 -19240 59137 -19210
rect 59137 -19240 59166 -19210
rect 59076 -19280 59166 -19240
rect 59576 -18898 59636 -18870
rect 59576 -18930 59580 -18898
rect 59580 -18930 59636 -18898
rect 59476 -19120 59502 -19050
rect 59502 -19120 59536 -19050
rect 59576 -19158 59590 -18990
rect 59590 -19158 59624 -18990
rect 59624 -19158 59636 -18990
rect 59576 -19160 59636 -19158
rect 59076 -19408 59166 -19370
rect 59076 -19440 59103 -19408
rect 59103 -19440 59137 -19408
rect 59137 -19440 59166 -19408
rect 59206 -19440 59266 -19370
rect 61206 -18900 61346 -18720
rect 59806 -19140 59818 -19000
rect 59818 -19140 59852 -19000
rect 59852 -19140 59866 -19000
rect 59916 -18982 60006 -18980
rect 59916 -19158 59940 -18982
rect 59940 -19158 60006 -18982
rect 59916 -19160 60006 -19158
rect 60306 -19090 60456 -18950
rect 59826 -19242 59862 -19210
rect 59862 -19242 59896 -19210
rect 59896 -19242 59916 -19210
rect 59826 -19280 59916 -19242
rect 59166 -19610 59196 -19530
rect 59196 -19610 59226 -19530
rect 59166 -19840 59196 -19760
rect 59196 -19840 59226 -19760
rect 59466 -19610 59501 -19530
rect 59501 -19610 59526 -19530
rect 59586 -19650 59589 -19510
rect 59589 -19650 59623 -19510
rect 59623 -19650 59646 -19510
rect 59516 -19721 59596 -19720
rect 59516 -19755 59545 -19721
rect 59545 -19755 59579 -19721
rect 59579 -19755 59596 -19721
rect 59516 -19780 59596 -19755
rect 59826 -19411 59926 -19370
rect 59826 -19440 59861 -19411
rect 59861 -19440 59895 -19411
rect 59895 -19440 59926 -19411
rect 60096 -19283 60127 -19280
rect 60127 -19283 60161 -19280
rect 60161 -19283 60176 -19280
rect 60096 -19341 60176 -19283
rect 60096 -19375 60127 -19341
rect 60127 -19375 60161 -19341
rect 60161 -19375 60176 -19341
rect 60096 -19433 60176 -19375
rect 60096 -19440 60127 -19433
rect 60127 -19440 60161 -19433
rect 60161 -19440 60176 -19433
rect 59796 -19495 59856 -19490
rect 59796 -19670 59817 -19495
rect 59817 -19670 59851 -19495
rect 59851 -19670 59856 -19495
rect 59916 -19495 60006 -19490
rect 59916 -19671 59939 -19495
rect 59939 -19671 60006 -19495
rect 59916 -19680 60006 -19671
rect 60476 -19525 60536 -19510
rect 60476 -19559 60484 -19525
rect 60484 -19559 60536 -19525
rect 60476 -19570 60536 -19559
rect 61036 -19130 61126 -19020
rect 61276 -19283 61291 -19250
rect 61291 -19283 61325 -19250
rect 61325 -19283 61356 -19250
rect 61276 -19341 61356 -19283
rect 61276 -19375 61291 -19341
rect 61291 -19375 61325 -19341
rect 61325 -19375 61356 -19341
rect 61276 -19433 61356 -19375
rect 61276 -19460 61291 -19433
rect 61291 -19460 61325 -19433
rect 61325 -19460 61356 -19433
rect 60476 -19660 60536 -19650
rect 60476 -19700 60486 -19660
rect 60486 -19700 60526 -19660
rect 60526 -19700 60536 -19660
rect 60476 -19710 60536 -19700
rect 60616 -19660 60736 -19650
rect 60616 -19700 60626 -19660
rect 60626 -19700 60666 -19660
rect 60666 -19700 60736 -19660
rect 60616 -19710 60736 -19700
rect 60756 -19660 60816 -19650
rect 60756 -19700 60766 -19660
rect 60766 -19700 60806 -19660
rect 60806 -19700 60816 -19660
rect 60756 -19710 60816 -19700
rect 60896 -19660 60956 -19650
rect 60896 -19700 60906 -19660
rect 60906 -19700 60946 -19660
rect 60946 -19700 60956 -19660
rect 60896 -19710 60956 -19700
rect 56380 -20088 56440 -19968
rect 55880 -20280 55970 -20278
rect 55880 -20314 55882 -20280
rect 55882 -20314 55970 -20280
rect 55880 -20358 55970 -20314
rect 55220 -20728 55330 -20618
rect 55530 -20802 55610 -20778
rect 55530 -20836 55560 -20802
rect 55560 -20836 55610 -20802
rect 55530 -20868 55610 -20836
rect 54140 -20908 54150 -20888
rect 54150 -20908 54840 -20888
rect 54840 -20908 54850 -20888
rect 54140 -21148 54850 -20908
rect 55320 -20948 55470 -20928
rect 55320 -21008 55470 -20948
rect 55320 -21068 55470 -21008
rect 56020 -20608 56080 -20458
rect 56170 -20608 56390 -20408
rect 56654 -20686 56998 -20468
rect 59076 -19970 59103 -19940
rect 59103 -19970 59137 -19940
rect 59137 -19970 59166 -19940
rect 59076 -20000 59166 -19970
rect 58926 -20110 58986 -20060
rect 58926 -20130 58966 -20110
rect 58966 -20130 58986 -20110
rect 59146 -20130 59226 -20060
rect 59276 -20130 59356 -20060
rect 59396 -20130 59476 -20060
rect 59646 -20120 59706 -20060
rect 59546 -20208 59606 -20200
rect 59256 -20262 59366 -20230
rect 59546 -20242 59560 -20208
rect 59560 -20242 59594 -20208
rect 59594 -20242 59606 -20208
rect 59016 -20316 59076 -20300
rect 59256 -20290 59366 -20262
rect 59546 -20260 59606 -20242
rect 59016 -20350 59032 -20316
rect 59032 -20350 59066 -20316
rect 59066 -20350 59076 -20316
rect 59016 -20360 59076 -20350
rect 58906 -20500 58926 -20430
rect 58926 -20500 58966 -20430
rect 58966 -20500 58986 -20430
rect 59146 -20500 59226 -20430
rect 59276 -20500 59356 -20430
rect 59396 -20500 59476 -20430
rect 59966 -19940 60326 -19920
rect 59966 -19974 60326 -19940
rect 59966 -19980 60326 -19974
rect 59856 -19994 59916 -19980
rect 59856 -20028 59874 -19994
rect 59874 -20028 59908 -19994
rect 59908 -20028 59916 -19994
rect 59856 -20040 59916 -20028
rect 60376 -19994 60436 -19980
rect 60376 -20028 60384 -19994
rect 60384 -20028 60418 -19994
rect 60418 -20028 60436 -19994
rect 60376 -20040 60436 -20028
rect 61056 -20040 61126 -19940
rect 59806 -20320 59916 -20210
rect 60446 -20350 60526 -20230
rect 59646 -20500 59706 -20440
rect 58986 -20960 59126 -20820
rect 59996 -20900 60106 -20790
rect 59800 -21300 60300 -21000
rect 55500 -21900 56100 -21500
rect 55440 -22760 55720 -22480
rect 53480 -23340 53780 -23140
rect 54150 -23108 54860 -22938
rect 54150 -23178 54850 -23108
rect 54850 -23178 54860 -23108
rect 53520 -23568 53640 -23458
rect 54750 -23508 54850 -23438
rect 54750 -23518 54840 -23508
rect 55430 -23488 55520 -23418
rect 55290 -23598 55390 -23528
rect 53050 -25508 53250 -23758
rect 53950 -23728 53998 -23698
rect 53998 -23728 54020 -23698
rect 53950 -23798 54020 -23728
rect 54920 -23690 54990 -23678
rect 54920 -23728 54926 -23690
rect 54926 -23728 54960 -23690
rect 54960 -23728 54990 -23690
rect 54920 -23768 54990 -23728
rect 53860 -24238 53920 -24128
rect 55230 -24028 55290 -23858
rect 55290 -24028 55320 -23858
rect 55430 -24018 55510 -23848
rect 55960 -23488 56040 -23338
rect 56190 -23568 56390 -23358
rect 56506 -23430 57016 -23180
rect 58966 -23230 59126 -23070
rect 59956 -23260 60166 -23100
rect 55880 -23656 55970 -23618
rect 55880 -23690 55882 -23656
rect 55882 -23690 55970 -23656
rect 55880 -23698 55970 -23690
rect 55000 -24238 55090 -24138
rect 54770 -24440 54840 -24438
rect 54770 -24528 54802 -24440
rect 54802 -24528 54840 -24440
rect 55540 -24238 55630 -24138
rect 56590 -23998 56660 -23868
rect 58906 -23620 58966 -23570
rect 58906 -23630 58926 -23620
rect 58926 -23630 58966 -23620
rect 59216 -23630 59276 -23570
rect 59326 -23630 59386 -23570
rect 59436 -23630 59496 -23570
rect 59636 -23630 59696 -23570
rect 59546 -23701 59606 -23690
rect 59286 -23755 59346 -23730
rect 59546 -23735 59560 -23701
rect 59560 -23735 59594 -23701
rect 59594 -23735 59606 -23701
rect 59286 -23789 59346 -23755
rect 59546 -23750 59606 -23735
rect 59286 -23790 59346 -23789
rect 59016 -23809 59076 -23800
rect 59016 -23843 59032 -23809
rect 59032 -23843 59066 -23809
rect 59066 -23843 59076 -23809
rect 59016 -23860 59076 -23843
rect 59546 -23870 59606 -23810
rect 58906 -23990 58966 -23930
rect 59216 -23980 59276 -23920
rect 59336 -23980 59396 -23920
rect 59436 -23980 59496 -23920
rect 55140 -24608 55200 -24538
rect 55030 -24728 55110 -24648
rect 55740 -24728 55810 -24648
rect 55880 -24728 55970 -24638
rect 56480 -24206 56550 -24188
rect 56480 -24240 56492 -24206
rect 56492 -24240 56530 -24206
rect 56530 -24240 56550 -24206
rect 56480 -24248 56550 -24240
rect 59866 -23830 59966 -23740
rect 60446 -23820 60526 -23720
rect 59636 -23990 59696 -23930
rect 59076 -24078 59166 -24040
rect 59076 -24110 59103 -24078
rect 59103 -24110 59137 -24078
rect 59137 -24110 59166 -24078
rect 60046 -23974 60126 -23940
rect 59856 -24028 59916 -24010
rect 60046 -24000 60126 -23974
rect 59856 -24062 59874 -24028
rect 59874 -24062 59908 -24028
rect 59908 -24062 59916 -24028
rect 59856 -24080 59916 -24062
rect 60376 -24028 60446 -24020
rect 60376 -24062 60384 -24028
rect 60384 -24062 60418 -24028
rect 60418 -24062 60446 -24028
rect 59976 -24116 60316 -24100
rect 60376 -24080 60446 -24062
rect 57098 -24189 57368 -24164
rect 57098 -24223 57125 -24189
rect 57125 -24223 57159 -24189
rect 57159 -24223 57217 -24189
rect 57217 -24223 57251 -24189
rect 57251 -24223 57309 -24189
rect 57309 -24223 57343 -24189
rect 57343 -24223 57368 -24189
rect 54770 -24928 54802 -24848
rect 54802 -24928 54840 -24848
rect 53850 -25248 53920 -25138
rect 54920 -25068 54980 -24998
rect 55000 -25238 55090 -25138
rect 55540 -25238 55630 -25138
rect 55220 -25518 55280 -25348
rect 55280 -25518 55310 -25348
rect 55410 -25528 55500 -25358
rect 53950 -25650 54010 -25608
rect 53950 -25688 53988 -25650
rect 53988 -25688 54010 -25650
rect 54910 -25650 54980 -25598
rect 54910 -25688 54916 -25650
rect 54916 -25688 54950 -25650
rect 54950 -25688 54980 -25650
rect 54910 -25698 54980 -25688
rect 15000 -31200 19400 -26400
rect 53510 -25848 53630 -25728
rect 54740 -25944 54850 -25868
rect 54740 -25958 54850 -25944
rect 55240 -25818 55370 -25758
rect 55410 -25938 55510 -25848
rect 57098 -24280 57368 -24223
rect 57098 -24304 57368 -24280
rect 56900 -24748 57020 -24618
rect 58576 -24840 58736 -24680
rect 57098 -25080 57368 -25074
rect 56480 -25134 56550 -25128
rect 56480 -25168 56492 -25134
rect 56492 -25168 56530 -25134
rect 56530 -25168 56550 -25134
rect 56480 -25188 56550 -25168
rect 57098 -25165 57368 -25080
rect 57098 -25199 57125 -25165
rect 57125 -25199 57159 -25165
rect 57159 -25199 57217 -25165
rect 57217 -25199 57251 -25165
rect 57251 -25199 57309 -25165
rect 57309 -25199 57343 -25165
rect 57343 -25199 57368 -25165
rect 57098 -25214 57368 -25199
rect 59976 -24152 60316 -24116
rect 59176 -24320 59196 -24240
rect 59196 -24320 59236 -24240
rect 59176 -24520 59196 -24440
rect 59196 -24520 59236 -24440
rect 59076 -24640 59103 -24610
rect 59103 -24640 59137 -24610
rect 59137 -24640 59166 -24610
rect 59076 -24680 59166 -24640
rect 59576 -24298 59636 -24270
rect 59576 -24330 59580 -24298
rect 59580 -24330 59636 -24298
rect 59476 -24520 59502 -24450
rect 59502 -24520 59536 -24450
rect 59576 -24558 59590 -24390
rect 59590 -24558 59624 -24390
rect 59624 -24558 59636 -24390
rect 59576 -24560 59636 -24558
rect 59076 -24808 59166 -24770
rect 59076 -24840 59103 -24808
rect 59103 -24840 59137 -24808
rect 59137 -24840 59166 -24808
rect 59206 -24840 59266 -24770
rect 61206 -24300 61346 -24120
rect 59806 -24540 59818 -24400
rect 59818 -24540 59852 -24400
rect 59852 -24540 59866 -24400
rect 59916 -24382 60006 -24380
rect 59916 -24558 59940 -24382
rect 59940 -24558 60006 -24382
rect 59916 -24560 60006 -24558
rect 60306 -24490 60456 -24350
rect 59826 -24642 59862 -24610
rect 59862 -24642 59896 -24610
rect 59896 -24642 59916 -24610
rect 59826 -24680 59916 -24642
rect 59166 -25010 59196 -24930
rect 59196 -25010 59226 -24930
rect 59166 -25240 59196 -25160
rect 59196 -25240 59226 -25160
rect 59466 -25010 59501 -24930
rect 59501 -25010 59526 -24930
rect 59586 -25050 59589 -24910
rect 59589 -25050 59623 -24910
rect 59623 -25050 59646 -24910
rect 59516 -25121 59596 -25120
rect 59516 -25155 59545 -25121
rect 59545 -25155 59579 -25121
rect 59579 -25155 59596 -25121
rect 59516 -25180 59596 -25155
rect 59826 -24811 59926 -24770
rect 59826 -24840 59861 -24811
rect 59861 -24840 59895 -24811
rect 59895 -24840 59926 -24811
rect 60096 -24683 60127 -24680
rect 60127 -24683 60161 -24680
rect 60161 -24683 60176 -24680
rect 60096 -24741 60176 -24683
rect 60096 -24775 60127 -24741
rect 60127 -24775 60161 -24741
rect 60161 -24775 60176 -24741
rect 60096 -24833 60176 -24775
rect 60096 -24840 60127 -24833
rect 60127 -24840 60161 -24833
rect 60161 -24840 60176 -24833
rect 59796 -24895 59856 -24890
rect 59796 -25070 59817 -24895
rect 59817 -25070 59851 -24895
rect 59851 -25070 59856 -24895
rect 59916 -24895 60006 -24890
rect 59916 -25071 59939 -24895
rect 59939 -25071 60006 -24895
rect 59916 -25080 60006 -25071
rect 60476 -24925 60536 -24910
rect 60476 -24959 60484 -24925
rect 60484 -24959 60536 -24925
rect 60476 -24970 60536 -24959
rect 61036 -24530 61126 -24420
rect 61276 -24683 61291 -24650
rect 61291 -24683 61325 -24650
rect 61325 -24683 61356 -24650
rect 61276 -24741 61356 -24683
rect 61276 -24775 61291 -24741
rect 61291 -24775 61325 -24741
rect 61325 -24775 61356 -24741
rect 61276 -24833 61356 -24775
rect 61276 -24860 61291 -24833
rect 61291 -24860 61325 -24833
rect 61325 -24860 61356 -24833
rect 60476 -25060 60536 -25050
rect 60476 -25100 60486 -25060
rect 60486 -25100 60526 -25060
rect 60526 -25100 60536 -25060
rect 60476 -25110 60536 -25100
rect 60616 -25060 60736 -25050
rect 60616 -25100 60626 -25060
rect 60626 -25100 60666 -25060
rect 60666 -25100 60736 -25060
rect 60616 -25110 60736 -25100
rect 60756 -25060 60816 -25050
rect 60756 -25100 60766 -25060
rect 60766 -25100 60806 -25060
rect 60806 -25100 60816 -25060
rect 60756 -25110 60816 -25100
rect 60896 -25060 60956 -25050
rect 60896 -25100 60906 -25060
rect 60906 -25100 60946 -25060
rect 60946 -25100 60956 -25060
rect 60896 -25110 60956 -25100
rect 56380 -25488 56440 -25368
rect 55880 -25680 55970 -25678
rect 55880 -25714 55882 -25680
rect 55882 -25714 55970 -25680
rect 55880 -25758 55970 -25714
rect 55220 -26128 55330 -26018
rect 55530 -26202 55610 -26178
rect 55530 -26236 55560 -26202
rect 55560 -26236 55610 -26202
rect 55530 -26268 55610 -26236
rect 54140 -26308 54150 -26288
rect 54150 -26308 54840 -26288
rect 54840 -26308 54850 -26288
rect 26600 -30400 35200 -26400
rect 54140 -26548 54850 -26308
rect 55320 -26348 55470 -26328
rect 55320 -26408 55470 -26348
rect 55320 -26468 55470 -26408
rect 56020 -26008 56080 -25858
rect 56170 -26008 56390 -25808
rect 56654 -26086 56998 -25868
rect 59076 -25370 59103 -25340
rect 59103 -25370 59137 -25340
rect 59137 -25370 59166 -25340
rect 59076 -25400 59166 -25370
rect 58926 -25510 58986 -25460
rect 58926 -25530 58966 -25510
rect 58966 -25530 58986 -25510
rect 59146 -25530 59226 -25460
rect 59276 -25530 59356 -25460
rect 59396 -25530 59476 -25460
rect 59646 -25520 59706 -25460
rect 59546 -25608 59606 -25600
rect 59256 -25662 59366 -25630
rect 59546 -25642 59560 -25608
rect 59560 -25642 59594 -25608
rect 59594 -25642 59606 -25608
rect 59016 -25716 59076 -25700
rect 59256 -25690 59366 -25662
rect 59546 -25660 59606 -25642
rect 59016 -25750 59032 -25716
rect 59032 -25750 59066 -25716
rect 59066 -25750 59076 -25716
rect 59016 -25760 59076 -25750
rect 58906 -25900 58926 -25830
rect 58926 -25900 58966 -25830
rect 58966 -25900 58986 -25830
rect 59146 -25900 59226 -25830
rect 59276 -25900 59356 -25830
rect 59396 -25900 59476 -25830
rect 59966 -25340 60326 -25320
rect 59966 -25374 60326 -25340
rect 59966 -25380 60326 -25374
rect 59856 -25394 59916 -25380
rect 59856 -25428 59874 -25394
rect 59874 -25428 59908 -25394
rect 59908 -25428 59916 -25394
rect 59856 -25440 59916 -25428
rect 60376 -25394 60436 -25380
rect 60376 -25428 60384 -25394
rect 60384 -25428 60418 -25394
rect 60418 -25428 60436 -25394
rect 60376 -25440 60436 -25428
rect 61056 -25440 61126 -25340
rect 59806 -25720 59916 -25610
rect 60446 -25750 60526 -25630
rect 59646 -25900 59706 -25840
rect 58986 -26360 59126 -26220
rect 59996 -26300 60106 -26190
rect 59700 -26800 60400 -26400
rect 55500 -27300 56100 -26900
rect 55460 -28160 55720 -27880
rect 53480 -28740 53780 -28540
rect 54150 -28508 54860 -28338
rect 54150 -28578 54850 -28508
rect 54850 -28578 54860 -28508
rect 53520 -28968 53640 -28858
rect 54750 -28908 54850 -28838
rect 54750 -28918 54840 -28908
rect 55430 -28888 55520 -28818
rect 55290 -28998 55390 -28928
rect 15000 -49000 24000 -38000
rect 53050 -30908 53250 -29158
rect 53950 -29128 53998 -29098
rect 53998 -29128 54020 -29098
rect 53950 -29198 54020 -29128
rect 54920 -29090 54990 -29078
rect 54920 -29128 54926 -29090
rect 54926 -29128 54960 -29090
rect 54960 -29128 54990 -29090
rect 54920 -29168 54990 -29128
rect 53860 -29638 53920 -29528
rect 55230 -29428 55290 -29258
rect 55290 -29428 55320 -29258
rect 55430 -29418 55510 -29248
rect 55960 -28888 56040 -28738
rect 56190 -28968 56390 -28758
rect 56506 -28830 57016 -28580
rect 58966 -28630 59126 -28470
rect 59956 -28660 60166 -28500
rect 55880 -29056 55970 -29018
rect 55880 -29090 55882 -29056
rect 55882 -29090 55970 -29056
rect 55880 -29098 55970 -29090
rect 55000 -29638 55090 -29538
rect 54770 -29840 54840 -29838
rect 54770 -29928 54802 -29840
rect 54802 -29928 54840 -29840
rect 55540 -29638 55630 -29538
rect 56590 -29398 56660 -29268
rect 58906 -29020 58966 -28970
rect 58906 -29030 58926 -29020
rect 58926 -29030 58966 -29020
rect 59216 -29030 59276 -28970
rect 59326 -29030 59386 -28970
rect 59436 -29030 59496 -28970
rect 59636 -29030 59696 -28970
rect 59546 -29101 59606 -29090
rect 59286 -29155 59346 -29130
rect 59546 -29135 59560 -29101
rect 59560 -29135 59594 -29101
rect 59594 -29135 59606 -29101
rect 59286 -29189 59346 -29155
rect 59546 -29150 59606 -29135
rect 59286 -29190 59346 -29189
rect 59016 -29209 59076 -29200
rect 59016 -29243 59032 -29209
rect 59032 -29243 59066 -29209
rect 59066 -29243 59076 -29209
rect 59016 -29260 59076 -29243
rect 59546 -29270 59606 -29210
rect 58906 -29390 58966 -29330
rect 59216 -29380 59276 -29320
rect 59336 -29380 59396 -29320
rect 59436 -29380 59496 -29320
rect 55140 -30008 55200 -29938
rect 55030 -30128 55110 -30048
rect 55740 -30128 55810 -30048
rect 55880 -30128 55970 -30038
rect 56480 -29606 56550 -29588
rect 56480 -29640 56492 -29606
rect 56492 -29640 56530 -29606
rect 56530 -29640 56550 -29606
rect 56480 -29648 56550 -29640
rect 59866 -29230 59966 -29140
rect 60446 -29220 60526 -29120
rect 59636 -29390 59696 -29330
rect 59076 -29478 59166 -29440
rect 59076 -29510 59103 -29478
rect 59103 -29510 59137 -29478
rect 59137 -29510 59166 -29478
rect 60046 -29374 60126 -29340
rect 59856 -29428 59916 -29410
rect 60046 -29400 60126 -29374
rect 59856 -29462 59874 -29428
rect 59874 -29462 59908 -29428
rect 59908 -29462 59916 -29428
rect 59856 -29480 59916 -29462
rect 60376 -29428 60446 -29420
rect 60376 -29462 60384 -29428
rect 60384 -29462 60418 -29428
rect 60418 -29462 60446 -29428
rect 59976 -29516 60316 -29500
rect 60376 -29480 60446 -29462
rect 57098 -29589 57368 -29564
rect 57098 -29623 57125 -29589
rect 57125 -29623 57159 -29589
rect 57159 -29623 57217 -29589
rect 57217 -29623 57251 -29589
rect 57251 -29623 57309 -29589
rect 57309 -29623 57343 -29589
rect 57343 -29623 57368 -29589
rect 54770 -30328 54802 -30248
rect 54802 -30328 54840 -30248
rect 53850 -30648 53920 -30538
rect 54920 -30468 54980 -30398
rect 55000 -30638 55090 -30538
rect 55540 -30638 55630 -30538
rect 55220 -30918 55280 -30748
rect 55280 -30918 55310 -30748
rect 55410 -30928 55500 -30758
rect 53950 -31050 54010 -31008
rect 53950 -31088 53988 -31050
rect 53988 -31088 54010 -31050
rect 54910 -31050 54980 -30998
rect 54910 -31088 54916 -31050
rect 54916 -31088 54950 -31050
rect 54950 -31088 54980 -31050
rect 54910 -31098 54980 -31088
rect 53510 -31248 53630 -31128
rect 54740 -31344 54850 -31268
rect 54740 -31358 54850 -31344
rect 55240 -31218 55370 -31158
rect 55410 -31338 55510 -31248
rect 57098 -29680 57368 -29623
rect 57098 -29704 57368 -29680
rect 56900 -30148 57020 -30018
rect 58576 -30240 58736 -30080
rect 57098 -30480 57368 -30474
rect 56480 -30534 56550 -30528
rect 56480 -30568 56492 -30534
rect 56492 -30568 56530 -30534
rect 56530 -30568 56550 -30534
rect 56480 -30588 56550 -30568
rect 57098 -30565 57368 -30480
rect 57098 -30599 57125 -30565
rect 57125 -30599 57159 -30565
rect 57159 -30599 57217 -30565
rect 57217 -30599 57251 -30565
rect 57251 -30599 57309 -30565
rect 57309 -30599 57343 -30565
rect 57343 -30599 57368 -30565
rect 57098 -30614 57368 -30599
rect 59976 -29552 60316 -29516
rect 59176 -29720 59196 -29640
rect 59196 -29720 59236 -29640
rect 59176 -29920 59196 -29840
rect 59196 -29920 59236 -29840
rect 59076 -30040 59103 -30010
rect 59103 -30040 59137 -30010
rect 59137 -30040 59166 -30010
rect 59076 -30080 59166 -30040
rect 59576 -29698 59636 -29670
rect 59576 -29730 59580 -29698
rect 59580 -29730 59636 -29698
rect 59476 -29920 59502 -29850
rect 59502 -29920 59536 -29850
rect 59576 -29958 59590 -29790
rect 59590 -29958 59624 -29790
rect 59624 -29958 59636 -29790
rect 59576 -29960 59636 -29958
rect 59076 -30208 59166 -30170
rect 59076 -30240 59103 -30208
rect 59103 -30240 59137 -30208
rect 59137 -30240 59166 -30208
rect 59206 -30240 59266 -30170
rect 61206 -29700 61346 -29520
rect 59806 -29940 59818 -29800
rect 59818 -29940 59852 -29800
rect 59852 -29940 59866 -29800
rect 59916 -29782 60006 -29780
rect 59916 -29958 59940 -29782
rect 59940 -29958 60006 -29782
rect 59916 -29960 60006 -29958
rect 60306 -29890 60456 -29750
rect 59826 -30042 59862 -30010
rect 59862 -30042 59896 -30010
rect 59896 -30042 59916 -30010
rect 59826 -30080 59916 -30042
rect 59166 -30410 59196 -30330
rect 59196 -30410 59226 -30330
rect 59166 -30640 59196 -30560
rect 59196 -30640 59226 -30560
rect 59466 -30410 59501 -30330
rect 59501 -30410 59526 -30330
rect 59586 -30450 59589 -30310
rect 59589 -30450 59623 -30310
rect 59623 -30450 59646 -30310
rect 59516 -30521 59596 -30520
rect 59516 -30555 59545 -30521
rect 59545 -30555 59579 -30521
rect 59579 -30555 59596 -30521
rect 59516 -30580 59596 -30555
rect 59826 -30211 59926 -30170
rect 59826 -30240 59861 -30211
rect 59861 -30240 59895 -30211
rect 59895 -30240 59926 -30211
rect 60096 -30083 60127 -30080
rect 60127 -30083 60161 -30080
rect 60161 -30083 60176 -30080
rect 60096 -30141 60176 -30083
rect 60096 -30175 60127 -30141
rect 60127 -30175 60161 -30141
rect 60161 -30175 60176 -30141
rect 60096 -30233 60176 -30175
rect 60096 -30240 60127 -30233
rect 60127 -30240 60161 -30233
rect 60161 -30240 60176 -30233
rect 59796 -30295 59856 -30290
rect 59796 -30470 59817 -30295
rect 59817 -30470 59851 -30295
rect 59851 -30470 59856 -30295
rect 59916 -30295 60006 -30290
rect 59916 -30471 59939 -30295
rect 59939 -30471 60006 -30295
rect 59916 -30480 60006 -30471
rect 60476 -30325 60536 -30310
rect 60476 -30359 60484 -30325
rect 60484 -30359 60536 -30325
rect 60476 -30370 60536 -30359
rect 61036 -29930 61126 -29820
rect 61276 -30083 61291 -30050
rect 61291 -30083 61325 -30050
rect 61325 -30083 61356 -30050
rect 61276 -30141 61356 -30083
rect 61276 -30175 61291 -30141
rect 61291 -30175 61325 -30141
rect 61325 -30175 61356 -30141
rect 61276 -30233 61356 -30175
rect 61276 -30260 61291 -30233
rect 61291 -30260 61325 -30233
rect 61325 -30260 61356 -30233
rect 60476 -30460 60536 -30450
rect 60476 -30500 60486 -30460
rect 60486 -30500 60526 -30460
rect 60526 -30500 60536 -30460
rect 60476 -30510 60536 -30500
rect 60616 -30460 60736 -30450
rect 60616 -30500 60626 -30460
rect 60626 -30500 60666 -30460
rect 60666 -30500 60736 -30460
rect 60616 -30510 60736 -30500
rect 60756 -30460 60816 -30450
rect 60756 -30500 60766 -30460
rect 60766 -30500 60806 -30460
rect 60806 -30500 60816 -30460
rect 60756 -30510 60816 -30500
rect 60896 -30460 60956 -30450
rect 60896 -30500 60906 -30460
rect 60906 -30500 60946 -30460
rect 60946 -30500 60956 -30460
rect 60896 -30510 60956 -30500
rect 56380 -30888 56440 -30768
rect 55880 -31080 55970 -31078
rect 55880 -31114 55882 -31080
rect 55882 -31114 55970 -31080
rect 55880 -31158 55970 -31114
rect 55220 -31528 55330 -31418
rect 55530 -31602 55610 -31578
rect 55530 -31636 55560 -31602
rect 55560 -31636 55610 -31602
rect 55530 -31668 55610 -31636
rect 54140 -31708 54150 -31688
rect 54150 -31708 54840 -31688
rect 54840 -31708 54850 -31688
rect 54140 -31948 54850 -31708
rect 55320 -31748 55470 -31728
rect 55320 -31808 55470 -31748
rect 55320 -31868 55470 -31808
rect 56020 -31408 56080 -31258
rect 56170 -31408 56390 -31208
rect 56654 -31486 56998 -31268
rect 59076 -30770 59103 -30740
rect 59103 -30770 59137 -30740
rect 59137 -30770 59166 -30740
rect 59076 -30800 59166 -30770
rect 58926 -30910 58986 -30860
rect 58926 -30930 58966 -30910
rect 58966 -30930 58986 -30910
rect 59146 -30930 59226 -30860
rect 59276 -30930 59356 -30860
rect 59396 -30930 59476 -30860
rect 59646 -30920 59706 -30860
rect 59546 -31008 59606 -31000
rect 59256 -31062 59366 -31030
rect 59546 -31042 59560 -31008
rect 59560 -31042 59594 -31008
rect 59594 -31042 59606 -31008
rect 59016 -31116 59076 -31100
rect 59256 -31090 59366 -31062
rect 59546 -31060 59606 -31042
rect 59016 -31150 59032 -31116
rect 59032 -31150 59066 -31116
rect 59066 -31150 59076 -31116
rect 59016 -31160 59076 -31150
rect 58906 -31300 58926 -31230
rect 58926 -31300 58966 -31230
rect 58966 -31300 58986 -31230
rect 59146 -31300 59226 -31230
rect 59276 -31300 59356 -31230
rect 59396 -31300 59476 -31230
rect 59966 -30740 60326 -30720
rect 59966 -30774 60326 -30740
rect 59966 -30780 60326 -30774
rect 59856 -30794 59916 -30780
rect 59856 -30828 59874 -30794
rect 59874 -30828 59908 -30794
rect 59908 -30828 59916 -30794
rect 59856 -30840 59916 -30828
rect 60376 -30794 60436 -30780
rect 60376 -30828 60384 -30794
rect 60384 -30828 60418 -30794
rect 60418 -30828 60436 -30794
rect 60376 -30840 60436 -30828
rect 61056 -30840 61126 -30740
rect 59806 -31120 59916 -31010
rect 60446 -31150 60526 -31030
rect 59646 -31300 59706 -31240
rect 58986 -31760 59126 -31620
rect 59996 -31700 60106 -31590
rect 59800 -32100 60300 -31800
rect 36200 -33000 36800 -32200
rect 55500 -32700 56100 -32300
rect 55460 -33560 55720 -33280
rect 36000 -34700 38100 -33700
rect 53480 -34140 53780 -33940
rect 54150 -33908 54860 -33738
rect 54150 -33978 54850 -33908
rect 54850 -33978 54860 -33908
rect 53520 -34368 53640 -34258
rect 54750 -34308 54850 -34238
rect 54750 -34318 54840 -34308
rect 55430 -34288 55520 -34218
rect 55290 -34398 55390 -34328
rect 36000 -36300 39000 -35300
rect 53050 -36308 53250 -34558
rect 53950 -34528 53998 -34498
rect 53998 -34528 54020 -34498
rect 53950 -34598 54020 -34528
rect 54920 -34490 54990 -34478
rect 54920 -34528 54926 -34490
rect 54926 -34528 54960 -34490
rect 54960 -34528 54990 -34490
rect 54920 -34568 54990 -34528
rect 53860 -35038 53920 -34928
rect 55230 -34828 55290 -34658
rect 55290 -34828 55320 -34658
rect 55430 -34818 55510 -34648
rect 55960 -34288 56040 -34138
rect 56190 -34368 56390 -34158
rect 56506 -34230 57016 -33980
rect 58966 -34030 59126 -33870
rect 59956 -34060 60166 -33900
rect 55880 -34456 55970 -34418
rect 55880 -34490 55882 -34456
rect 55882 -34490 55970 -34456
rect 55880 -34498 55970 -34490
rect 55000 -35038 55090 -34938
rect 54770 -35240 54840 -35238
rect 54770 -35328 54802 -35240
rect 54802 -35328 54840 -35240
rect 55540 -35038 55630 -34938
rect 56590 -34798 56660 -34668
rect 58906 -34420 58966 -34370
rect 58906 -34430 58926 -34420
rect 58926 -34430 58966 -34420
rect 59216 -34430 59276 -34370
rect 59326 -34430 59386 -34370
rect 59436 -34430 59496 -34370
rect 59636 -34430 59696 -34370
rect 59546 -34501 59606 -34490
rect 59286 -34555 59346 -34530
rect 59546 -34535 59560 -34501
rect 59560 -34535 59594 -34501
rect 59594 -34535 59606 -34501
rect 59286 -34589 59346 -34555
rect 59546 -34550 59606 -34535
rect 59286 -34590 59346 -34589
rect 59016 -34609 59076 -34600
rect 59016 -34643 59032 -34609
rect 59032 -34643 59066 -34609
rect 59066 -34643 59076 -34609
rect 59016 -34660 59076 -34643
rect 59546 -34670 59606 -34610
rect 58906 -34790 58966 -34730
rect 59216 -34780 59276 -34720
rect 59336 -34780 59396 -34720
rect 59436 -34780 59496 -34720
rect 55140 -35408 55200 -35338
rect 55030 -35528 55110 -35448
rect 55740 -35528 55810 -35448
rect 55880 -35528 55970 -35438
rect 56480 -35006 56550 -34988
rect 56480 -35040 56492 -35006
rect 56492 -35040 56530 -35006
rect 56530 -35040 56550 -35006
rect 56480 -35048 56550 -35040
rect 59866 -34630 59966 -34540
rect 60446 -34620 60526 -34520
rect 59636 -34790 59696 -34730
rect 59076 -34878 59166 -34840
rect 59076 -34910 59103 -34878
rect 59103 -34910 59137 -34878
rect 59137 -34910 59166 -34878
rect 60046 -34774 60126 -34740
rect 59856 -34828 59916 -34810
rect 60046 -34800 60126 -34774
rect 59856 -34862 59874 -34828
rect 59874 -34862 59908 -34828
rect 59908 -34862 59916 -34828
rect 59856 -34880 59916 -34862
rect 60376 -34828 60446 -34820
rect 60376 -34862 60384 -34828
rect 60384 -34862 60418 -34828
rect 60418 -34862 60446 -34828
rect 59976 -34916 60316 -34900
rect 60376 -34880 60446 -34862
rect 57098 -34989 57368 -34964
rect 57098 -35023 57125 -34989
rect 57125 -35023 57159 -34989
rect 57159 -35023 57217 -34989
rect 57217 -35023 57251 -34989
rect 57251 -35023 57309 -34989
rect 57309 -35023 57343 -34989
rect 57343 -35023 57368 -34989
rect 54770 -35728 54802 -35648
rect 54802 -35728 54840 -35648
rect 53850 -36048 53920 -35938
rect 54920 -35868 54980 -35798
rect 55000 -36038 55090 -35938
rect 55540 -36038 55630 -35938
rect 55220 -36318 55280 -36148
rect 55280 -36318 55310 -36148
rect 55410 -36328 55500 -36158
rect 53950 -36450 54010 -36408
rect 53950 -36488 53988 -36450
rect 53988 -36488 54010 -36450
rect 54910 -36450 54980 -36398
rect 54910 -36488 54916 -36450
rect 54916 -36488 54950 -36450
rect 54950 -36488 54980 -36450
rect 54910 -36498 54980 -36488
rect 53510 -36648 53630 -36528
rect 54740 -36744 54850 -36668
rect 54740 -36758 54850 -36744
rect 55240 -36618 55370 -36558
rect 55410 -36738 55510 -36648
rect 57098 -35080 57368 -35023
rect 57098 -35104 57368 -35080
rect 56900 -35548 57020 -35418
rect 58576 -35640 58736 -35480
rect 57098 -35880 57368 -35874
rect 56480 -35934 56550 -35928
rect 56480 -35968 56492 -35934
rect 56492 -35968 56530 -35934
rect 56530 -35968 56550 -35934
rect 56480 -35988 56550 -35968
rect 57098 -35965 57368 -35880
rect 57098 -35999 57125 -35965
rect 57125 -35999 57159 -35965
rect 57159 -35999 57217 -35965
rect 57217 -35999 57251 -35965
rect 57251 -35999 57309 -35965
rect 57309 -35999 57343 -35965
rect 57343 -35999 57368 -35965
rect 57098 -36014 57368 -35999
rect 59976 -34952 60316 -34916
rect 59176 -35120 59196 -35040
rect 59196 -35120 59236 -35040
rect 59176 -35320 59196 -35240
rect 59196 -35320 59236 -35240
rect 59076 -35440 59103 -35410
rect 59103 -35440 59137 -35410
rect 59137 -35440 59166 -35410
rect 59076 -35480 59166 -35440
rect 59576 -35098 59636 -35070
rect 59576 -35130 59580 -35098
rect 59580 -35130 59636 -35098
rect 59476 -35320 59502 -35250
rect 59502 -35320 59536 -35250
rect 59576 -35358 59590 -35190
rect 59590 -35358 59624 -35190
rect 59624 -35358 59636 -35190
rect 59576 -35360 59636 -35358
rect 59076 -35608 59166 -35570
rect 59076 -35640 59103 -35608
rect 59103 -35640 59137 -35608
rect 59137 -35640 59166 -35608
rect 59206 -35640 59266 -35570
rect 61206 -35100 61346 -34920
rect 59806 -35340 59818 -35200
rect 59818 -35340 59852 -35200
rect 59852 -35340 59866 -35200
rect 59916 -35182 60006 -35180
rect 59916 -35358 59940 -35182
rect 59940 -35358 60006 -35182
rect 59916 -35360 60006 -35358
rect 60306 -35290 60456 -35150
rect 59826 -35442 59862 -35410
rect 59862 -35442 59896 -35410
rect 59896 -35442 59916 -35410
rect 59826 -35480 59916 -35442
rect 59166 -35810 59196 -35730
rect 59196 -35810 59226 -35730
rect 59166 -36040 59196 -35960
rect 59196 -36040 59226 -35960
rect 59466 -35810 59501 -35730
rect 59501 -35810 59526 -35730
rect 59586 -35850 59589 -35710
rect 59589 -35850 59623 -35710
rect 59623 -35850 59646 -35710
rect 59516 -35921 59596 -35920
rect 59516 -35955 59545 -35921
rect 59545 -35955 59579 -35921
rect 59579 -35955 59596 -35921
rect 59516 -35980 59596 -35955
rect 59826 -35611 59926 -35570
rect 59826 -35640 59861 -35611
rect 59861 -35640 59895 -35611
rect 59895 -35640 59926 -35611
rect 60096 -35483 60127 -35480
rect 60127 -35483 60161 -35480
rect 60161 -35483 60176 -35480
rect 60096 -35541 60176 -35483
rect 60096 -35575 60127 -35541
rect 60127 -35575 60161 -35541
rect 60161 -35575 60176 -35541
rect 60096 -35633 60176 -35575
rect 60096 -35640 60127 -35633
rect 60127 -35640 60161 -35633
rect 60161 -35640 60176 -35633
rect 59796 -35695 59856 -35690
rect 59796 -35870 59817 -35695
rect 59817 -35870 59851 -35695
rect 59851 -35870 59856 -35695
rect 59916 -35695 60006 -35690
rect 59916 -35871 59939 -35695
rect 59939 -35871 60006 -35695
rect 59916 -35880 60006 -35871
rect 60476 -35725 60536 -35710
rect 60476 -35759 60484 -35725
rect 60484 -35759 60536 -35725
rect 60476 -35770 60536 -35759
rect 61036 -35330 61126 -35220
rect 61276 -35483 61291 -35450
rect 61291 -35483 61325 -35450
rect 61325 -35483 61356 -35450
rect 61276 -35541 61356 -35483
rect 61276 -35575 61291 -35541
rect 61291 -35575 61325 -35541
rect 61325 -35575 61356 -35541
rect 61276 -35633 61356 -35575
rect 61276 -35660 61291 -35633
rect 61291 -35660 61325 -35633
rect 61325 -35660 61356 -35633
rect 72000 -35500 74000 -34100
rect 60476 -35860 60536 -35850
rect 60476 -35900 60486 -35860
rect 60486 -35900 60526 -35860
rect 60526 -35900 60536 -35860
rect 60476 -35910 60536 -35900
rect 60616 -35860 60736 -35850
rect 60616 -35900 60626 -35860
rect 60626 -35900 60666 -35860
rect 60666 -35900 60736 -35860
rect 60616 -35910 60736 -35900
rect 60756 -35860 60816 -35850
rect 60756 -35900 60766 -35860
rect 60766 -35900 60806 -35860
rect 60806 -35900 60816 -35860
rect 60756 -35910 60816 -35900
rect 60896 -35860 60956 -35850
rect 60896 -35900 60906 -35860
rect 60906 -35900 60946 -35860
rect 60946 -35900 60956 -35860
rect 60896 -35910 60956 -35900
rect 56380 -36288 56440 -36168
rect 55880 -36480 55970 -36478
rect 55880 -36514 55882 -36480
rect 55882 -36514 55970 -36480
rect 55880 -36558 55970 -36514
rect 36000 -37900 40000 -36900
rect 55220 -36928 55330 -36818
rect 55530 -37002 55610 -36978
rect 55530 -37036 55560 -37002
rect 55560 -37036 55610 -37002
rect 55530 -37068 55610 -37036
rect 54140 -37108 54150 -37088
rect 54150 -37108 54840 -37088
rect 54840 -37108 54850 -37088
rect 54140 -37348 54850 -37108
rect 55320 -37148 55470 -37128
rect 55320 -37208 55470 -37148
rect 55320 -37268 55470 -37208
rect 56020 -36808 56080 -36658
rect 56170 -36808 56390 -36608
rect 56654 -36886 56998 -36668
rect 59076 -36170 59103 -36140
rect 59103 -36170 59137 -36140
rect 59137 -36170 59166 -36140
rect 59076 -36200 59166 -36170
rect 58926 -36310 58986 -36260
rect 58926 -36330 58966 -36310
rect 58966 -36330 58986 -36310
rect 59146 -36330 59226 -36260
rect 59276 -36330 59356 -36260
rect 59396 -36330 59476 -36260
rect 59646 -36320 59706 -36260
rect 59546 -36408 59606 -36400
rect 59256 -36462 59366 -36430
rect 59546 -36442 59560 -36408
rect 59560 -36442 59594 -36408
rect 59594 -36442 59606 -36408
rect 59016 -36516 59076 -36500
rect 59256 -36490 59366 -36462
rect 59546 -36460 59606 -36442
rect 59016 -36550 59032 -36516
rect 59032 -36550 59066 -36516
rect 59066 -36550 59076 -36516
rect 59016 -36560 59076 -36550
rect 58906 -36700 58926 -36630
rect 58926 -36700 58966 -36630
rect 58966 -36700 58986 -36630
rect 59146 -36700 59226 -36630
rect 59276 -36700 59356 -36630
rect 59396 -36700 59476 -36630
rect 59966 -36140 60326 -36120
rect 59966 -36174 60326 -36140
rect 59966 -36180 60326 -36174
rect 59856 -36194 59916 -36180
rect 59856 -36228 59874 -36194
rect 59874 -36228 59908 -36194
rect 59908 -36228 59916 -36194
rect 59856 -36240 59916 -36228
rect 60376 -36194 60436 -36180
rect 60376 -36228 60384 -36194
rect 60384 -36228 60418 -36194
rect 60418 -36228 60436 -36194
rect 60376 -36240 60436 -36228
rect 61056 -36240 61126 -36140
rect 59806 -36520 59916 -36410
rect 60446 -36550 60526 -36430
rect 59646 -36700 59706 -36640
rect 58986 -37160 59126 -37020
rect 59996 -37100 60106 -36990
rect 59900 -37400 60200 -37200
rect 55400 -38100 56100 -37700
rect 36000 -39500 41000 -38500
rect 73220 -38550 73340 -38360
rect 73470 -38550 73590 -38360
rect 73720 -38550 73840 -38360
rect 73970 -38550 74090 -38360
rect 74220 -38550 74340 -38360
rect 74470 -38550 74590 -38360
rect 74720 -38550 74840 -38360
rect 74970 -38550 75090 -38360
rect 75390 -38270 75550 -38150
rect 75220 -38550 75340 -38360
rect 73723 -38648 73840 -38596
rect 75410 -38650 75470 -38590
rect 75673 -38609 75751 -38583
rect 75673 -38643 75704 -38609
rect 75704 -38643 75751 -38609
rect 75673 -38661 75751 -38643
rect 55460 -38960 55720 -38680
rect 75946 -38609 76024 -38583
rect 75946 -38643 75947 -38609
rect 75947 -38643 75981 -38609
rect 75981 -38643 76024 -38609
rect 75946 -38661 76024 -38643
rect 72820 -38920 73040 -38740
rect 74220 -38840 74340 -38760
rect 76102 -38610 76167 -38583
rect 76920 -38530 77060 -38410
rect 84960 -38480 85400 -38050
rect 76102 -38644 76128 -38610
rect 76128 -38644 76162 -38610
rect 76162 -38644 76167 -38610
rect 76102 -38661 76167 -38644
rect 76232 -38610 76310 -38583
rect 76232 -38644 76258 -38610
rect 76258 -38644 76310 -38610
rect 76232 -38661 76310 -38644
rect 76380 -38609 76440 -38600
rect 76380 -38643 76404 -38609
rect 76404 -38643 76438 -38609
rect 76438 -38643 76440 -38609
rect 76380 -38660 76440 -38643
rect 76505 -38609 76583 -38596
rect 76505 -38643 76531 -38609
rect 76531 -38643 76583 -38609
rect 76505 -38661 76583 -38643
rect 76648 -38609 76726 -38596
rect 76648 -38643 76680 -38609
rect 76680 -38643 76714 -38609
rect 76714 -38643 76726 -38609
rect 76648 -38674 76726 -38643
rect 76791 -38610 76843 -38596
rect 76791 -38644 76806 -38610
rect 76806 -38644 76843 -38610
rect 76791 -38674 76843 -38644
rect 77170 -39040 77430 -38790
rect 53480 -39540 53780 -39340
rect 54150 -39308 54860 -39138
rect 54150 -39378 54850 -39308
rect 54850 -39378 54860 -39308
rect 53520 -39768 53640 -39658
rect 54750 -39708 54850 -39638
rect 54750 -39718 54840 -39708
rect 55430 -39688 55520 -39618
rect 55290 -39798 55390 -39728
rect 36000 -41100 42100 -40100
rect 36000 -42700 43100 -41700
rect 53050 -41708 53250 -39958
rect 53950 -39928 53998 -39898
rect 53998 -39928 54020 -39898
rect 53950 -39998 54020 -39928
rect 54920 -39890 54990 -39878
rect 54920 -39928 54926 -39890
rect 54926 -39928 54960 -39890
rect 54960 -39928 54990 -39890
rect 54920 -39968 54990 -39928
rect 53860 -40438 53920 -40328
rect 55230 -40228 55290 -40058
rect 55290 -40228 55320 -40058
rect 55430 -40218 55510 -40048
rect 55960 -39688 56040 -39538
rect 56190 -39768 56390 -39558
rect 56506 -39630 57016 -39380
rect 58966 -39430 59126 -39270
rect 72820 -39250 73040 -39070
rect 73480 -39180 73580 -39120
rect 88150 -38820 88590 -38390
rect 73730 -39290 73830 -39230
rect 59956 -39460 60166 -39300
rect 73230 -39400 73330 -39340
rect 78150 -39350 78210 -39340
rect 78150 -39390 78160 -39350
rect 78160 -39390 78200 -39350
rect 78200 -39390 78210 -39350
rect 78150 -39400 78210 -39390
rect 78280 -39350 78340 -39340
rect 78280 -39390 78290 -39350
rect 78290 -39390 78330 -39350
rect 78330 -39390 78340 -39350
rect 78580 -39330 78640 -39320
rect 78580 -39370 78590 -39330
rect 78590 -39370 78630 -39330
rect 78630 -39370 78640 -39330
rect 78580 -39380 78640 -39370
rect 78800 -39340 78860 -39330
rect 78800 -39380 78850 -39340
rect 78850 -39380 78860 -39340
rect 78800 -39390 78860 -39380
rect 78280 -39400 78340 -39390
rect 55880 -39856 55970 -39818
rect 55880 -39890 55882 -39856
rect 55882 -39890 55970 -39856
rect 55880 -39898 55970 -39890
rect 55000 -40438 55090 -40338
rect 54770 -40640 54840 -40638
rect 54770 -40728 54802 -40640
rect 54802 -40728 54840 -40640
rect 55540 -40438 55630 -40338
rect 56590 -40198 56660 -40068
rect 77230 -39450 77310 -39440
rect 77230 -39490 77240 -39450
rect 77240 -39490 77300 -39450
rect 77300 -39490 77310 -39450
rect 77230 -39500 77310 -39490
rect 58906 -39820 58966 -39770
rect 58906 -39830 58926 -39820
rect 58926 -39830 58966 -39820
rect 59216 -39830 59276 -39770
rect 59326 -39830 59386 -39770
rect 59436 -39830 59496 -39770
rect 72820 -39740 73040 -39560
rect 76920 -39720 77060 -39570
rect 79080 -39400 79140 -39350
rect 79140 -39400 79250 -39350
rect 79080 -39450 79250 -39400
rect 79080 -39510 79140 -39450
rect 79140 -39510 79250 -39450
rect 80080 -39580 80430 -39270
rect 82780 -39280 82820 -39270
rect 82820 -39280 82890 -39270
rect 82780 -39320 82890 -39280
rect 82780 -39360 82820 -39320
rect 82820 -39360 82890 -39320
rect 82780 -39400 82890 -39360
rect 82780 -39440 82820 -39400
rect 82820 -39440 82890 -39400
rect 82780 -39490 82890 -39440
rect 82780 -39520 82820 -39490
rect 82820 -39520 82890 -39490
rect 83370 -39394 83770 -39380
rect 83370 -39434 83770 -39394
rect 83370 -39450 83770 -39434
rect 84230 -39260 84310 -39250
rect 84230 -39530 84250 -39260
rect 84250 -39530 84290 -39260
rect 84290 -39530 84310 -39260
rect 84230 -39540 84310 -39530
rect 84870 -39397 85240 -39380
rect 84870 -39437 85240 -39397
rect 84870 -39450 85240 -39437
rect 85710 -39270 85790 -39260
rect 85710 -39540 85730 -39270
rect 85730 -39540 85770 -39270
rect 85770 -39540 85790 -39270
rect 85710 -39550 85790 -39540
rect 86320 -39394 86710 -39380
rect 86320 -39434 86329 -39394
rect 86329 -39434 86699 -39394
rect 86699 -39434 86710 -39394
rect 86320 -39450 86710 -39434
rect 87180 -39510 87200 -39240
rect 87200 -39510 87240 -39240
rect 87240 -39510 87260 -39240
rect 87450 -39395 87760 -39380
rect 87450 -39435 87469 -39395
rect 87469 -39435 87749 -39395
rect 87749 -39435 87760 -39395
rect 87450 -39450 87760 -39435
rect 88650 -39260 88730 -39250
rect 88650 -39530 88670 -39260
rect 88670 -39530 88710 -39260
rect 88710 -39530 88730 -39260
rect 88650 -39540 88730 -39530
rect 59636 -39830 59696 -39770
rect 59546 -39901 59606 -39890
rect 59286 -39955 59346 -39930
rect 59546 -39935 59560 -39901
rect 59560 -39935 59594 -39901
rect 59594 -39935 59606 -39901
rect 59286 -39989 59346 -39955
rect 59546 -39950 59606 -39935
rect 59286 -39990 59346 -39989
rect 59016 -40009 59076 -40000
rect 59016 -40043 59032 -40009
rect 59032 -40043 59066 -40009
rect 59066 -40043 59076 -40009
rect 59016 -40060 59076 -40043
rect 59546 -40070 59606 -40010
rect 58906 -40190 58966 -40130
rect 59216 -40180 59276 -40120
rect 59336 -40180 59396 -40120
rect 59436 -40180 59496 -40120
rect 55140 -40808 55200 -40738
rect 55030 -40928 55110 -40848
rect 55740 -40928 55810 -40848
rect 55880 -40928 55970 -40838
rect 56480 -40406 56550 -40388
rect 56480 -40440 56492 -40406
rect 56492 -40440 56530 -40406
rect 56530 -40440 56550 -40406
rect 56480 -40448 56550 -40440
rect 59866 -40030 59966 -39940
rect 60446 -40020 60526 -39920
rect 72820 -40020 73040 -39840
rect 77170 -39790 77260 -39780
rect 77170 -39840 77260 -39790
rect 77170 -39850 77260 -39840
rect 74230 -39950 74330 -39890
rect 74730 -40040 74830 -39980
rect 59636 -40190 59696 -40130
rect 78150 -39830 78160 -39790
rect 78160 -39830 78200 -39790
rect 78200 -39830 78210 -39790
rect 78150 -39900 78210 -39830
rect 78150 -39940 78160 -39900
rect 78160 -39940 78200 -39900
rect 78200 -39940 78210 -39900
rect 78150 -40020 78210 -39940
rect 78150 -40060 78160 -40020
rect 78160 -40060 78200 -40020
rect 78200 -40060 78210 -40020
rect 78150 -40080 78210 -40060
rect 80080 -40060 80430 -39680
rect 59076 -40278 59166 -40240
rect 59076 -40310 59103 -40278
rect 59103 -40310 59137 -40278
rect 59137 -40310 59166 -40278
rect 60046 -40174 60126 -40140
rect 59856 -40228 59916 -40210
rect 60046 -40200 60126 -40174
rect 77410 -40120 77480 -40110
rect 77410 -40170 77420 -40120
rect 77420 -40170 77470 -40120
rect 77470 -40170 77480 -40120
rect 77410 -40180 77480 -40170
rect 59856 -40262 59874 -40228
rect 59874 -40262 59908 -40228
rect 59908 -40262 59916 -40228
rect 59856 -40280 59916 -40262
rect 60376 -40228 60446 -40220
rect 60376 -40262 60384 -40228
rect 60384 -40262 60418 -40228
rect 60418 -40262 60446 -40228
rect 59976 -40316 60316 -40300
rect 60376 -40280 60446 -40262
rect 57098 -40389 57368 -40364
rect 57098 -40423 57125 -40389
rect 57125 -40423 57159 -40389
rect 57159 -40423 57217 -40389
rect 57217 -40423 57251 -40389
rect 57251 -40423 57309 -40389
rect 57309 -40423 57343 -40389
rect 57343 -40423 57368 -40389
rect 54770 -41128 54802 -41048
rect 54802 -41128 54840 -41048
rect 53850 -41448 53920 -41338
rect 54920 -41268 54980 -41198
rect 55000 -41438 55090 -41338
rect 55540 -41438 55630 -41338
rect 55220 -41718 55280 -41548
rect 55280 -41718 55310 -41548
rect 55410 -41728 55500 -41558
rect 53950 -41850 54010 -41808
rect 53950 -41888 53988 -41850
rect 53988 -41888 54010 -41850
rect 54910 -41850 54980 -41798
rect 54910 -41888 54916 -41850
rect 54916 -41888 54950 -41850
rect 54950 -41888 54980 -41850
rect 54910 -41898 54980 -41888
rect 53510 -42048 53630 -41928
rect 54740 -42144 54850 -42068
rect 54740 -42158 54850 -42144
rect 55240 -42018 55370 -41958
rect 55410 -42138 55510 -42048
rect 57098 -40480 57368 -40423
rect 57098 -40504 57368 -40480
rect 56900 -40948 57020 -40818
rect 58576 -41040 58736 -40880
rect 57098 -41280 57368 -41274
rect 56480 -41334 56550 -41328
rect 56480 -41368 56492 -41334
rect 56492 -41368 56530 -41334
rect 56530 -41368 56550 -41334
rect 56480 -41388 56550 -41368
rect 57098 -41365 57368 -41280
rect 57098 -41399 57125 -41365
rect 57125 -41399 57159 -41365
rect 57159 -41399 57217 -41365
rect 57217 -41399 57251 -41365
rect 57251 -41399 57309 -41365
rect 57309 -41399 57343 -41365
rect 57343 -41399 57368 -41365
rect 57098 -41414 57368 -41399
rect 59976 -40352 60316 -40316
rect 59176 -40520 59196 -40440
rect 59196 -40520 59236 -40440
rect 59176 -40720 59196 -40640
rect 59196 -40720 59236 -40640
rect 59076 -40840 59103 -40810
rect 59103 -40840 59137 -40810
rect 59137 -40840 59166 -40810
rect 59076 -40880 59166 -40840
rect 59576 -40498 59636 -40470
rect 59576 -40530 59580 -40498
rect 59580 -40530 59636 -40498
rect 59476 -40720 59502 -40650
rect 59502 -40720 59536 -40650
rect 59576 -40758 59590 -40590
rect 59590 -40758 59624 -40590
rect 59624 -40758 59636 -40590
rect 59576 -40760 59636 -40758
rect 59076 -41008 59166 -40970
rect 59076 -41040 59103 -41008
rect 59103 -41040 59137 -41008
rect 59137 -41040 59166 -41008
rect 59206 -41040 59266 -40970
rect 61206 -40500 61346 -40320
rect 72820 -40480 73040 -40300
rect 79410 -40390 79680 -40150
rect 79780 -40370 79910 -40130
rect 83150 -40180 83510 -39830
rect 81140 -40510 81570 -40250
rect 91780 -39960 92130 -39580
rect 59806 -40740 59818 -40600
rect 59818 -40740 59852 -40600
rect 59852 -40740 59866 -40600
rect 59916 -40582 60006 -40580
rect 59916 -40758 59940 -40582
rect 59940 -40758 60006 -40582
rect 59916 -40760 60006 -40758
rect 60306 -40690 60456 -40550
rect 59826 -40842 59862 -40810
rect 59862 -40842 59896 -40810
rect 59896 -40842 59916 -40810
rect 59826 -40880 59916 -40842
rect 59166 -41210 59196 -41130
rect 59196 -41210 59226 -41130
rect 59166 -41440 59196 -41360
rect 59196 -41440 59226 -41360
rect 59466 -41210 59501 -41130
rect 59501 -41210 59526 -41130
rect 59586 -41250 59589 -41110
rect 59589 -41250 59623 -41110
rect 59623 -41250 59646 -41110
rect 59516 -41321 59596 -41320
rect 59516 -41355 59545 -41321
rect 59545 -41355 59579 -41321
rect 59579 -41355 59596 -41321
rect 59516 -41380 59596 -41355
rect 59826 -41011 59926 -40970
rect 59826 -41040 59861 -41011
rect 59861 -41040 59895 -41011
rect 59895 -41040 59926 -41011
rect 60096 -40883 60127 -40880
rect 60127 -40883 60161 -40880
rect 60161 -40883 60176 -40880
rect 60096 -40941 60176 -40883
rect 60096 -40975 60127 -40941
rect 60127 -40975 60161 -40941
rect 60161 -40975 60176 -40941
rect 60096 -41033 60176 -40975
rect 60096 -41040 60127 -41033
rect 60127 -41040 60161 -41033
rect 60161 -41040 60176 -41033
rect 59796 -41095 59856 -41090
rect 59796 -41270 59817 -41095
rect 59817 -41270 59851 -41095
rect 59851 -41270 59856 -41095
rect 59916 -41095 60006 -41090
rect 59916 -41271 59939 -41095
rect 59939 -41271 60006 -41095
rect 59916 -41280 60006 -41271
rect 60476 -41125 60536 -41110
rect 60476 -41159 60484 -41125
rect 60484 -41159 60536 -41125
rect 60476 -41170 60536 -41159
rect 61036 -40730 61126 -40620
rect 77450 -40550 77520 -40540
rect 77450 -40600 77460 -40550
rect 77460 -40600 77510 -40550
rect 77510 -40600 77520 -40550
rect 77450 -40610 77520 -40600
rect 77780 -40590 77840 -40570
rect 77780 -40630 77790 -40590
rect 77790 -40630 77830 -40590
rect 77830 -40630 77840 -40590
rect 72820 -40840 73040 -40660
rect 78310 -40760 78410 -40650
rect 87830 -40590 88190 -40240
rect 61276 -40883 61291 -40850
rect 61291 -40883 61325 -40850
rect 61325 -40883 61356 -40850
rect 61276 -40941 61356 -40883
rect 61276 -40975 61291 -40941
rect 61291 -40975 61325 -40941
rect 61325 -40975 61356 -40941
rect 61276 -41033 61356 -40975
rect 61276 -41060 61291 -41033
rect 61291 -41060 61325 -41033
rect 61325 -41060 61356 -41033
rect 76920 -40960 77060 -40820
rect 60476 -41260 60536 -41250
rect 60476 -41300 60486 -41260
rect 60486 -41300 60526 -41260
rect 60526 -41300 60536 -41260
rect 60476 -41310 60536 -41300
rect 60616 -41260 60736 -41250
rect 60616 -41300 60626 -41260
rect 60626 -41300 60666 -41260
rect 60666 -41300 60736 -41260
rect 60616 -41310 60736 -41300
rect 60756 -41260 60816 -41250
rect 60756 -41300 60766 -41260
rect 60766 -41300 60806 -41260
rect 60806 -41300 60816 -41260
rect 60756 -41310 60816 -41300
rect 60896 -41260 60956 -41250
rect 60896 -41300 60906 -41260
rect 60906 -41300 60946 -41260
rect 60946 -41300 60956 -41260
rect 60896 -41310 60956 -41300
rect 56380 -41688 56440 -41568
rect 55880 -41880 55970 -41878
rect 55880 -41914 55882 -41880
rect 55882 -41914 55970 -41880
rect 55880 -41958 55970 -41914
rect 55220 -42328 55330 -42218
rect 55530 -42402 55610 -42378
rect 55530 -42436 55560 -42402
rect 55560 -42436 55610 -42402
rect 55530 -42468 55610 -42436
rect 54140 -42508 54150 -42488
rect 54150 -42508 54840 -42488
rect 54840 -42508 54850 -42488
rect 54140 -42748 54850 -42508
rect 55320 -42548 55470 -42528
rect 55320 -42608 55470 -42548
rect 55320 -42668 55470 -42608
rect 56020 -42208 56080 -42058
rect 56170 -42208 56390 -42008
rect 56654 -42286 56998 -42068
rect 59076 -41570 59103 -41540
rect 59103 -41570 59137 -41540
rect 59137 -41570 59166 -41540
rect 59076 -41600 59166 -41570
rect 58926 -41710 58986 -41660
rect 58926 -41730 58966 -41710
rect 58966 -41730 58986 -41710
rect 59146 -41730 59226 -41660
rect 59276 -41730 59356 -41660
rect 59396 -41730 59476 -41660
rect 59646 -41720 59706 -41660
rect 59546 -41808 59606 -41800
rect 59256 -41862 59366 -41830
rect 59546 -41842 59560 -41808
rect 59560 -41842 59594 -41808
rect 59594 -41842 59606 -41808
rect 59016 -41916 59076 -41900
rect 59256 -41890 59366 -41862
rect 59546 -41860 59606 -41842
rect 59016 -41950 59032 -41916
rect 59032 -41950 59066 -41916
rect 59066 -41950 59076 -41916
rect 59016 -41960 59076 -41950
rect 58906 -42100 58926 -42030
rect 58926 -42100 58966 -42030
rect 58966 -42100 58986 -42030
rect 59146 -42100 59226 -42030
rect 59276 -42100 59356 -42030
rect 59396 -42100 59476 -42030
rect 59966 -41540 60326 -41520
rect 59966 -41574 60326 -41540
rect 72820 -41240 73040 -41060
rect 77450 -41180 77530 -41160
rect 77450 -41220 77470 -41180
rect 77470 -41220 77510 -41180
rect 77510 -41220 77530 -41180
rect 77450 -41240 77530 -41220
rect 77780 -41150 77840 -41140
rect 77780 -41190 77790 -41150
rect 77790 -41190 77830 -41150
rect 77830 -41190 77840 -41150
rect 77780 -41200 77840 -41190
rect 78060 -41180 78070 -41090
rect 78070 -41180 78110 -41090
rect 78110 -41180 78120 -41090
rect 78180 -41230 78190 -41140
rect 78190 -41230 78280 -41140
rect 78280 -41230 78290 -41140
rect 78180 -41240 78290 -41230
rect 78350 -41140 78410 -41130
rect 78350 -41180 78360 -41140
rect 78360 -41180 78400 -41140
rect 78400 -41180 78410 -41140
rect 78350 -41190 78410 -41180
rect 78670 -41380 78780 -41030
rect 80080 -41290 80430 -40910
rect 59966 -41580 60326 -41574
rect 59856 -41594 59916 -41580
rect 59856 -41628 59874 -41594
rect 59874 -41628 59908 -41594
rect 59908 -41628 59916 -41594
rect 59856 -41640 59916 -41628
rect 60376 -41594 60436 -41580
rect 60376 -41628 60384 -41594
rect 60384 -41628 60418 -41594
rect 60418 -41628 60436 -41594
rect 60376 -41640 60436 -41628
rect 61056 -41640 61126 -41540
rect 72820 -41690 73040 -41510
rect 79410 -41620 79680 -41380
rect 59806 -41920 59916 -41810
rect 60446 -41950 60526 -41830
rect 77490 -41790 77580 -41770
rect 77490 -41840 77510 -41790
rect 77510 -41840 77560 -41790
rect 77560 -41840 77580 -41790
rect 77490 -41860 77580 -41840
rect 77780 -41830 77840 -41810
rect 77780 -41870 77790 -41830
rect 77790 -41870 77830 -41830
rect 77830 -41870 77840 -41830
rect 59646 -42100 59706 -42040
rect 72820 -42060 73040 -41880
rect 76920 -42220 77060 -42060
rect 78170 -42000 78290 -41730
rect 78530 -42000 78590 -41730
rect 58986 -42560 59126 -42420
rect 59996 -42500 60106 -42390
rect 77470 -42430 77560 -42410
rect 77470 -42480 77490 -42430
rect 77490 -42480 77540 -42430
rect 77540 -42480 77560 -42430
rect 77470 -42500 77560 -42480
rect 77780 -42400 77840 -42380
rect 77780 -42440 77790 -42400
rect 77790 -42440 77830 -42400
rect 77830 -42440 77840 -42400
rect 78060 -42640 78120 -42340
rect 36000 -44300 44300 -43300
rect 55500 -43500 56100 -43100
rect 59800 -43400 60400 -42800
rect 77470 -43000 77540 -42930
rect 78240 -42889 78300 -42880
rect 78240 -42923 78250 -42889
rect 78250 -42923 78290 -42889
rect 78290 -42923 78300 -42889
rect 78240 -42940 78300 -42923
rect 79410 -42880 79680 -42640
rect 78860 -42970 78900 -42920
rect 78900 -42970 78980 -42920
rect 75940 -43140 76050 -43080
rect 77200 -43140 77260 -43080
rect 77860 -43110 77920 -43050
rect 76920 -43450 77060 -43310
rect 78860 -43040 78980 -42970
rect 78630 -43090 78700 -43080
rect 78630 -43130 78640 -43090
rect 78640 -43130 78690 -43090
rect 78690 -43130 78700 -43090
rect 78630 -43140 78700 -43130
rect 77960 -43210 78020 -43190
rect 77960 -43250 77970 -43210
rect 77970 -43250 78010 -43210
rect 78010 -43250 78020 -43210
rect 78340 -43180 78350 -43140
rect 78350 -43180 78400 -43140
rect 78400 -43180 78410 -43140
rect 78340 -43200 78410 -43180
rect 78860 -43090 78900 -43040
rect 78900 -43090 78980 -43040
rect 78860 -43160 78980 -43090
rect 78860 -43210 78900 -43160
rect 78900 -43210 78980 -43160
rect 80010 -43290 80360 -42910
rect 82820 -43310 91410 -42740
rect 77200 -43590 77260 -43530
rect 77860 -43540 77920 -43500
rect 77860 -43580 77870 -43540
rect 77870 -43580 77910 -43540
rect 77910 -43580 77920 -43540
rect 77860 -43620 77920 -43580
rect 77860 -43660 77870 -43620
rect 77870 -43660 77910 -43620
rect 77910 -43660 77920 -43620
rect 77860 -43670 77920 -43660
rect 78240 -43510 78300 -43500
rect 78240 -43560 78280 -43510
rect 78280 -43560 78300 -43510
rect 77970 -43630 78030 -43620
rect 77970 -43670 78010 -43630
rect 78010 -43670 78030 -43630
rect 77970 -43680 78030 -43670
rect 78240 -43650 78300 -43560
rect 78240 -43700 78280 -43650
rect 78280 -43700 78300 -43650
rect 77430 -43770 77500 -43760
rect 77430 -43820 77440 -43770
rect 77440 -43820 77490 -43770
rect 77490 -43820 77500 -43770
rect 77430 -43830 77500 -43820
rect 78240 -43790 78300 -43700
rect 78240 -43840 78280 -43790
rect 78280 -43840 78300 -43790
rect 78240 -43870 78300 -43840
rect 55500 -44360 55720 -44080
rect 79410 -44100 79680 -43860
rect 82470 -44000 82550 -43890
rect 83040 -43910 83100 -43890
rect 83040 -43990 83050 -43910
rect 83050 -43990 83090 -43910
rect 83090 -43990 83100 -43910
rect 83040 -44000 83100 -43990
rect 85320 -43820 85390 -43810
rect 85320 -43990 85330 -43820
rect 85330 -43990 85380 -43820
rect 85380 -43990 85390 -43820
rect 85320 -44000 85390 -43990
rect 85590 -43897 86480 -43870
rect 85590 -43931 85610 -43897
rect 85610 -43931 86471 -43897
rect 86471 -43931 86480 -43897
rect 85590 -43950 86480 -43931
rect 86800 -43800 86870 -43790
rect 86800 -43990 86810 -43800
rect 86810 -43990 86860 -43800
rect 86860 -43990 86870 -43800
rect 86800 -44000 86870 -43990
rect 87040 -43896 87920 -43870
rect 87040 -43930 87044 -43896
rect 87044 -43930 87905 -43896
rect 87905 -43930 87920 -43896
rect 87040 -43950 87920 -43930
rect 88270 -43810 88340 -43800
rect 88270 -43990 88280 -43810
rect 88280 -43990 88330 -43810
rect 88330 -43990 88340 -43810
rect 88270 -44000 88340 -43990
rect 88510 -43896 89390 -43880
rect 88510 -43930 88523 -43896
rect 88523 -43930 89384 -43896
rect 89384 -43930 89390 -43896
rect 88510 -43950 89390 -43930
rect 89740 -43810 89810 -43800
rect 89740 -44000 89750 -43810
rect 89750 -44000 89800 -43810
rect 89800 -44000 89810 -43810
rect 89740 -44010 89810 -44000
rect 89982 -43897 90762 -43879
rect 89982 -43899 90747 -43897
rect 90747 -43899 90762 -43897
rect 89982 -43933 90748 -43899
rect 90748 -43933 90762 -43899
rect 89982 -43951 90762 -43933
rect 91210 -43810 91280 -43800
rect 91210 -44000 91220 -43810
rect 91220 -44000 91270 -43810
rect 91270 -44000 91280 -43810
rect 91210 -44010 91280 -44000
rect 75940 -44240 76050 -44150
rect 75660 -44330 75760 -44270
rect 36000 -45900 44300 -44900
rect 53480 -44940 53780 -44740
rect 54150 -44708 54860 -44538
rect 54150 -44778 54850 -44708
rect 54850 -44778 54860 -44708
rect 53520 -45168 53640 -45058
rect 54750 -45108 54850 -45038
rect 54750 -45118 54840 -45108
rect 55430 -45088 55520 -45018
rect 55290 -45198 55390 -45128
rect 36000 -47500 43400 -46500
rect 53050 -47108 53250 -45358
rect 53950 -45328 53998 -45298
rect 53998 -45328 54020 -45298
rect 53950 -45398 54020 -45328
rect 54920 -45290 54990 -45278
rect 54920 -45328 54926 -45290
rect 54926 -45328 54960 -45290
rect 54960 -45328 54990 -45290
rect 54920 -45368 54990 -45328
rect 53860 -45838 53920 -45728
rect 55230 -45628 55290 -45458
rect 55290 -45628 55320 -45458
rect 55430 -45618 55510 -45448
rect 77760 -44440 77820 -44420
rect 77760 -44480 77770 -44440
rect 77770 -44480 77810 -44440
rect 77810 -44480 77820 -44440
rect 77970 -44360 78030 -44350
rect 77970 -44460 78010 -44360
rect 78010 -44460 78030 -44360
rect 77970 -44470 78030 -44460
rect 78180 -44140 78300 -44130
rect 78180 -44460 78290 -44140
rect 78290 -44460 78300 -44140
rect 78180 -44470 78300 -44460
rect 55960 -45088 56040 -44938
rect 56190 -45168 56390 -44958
rect 56506 -45030 57016 -44780
rect 58966 -44830 59126 -44670
rect 76920 -44610 77060 -44520
rect 59956 -44860 60166 -44700
rect 77760 -44780 77770 -44740
rect 77770 -44780 77810 -44740
rect 77810 -44780 77820 -44740
rect 77760 -44800 77820 -44780
rect 55880 -45256 55970 -45218
rect 55880 -45290 55882 -45256
rect 55882 -45290 55970 -45256
rect 55880 -45298 55970 -45290
rect 55000 -45838 55090 -45738
rect 54770 -46040 54840 -46038
rect 54770 -46128 54802 -46040
rect 54802 -46128 54840 -46040
rect 55540 -45838 55630 -45738
rect 56590 -45598 56660 -45468
rect 75940 -44900 76050 -44840
rect 77960 -44860 78020 -44850
rect 77960 -44910 78010 -44860
rect 78010 -44910 78020 -44860
rect 77960 -44920 78020 -44910
rect 75230 -45060 75330 -44970
rect 78640 -45090 78750 -44950
rect 82820 -45010 91410 -44440
rect 91780 -44460 92130 -44080
rect 58906 -45220 58966 -45170
rect 58906 -45230 58926 -45220
rect 58926 -45230 58966 -45220
rect 59216 -45230 59276 -45170
rect 59326 -45230 59386 -45170
rect 59436 -45230 59496 -45170
rect 59636 -45230 59696 -45170
rect 59546 -45301 59606 -45290
rect 59286 -45355 59346 -45330
rect 59546 -45335 59560 -45301
rect 59560 -45335 59594 -45301
rect 59594 -45335 59606 -45301
rect 59286 -45389 59346 -45355
rect 59546 -45350 59606 -45335
rect 59286 -45390 59346 -45389
rect 59016 -45409 59076 -45400
rect 59016 -45443 59032 -45409
rect 59032 -45443 59066 -45409
rect 59066 -45443 59076 -45409
rect 59016 -45460 59076 -45443
rect 59546 -45470 59606 -45410
rect 58906 -45590 58966 -45530
rect 59216 -45580 59276 -45520
rect 59336 -45580 59396 -45520
rect 59436 -45580 59496 -45520
rect 55140 -46208 55200 -46138
rect 55030 -46328 55110 -46248
rect 55740 -46328 55810 -46248
rect 55880 -46328 55970 -46238
rect 56480 -45806 56550 -45788
rect 56480 -45840 56492 -45806
rect 56492 -45840 56530 -45806
rect 56530 -45840 56550 -45806
rect 56480 -45848 56550 -45840
rect 59866 -45430 59966 -45340
rect 60446 -45420 60526 -45320
rect 76500 -45420 76600 -45350
rect 79410 -45360 79680 -45120
rect 59636 -45590 59696 -45530
rect 59076 -45678 59166 -45640
rect 59076 -45710 59103 -45678
rect 59103 -45710 59137 -45678
rect 59137 -45710 59166 -45678
rect 60046 -45574 60126 -45540
rect 75230 -45570 75330 -45500
rect 59856 -45628 59916 -45610
rect 60046 -45600 60126 -45574
rect 59856 -45662 59874 -45628
rect 59874 -45662 59908 -45628
rect 59908 -45662 59916 -45628
rect 59856 -45680 59916 -45662
rect 60376 -45628 60446 -45620
rect 60376 -45662 60384 -45628
rect 60384 -45662 60418 -45628
rect 60418 -45662 60446 -45628
rect 59976 -45716 60316 -45700
rect 60376 -45680 60446 -45662
rect 57098 -45789 57368 -45764
rect 57098 -45823 57125 -45789
rect 57125 -45823 57159 -45789
rect 57159 -45823 57217 -45789
rect 57217 -45823 57251 -45789
rect 57251 -45823 57309 -45789
rect 57309 -45823 57343 -45789
rect 57343 -45823 57368 -45789
rect 54770 -46528 54802 -46448
rect 54802 -46528 54840 -46448
rect 53850 -46848 53920 -46738
rect 54920 -46668 54980 -46598
rect 55000 -46838 55090 -46738
rect 55540 -46838 55630 -46738
rect 55220 -47118 55280 -46948
rect 55280 -47118 55310 -46948
rect 55410 -47128 55500 -46958
rect 53950 -47250 54010 -47208
rect 53950 -47288 53988 -47250
rect 53988 -47288 54010 -47250
rect 54910 -47250 54980 -47198
rect 54910 -47288 54916 -47250
rect 54916 -47288 54950 -47250
rect 54950 -47288 54980 -47250
rect 54910 -47298 54980 -47288
rect 53510 -47448 53630 -47328
rect 54740 -47544 54850 -47468
rect 54740 -47558 54850 -47544
rect 55240 -47418 55370 -47358
rect 55410 -47538 55510 -47448
rect 57098 -45880 57368 -45823
rect 57098 -45904 57368 -45880
rect 56900 -46348 57020 -46218
rect 58576 -46440 58736 -46280
rect 57098 -46680 57368 -46674
rect 56480 -46734 56550 -46728
rect 56480 -46768 56492 -46734
rect 56492 -46768 56530 -46734
rect 56530 -46768 56550 -46734
rect 56480 -46788 56550 -46768
rect 57098 -46765 57368 -46680
rect 57098 -46799 57125 -46765
rect 57125 -46799 57159 -46765
rect 57159 -46799 57217 -46765
rect 57217 -46799 57251 -46765
rect 57251 -46799 57309 -46765
rect 57309 -46799 57343 -46765
rect 57343 -46799 57368 -46765
rect 57098 -46814 57368 -46799
rect 59976 -45752 60316 -45716
rect 59176 -45920 59196 -45840
rect 59196 -45920 59236 -45840
rect 59176 -46120 59196 -46040
rect 59196 -46120 59236 -46040
rect 59076 -46240 59103 -46210
rect 59103 -46240 59137 -46210
rect 59137 -46240 59166 -46210
rect 59076 -46280 59166 -46240
rect 59576 -45898 59636 -45870
rect 59576 -45930 59580 -45898
rect 59580 -45930 59636 -45898
rect 59476 -46120 59502 -46050
rect 59502 -46120 59536 -46050
rect 59576 -46158 59590 -45990
rect 59590 -46158 59624 -45990
rect 59624 -46158 59636 -45990
rect 59576 -46160 59636 -46158
rect 59076 -46408 59166 -46370
rect 59076 -46440 59103 -46408
rect 59103 -46440 59137 -46408
rect 59137 -46440 59166 -46408
rect 59206 -46440 59266 -46370
rect 61206 -45900 61346 -45720
rect 76920 -45740 77060 -45640
rect 77600 -45620 77710 -45610
rect 77600 -45670 77620 -45620
rect 77620 -45670 77690 -45620
rect 77690 -45670 77710 -45620
rect 77600 -45680 77710 -45670
rect 78070 -45490 78140 -45480
rect 78070 -45580 78080 -45490
rect 78080 -45580 78130 -45490
rect 78130 -45580 78140 -45490
rect 78070 -45590 78140 -45580
rect 78240 -45550 78300 -45530
rect 78240 -45590 78250 -45550
rect 78250 -45590 78290 -45550
rect 78290 -45590 78300 -45550
rect 78640 -45520 78740 -45510
rect 78640 -45590 78650 -45520
rect 78650 -45590 78730 -45520
rect 78730 -45590 78740 -45520
rect 78640 -45600 78740 -45590
rect 78810 -45560 78870 -45550
rect 78810 -45600 78820 -45560
rect 78820 -45600 78860 -45560
rect 78860 -45600 78870 -45560
rect 78810 -45610 78870 -45600
rect 79080 -45680 79190 -45380
rect 80010 -45810 80360 -45430
rect 59806 -46140 59818 -46000
rect 59818 -46140 59852 -46000
rect 59852 -46140 59866 -46000
rect 59916 -45982 60006 -45980
rect 59916 -46158 59940 -45982
rect 59940 -46158 60006 -45982
rect 59916 -46160 60006 -46158
rect 60306 -46090 60456 -45950
rect 59826 -46242 59862 -46210
rect 59862 -46242 59896 -46210
rect 59896 -46242 59916 -46210
rect 59826 -46280 59916 -46242
rect 59166 -46610 59196 -46530
rect 59196 -46610 59226 -46530
rect 59166 -46840 59196 -46760
rect 59196 -46840 59226 -46760
rect 59466 -46610 59501 -46530
rect 59501 -46610 59526 -46530
rect 59586 -46650 59589 -46510
rect 59589 -46650 59623 -46510
rect 59623 -46650 59646 -46510
rect 59516 -46721 59596 -46720
rect 59516 -46755 59545 -46721
rect 59545 -46755 59579 -46721
rect 59579 -46755 59596 -46721
rect 59516 -46780 59596 -46755
rect 59826 -46411 59926 -46370
rect 59826 -46440 59861 -46411
rect 59861 -46440 59895 -46411
rect 59895 -46440 59926 -46411
rect 60096 -46283 60127 -46280
rect 60127 -46283 60161 -46280
rect 60161 -46283 60176 -46280
rect 60096 -46341 60176 -46283
rect 60096 -46375 60127 -46341
rect 60127 -46375 60161 -46341
rect 60161 -46375 60176 -46341
rect 60096 -46433 60176 -46375
rect 60096 -46440 60127 -46433
rect 60127 -46440 60161 -46433
rect 60161 -46440 60176 -46433
rect 59796 -46495 59856 -46490
rect 59796 -46670 59817 -46495
rect 59817 -46670 59851 -46495
rect 59851 -46670 59856 -46495
rect 59916 -46495 60006 -46490
rect 59916 -46671 59939 -46495
rect 59939 -46671 60006 -46495
rect 59916 -46680 60006 -46671
rect 60476 -46525 60536 -46510
rect 60476 -46559 60484 -46525
rect 60484 -46559 60536 -46525
rect 60476 -46570 60536 -46559
rect 61036 -46130 61126 -46020
rect 61276 -46283 61291 -46250
rect 61291 -46283 61325 -46250
rect 61325 -46283 61356 -46250
rect 61276 -46341 61356 -46283
rect 61276 -46375 61291 -46341
rect 61291 -46375 61325 -46341
rect 61325 -46375 61356 -46341
rect 61276 -46433 61356 -46375
rect 61276 -46460 61291 -46433
rect 61291 -46460 61325 -46433
rect 61325 -46460 61356 -46433
rect 73220 -46590 73340 -46400
rect 60476 -46660 60536 -46650
rect 60476 -46700 60486 -46660
rect 60486 -46700 60526 -46660
rect 60526 -46700 60536 -46660
rect 60476 -46710 60536 -46700
rect 60616 -46660 60736 -46650
rect 60616 -46700 60626 -46660
rect 60626 -46700 60666 -46660
rect 60666 -46700 60736 -46660
rect 60616 -46710 60736 -46700
rect 60756 -46660 60816 -46650
rect 60756 -46700 60766 -46660
rect 60766 -46700 60806 -46660
rect 60806 -46700 60816 -46660
rect 60756 -46710 60816 -46700
rect 60896 -46660 60956 -46650
rect 60896 -46700 60906 -46660
rect 60906 -46700 60946 -46660
rect 60946 -46700 60956 -46660
rect 60896 -46710 60956 -46700
rect 56380 -47088 56440 -46968
rect 55880 -47280 55970 -47278
rect 55880 -47314 55882 -47280
rect 55882 -47314 55970 -47280
rect 55880 -47358 55970 -47314
rect 55220 -47728 55330 -47618
rect 55530 -47802 55610 -47778
rect 55530 -47836 55560 -47802
rect 55560 -47836 55610 -47802
rect 55530 -47868 55610 -47836
rect 54140 -47908 54150 -47888
rect 54150 -47908 54840 -47888
rect 54840 -47908 54850 -47888
rect 36000 -49100 42500 -48100
rect 54140 -48148 54850 -47908
rect 55320 -47948 55470 -47928
rect 55320 -48008 55470 -47948
rect 55320 -48068 55470 -48008
rect 56020 -47608 56080 -47458
rect 56170 -47608 56390 -47408
rect 56654 -47686 56998 -47468
rect 59076 -46970 59103 -46940
rect 59103 -46970 59137 -46940
rect 59137 -46970 59166 -46940
rect 59076 -47000 59166 -46970
rect 58926 -47110 58986 -47060
rect 58926 -47130 58966 -47110
rect 58966 -47130 58986 -47110
rect 59146 -47130 59226 -47060
rect 59276 -47130 59356 -47060
rect 59396 -47130 59476 -47060
rect 59646 -47120 59706 -47060
rect 59546 -47208 59606 -47200
rect 59256 -47262 59366 -47230
rect 59546 -47242 59560 -47208
rect 59560 -47242 59594 -47208
rect 59594 -47242 59606 -47208
rect 59016 -47316 59076 -47300
rect 59256 -47290 59366 -47262
rect 59546 -47260 59606 -47242
rect 59016 -47350 59032 -47316
rect 59032 -47350 59066 -47316
rect 59066 -47350 59076 -47316
rect 59016 -47360 59076 -47350
rect 58906 -47500 58926 -47430
rect 58926 -47500 58966 -47430
rect 58966 -47500 58986 -47430
rect 59146 -47500 59226 -47430
rect 59276 -47500 59356 -47430
rect 59396 -47500 59476 -47430
rect 59966 -46940 60326 -46920
rect 59966 -46974 60326 -46940
rect 73470 -46590 73590 -46400
rect 73720 -46590 73840 -46400
rect 73970 -46590 74090 -46400
rect 74220 -46590 74340 -46400
rect 74470 -46590 74590 -46400
rect 74720 -46590 74840 -46400
rect 74970 -46590 75090 -46400
rect 75390 -46310 75550 -46190
rect 75220 -46590 75340 -46400
rect 73723 -46688 73840 -46636
rect 75410 -46690 75470 -46630
rect 75673 -46649 75751 -46623
rect 75673 -46683 75704 -46649
rect 75704 -46683 75751 -46649
rect 75673 -46701 75751 -46683
rect 75946 -46649 76024 -46623
rect 75946 -46683 75947 -46649
rect 75947 -46683 75981 -46649
rect 75981 -46683 76024 -46649
rect 75946 -46701 76024 -46683
rect 74220 -46880 74340 -46800
rect 76102 -46650 76167 -46623
rect 76920 -46570 77060 -46450
rect 76102 -46684 76128 -46650
rect 76128 -46684 76162 -46650
rect 76162 -46684 76167 -46650
rect 76102 -46701 76167 -46684
rect 76232 -46650 76310 -46623
rect 76232 -46684 76258 -46650
rect 76258 -46684 76310 -46650
rect 76232 -46701 76310 -46684
rect 76380 -46649 76440 -46640
rect 76380 -46683 76404 -46649
rect 76404 -46683 76438 -46649
rect 76438 -46683 76440 -46649
rect 76380 -46700 76440 -46683
rect 76505 -46649 76583 -46636
rect 76505 -46683 76531 -46649
rect 76531 -46683 76583 -46649
rect 76505 -46701 76583 -46683
rect 76648 -46649 76726 -46636
rect 76648 -46683 76680 -46649
rect 76680 -46683 76714 -46649
rect 76714 -46683 76726 -46649
rect 76648 -46714 76726 -46683
rect 76791 -46650 76843 -46636
rect 76791 -46684 76806 -46650
rect 76806 -46684 76843 -46650
rect 76791 -46714 76843 -46684
rect 59966 -46980 60326 -46974
rect 59856 -46994 59916 -46980
rect 59856 -47028 59874 -46994
rect 59874 -47028 59908 -46994
rect 59908 -47028 59916 -46994
rect 59856 -47040 59916 -47028
rect 60376 -46994 60436 -46980
rect 60376 -47028 60384 -46994
rect 60384 -47028 60418 -46994
rect 60418 -47028 60436 -46994
rect 60376 -47040 60436 -47028
rect 61056 -47040 61126 -46940
rect 72820 -47080 73040 -46900
rect 77170 -47080 77430 -46830
rect 59806 -47320 59916 -47210
rect 73480 -47220 73580 -47160
rect 60446 -47350 60526 -47230
rect 72820 -47410 73040 -47230
rect 73730 -47330 73830 -47270
rect 59646 -47500 59706 -47440
rect 73230 -47440 73330 -47380
rect 78150 -47390 78210 -47380
rect 78150 -47430 78160 -47390
rect 78160 -47430 78200 -47390
rect 78200 -47430 78210 -47390
rect 78150 -47440 78210 -47430
rect 78280 -47390 78340 -47380
rect 78280 -47430 78290 -47390
rect 78290 -47430 78330 -47390
rect 78330 -47430 78340 -47390
rect 78580 -47370 78640 -47360
rect 78580 -47410 78590 -47370
rect 78590 -47410 78630 -47370
rect 78630 -47410 78640 -47370
rect 78580 -47420 78640 -47410
rect 78800 -47380 78860 -47370
rect 78800 -47420 78850 -47380
rect 78850 -47420 78860 -47380
rect 78800 -47430 78860 -47420
rect 78280 -47440 78340 -47430
rect 77230 -47490 77310 -47480
rect 77230 -47530 77240 -47490
rect 77240 -47530 77300 -47490
rect 77300 -47530 77310 -47490
rect 77230 -47540 77310 -47530
rect 58986 -47960 59126 -47820
rect 59996 -47900 60106 -47790
rect 72820 -47900 73040 -47720
rect 76920 -47760 77060 -47610
rect 79080 -47440 79140 -47390
rect 79140 -47440 79250 -47390
rect 79080 -47490 79250 -47440
rect 79080 -47550 79140 -47490
rect 79140 -47550 79250 -47490
rect 80080 -47620 80430 -47310
rect 82824 -47448 91414 -46878
rect 77170 -47830 77260 -47820
rect 77170 -47880 77260 -47830
rect 77170 -47890 77260 -47880
rect 74230 -47990 74330 -47930
rect 72820 -48180 73040 -48000
rect 74730 -48080 74830 -48020
rect 78150 -47870 78160 -47830
rect 78160 -47870 78200 -47830
rect 78200 -47870 78210 -47830
rect 78150 -47940 78210 -47870
rect 78150 -47980 78160 -47940
rect 78160 -47980 78200 -47940
rect 78200 -47980 78210 -47940
rect 78150 -48060 78210 -47980
rect 78150 -48100 78160 -48060
rect 78160 -48100 78200 -48060
rect 78200 -48100 78210 -48060
rect 78150 -48120 78210 -48100
rect 80080 -48100 80430 -47720
rect 81950 -48140 82070 -48020
rect 83040 -48040 83100 -48020
rect 83040 -48130 83050 -48040
rect 83050 -48130 83090 -48040
rect 83090 -48130 83100 -48040
rect 83040 -48140 83100 -48130
rect 85324 -47958 85394 -47948
rect 85324 -48128 85334 -47958
rect 85334 -48128 85384 -47958
rect 85384 -48128 85394 -47958
rect 85324 -48138 85394 -48128
rect 85594 -48035 86484 -48008
rect 85594 -48069 85614 -48035
rect 85614 -48069 86475 -48035
rect 86475 -48069 86484 -48035
rect 85594 -48088 86484 -48069
rect 86804 -47938 86874 -47928
rect 86804 -48128 86814 -47938
rect 86814 -48128 86864 -47938
rect 86864 -48128 86874 -47938
rect 86804 -48138 86874 -48128
rect 87044 -48034 87924 -48008
rect 87044 -48068 87048 -48034
rect 87048 -48068 87909 -48034
rect 87909 -48068 87924 -48034
rect 87044 -48088 87924 -48068
rect 88274 -47948 88344 -47938
rect 88274 -48128 88284 -47948
rect 88284 -48128 88334 -47948
rect 88334 -48128 88344 -47948
rect 88274 -48138 88344 -48128
rect 88514 -48034 89394 -48018
rect 88514 -48068 88527 -48034
rect 88527 -48068 89388 -48034
rect 89388 -48068 89394 -48034
rect 88514 -48088 89394 -48068
rect 89744 -47948 89814 -47938
rect 89744 -48138 89754 -47948
rect 89754 -48138 89804 -47948
rect 89804 -48138 89814 -47948
rect 89744 -48148 89814 -48138
rect 89986 -48035 90766 -48017
rect 89986 -48037 90751 -48035
rect 90751 -48037 90766 -48035
rect 89986 -48071 90752 -48037
rect 90752 -48071 90766 -48037
rect 89986 -48089 90766 -48071
rect 77410 -48160 77480 -48150
rect 77410 -48210 77420 -48160
rect 77420 -48210 77470 -48160
rect 77470 -48210 77480 -48160
rect 77410 -48220 77480 -48210
rect 91214 -47948 91284 -47938
rect 91214 -48138 91224 -47948
rect 91224 -48138 91274 -47948
rect 91274 -48138 91284 -47948
rect 91214 -48148 91284 -48138
rect 79410 -48430 79680 -48190
rect 55500 -48900 56100 -48500
rect 72820 -48640 73040 -48460
rect 77450 -48590 77520 -48580
rect 77450 -48640 77460 -48590
rect 77460 -48640 77510 -48590
rect 77510 -48640 77520 -48590
rect 77450 -48650 77520 -48640
rect 77780 -48630 77840 -48610
rect 77780 -48670 77790 -48630
rect 77790 -48670 77830 -48630
rect 77830 -48670 77840 -48630
rect 72820 -49000 73040 -48820
rect 78310 -48800 78410 -48690
rect 76920 -49000 77060 -48860
rect 72820 -49400 73040 -49220
rect 77450 -49220 77530 -49200
rect 77450 -49260 77470 -49220
rect 77470 -49260 77510 -49220
rect 77510 -49260 77530 -49220
rect 77450 -49280 77530 -49260
rect 77780 -49190 77840 -49180
rect 77780 -49230 77790 -49190
rect 77790 -49230 77830 -49190
rect 77830 -49230 77840 -49190
rect 77780 -49240 77840 -49230
rect 78060 -49220 78070 -49130
rect 78070 -49220 78110 -49130
rect 78110 -49220 78120 -49130
rect 78180 -49270 78190 -49180
rect 78190 -49270 78280 -49180
rect 78280 -49270 78290 -49180
rect 78180 -49280 78290 -49270
rect 78350 -49180 78410 -49170
rect 78350 -49220 78360 -49180
rect 78360 -49220 78400 -49180
rect 78400 -49220 78410 -49180
rect 78350 -49230 78410 -49220
rect 78670 -49420 78780 -49070
rect 80080 -49330 80430 -48950
rect 82824 -49148 91414 -48578
rect 91780 -48620 92130 -48240
rect 36000 -50700 41600 -49700
rect 55460 -49760 55720 -49480
rect 79410 -49660 79680 -49420
rect 53460 -50340 53780 -50140
rect 54150 -50108 54860 -49938
rect 54150 -50178 54850 -50108
rect 54850 -50178 54860 -50108
rect 53520 -50568 53640 -50458
rect 54750 -50508 54850 -50438
rect 54750 -50518 54840 -50508
rect 55430 -50488 55520 -50418
rect 55290 -50598 55390 -50528
rect 36000 -52300 40700 -51300
rect 53050 -52508 53250 -50758
rect 53950 -50728 53998 -50698
rect 53998 -50728 54020 -50698
rect 53950 -50798 54020 -50728
rect 54920 -50690 54990 -50678
rect 54920 -50728 54926 -50690
rect 54926 -50728 54960 -50690
rect 54960 -50728 54990 -50690
rect 54920 -50768 54990 -50728
rect 53860 -51238 53920 -51128
rect 55230 -51028 55290 -50858
rect 55290 -51028 55320 -50858
rect 55430 -51018 55510 -50848
rect 72820 -49850 73040 -49670
rect 77490 -49830 77580 -49810
rect 77490 -49880 77510 -49830
rect 77510 -49880 77560 -49830
rect 77560 -49880 77580 -49830
rect 77490 -49900 77580 -49880
rect 77780 -49870 77840 -49850
rect 77780 -49910 77790 -49870
rect 77790 -49910 77830 -49870
rect 77830 -49910 77840 -49870
rect 55960 -50488 56040 -50338
rect 56190 -50568 56390 -50358
rect 56506 -50430 57016 -50180
rect 58966 -50230 59126 -50070
rect 59956 -50260 60166 -50100
rect 72820 -50220 73040 -50040
rect 55880 -50656 55970 -50618
rect 55880 -50690 55882 -50656
rect 55882 -50690 55970 -50656
rect 55880 -50698 55970 -50690
rect 55000 -51238 55090 -51138
rect 54770 -51440 54840 -51438
rect 54770 -51528 54802 -51440
rect 54802 -51528 54840 -51440
rect 55540 -51238 55630 -51138
rect 56590 -50998 56660 -50868
rect 76920 -50260 77060 -50100
rect 78170 -50040 78290 -49770
rect 78530 -50040 78590 -49770
rect 58906 -50620 58966 -50570
rect 58906 -50630 58926 -50620
rect 58926 -50630 58966 -50620
rect 59216 -50630 59276 -50570
rect 59326 -50630 59386 -50570
rect 59436 -50630 59496 -50570
rect 77470 -50470 77560 -50450
rect 77470 -50520 77490 -50470
rect 77490 -50520 77540 -50470
rect 77540 -50520 77560 -50470
rect 77470 -50540 77560 -50520
rect 77780 -50440 77840 -50420
rect 77780 -50480 77790 -50440
rect 77790 -50480 77830 -50440
rect 77830 -50480 77840 -50440
rect 59636 -50630 59696 -50570
rect 59546 -50701 59606 -50690
rect 59286 -50755 59346 -50730
rect 59546 -50735 59560 -50701
rect 59560 -50735 59594 -50701
rect 59594 -50735 59606 -50701
rect 59286 -50789 59346 -50755
rect 59546 -50750 59606 -50735
rect 59286 -50790 59346 -50789
rect 59016 -50809 59076 -50800
rect 59016 -50843 59032 -50809
rect 59032 -50843 59066 -50809
rect 59066 -50843 59076 -50809
rect 59016 -50860 59076 -50843
rect 59546 -50870 59606 -50810
rect 58906 -50990 58966 -50930
rect 59216 -50980 59276 -50920
rect 59336 -50980 59396 -50920
rect 59436 -50980 59496 -50920
rect 55140 -51608 55200 -51538
rect 55030 -51728 55110 -51648
rect 55740 -51728 55810 -51648
rect 55880 -51728 55970 -51638
rect 56480 -51206 56550 -51188
rect 56480 -51240 56492 -51206
rect 56492 -51240 56530 -51206
rect 56530 -51240 56550 -51206
rect 56480 -51248 56550 -51240
rect 78060 -50680 78120 -50380
rect 59866 -50830 59966 -50740
rect 60446 -50820 60526 -50720
rect 59636 -50990 59696 -50930
rect 59076 -51078 59166 -51040
rect 59076 -51110 59103 -51078
rect 59103 -51110 59137 -51078
rect 59137 -51110 59166 -51078
rect 60046 -50974 60126 -50940
rect 59856 -51028 59916 -51010
rect 60046 -51000 60126 -50974
rect 59856 -51062 59874 -51028
rect 59874 -51062 59908 -51028
rect 59908 -51062 59916 -51028
rect 59856 -51080 59916 -51062
rect 60376 -51028 60446 -51020
rect 60376 -51062 60384 -51028
rect 60384 -51062 60418 -51028
rect 60418 -51062 60446 -51028
rect 77470 -51040 77540 -50970
rect 78240 -50929 78300 -50920
rect 78240 -50963 78250 -50929
rect 78250 -50963 78290 -50929
rect 78290 -50963 78300 -50929
rect 78240 -50980 78300 -50963
rect 79410 -50920 79680 -50680
rect 78860 -51010 78900 -50960
rect 78900 -51010 78980 -50960
rect 59976 -51116 60316 -51100
rect 60376 -51080 60446 -51062
rect 57098 -51189 57368 -51164
rect 57098 -51223 57125 -51189
rect 57125 -51223 57159 -51189
rect 57159 -51223 57217 -51189
rect 57217 -51223 57251 -51189
rect 57251 -51223 57309 -51189
rect 57309 -51223 57343 -51189
rect 57343 -51223 57368 -51189
rect 54770 -51928 54802 -51848
rect 54802 -51928 54840 -51848
rect 53850 -52248 53920 -52138
rect 54920 -52068 54980 -51998
rect 55000 -52238 55090 -52138
rect 55540 -52238 55630 -52138
rect 55220 -52518 55280 -52348
rect 55280 -52518 55310 -52348
rect 55410 -52528 55500 -52358
rect 53950 -52650 54010 -52608
rect 53950 -52688 53988 -52650
rect 53988 -52688 54010 -52650
rect 54910 -52650 54980 -52598
rect 54910 -52688 54916 -52650
rect 54916 -52688 54950 -52650
rect 54950 -52688 54980 -52650
rect 54910 -52698 54980 -52688
rect 53510 -52848 53630 -52728
rect 36000 -53900 39800 -52900
rect 54740 -52944 54850 -52868
rect 54740 -52958 54850 -52944
rect 55240 -52818 55370 -52758
rect 55410 -52938 55510 -52848
rect 57098 -51280 57368 -51223
rect 57098 -51304 57368 -51280
rect 56900 -51748 57020 -51618
rect 58576 -51840 58736 -51680
rect 57098 -52080 57368 -52074
rect 56480 -52134 56550 -52128
rect 56480 -52168 56492 -52134
rect 56492 -52168 56530 -52134
rect 56530 -52168 56550 -52134
rect 56480 -52188 56550 -52168
rect 57098 -52165 57368 -52080
rect 57098 -52199 57125 -52165
rect 57125 -52199 57159 -52165
rect 57159 -52199 57217 -52165
rect 57217 -52199 57251 -52165
rect 57251 -52199 57309 -52165
rect 57309 -52199 57343 -52165
rect 57343 -52199 57368 -52165
rect 57098 -52214 57368 -52199
rect 59976 -51152 60316 -51116
rect 59176 -51320 59196 -51240
rect 59196 -51320 59236 -51240
rect 59176 -51520 59196 -51440
rect 59196 -51520 59236 -51440
rect 59076 -51640 59103 -51610
rect 59103 -51640 59137 -51610
rect 59137 -51640 59166 -51610
rect 59076 -51680 59166 -51640
rect 59576 -51298 59636 -51270
rect 59576 -51330 59580 -51298
rect 59580 -51330 59636 -51298
rect 59476 -51520 59502 -51450
rect 59502 -51520 59536 -51450
rect 59576 -51558 59590 -51390
rect 59590 -51558 59624 -51390
rect 59624 -51558 59636 -51390
rect 59576 -51560 59636 -51558
rect 59076 -51808 59166 -51770
rect 59076 -51840 59103 -51808
rect 59103 -51840 59137 -51808
rect 59137 -51840 59166 -51808
rect 59206 -51840 59266 -51770
rect 61206 -51300 61346 -51120
rect 75940 -51180 76050 -51120
rect 77200 -51180 77260 -51120
rect 77860 -51150 77920 -51090
rect 59806 -51540 59818 -51400
rect 59818 -51540 59852 -51400
rect 59852 -51540 59866 -51400
rect 59916 -51382 60006 -51380
rect 59916 -51558 59940 -51382
rect 59940 -51558 60006 -51382
rect 59916 -51560 60006 -51558
rect 60306 -51490 60456 -51350
rect 59826 -51642 59862 -51610
rect 59862 -51642 59896 -51610
rect 59896 -51642 59916 -51610
rect 59826 -51680 59916 -51642
rect 59166 -52010 59196 -51930
rect 59196 -52010 59226 -51930
rect 59166 -52240 59196 -52160
rect 59196 -52240 59226 -52160
rect 59466 -52010 59501 -51930
rect 59501 -52010 59526 -51930
rect 59586 -52050 59589 -51910
rect 59589 -52050 59623 -51910
rect 59623 -52050 59646 -51910
rect 59516 -52121 59596 -52120
rect 59516 -52155 59545 -52121
rect 59545 -52155 59579 -52121
rect 59579 -52155 59596 -52121
rect 59516 -52180 59596 -52155
rect 59826 -51811 59926 -51770
rect 59826 -51840 59861 -51811
rect 59861 -51840 59895 -51811
rect 59895 -51840 59926 -51811
rect 60096 -51683 60127 -51680
rect 60127 -51683 60161 -51680
rect 60161 -51683 60176 -51680
rect 60096 -51741 60176 -51683
rect 60096 -51775 60127 -51741
rect 60127 -51775 60161 -51741
rect 60161 -51775 60176 -51741
rect 60096 -51833 60176 -51775
rect 60096 -51840 60127 -51833
rect 60127 -51840 60161 -51833
rect 60161 -51840 60176 -51833
rect 59796 -51895 59856 -51890
rect 59796 -52070 59817 -51895
rect 59817 -52070 59851 -51895
rect 59851 -52070 59856 -51895
rect 59916 -51895 60006 -51890
rect 59916 -52071 59939 -51895
rect 59939 -52071 60006 -51895
rect 59916 -52080 60006 -52071
rect 60476 -51925 60536 -51910
rect 60476 -51959 60484 -51925
rect 60484 -51959 60536 -51925
rect 60476 -51970 60536 -51959
rect 61036 -51530 61126 -51420
rect 76920 -51490 77060 -51350
rect 78860 -51080 78980 -51010
rect 78630 -51130 78700 -51120
rect 78630 -51170 78640 -51130
rect 78640 -51170 78690 -51130
rect 78690 -51170 78700 -51130
rect 78630 -51180 78700 -51170
rect 77960 -51250 78020 -51230
rect 77960 -51290 77970 -51250
rect 77970 -51290 78010 -51250
rect 78010 -51290 78020 -51250
rect 78340 -51220 78350 -51180
rect 78350 -51220 78400 -51180
rect 78400 -51220 78410 -51180
rect 78340 -51240 78410 -51220
rect 78860 -51130 78900 -51080
rect 78900 -51130 78980 -51080
rect 78860 -51200 78980 -51130
rect 78860 -51250 78900 -51200
rect 78900 -51250 78980 -51200
rect 80010 -51330 80360 -50950
rect 82820 -51100 91410 -50530
rect 77200 -51630 77260 -51570
rect 61276 -51683 61291 -51650
rect 61291 -51683 61325 -51650
rect 61325 -51683 61356 -51650
rect 61276 -51741 61356 -51683
rect 61276 -51775 61291 -51741
rect 61291 -51775 61325 -51741
rect 61325 -51775 61356 -51741
rect 61276 -51833 61356 -51775
rect 61276 -51860 61291 -51833
rect 61291 -51860 61325 -51833
rect 61325 -51860 61356 -51833
rect 77860 -51580 77920 -51540
rect 77860 -51620 77870 -51580
rect 77870 -51620 77910 -51580
rect 77910 -51620 77920 -51580
rect 77860 -51660 77920 -51620
rect 77860 -51700 77870 -51660
rect 77870 -51700 77910 -51660
rect 77910 -51700 77920 -51660
rect 77860 -51710 77920 -51700
rect 78240 -51550 78300 -51540
rect 78240 -51600 78280 -51550
rect 78280 -51600 78300 -51550
rect 77970 -51670 78030 -51660
rect 77970 -51710 78010 -51670
rect 78010 -51710 78030 -51670
rect 77970 -51720 78030 -51710
rect 78240 -51690 78300 -51600
rect 78240 -51740 78280 -51690
rect 78280 -51740 78300 -51690
rect 77430 -51810 77500 -51800
rect 77430 -51860 77440 -51810
rect 77440 -51860 77490 -51810
rect 77490 -51860 77500 -51810
rect 77430 -51870 77500 -51860
rect 78240 -51830 78300 -51740
rect 78240 -51880 78280 -51830
rect 78280 -51880 78300 -51830
rect 78240 -51910 78300 -51880
rect 82290 -51790 82440 -51680
rect 83030 -51690 83100 -51680
rect 83030 -51780 83040 -51690
rect 83040 -51780 83090 -51690
rect 83090 -51780 83100 -51690
rect 83030 -51790 83100 -51780
rect 85320 -51610 85390 -51600
rect 85320 -51780 85330 -51610
rect 85330 -51780 85380 -51610
rect 85380 -51780 85390 -51610
rect 85320 -51790 85390 -51780
rect 85590 -51687 86480 -51660
rect 85590 -51721 85610 -51687
rect 85610 -51721 86471 -51687
rect 86471 -51721 86480 -51687
rect 85590 -51740 86480 -51721
rect 86800 -51590 86870 -51580
rect 86800 -51780 86810 -51590
rect 86810 -51780 86860 -51590
rect 86860 -51780 86870 -51590
rect 86800 -51790 86870 -51780
rect 87040 -51686 87920 -51660
rect 87040 -51720 87044 -51686
rect 87044 -51720 87905 -51686
rect 87905 -51720 87920 -51686
rect 87040 -51740 87920 -51720
rect 88270 -51600 88340 -51590
rect 88270 -51780 88280 -51600
rect 88280 -51780 88330 -51600
rect 88330 -51780 88340 -51600
rect 88270 -51790 88340 -51780
rect 88510 -51686 89390 -51670
rect 88510 -51720 88523 -51686
rect 88523 -51720 89384 -51686
rect 89384 -51720 89390 -51686
rect 88510 -51740 89390 -51720
rect 89740 -51600 89810 -51590
rect 89740 -51790 89750 -51600
rect 89750 -51790 89800 -51600
rect 89800 -51790 89810 -51600
rect 89740 -51800 89810 -51790
rect 89982 -51687 90762 -51669
rect 89982 -51689 90747 -51687
rect 90747 -51689 90762 -51687
rect 89982 -51723 90748 -51689
rect 90748 -51723 90762 -51689
rect 89982 -51741 90762 -51723
rect 91210 -51600 91280 -51590
rect 91210 -51790 91220 -51600
rect 91220 -51790 91270 -51600
rect 91270 -51790 91280 -51600
rect 91210 -51800 91280 -51790
rect 60476 -52060 60536 -52050
rect 60476 -52100 60486 -52060
rect 60486 -52100 60526 -52060
rect 60526 -52100 60536 -52060
rect 60476 -52110 60536 -52100
rect 60616 -52060 60736 -52050
rect 60616 -52100 60626 -52060
rect 60626 -52100 60666 -52060
rect 60666 -52100 60736 -52060
rect 60616 -52110 60736 -52100
rect 60756 -52060 60816 -52050
rect 60756 -52100 60766 -52060
rect 60766 -52100 60806 -52060
rect 60806 -52100 60816 -52060
rect 60756 -52110 60816 -52100
rect 60896 -52060 60956 -52050
rect 60896 -52100 60906 -52060
rect 60906 -52100 60946 -52060
rect 60946 -52100 60956 -52060
rect 60896 -52110 60956 -52100
rect 56380 -52488 56440 -52368
rect 55880 -52680 55970 -52678
rect 55880 -52714 55882 -52680
rect 55882 -52714 55970 -52680
rect 55880 -52758 55970 -52714
rect 55220 -53128 55330 -53018
rect 55530 -53202 55610 -53178
rect 55530 -53236 55560 -53202
rect 55560 -53236 55610 -53202
rect 55530 -53268 55610 -53236
rect 54140 -53308 54150 -53288
rect 54150 -53308 54840 -53288
rect 54840 -53308 54850 -53288
rect 54140 -53548 54850 -53308
rect 55320 -53348 55470 -53328
rect 55320 -53408 55470 -53348
rect 55320 -53468 55470 -53408
rect 56020 -53008 56080 -52858
rect 56170 -53008 56390 -52808
rect 56654 -53086 56998 -52868
rect 59076 -52370 59103 -52340
rect 59103 -52370 59137 -52340
rect 59137 -52370 59166 -52340
rect 59076 -52400 59166 -52370
rect 58926 -52510 58986 -52460
rect 58926 -52530 58966 -52510
rect 58966 -52530 58986 -52510
rect 59146 -52530 59226 -52460
rect 59276 -52530 59356 -52460
rect 59396 -52530 59476 -52460
rect 59646 -52520 59706 -52460
rect 59546 -52608 59606 -52600
rect 59256 -52662 59366 -52630
rect 59546 -52642 59560 -52608
rect 59560 -52642 59594 -52608
rect 59594 -52642 59606 -52608
rect 59016 -52716 59076 -52700
rect 59256 -52690 59366 -52662
rect 59546 -52660 59606 -52642
rect 59016 -52750 59032 -52716
rect 59032 -52750 59066 -52716
rect 59066 -52750 59076 -52716
rect 59016 -52760 59076 -52750
rect 58906 -52900 58926 -52830
rect 58926 -52900 58966 -52830
rect 58966 -52900 58986 -52830
rect 59146 -52900 59226 -52830
rect 59276 -52900 59356 -52830
rect 59396 -52900 59476 -52830
rect 59966 -52340 60326 -52320
rect 59966 -52374 60326 -52340
rect 79410 -52140 79680 -51900
rect 75940 -52280 76050 -52190
rect 59966 -52380 60326 -52374
rect 59856 -52394 59916 -52380
rect 59856 -52428 59874 -52394
rect 59874 -52428 59908 -52394
rect 59908 -52428 59916 -52394
rect 59856 -52440 59916 -52428
rect 60376 -52394 60436 -52380
rect 60376 -52428 60384 -52394
rect 60384 -52428 60418 -52394
rect 60418 -52428 60436 -52394
rect 60376 -52440 60436 -52428
rect 61056 -52440 61126 -52340
rect 75660 -52370 75760 -52310
rect 77760 -52480 77820 -52460
rect 77760 -52520 77770 -52480
rect 77770 -52520 77810 -52480
rect 77810 -52520 77820 -52480
rect 77970 -52400 78030 -52390
rect 77970 -52500 78010 -52400
rect 78010 -52500 78030 -52400
rect 77970 -52510 78030 -52500
rect 78180 -52180 78300 -52170
rect 78180 -52500 78290 -52180
rect 78290 -52500 78300 -52180
rect 78180 -52510 78300 -52500
rect 59806 -52720 59916 -52610
rect 60446 -52750 60526 -52630
rect 76920 -52650 77060 -52560
rect 59646 -52900 59706 -52840
rect 77760 -52820 77770 -52780
rect 77770 -52820 77810 -52780
rect 77810 -52820 77820 -52780
rect 77760 -52840 77820 -52820
rect 82820 -52800 91410 -52230
rect 91780 -52250 92130 -51870
rect 75940 -52940 76050 -52880
rect 77960 -52900 78020 -52890
rect 77960 -52950 78010 -52900
rect 78010 -52950 78020 -52900
rect 77960 -52960 78020 -52950
rect 75230 -53100 75330 -53010
rect 78640 -53130 78750 -52990
rect 58986 -53360 59126 -53220
rect 59996 -53300 60106 -53190
rect 76500 -53460 76600 -53390
rect 79410 -53400 79680 -53160
rect 75230 -53610 75330 -53540
rect 76920 -53780 77060 -53680
rect 77600 -53660 77710 -53650
rect 77600 -53710 77620 -53660
rect 77620 -53710 77690 -53660
rect 77690 -53710 77710 -53660
rect 77600 -53720 77710 -53710
rect 78070 -53530 78140 -53520
rect 78070 -53620 78080 -53530
rect 78080 -53620 78130 -53530
rect 78130 -53620 78140 -53530
rect 78070 -53630 78140 -53620
rect 78240 -53590 78300 -53570
rect 78240 -53630 78250 -53590
rect 78250 -53630 78290 -53590
rect 78290 -53630 78300 -53590
rect 78640 -53560 78740 -53550
rect 78640 -53630 78650 -53560
rect 78650 -53630 78730 -53560
rect 78730 -53630 78740 -53560
rect 78640 -53640 78740 -53630
rect 78810 -53600 78870 -53590
rect 78810 -53640 78820 -53600
rect 78820 -53640 78860 -53600
rect 78860 -53640 78870 -53600
rect 78810 -53650 78870 -53640
rect 79080 -53720 79190 -53420
rect 55400 -54300 56100 -53900
rect 80010 -53850 80360 -53470
rect 36000 -55500 38800 -54500
rect 55460 -55160 55720 -54880
rect 53480 -55740 53780 -55540
rect 54150 -55508 54860 -55338
rect 54150 -55578 54850 -55508
rect 54850 -55578 54860 -55508
rect 36000 -57100 37700 -56100
rect 53520 -55968 53640 -55858
rect 54750 -55908 54850 -55838
rect 54750 -55918 54840 -55908
rect 55430 -55888 55520 -55818
rect 55290 -55998 55390 -55928
rect 53050 -57908 53250 -56158
rect 53950 -56128 53998 -56098
rect 53998 -56128 54020 -56098
rect 53950 -56198 54020 -56128
rect 54920 -56090 54990 -56078
rect 54920 -56128 54926 -56090
rect 54926 -56128 54960 -56090
rect 54960 -56128 54990 -56090
rect 54920 -56168 54990 -56128
rect 53860 -56638 53920 -56528
rect 55230 -56428 55290 -56258
rect 55290 -56428 55320 -56258
rect 55430 -56418 55510 -56248
rect 55960 -55888 56040 -55738
rect 56190 -55968 56390 -55758
rect 56506 -55830 57016 -55580
rect 58966 -55630 59126 -55470
rect 59956 -55660 60166 -55500
rect 55880 -56056 55970 -56018
rect 55880 -56090 55882 -56056
rect 55882 -56090 55970 -56056
rect 55880 -56098 55970 -56090
rect 55000 -56638 55090 -56538
rect 54770 -56840 54840 -56838
rect 54770 -56928 54802 -56840
rect 54802 -56928 54840 -56840
rect 55540 -56638 55630 -56538
rect 56590 -56398 56660 -56268
rect 58906 -56020 58966 -55970
rect 58906 -56030 58926 -56020
rect 58926 -56030 58966 -56020
rect 59216 -56030 59276 -55970
rect 59326 -56030 59386 -55970
rect 59436 -56030 59496 -55970
rect 59636 -56030 59696 -55970
rect 59546 -56101 59606 -56090
rect 59286 -56155 59346 -56130
rect 59546 -56135 59560 -56101
rect 59560 -56135 59594 -56101
rect 59594 -56135 59606 -56101
rect 59286 -56189 59346 -56155
rect 59546 -56150 59606 -56135
rect 59286 -56190 59346 -56189
rect 59016 -56209 59076 -56200
rect 59016 -56243 59032 -56209
rect 59032 -56243 59066 -56209
rect 59066 -56243 59076 -56209
rect 59016 -56260 59076 -56243
rect 59546 -56270 59606 -56210
rect 58906 -56390 58966 -56330
rect 59216 -56380 59276 -56320
rect 59336 -56380 59396 -56320
rect 59436 -56380 59496 -56320
rect 55140 -57008 55200 -56938
rect 55030 -57128 55110 -57048
rect 55740 -57128 55810 -57048
rect 55880 -57128 55970 -57038
rect 56480 -56606 56550 -56588
rect 56480 -56640 56492 -56606
rect 56492 -56640 56530 -56606
rect 56530 -56640 56550 -56606
rect 56480 -56648 56550 -56640
rect 59866 -56230 59966 -56140
rect 60446 -56220 60526 -56120
rect 59636 -56390 59696 -56330
rect 59076 -56478 59166 -56440
rect 59076 -56510 59103 -56478
rect 59103 -56510 59137 -56478
rect 59137 -56510 59166 -56478
rect 60046 -56374 60126 -56340
rect 59856 -56428 59916 -56410
rect 60046 -56400 60126 -56374
rect 59856 -56462 59874 -56428
rect 59874 -56462 59908 -56428
rect 59908 -56462 59916 -56428
rect 59856 -56480 59916 -56462
rect 60376 -56428 60446 -56420
rect 60376 -56462 60384 -56428
rect 60384 -56462 60418 -56428
rect 60418 -56462 60446 -56428
rect 59976 -56516 60316 -56500
rect 60376 -56480 60446 -56462
rect 57098 -56589 57368 -56564
rect 57098 -56623 57125 -56589
rect 57125 -56623 57159 -56589
rect 57159 -56623 57217 -56589
rect 57217 -56623 57251 -56589
rect 57251 -56623 57309 -56589
rect 57309 -56623 57343 -56589
rect 57343 -56623 57368 -56589
rect 54770 -57328 54802 -57248
rect 54802 -57328 54840 -57248
rect 53850 -57648 53920 -57538
rect 54920 -57468 54980 -57398
rect 55000 -57638 55090 -57538
rect 55540 -57638 55630 -57538
rect 55220 -57918 55280 -57748
rect 55280 -57918 55310 -57748
rect 55410 -57928 55500 -57758
rect 53950 -58050 54010 -58008
rect 53950 -58088 53988 -58050
rect 53988 -58088 54010 -58050
rect 54910 -58050 54980 -57998
rect 54910 -58088 54916 -58050
rect 54916 -58088 54950 -58050
rect 54950 -58088 54980 -58050
rect 54910 -58098 54980 -58088
rect 53510 -58248 53630 -58128
rect 54740 -58344 54850 -58268
rect 54740 -58358 54850 -58344
rect 55240 -58218 55370 -58158
rect 55410 -58338 55510 -58248
rect 57098 -56680 57368 -56623
rect 57098 -56704 57368 -56680
rect 56900 -57148 57020 -57018
rect 58576 -57240 58736 -57080
rect 57098 -57480 57368 -57474
rect 56480 -57534 56550 -57528
rect 56480 -57568 56492 -57534
rect 56492 -57568 56530 -57534
rect 56530 -57568 56550 -57534
rect 56480 -57588 56550 -57568
rect 57098 -57565 57368 -57480
rect 57098 -57599 57125 -57565
rect 57125 -57599 57159 -57565
rect 57159 -57599 57217 -57565
rect 57217 -57599 57251 -57565
rect 57251 -57599 57309 -57565
rect 57309 -57599 57343 -57565
rect 57343 -57599 57368 -57565
rect 57098 -57614 57368 -57599
rect 59976 -56552 60316 -56516
rect 59176 -56720 59196 -56640
rect 59196 -56720 59236 -56640
rect 59176 -56920 59196 -56840
rect 59196 -56920 59236 -56840
rect 59076 -57040 59103 -57010
rect 59103 -57040 59137 -57010
rect 59137 -57040 59166 -57010
rect 59076 -57080 59166 -57040
rect 59576 -56698 59636 -56670
rect 59576 -56730 59580 -56698
rect 59580 -56730 59636 -56698
rect 59476 -56920 59502 -56850
rect 59502 -56920 59536 -56850
rect 59576 -56958 59590 -56790
rect 59590 -56958 59624 -56790
rect 59624 -56958 59636 -56790
rect 59576 -56960 59636 -56958
rect 59076 -57208 59166 -57170
rect 59076 -57240 59103 -57208
rect 59103 -57240 59137 -57208
rect 59137 -57240 59166 -57208
rect 59206 -57240 59266 -57170
rect 61206 -56700 61346 -56520
rect 59806 -56940 59818 -56800
rect 59818 -56940 59852 -56800
rect 59852 -56940 59866 -56800
rect 59916 -56782 60006 -56780
rect 59916 -56958 59940 -56782
rect 59940 -56958 60006 -56782
rect 59916 -56960 60006 -56958
rect 60306 -56890 60456 -56750
rect 59826 -57042 59862 -57010
rect 59862 -57042 59896 -57010
rect 59896 -57042 59916 -57010
rect 59826 -57080 59916 -57042
rect 59166 -57410 59196 -57330
rect 59196 -57410 59226 -57330
rect 59166 -57640 59196 -57560
rect 59196 -57640 59226 -57560
rect 59466 -57410 59501 -57330
rect 59501 -57410 59526 -57330
rect 59586 -57450 59589 -57310
rect 59589 -57450 59623 -57310
rect 59623 -57450 59646 -57310
rect 59516 -57521 59596 -57520
rect 59516 -57555 59545 -57521
rect 59545 -57555 59579 -57521
rect 59579 -57555 59596 -57521
rect 59516 -57580 59596 -57555
rect 59826 -57211 59926 -57170
rect 59826 -57240 59861 -57211
rect 59861 -57240 59895 -57211
rect 59895 -57240 59926 -57211
rect 60096 -57083 60127 -57080
rect 60127 -57083 60161 -57080
rect 60161 -57083 60176 -57080
rect 60096 -57141 60176 -57083
rect 60096 -57175 60127 -57141
rect 60127 -57175 60161 -57141
rect 60161 -57175 60176 -57141
rect 60096 -57233 60176 -57175
rect 60096 -57240 60127 -57233
rect 60127 -57240 60161 -57233
rect 60161 -57240 60176 -57233
rect 59796 -57295 59856 -57290
rect 59796 -57470 59817 -57295
rect 59817 -57470 59851 -57295
rect 59851 -57470 59856 -57295
rect 59916 -57295 60006 -57290
rect 59916 -57471 59939 -57295
rect 59939 -57471 60006 -57295
rect 59916 -57480 60006 -57471
rect 60476 -57325 60536 -57310
rect 60476 -57359 60484 -57325
rect 60484 -57359 60536 -57325
rect 60476 -57370 60536 -57359
rect 61036 -56930 61126 -56820
rect 61276 -57083 61291 -57050
rect 61291 -57083 61325 -57050
rect 61325 -57083 61356 -57050
rect 61276 -57141 61356 -57083
rect 61276 -57175 61291 -57141
rect 61291 -57175 61325 -57141
rect 61325 -57175 61356 -57141
rect 61276 -57233 61356 -57175
rect 61276 -57260 61291 -57233
rect 61291 -57260 61325 -57233
rect 61325 -57260 61356 -57233
rect 60476 -57460 60536 -57450
rect 60476 -57500 60486 -57460
rect 60486 -57500 60526 -57460
rect 60526 -57500 60536 -57460
rect 60476 -57510 60536 -57500
rect 60616 -57460 60736 -57450
rect 60616 -57500 60626 -57460
rect 60626 -57500 60666 -57460
rect 60666 -57500 60736 -57460
rect 60616 -57510 60736 -57500
rect 60756 -57460 60816 -57450
rect 60756 -57500 60766 -57460
rect 60766 -57500 60806 -57460
rect 60806 -57500 60816 -57460
rect 60756 -57510 60816 -57500
rect 60896 -57460 60956 -57450
rect 60896 -57500 60906 -57460
rect 60906 -57500 60946 -57460
rect 60946 -57500 60956 -57460
rect 60896 -57510 60956 -57500
rect 56380 -57888 56440 -57768
rect 55880 -58080 55970 -58078
rect 55880 -58114 55882 -58080
rect 55882 -58114 55970 -58080
rect 55880 -58158 55970 -58114
rect 55220 -58528 55330 -58418
rect 55530 -58602 55610 -58578
rect 55530 -58636 55560 -58602
rect 55560 -58636 55610 -58602
rect 55530 -58668 55610 -58636
rect 54140 -58708 54150 -58688
rect 54150 -58708 54840 -58688
rect 54840 -58708 54850 -58688
rect 15200 -64800 19600 -60000
rect 25000 -64800 35400 -58800
rect 54140 -58948 54850 -58708
rect 55320 -58748 55470 -58728
rect 55320 -58808 55470 -58748
rect 55320 -58868 55470 -58808
rect 56020 -58408 56080 -58258
rect 56170 -58408 56390 -58208
rect 56654 -58486 56998 -58268
rect 59076 -57770 59103 -57740
rect 59103 -57770 59137 -57740
rect 59137 -57770 59166 -57740
rect 59076 -57800 59166 -57770
rect 58926 -57910 58986 -57860
rect 58926 -57930 58966 -57910
rect 58966 -57930 58986 -57910
rect 59146 -57930 59226 -57860
rect 59276 -57930 59356 -57860
rect 59396 -57930 59476 -57860
rect 59646 -57920 59706 -57860
rect 59546 -58008 59606 -58000
rect 59256 -58062 59366 -58030
rect 59546 -58042 59560 -58008
rect 59560 -58042 59594 -58008
rect 59594 -58042 59606 -58008
rect 59016 -58116 59076 -58100
rect 59256 -58090 59366 -58062
rect 59546 -58060 59606 -58042
rect 59016 -58150 59032 -58116
rect 59032 -58150 59066 -58116
rect 59066 -58150 59076 -58116
rect 59016 -58160 59076 -58150
rect 58906 -58300 58926 -58230
rect 58926 -58300 58966 -58230
rect 58966 -58300 58986 -58230
rect 59146 -58300 59226 -58230
rect 59276 -58300 59356 -58230
rect 59396 -58300 59476 -58230
rect 59966 -57740 60326 -57720
rect 59966 -57774 60326 -57740
rect 59966 -57780 60326 -57774
rect 59856 -57794 59916 -57780
rect 59856 -57828 59874 -57794
rect 59874 -57828 59908 -57794
rect 59908 -57828 59916 -57794
rect 59856 -57840 59916 -57828
rect 60376 -57794 60436 -57780
rect 60376 -57828 60384 -57794
rect 60384 -57828 60418 -57794
rect 60418 -57828 60436 -57794
rect 60376 -57840 60436 -57828
rect 61056 -57840 61126 -57740
rect 59806 -58120 59916 -58010
rect 60446 -58150 60526 -58030
rect 59646 -58300 59706 -58240
rect 58986 -58760 59126 -58620
rect 59996 -58700 60106 -58590
rect 55500 -59700 56100 -59300
rect 55460 -60560 55720 -60280
rect 53480 -61140 53780 -60940
rect 54150 -60908 54860 -60738
rect 54150 -60978 54850 -60908
rect 54850 -60978 54860 -60908
rect 53520 -61368 53640 -61258
rect 54750 -61308 54850 -61238
rect 54750 -61318 54840 -61308
rect 55430 -61288 55520 -61218
rect 55290 -61398 55390 -61328
rect 53050 -63308 53250 -61558
rect 53950 -61528 53998 -61498
rect 53998 -61528 54020 -61498
rect 53950 -61598 54020 -61528
rect 54920 -61490 54990 -61478
rect 54920 -61528 54926 -61490
rect 54926 -61528 54960 -61490
rect 54960 -61528 54990 -61490
rect 54920 -61568 54990 -61528
rect 53860 -62038 53920 -61928
rect 55230 -61828 55290 -61658
rect 55290 -61828 55320 -61658
rect 55430 -61818 55510 -61648
rect 55960 -61288 56040 -61138
rect 56190 -61368 56390 -61158
rect 56506 -61230 57016 -60980
rect 58966 -61030 59126 -60870
rect 59956 -61060 60166 -60900
rect 55880 -61456 55970 -61418
rect 55880 -61490 55882 -61456
rect 55882 -61490 55970 -61456
rect 55880 -61498 55970 -61490
rect 55000 -62038 55090 -61938
rect 54770 -62240 54840 -62238
rect 54770 -62328 54802 -62240
rect 54802 -62328 54840 -62240
rect 55540 -62038 55630 -61938
rect 56590 -61798 56660 -61668
rect 58906 -61420 58966 -61370
rect 58906 -61430 58926 -61420
rect 58926 -61430 58966 -61420
rect 59216 -61430 59276 -61370
rect 59326 -61430 59386 -61370
rect 59436 -61430 59496 -61370
rect 59636 -61430 59696 -61370
rect 59546 -61501 59606 -61490
rect 59286 -61555 59346 -61530
rect 59546 -61535 59560 -61501
rect 59560 -61535 59594 -61501
rect 59594 -61535 59606 -61501
rect 59286 -61589 59346 -61555
rect 59546 -61550 59606 -61535
rect 59286 -61590 59346 -61589
rect 59016 -61609 59076 -61600
rect 59016 -61643 59032 -61609
rect 59032 -61643 59066 -61609
rect 59066 -61643 59076 -61609
rect 59016 -61660 59076 -61643
rect 59546 -61670 59606 -61610
rect 58906 -61790 58966 -61730
rect 59216 -61780 59276 -61720
rect 59336 -61780 59396 -61720
rect 59436 -61780 59496 -61720
rect 55140 -62408 55200 -62338
rect 55030 -62528 55110 -62448
rect 55740 -62528 55810 -62448
rect 55880 -62528 55970 -62438
rect 56480 -62006 56550 -61988
rect 56480 -62040 56492 -62006
rect 56492 -62040 56530 -62006
rect 56530 -62040 56550 -62006
rect 56480 -62048 56550 -62040
rect 59866 -61630 59966 -61540
rect 60446 -61620 60526 -61520
rect 59636 -61790 59696 -61730
rect 59076 -61878 59166 -61840
rect 59076 -61910 59103 -61878
rect 59103 -61910 59137 -61878
rect 59137 -61910 59166 -61878
rect 60046 -61774 60126 -61740
rect 59856 -61828 59916 -61810
rect 60046 -61800 60126 -61774
rect 59856 -61862 59874 -61828
rect 59874 -61862 59908 -61828
rect 59908 -61862 59916 -61828
rect 59856 -61880 59916 -61862
rect 60376 -61828 60446 -61820
rect 60376 -61862 60384 -61828
rect 60384 -61862 60418 -61828
rect 60418 -61862 60446 -61828
rect 59976 -61916 60316 -61900
rect 60376 -61880 60446 -61862
rect 57098 -61989 57368 -61964
rect 57098 -62023 57125 -61989
rect 57125 -62023 57159 -61989
rect 57159 -62023 57217 -61989
rect 57217 -62023 57251 -61989
rect 57251 -62023 57309 -61989
rect 57309 -62023 57343 -61989
rect 57343 -62023 57368 -61989
rect 54770 -62728 54802 -62648
rect 54802 -62728 54840 -62648
rect 53850 -63048 53920 -62938
rect 54920 -62868 54980 -62798
rect 55000 -63038 55090 -62938
rect 55540 -63038 55630 -62938
rect 55220 -63318 55280 -63148
rect 55280 -63318 55310 -63148
rect 55410 -63328 55500 -63158
rect 53950 -63450 54010 -63408
rect 53950 -63488 53988 -63450
rect 53988 -63488 54010 -63450
rect 54910 -63450 54980 -63398
rect 54910 -63488 54916 -63450
rect 54916 -63488 54950 -63450
rect 54950 -63488 54980 -63450
rect 54910 -63498 54980 -63488
rect 53510 -63648 53630 -63528
rect 54740 -63744 54850 -63668
rect 54740 -63758 54850 -63744
rect 55240 -63618 55370 -63558
rect 55410 -63738 55510 -63648
rect 57098 -62080 57368 -62023
rect 57098 -62104 57368 -62080
rect 56900 -62548 57020 -62418
rect 58576 -62640 58736 -62480
rect 57098 -62880 57368 -62874
rect 56480 -62934 56550 -62928
rect 56480 -62968 56492 -62934
rect 56492 -62968 56530 -62934
rect 56530 -62968 56550 -62934
rect 56480 -62988 56550 -62968
rect 57098 -62965 57368 -62880
rect 57098 -62999 57125 -62965
rect 57125 -62999 57159 -62965
rect 57159 -62999 57217 -62965
rect 57217 -62999 57251 -62965
rect 57251 -62999 57309 -62965
rect 57309 -62999 57343 -62965
rect 57343 -62999 57368 -62965
rect 57098 -63014 57368 -62999
rect 59976 -61952 60316 -61916
rect 59176 -62120 59196 -62040
rect 59196 -62120 59236 -62040
rect 59176 -62320 59196 -62240
rect 59196 -62320 59236 -62240
rect 59076 -62440 59103 -62410
rect 59103 -62440 59137 -62410
rect 59137 -62440 59166 -62410
rect 59076 -62480 59166 -62440
rect 59576 -62098 59636 -62070
rect 59576 -62130 59580 -62098
rect 59580 -62130 59636 -62098
rect 59476 -62320 59502 -62250
rect 59502 -62320 59536 -62250
rect 59576 -62358 59590 -62190
rect 59590 -62358 59624 -62190
rect 59624 -62358 59636 -62190
rect 59576 -62360 59636 -62358
rect 59076 -62608 59166 -62570
rect 59076 -62640 59103 -62608
rect 59103 -62640 59137 -62608
rect 59137 -62640 59166 -62608
rect 59206 -62640 59266 -62570
rect 61206 -62100 61346 -61920
rect 59806 -62340 59818 -62200
rect 59818 -62340 59852 -62200
rect 59852 -62340 59866 -62200
rect 59916 -62182 60006 -62180
rect 59916 -62358 59940 -62182
rect 59940 -62358 60006 -62182
rect 59916 -62360 60006 -62358
rect 60306 -62290 60456 -62150
rect 59826 -62442 59862 -62410
rect 59862 -62442 59896 -62410
rect 59896 -62442 59916 -62410
rect 59826 -62480 59916 -62442
rect 59166 -62810 59196 -62730
rect 59196 -62810 59226 -62730
rect 59166 -63040 59196 -62960
rect 59196 -63040 59226 -62960
rect 59466 -62810 59501 -62730
rect 59501 -62810 59526 -62730
rect 59586 -62850 59589 -62710
rect 59589 -62850 59623 -62710
rect 59623 -62850 59646 -62710
rect 59516 -62921 59596 -62920
rect 59516 -62955 59545 -62921
rect 59545 -62955 59579 -62921
rect 59579 -62955 59596 -62921
rect 59516 -62980 59596 -62955
rect 59826 -62611 59926 -62570
rect 59826 -62640 59861 -62611
rect 59861 -62640 59895 -62611
rect 59895 -62640 59926 -62611
rect 60096 -62483 60127 -62480
rect 60127 -62483 60161 -62480
rect 60161 -62483 60176 -62480
rect 60096 -62541 60176 -62483
rect 60096 -62575 60127 -62541
rect 60127 -62575 60161 -62541
rect 60161 -62575 60176 -62541
rect 60096 -62633 60176 -62575
rect 60096 -62640 60127 -62633
rect 60127 -62640 60161 -62633
rect 60161 -62640 60176 -62633
rect 59796 -62695 59856 -62690
rect 59796 -62870 59817 -62695
rect 59817 -62870 59851 -62695
rect 59851 -62870 59856 -62695
rect 59916 -62695 60006 -62690
rect 59916 -62871 59939 -62695
rect 59939 -62871 60006 -62695
rect 59916 -62880 60006 -62871
rect 60476 -62725 60536 -62710
rect 60476 -62759 60484 -62725
rect 60484 -62759 60536 -62725
rect 60476 -62770 60536 -62759
rect 61036 -62330 61126 -62220
rect 61276 -62483 61291 -62450
rect 61291 -62483 61325 -62450
rect 61325 -62483 61356 -62450
rect 61276 -62541 61356 -62483
rect 61276 -62575 61291 -62541
rect 61291 -62575 61325 -62541
rect 61325 -62575 61356 -62541
rect 61276 -62633 61356 -62575
rect 61276 -62660 61291 -62633
rect 61291 -62660 61325 -62633
rect 61325 -62660 61356 -62633
rect 60476 -62860 60536 -62850
rect 60476 -62900 60486 -62860
rect 60486 -62900 60526 -62860
rect 60526 -62900 60536 -62860
rect 60476 -62910 60536 -62900
rect 60616 -62860 60736 -62850
rect 60616 -62900 60626 -62860
rect 60626 -62900 60666 -62860
rect 60666 -62900 60736 -62860
rect 60616 -62910 60736 -62900
rect 60756 -62860 60816 -62850
rect 60756 -62900 60766 -62860
rect 60766 -62900 60806 -62860
rect 60806 -62900 60816 -62860
rect 60756 -62910 60816 -62900
rect 60896 -62860 60956 -62850
rect 60896 -62900 60906 -62860
rect 60906 -62900 60946 -62860
rect 60946 -62900 60956 -62860
rect 60896 -62910 60956 -62900
rect 56380 -63288 56440 -63168
rect 55880 -63480 55970 -63478
rect 55880 -63514 55882 -63480
rect 55882 -63514 55970 -63480
rect 55880 -63558 55970 -63514
rect 55220 -63928 55330 -63818
rect 55530 -64002 55610 -63978
rect 55530 -64036 55560 -64002
rect 55560 -64036 55610 -64002
rect 55530 -64068 55610 -64036
rect 54140 -64108 54150 -64088
rect 54150 -64108 54840 -64088
rect 54840 -64108 54850 -64088
rect 54140 -64348 54850 -64108
rect 55320 -64148 55470 -64128
rect 55320 -64208 55470 -64148
rect 55320 -64268 55470 -64208
rect 56020 -63808 56080 -63658
rect 56170 -63808 56390 -63608
rect 56654 -63886 56998 -63668
rect 59076 -63170 59103 -63140
rect 59103 -63170 59137 -63140
rect 59137 -63170 59166 -63140
rect 59076 -63200 59166 -63170
rect 58926 -63310 58986 -63260
rect 58926 -63330 58966 -63310
rect 58966 -63330 58986 -63310
rect 59146 -63330 59226 -63260
rect 59276 -63330 59356 -63260
rect 59396 -63330 59476 -63260
rect 59646 -63320 59706 -63260
rect 59546 -63408 59606 -63400
rect 59256 -63462 59366 -63430
rect 59546 -63442 59560 -63408
rect 59560 -63442 59594 -63408
rect 59594 -63442 59606 -63408
rect 59016 -63516 59076 -63500
rect 59256 -63490 59366 -63462
rect 59546 -63460 59606 -63442
rect 59016 -63550 59032 -63516
rect 59032 -63550 59066 -63516
rect 59066 -63550 59076 -63516
rect 59016 -63560 59076 -63550
rect 58906 -63700 58926 -63630
rect 58926 -63700 58966 -63630
rect 58966 -63700 58986 -63630
rect 59146 -63700 59226 -63630
rect 59276 -63700 59356 -63630
rect 59396 -63700 59476 -63630
rect 59966 -63140 60326 -63120
rect 59966 -63174 60326 -63140
rect 59966 -63180 60326 -63174
rect 59856 -63194 59916 -63180
rect 59856 -63228 59874 -63194
rect 59874 -63228 59908 -63194
rect 59908 -63228 59916 -63194
rect 59856 -63240 59916 -63228
rect 60376 -63194 60436 -63180
rect 60376 -63228 60384 -63194
rect 60384 -63228 60418 -63194
rect 60418 -63228 60436 -63194
rect 60376 -63240 60436 -63228
rect 61056 -63240 61126 -63140
rect 59806 -63520 59916 -63410
rect 60446 -63550 60526 -63430
rect 59646 -63700 59706 -63640
rect 58986 -64160 59126 -64020
rect 59996 -64100 60106 -63990
rect 55500 -65100 56100 -64700
rect 55440 -65960 55720 -65680
rect 53480 -66540 53780 -66340
rect 54150 -66308 54860 -66138
rect 54150 -66378 54850 -66308
rect 54850 -66378 54860 -66308
rect 53520 -66768 53640 -66658
rect 54750 -66708 54850 -66638
rect 54750 -66718 54840 -66708
rect 55430 -66688 55520 -66618
rect 55290 -66798 55390 -66728
rect 53050 -68708 53250 -66958
rect 53950 -66928 53998 -66898
rect 53998 -66928 54020 -66898
rect 53950 -66998 54020 -66928
rect 54920 -66890 54990 -66878
rect 54920 -66928 54926 -66890
rect 54926 -66928 54960 -66890
rect 54960 -66928 54990 -66890
rect 54920 -66968 54990 -66928
rect 53860 -67438 53920 -67328
rect 55230 -67228 55290 -67058
rect 55290 -67228 55320 -67058
rect 55430 -67218 55510 -67048
rect 55960 -66688 56040 -66538
rect 56190 -66768 56390 -66558
rect 56506 -66630 57016 -66380
rect 58966 -66430 59126 -66270
rect 59956 -66460 60166 -66300
rect 55880 -66856 55970 -66818
rect 55880 -66890 55882 -66856
rect 55882 -66890 55970 -66856
rect 55880 -66898 55970 -66890
rect 55000 -67438 55090 -67338
rect 54770 -67640 54840 -67638
rect 54770 -67728 54802 -67640
rect 54802 -67728 54840 -67640
rect 55540 -67438 55630 -67338
rect 56590 -67198 56660 -67068
rect 58906 -66820 58966 -66770
rect 58906 -66830 58926 -66820
rect 58926 -66830 58966 -66820
rect 59216 -66830 59276 -66770
rect 59326 -66830 59386 -66770
rect 59436 -66830 59496 -66770
rect 59636 -66830 59696 -66770
rect 59546 -66901 59606 -66890
rect 59286 -66955 59346 -66930
rect 59546 -66935 59560 -66901
rect 59560 -66935 59594 -66901
rect 59594 -66935 59606 -66901
rect 59286 -66989 59346 -66955
rect 59546 -66950 59606 -66935
rect 59286 -66990 59346 -66989
rect 59016 -67009 59076 -67000
rect 59016 -67043 59032 -67009
rect 59032 -67043 59066 -67009
rect 59066 -67043 59076 -67009
rect 59016 -67060 59076 -67043
rect 59546 -67070 59606 -67010
rect 58906 -67190 58966 -67130
rect 59216 -67180 59276 -67120
rect 59336 -67180 59396 -67120
rect 59436 -67180 59496 -67120
rect 55140 -67808 55200 -67738
rect 55030 -67928 55110 -67848
rect 55740 -67928 55810 -67848
rect 55880 -67928 55970 -67838
rect 56480 -67406 56550 -67388
rect 56480 -67440 56492 -67406
rect 56492 -67440 56530 -67406
rect 56530 -67440 56550 -67406
rect 56480 -67448 56550 -67440
rect 59866 -67030 59966 -66940
rect 60446 -67020 60526 -66920
rect 59636 -67190 59696 -67130
rect 59076 -67278 59166 -67240
rect 59076 -67310 59103 -67278
rect 59103 -67310 59137 -67278
rect 59137 -67310 59166 -67278
rect 60046 -67174 60126 -67140
rect 59856 -67228 59916 -67210
rect 60046 -67200 60126 -67174
rect 59856 -67262 59874 -67228
rect 59874 -67262 59908 -67228
rect 59908 -67262 59916 -67228
rect 59856 -67280 59916 -67262
rect 60376 -67228 60446 -67220
rect 60376 -67262 60384 -67228
rect 60384 -67262 60418 -67228
rect 60418 -67262 60446 -67228
rect 59976 -67316 60316 -67300
rect 60376 -67280 60446 -67262
rect 57098 -67389 57368 -67364
rect 57098 -67423 57125 -67389
rect 57125 -67423 57159 -67389
rect 57159 -67423 57217 -67389
rect 57217 -67423 57251 -67389
rect 57251 -67423 57309 -67389
rect 57309 -67423 57343 -67389
rect 57343 -67423 57368 -67389
rect 54770 -68128 54802 -68048
rect 54802 -68128 54840 -68048
rect 53850 -68448 53920 -68338
rect 54920 -68268 54980 -68198
rect 55000 -68438 55090 -68338
rect 55540 -68438 55630 -68338
rect 55220 -68718 55280 -68548
rect 55280 -68718 55310 -68548
rect 55410 -68728 55500 -68558
rect 53950 -68850 54010 -68808
rect 53950 -68888 53988 -68850
rect 53988 -68888 54010 -68850
rect 54910 -68850 54980 -68798
rect 54910 -68888 54916 -68850
rect 54916 -68888 54950 -68850
rect 54950 -68888 54980 -68850
rect 54910 -68898 54980 -68888
rect 53510 -69048 53630 -68928
rect 54740 -69144 54850 -69068
rect 54740 -69158 54850 -69144
rect 55240 -69018 55370 -68958
rect 55410 -69138 55510 -69048
rect 57098 -67480 57368 -67423
rect 57098 -67504 57368 -67480
rect 56900 -67948 57020 -67818
rect 58576 -68040 58736 -67880
rect 57098 -68280 57368 -68274
rect 56480 -68334 56550 -68328
rect 56480 -68368 56492 -68334
rect 56492 -68368 56530 -68334
rect 56530 -68368 56550 -68334
rect 56480 -68388 56550 -68368
rect 57098 -68365 57368 -68280
rect 57098 -68399 57125 -68365
rect 57125 -68399 57159 -68365
rect 57159 -68399 57217 -68365
rect 57217 -68399 57251 -68365
rect 57251 -68399 57309 -68365
rect 57309 -68399 57343 -68365
rect 57343 -68399 57368 -68365
rect 57098 -68414 57368 -68399
rect 59976 -67352 60316 -67316
rect 59176 -67520 59196 -67440
rect 59196 -67520 59236 -67440
rect 59176 -67720 59196 -67640
rect 59196 -67720 59236 -67640
rect 59076 -67840 59103 -67810
rect 59103 -67840 59137 -67810
rect 59137 -67840 59166 -67810
rect 59076 -67880 59166 -67840
rect 59576 -67498 59636 -67470
rect 59576 -67530 59580 -67498
rect 59580 -67530 59636 -67498
rect 59476 -67720 59502 -67650
rect 59502 -67720 59536 -67650
rect 59576 -67758 59590 -67590
rect 59590 -67758 59624 -67590
rect 59624 -67758 59636 -67590
rect 59576 -67760 59636 -67758
rect 59076 -68008 59166 -67970
rect 59076 -68040 59103 -68008
rect 59103 -68040 59137 -68008
rect 59137 -68040 59166 -68008
rect 59206 -68040 59266 -67970
rect 61206 -67500 61346 -67320
rect 59806 -67740 59818 -67600
rect 59818 -67740 59852 -67600
rect 59852 -67740 59866 -67600
rect 59916 -67582 60006 -67580
rect 59916 -67758 59940 -67582
rect 59940 -67758 60006 -67582
rect 59916 -67760 60006 -67758
rect 60306 -67690 60456 -67550
rect 59826 -67842 59862 -67810
rect 59862 -67842 59896 -67810
rect 59896 -67842 59916 -67810
rect 59826 -67880 59916 -67842
rect 59166 -68210 59196 -68130
rect 59196 -68210 59226 -68130
rect 59166 -68440 59196 -68360
rect 59196 -68440 59226 -68360
rect 59466 -68210 59501 -68130
rect 59501 -68210 59526 -68130
rect 59586 -68250 59589 -68110
rect 59589 -68250 59623 -68110
rect 59623 -68250 59646 -68110
rect 59516 -68321 59596 -68320
rect 59516 -68355 59545 -68321
rect 59545 -68355 59579 -68321
rect 59579 -68355 59596 -68321
rect 59516 -68380 59596 -68355
rect 59826 -68011 59926 -67970
rect 59826 -68040 59861 -68011
rect 59861 -68040 59895 -68011
rect 59895 -68040 59926 -68011
rect 60096 -67883 60127 -67880
rect 60127 -67883 60161 -67880
rect 60161 -67883 60176 -67880
rect 60096 -67941 60176 -67883
rect 60096 -67975 60127 -67941
rect 60127 -67975 60161 -67941
rect 60161 -67975 60176 -67941
rect 60096 -68033 60176 -67975
rect 60096 -68040 60127 -68033
rect 60127 -68040 60161 -68033
rect 60161 -68040 60176 -68033
rect 59796 -68095 59856 -68090
rect 59796 -68270 59817 -68095
rect 59817 -68270 59851 -68095
rect 59851 -68270 59856 -68095
rect 59916 -68095 60006 -68090
rect 59916 -68271 59939 -68095
rect 59939 -68271 60006 -68095
rect 59916 -68280 60006 -68271
rect 60476 -68125 60536 -68110
rect 60476 -68159 60484 -68125
rect 60484 -68159 60536 -68125
rect 60476 -68170 60536 -68159
rect 61036 -67730 61126 -67620
rect 61276 -67883 61291 -67850
rect 61291 -67883 61325 -67850
rect 61325 -67883 61356 -67850
rect 61276 -67941 61356 -67883
rect 61276 -67975 61291 -67941
rect 61291 -67975 61325 -67941
rect 61325 -67975 61356 -67941
rect 61276 -68033 61356 -67975
rect 61276 -68060 61291 -68033
rect 61291 -68060 61325 -68033
rect 61325 -68060 61356 -68033
rect 60476 -68260 60536 -68250
rect 60476 -68300 60486 -68260
rect 60486 -68300 60526 -68260
rect 60526 -68300 60536 -68260
rect 60476 -68310 60536 -68300
rect 60616 -68260 60736 -68250
rect 60616 -68300 60626 -68260
rect 60626 -68300 60666 -68260
rect 60666 -68300 60736 -68260
rect 60616 -68310 60736 -68300
rect 60756 -68260 60816 -68250
rect 60756 -68300 60766 -68260
rect 60766 -68300 60806 -68260
rect 60806 -68300 60816 -68260
rect 60756 -68310 60816 -68300
rect 60896 -68260 60956 -68250
rect 60896 -68300 60906 -68260
rect 60906 -68300 60946 -68260
rect 60946 -68300 60956 -68260
rect 60896 -68310 60956 -68300
rect 56380 -68688 56440 -68568
rect 55880 -68880 55970 -68878
rect 55880 -68914 55882 -68880
rect 55882 -68914 55970 -68880
rect 55880 -68958 55970 -68914
rect 55220 -69328 55330 -69218
rect 55530 -69402 55610 -69378
rect 55530 -69436 55560 -69402
rect 55560 -69436 55610 -69402
rect 55530 -69468 55610 -69436
rect 54140 -69508 54150 -69488
rect 54150 -69508 54840 -69488
rect 54840 -69508 54850 -69488
rect 54140 -69748 54850 -69508
rect 55320 -69548 55470 -69528
rect 55320 -69608 55470 -69548
rect 55320 -69668 55470 -69608
rect 56020 -69208 56080 -69058
rect 56170 -69208 56390 -69008
rect 56654 -69286 56998 -69068
rect 59076 -68570 59103 -68540
rect 59103 -68570 59137 -68540
rect 59137 -68570 59166 -68540
rect 59076 -68600 59166 -68570
rect 58926 -68710 58986 -68660
rect 58926 -68730 58966 -68710
rect 58966 -68730 58986 -68710
rect 59146 -68730 59226 -68660
rect 59276 -68730 59356 -68660
rect 59396 -68730 59476 -68660
rect 59646 -68720 59706 -68660
rect 59546 -68808 59606 -68800
rect 59256 -68862 59366 -68830
rect 59546 -68842 59560 -68808
rect 59560 -68842 59594 -68808
rect 59594 -68842 59606 -68808
rect 59016 -68916 59076 -68900
rect 59256 -68890 59366 -68862
rect 59546 -68860 59606 -68842
rect 59016 -68950 59032 -68916
rect 59032 -68950 59066 -68916
rect 59066 -68950 59076 -68916
rect 59016 -68960 59076 -68950
rect 58906 -69100 58926 -69030
rect 58926 -69100 58966 -69030
rect 58966 -69100 58986 -69030
rect 59146 -69100 59226 -69030
rect 59276 -69100 59356 -69030
rect 59396 -69100 59476 -69030
rect 59966 -68540 60326 -68520
rect 59966 -68574 60326 -68540
rect 59966 -68580 60326 -68574
rect 59856 -68594 59916 -68580
rect 59856 -68628 59874 -68594
rect 59874 -68628 59908 -68594
rect 59908 -68628 59916 -68594
rect 59856 -68640 59916 -68628
rect 60376 -68594 60436 -68580
rect 60376 -68628 60384 -68594
rect 60384 -68628 60418 -68594
rect 60418 -68628 60436 -68594
rect 60376 -68640 60436 -68628
rect 61056 -68640 61126 -68540
rect 59806 -68920 59916 -68810
rect 60446 -68950 60526 -68830
rect 59646 -69100 59706 -69040
rect 58986 -69560 59126 -69420
rect 59996 -69500 60106 -69390
rect 55500 -70500 56100 -70100
rect 55460 -71360 55720 -71080
rect 53480 -71940 53780 -71740
rect 54150 -71708 54860 -71538
rect 54150 -71778 54850 -71708
rect 54850 -71778 54860 -71708
rect 53520 -72168 53640 -72058
rect 54750 -72108 54850 -72038
rect 54750 -72118 54840 -72108
rect 55430 -72088 55520 -72018
rect 55290 -72198 55390 -72128
rect 53050 -74108 53250 -72358
rect 53950 -72328 53998 -72298
rect 53998 -72328 54020 -72298
rect 53950 -72398 54020 -72328
rect 54920 -72290 54990 -72278
rect 54920 -72328 54926 -72290
rect 54926 -72328 54960 -72290
rect 54960 -72328 54990 -72290
rect 54920 -72368 54990 -72328
rect 53860 -72838 53920 -72728
rect 55230 -72628 55290 -72458
rect 55290 -72628 55320 -72458
rect 55430 -72618 55510 -72448
rect 55960 -72088 56040 -71938
rect 56190 -72168 56390 -71958
rect 56506 -72030 57016 -71780
rect 58966 -71830 59126 -71670
rect 59956 -71860 60166 -71700
rect 55880 -72256 55970 -72218
rect 55880 -72290 55882 -72256
rect 55882 -72290 55970 -72256
rect 55880 -72298 55970 -72290
rect 55000 -72838 55090 -72738
rect 54770 -73040 54840 -73038
rect 54770 -73128 54802 -73040
rect 54802 -73128 54840 -73040
rect 55540 -72838 55630 -72738
rect 56590 -72598 56660 -72468
rect 58906 -72220 58966 -72170
rect 58906 -72230 58926 -72220
rect 58926 -72230 58966 -72220
rect 59216 -72230 59276 -72170
rect 59326 -72230 59386 -72170
rect 59436 -72230 59496 -72170
rect 59636 -72230 59696 -72170
rect 59546 -72301 59606 -72290
rect 59286 -72355 59346 -72330
rect 59546 -72335 59560 -72301
rect 59560 -72335 59594 -72301
rect 59594 -72335 59606 -72301
rect 59286 -72389 59346 -72355
rect 59546 -72350 59606 -72335
rect 59286 -72390 59346 -72389
rect 59016 -72409 59076 -72400
rect 59016 -72443 59032 -72409
rect 59032 -72443 59066 -72409
rect 59066 -72443 59076 -72409
rect 59016 -72460 59076 -72443
rect 59546 -72470 59606 -72410
rect 58906 -72590 58966 -72530
rect 59216 -72580 59276 -72520
rect 59336 -72580 59396 -72520
rect 59436 -72580 59496 -72520
rect 55140 -73208 55200 -73138
rect 55030 -73328 55110 -73248
rect 55740 -73328 55810 -73248
rect 55880 -73328 55970 -73238
rect 56480 -72806 56550 -72788
rect 56480 -72840 56492 -72806
rect 56492 -72840 56530 -72806
rect 56530 -72840 56550 -72806
rect 56480 -72848 56550 -72840
rect 59866 -72430 59966 -72340
rect 60446 -72420 60526 -72320
rect 59636 -72590 59696 -72530
rect 59076 -72678 59166 -72640
rect 59076 -72710 59103 -72678
rect 59103 -72710 59137 -72678
rect 59137 -72710 59166 -72678
rect 60046 -72574 60126 -72540
rect 59856 -72628 59916 -72610
rect 60046 -72600 60126 -72574
rect 59856 -72662 59874 -72628
rect 59874 -72662 59908 -72628
rect 59908 -72662 59916 -72628
rect 59856 -72680 59916 -72662
rect 60376 -72628 60446 -72620
rect 60376 -72662 60384 -72628
rect 60384 -72662 60418 -72628
rect 60418 -72662 60446 -72628
rect 59976 -72716 60316 -72700
rect 60376 -72680 60446 -72662
rect 57098 -72789 57368 -72764
rect 57098 -72823 57125 -72789
rect 57125 -72823 57159 -72789
rect 57159 -72823 57217 -72789
rect 57217 -72823 57251 -72789
rect 57251 -72823 57309 -72789
rect 57309 -72823 57343 -72789
rect 57343 -72823 57368 -72789
rect 54770 -73528 54802 -73448
rect 54802 -73528 54840 -73448
rect 53850 -73848 53920 -73738
rect 54920 -73668 54980 -73598
rect 55000 -73838 55090 -73738
rect 55540 -73838 55630 -73738
rect 55220 -74118 55280 -73948
rect 55280 -74118 55310 -73948
rect 55410 -74128 55500 -73958
rect 53950 -74250 54010 -74208
rect 53950 -74288 53988 -74250
rect 53988 -74288 54010 -74250
rect 54910 -74250 54980 -74198
rect 54910 -74288 54916 -74250
rect 54916 -74288 54950 -74250
rect 54950 -74288 54980 -74250
rect 54910 -74298 54980 -74288
rect 53510 -74448 53630 -74328
rect 54740 -74544 54850 -74468
rect 54740 -74558 54850 -74544
rect 55240 -74418 55370 -74358
rect 55410 -74538 55510 -74448
rect 57098 -72880 57368 -72823
rect 57098 -72904 57368 -72880
rect 56900 -73348 57020 -73218
rect 58576 -73440 58736 -73280
rect 57098 -73680 57368 -73674
rect 56480 -73734 56550 -73728
rect 56480 -73768 56492 -73734
rect 56492 -73768 56530 -73734
rect 56530 -73768 56550 -73734
rect 56480 -73788 56550 -73768
rect 57098 -73765 57368 -73680
rect 57098 -73799 57125 -73765
rect 57125 -73799 57159 -73765
rect 57159 -73799 57217 -73765
rect 57217 -73799 57251 -73765
rect 57251 -73799 57309 -73765
rect 57309 -73799 57343 -73765
rect 57343 -73799 57368 -73765
rect 57098 -73814 57368 -73799
rect 59976 -72752 60316 -72716
rect 59176 -72920 59196 -72840
rect 59196 -72920 59236 -72840
rect 59176 -73120 59196 -73040
rect 59196 -73120 59236 -73040
rect 59076 -73240 59103 -73210
rect 59103 -73240 59137 -73210
rect 59137 -73240 59166 -73210
rect 59076 -73280 59166 -73240
rect 59576 -72898 59636 -72870
rect 59576 -72930 59580 -72898
rect 59580 -72930 59636 -72898
rect 59476 -73120 59502 -73050
rect 59502 -73120 59536 -73050
rect 59576 -73158 59590 -72990
rect 59590 -73158 59624 -72990
rect 59624 -73158 59636 -72990
rect 59576 -73160 59636 -73158
rect 59076 -73408 59166 -73370
rect 59076 -73440 59103 -73408
rect 59103 -73440 59137 -73408
rect 59137 -73440 59166 -73408
rect 59206 -73440 59266 -73370
rect 61206 -72900 61346 -72720
rect 59806 -73140 59818 -73000
rect 59818 -73140 59852 -73000
rect 59852 -73140 59866 -73000
rect 59916 -72982 60006 -72980
rect 59916 -73158 59940 -72982
rect 59940 -73158 60006 -72982
rect 59916 -73160 60006 -73158
rect 60306 -73090 60456 -72950
rect 59826 -73242 59862 -73210
rect 59862 -73242 59896 -73210
rect 59896 -73242 59916 -73210
rect 59826 -73280 59916 -73242
rect 59166 -73610 59196 -73530
rect 59196 -73610 59226 -73530
rect 59166 -73840 59196 -73760
rect 59196 -73840 59226 -73760
rect 59466 -73610 59501 -73530
rect 59501 -73610 59526 -73530
rect 59586 -73650 59589 -73510
rect 59589 -73650 59623 -73510
rect 59623 -73650 59646 -73510
rect 59516 -73721 59596 -73720
rect 59516 -73755 59545 -73721
rect 59545 -73755 59579 -73721
rect 59579 -73755 59596 -73721
rect 59516 -73780 59596 -73755
rect 59826 -73411 59926 -73370
rect 59826 -73440 59861 -73411
rect 59861 -73440 59895 -73411
rect 59895 -73440 59926 -73411
rect 60096 -73283 60127 -73280
rect 60127 -73283 60161 -73280
rect 60161 -73283 60176 -73280
rect 60096 -73341 60176 -73283
rect 60096 -73375 60127 -73341
rect 60127 -73375 60161 -73341
rect 60161 -73375 60176 -73341
rect 60096 -73433 60176 -73375
rect 60096 -73440 60127 -73433
rect 60127 -73440 60161 -73433
rect 60161 -73440 60176 -73433
rect 59796 -73495 59856 -73490
rect 59796 -73670 59817 -73495
rect 59817 -73670 59851 -73495
rect 59851 -73670 59856 -73495
rect 59916 -73495 60006 -73490
rect 59916 -73671 59939 -73495
rect 59939 -73671 60006 -73495
rect 59916 -73680 60006 -73671
rect 60476 -73525 60536 -73510
rect 60476 -73559 60484 -73525
rect 60484 -73559 60536 -73525
rect 60476 -73570 60536 -73559
rect 61036 -73130 61126 -73020
rect 61276 -73283 61291 -73250
rect 61291 -73283 61325 -73250
rect 61325 -73283 61356 -73250
rect 61276 -73341 61356 -73283
rect 61276 -73375 61291 -73341
rect 61291 -73375 61325 -73341
rect 61325 -73375 61356 -73341
rect 61276 -73433 61356 -73375
rect 61276 -73460 61291 -73433
rect 61291 -73460 61325 -73433
rect 61325 -73460 61356 -73433
rect 60476 -73660 60536 -73650
rect 60476 -73700 60486 -73660
rect 60486 -73700 60526 -73660
rect 60526 -73700 60536 -73660
rect 60476 -73710 60536 -73700
rect 60616 -73660 60736 -73650
rect 60616 -73700 60626 -73660
rect 60626 -73700 60666 -73660
rect 60666 -73700 60736 -73660
rect 60616 -73710 60736 -73700
rect 60756 -73660 60816 -73650
rect 60756 -73700 60766 -73660
rect 60766 -73700 60806 -73660
rect 60806 -73700 60816 -73660
rect 60756 -73710 60816 -73700
rect 60896 -73660 60956 -73650
rect 60896 -73700 60906 -73660
rect 60906 -73700 60946 -73660
rect 60946 -73700 60956 -73660
rect 60896 -73710 60956 -73700
rect 56380 -74088 56440 -73968
rect 55880 -74280 55970 -74278
rect 55880 -74314 55882 -74280
rect 55882 -74314 55970 -74280
rect 55880 -74358 55970 -74314
rect 55220 -74728 55330 -74618
rect 55530 -74802 55610 -74778
rect 55530 -74836 55560 -74802
rect 55560 -74836 55610 -74802
rect 55530 -74868 55610 -74836
rect 54140 -74908 54150 -74888
rect 54150 -74908 54840 -74888
rect 54840 -74908 54850 -74888
rect 54140 -75148 54850 -74908
rect 55320 -74948 55470 -74928
rect 55320 -75008 55470 -74948
rect 55320 -75068 55470 -75008
rect 56020 -74608 56080 -74458
rect 56170 -74608 56390 -74408
rect 56654 -74686 56998 -74468
rect 59076 -73970 59103 -73940
rect 59103 -73970 59137 -73940
rect 59137 -73970 59166 -73940
rect 59076 -74000 59166 -73970
rect 58926 -74110 58986 -74060
rect 58926 -74130 58966 -74110
rect 58966 -74130 58986 -74110
rect 59146 -74130 59226 -74060
rect 59276 -74130 59356 -74060
rect 59396 -74130 59476 -74060
rect 59646 -74120 59706 -74060
rect 59546 -74208 59606 -74200
rect 59256 -74262 59366 -74230
rect 59546 -74242 59560 -74208
rect 59560 -74242 59594 -74208
rect 59594 -74242 59606 -74208
rect 59016 -74316 59076 -74300
rect 59256 -74290 59366 -74262
rect 59546 -74260 59606 -74242
rect 59016 -74350 59032 -74316
rect 59032 -74350 59066 -74316
rect 59066 -74350 59076 -74316
rect 59016 -74360 59076 -74350
rect 58906 -74500 58926 -74430
rect 58926 -74500 58966 -74430
rect 58966 -74500 58986 -74430
rect 59146 -74500 59226 -74430
rect 59276 -74500 59356 -74430
rect 59396 -74500 59476 -74430
rect 59966 -73940 60326 -73920
rect 59966 -73974 60326 -73940
rect 59966 -73980 60326 -73974
rect 59856 -73994 59916 -73980
rect 59856 -74028 59874 -73994
rect 59874 -74028 59908 -73994
rect 59908 -74028 59916 -73994
rect 59856 -74040 59916 -74028
rect 60376 -73994 60436 -73980
rect 60376 -74028 60384 -73994
rect 60384 -74028 60418 -73994
rect 60418 -74028 60436 -73994
rect 60376 -74040 60436 -74028
rect 61056 -74040 61126 -73940
rect 59806 -74320 59916 -74210
rect 60446 -74350 60526 -74230
rect 59646 -74500 59706 -74440
rect 58986 -74960 59126 -74820
rect 59996 -74900 60106 -74790
rect 55500 -75900 56100 -75500
rect 55400 -76760 55720 -76480
rect 53480 -77340 53780 -77140
rect 54150 -77108 54860 -76938
rect 54150 -77178 54850 -77108
rect 54850 -77178 54860 -77108
rect 53520 -77568 53640 -77458
rect 54750 -77508 54850 -77438
rect 54750 -77518 54840 -77508
rect 55430 -77488 55520 -77418
rect 55290 -77598 55390 -77528
rect 53050 -79508 53250 -77758
rect 53950 -77728 53998 -77698
rect 53998 -77728 54020 -77698
rect 53950 -77798 54020 -77728
rect 54920 -77690 54990 -77678
rect 54920 -77728 54926 -77690
rect 54926 -77728 54960 -77690
rect 54960 -77728 54990 -77690
rect 54920 -77768 54990 -77728
rect 53860 -78238 53920 -78128
rect 55230 -78028 55290 -77858
rect 55290 -78028 55320 -77858
rect 55430 -78018 55510 -77848
rect 55960 -77488 56040 -77338
rect 56190 -77568 56390 -77358
rect 56506 -77430 57016 -77180
rect 58966 -77230 59126 -77070
rect 59956 -77260 60166 -77100
rect 55880 -77656 55970 -77618
rect 55880 -77690 55882 -77656
rect 55882 -77690 55970 -77656
rect 55880 -77698 55970 -77690
rect 55000 -78238 55090 -78138
rect 54770 -78440 54840 -78438
rect 54770 -78528 54802 -78440
rect 54802 -78528 54840 -78440
rect 55540 -78238 55630 -78138
rect 56590 -77998 56660 -77868
rect 58906 -77620 58966 -77570
rect 58906 -77630 58926 -77620
rect 58926 -77630 58966 -77620
rect 59216 -77630 59276 -77570
rect 59326 -77630 59386 -77570
rect 59436 -77630 59496 -77570
rect 59636 -77630 59696 -77570
rect 59546 -77701 59606 -77690
rect 59286 -77755 59346 -77730
rect 59546 -77735 59560 -77701
rect 59560 -77735 59594 -77701
rect 59594 -77735 59606 -77701
rect 59286 -77789 59346 -77755
rect 59546 -77750 59606 -77735
rect 59286 -77790 59346 -77789
rect 59016 -77809 59076 -77800
rect 59016 -77843 59032 -77809
rect 59032 -77843 59066 -77809
rect 59066 -77843 59076 -77809
rect 59016 -77860 59076 -77843
rect 59546 -77870 59606 -77810
rect 58906 -77990 58966 -77930
rect 59216 -77980 59276 -77920
rect 59336 -77980 59396 -77920
rect 59436 -77980 59496 -77920
rect 55140 -78608 55200 -78538
rect 55030 -78728 55110 -78648
rect 55740 -78728 55810 -78648
rect 55880 -78728 55970 -78638
rect 56480 -78206 56550 -78188
rect 56480 -78240 56492 -78206
rect 56492 -78240 56530 -78206
rect 56530 -78240 56550 -78206
rect 56480 -78248 56550 -78240
rect 59866 -77830 59966 -77740
rect 60446 -77820 60526 -77720
rect 59636 -77990 59696 -77930
rect 59076 -78078 59166 -78040
rect 59076 -78110 59103 -78078
rect 59103 -78110 59137 -78078
rect 59137 -78110 59166 -78078
rect 60046 -77974 60126 -77940
rect 59856 -78028 59916 -78010
rect 60046 -78000 60126 -77974
rect 59856 -78062 59874 -78028
rect 59874 -78062 59908 -78028
rect 59908 -78062 59916 -78028
rect 59856 -78080 59916 -78062
rect 60376 -78028 60446 -78020
rect 60376 -78062 60384 -78028
rect 60384 -78062 60418 -78028
rect 60418 -78062 60446 -78028
rect 59976 -78116 60316 -78100
rect 60376 -78080 60446 -78062
rect 57098 -78189 57368 -78164
rect 57098 -78223 57125 -78189
rect 57125 -78223 57159 -78189
rect 57159 -78223 57217 -78189
rect 57217 -78223 57251 -78189
rect 57251 -78223 57309 -78189
rect 57309 -78223 57343 -78189
rect 57343 -78223 57368 -78189
rect 54770 -78928 54802 -78848
rect 54802 -78928 54840 -78848
rect 53850 -79248 53920 -79138
rect 54920 -79068 54980 -78998
rect 55000 -79238 55090 -79138
rect 55540 -79238 55630 -79138
rect 55220 -79518 55280 -79348
rect 55280 -79518 55310 -79348
rect 55410 -79528 55500 -79358
rect 53950 -79650 54010 -79608
rect 53950 -79688 53988 -79650
rect 53988 -79688 54010 -79650
rect 54910 -79650 54980 -79598
rect 54910 -79688 54916 -79650
rect 54916 -79688 54950 -79650
rect 54950 -79688 54980 -79650
rect 54910 -79698 54980 -79688
rect 53510 -79848 53630 -79728
rect 54740 -79944 54850 -79868
rect 54740 -79958 54850 -79944
rect 55240 -79818 55370 -79758
rect 55410 -79938 55510 -79848
rect 57098 -78280 57368 -78223
rect 57098 -78304 57368 -78280
rect 56900 -78748 57020 -78618
rect 58576 -78840 58736 -78680
rect 57098 -79080 57368 -79074
rect 56480 -79134 56550 -79128
rect 56480 -79168 56492 -79134
rect 56492 -79168 56530 -79134
rect 56530 -79168 56550 -79134
rect 56480 -79188 56550 -79168
rect 57098 -79165 57368 -79080
rect 57098 -79199 57125 -79165
rect 57125 -79199 57159 -79165
rect 57159 -79199 57217 -79165
rect 57217 -79199 57251 -79165
rect 57251 -79199 57309 -79165
rect 57309 -79199 57343 -79165
rect 57343 -79199 57368 -79165
rect 57098 -79214 57368 -79199
rect 59976 -78152 60316 -78116
rect 59176 -78320 59196 -78240
rect 59196 -78320 59236 -78240
rect 59176 -78520 59196 -78440
rect 59196 -78520 59236 -78440
rect 59076 -78640 59103 -78610
rect 59103 -78640 59137 -78610
rect 59137 -78640 59166 -78610
rect 59076 -78680 59166 -78640
rect 59576 -78298 59636 -78270
rect 59576 -78330 59580 -78298
rect 59580 -78330 59636 -78298
rect 59476 -78520 59502 -78450
rect 59502 -78520 59536 -78450
rect 59576 -78558 59590 -78390
rect 59590 -78558 59624 -78390
rect 59624 -78558 59636 -78390
rect 59576 -78560 59636 -78558
rect 59076 -78808 59166 -78770
rect 59076 -78840 59103 -78808
rect 59103 -78840 59137 -78808
rect 59137 -78840 59166 -78808
rect 59206 -78840 59266 -78770
rect 61206 -78300 61346 -78120
rect 59806 -78540 59818 -78400
rect 59818 -78540 59852 -78400
rect 59852 -78540 59866 -78400
rect 59916 -78382 60006 -78380
rect 59916 -78558 59940 -78382
rect 59940 -78558 60006 -78382
rect 59916 -78560 60006 -78558
rect 60306 -78490 60456 -78350
rect 59826 -78642 59862 -78610
rect 59862 -78642 59896 -78610
rect 59896 -78642 59916 -78610
rect 59826 -78680 59916 -78642
rect 59166 -79010 59196 -78930
rect 59196 -79010 59226 -78930
rect 59166 -79240 59196 -79160
rect 59196 -79240 59226 -79160
rect 59466 -79010 59501 -78930
rect 59501 -79010 59526 -78930
rect 59586 -79050 59589 -78910
rect 59589 -79050 59623 -78910
rect 59623 -79050 59646 -78910
rect 59516 -79121 59596 -79120
rect 59516 -79155 59545 -79121
rect 59545 -79155 59579 -79121
rect 59579 -79155 59596 -79121
rect 59516 -79180 59596 -79155
rect 59826 -78811 59926 -78770
rect 59826 -78840 59861 -78811
rect 59861 -78840 59895 -78811
rect 59895 -78840 59926 -78811
rect 60096 -78683 60127 -78680
rect 60127 -78683 60161 -78680
rect 60161 -78683 60176 -78680
rect 60096 -78741 60176 -78683
rect 60096 -78775 60127 -78741
rect 60127 -78775 60161 -78741
rect 60161 -78775 60176 -78741
rect 60096 -78833 60176 -78775
rect 60096 -78840 60127 -78833
rect 60127 -78840 60161 -78833
rect 60161 -78840 60176 -78833
rect 59796 -78895 59856 -78890
rect 59796 -79070 59817 -78895
rect 59817 -79070 59851 -78895
rect 59851 -79070 59856 -78895
rect 59916 -78895 60006 -78890
rect 59916 -79071 59939 -78895
rect 59939 -79071 60006 -78895
rect 59916 -79080 60006 -79071
rect 60476 -78925 60536 -78910
rect 60476 -78959 60484 -78925
rect 60484 -78959 60536 -78925
rect 60476 -78970 60536 -78959
rect 61036 -78530 61126 -78420
rect 61276 -78683 61291 -78650
rect 61291 -78683 61325 -78650
rect 61325 -78683 61356 -78650
rect 61276 -78741 61356 -78683
rect 61276 -78775 61291 -78741
rect 61291 -78775 61325 -78741
rect 61325 -78775 61356 -78741
rect 61276 -78833 61356 -78775
rect 61276 -78860 61291 -78833
rect 61291 -78860 61325 -78833
rect 61325 -78860 61356 -78833
rect 60476 -79060 60536 -79050
rect 60476 -79100 60486 -79060
rect 60486 -79100 60526 -79060
rect 60526 -79100 60536 -79060
rect 60476 -79110 60536 -79100
rect 60616 -79060 60736 -79050
rect 60616 -79100 60626 -79060
rect 60626 -79100 60666 -79060
rect 60666 -79100 60736 -79060
rect 60616 -79110 60736 -79100
rect 60756 -79060 60816 -79050
rect 60756 -79100 60766 -79060
rect 60766 -79100 60806 -79060
rect 60806 -79100 60816 -79060
rect 60756 -79110 60816 -79100
rect 60896 -79060 60956 -79050
rect 60896 -79100 60906 -79060
rect 60906 -79100 60946 -79060
rect 60946 -79100 60956 -79060
rect 60896 -79110 60956 -79100
rect 56380 -79488 56440 -79368
rect 55880 -79680 55970 -79678
rect 55880 -79714 55882 -79680
rect 55882 -79714 55970 -79680
rect 55880 -79758 55970 -79714
rect 55220 -80128 55330 -80018
rect 55530 -80202 55610 -80178
rect 55530 -80236 55560 -80202
rect 55560 -80236 55610 -80202
rect 55530 -80268 55610 -80236
rect 54140 -80308 54150 -80288
rect 54150 -80308 54840 -80288
rect 54840 -80308 54850 -80288
rect 54140 -80548 54850 -80308
rect 55320 -80348 55470 -80328
rect 55320 -80408 55470 -80348
rect 55320 -80468 55470 -80408
rect 56020 -80008 56080 -79858
rect 56170 -80008 56390 -79808
rect 56654 -80086 56998 -79868
rect 59076 -79370 59103 -79340
rect 59103 -79370 59137 -79340
rect 59137 -79370 59166 -79340
rect 59076 -79400 59166 -79370
rect 58926 -79510 58986 -79460
rect 58926 -79530 58966 -79510
rect 58966 -79530 58986 -79510
rect 59146 -79530 59226 -79460
rect 59276 -79530 59356 -79460
rect 59396 -79530 59476 -79460
rect 59646 -79520 59706 -79460
rect 59546 -79608 59606 -79600
rect 59256 -79662 59366 -79630
rect 59546 -79642 59560 -79608
rect 59560 -79642 59594 -79608
rect 59594 -79642 59606 -79608
rect 59016 -79716 59076 -79700
rect 59256 -79690 59366 -79662
rect 59546 -79660 59606 -79642
rect 59016 -79750 59032 -79716
rect 59032 -79750 59066 -79716
rect 59066 -79750 59076 -79716
rect 59016 -79760 59076 -79750
rect 58906 -79900 58926 -79830
rect 58926 -79900 58966 -79830
rect 58966 -79900 58986 -79830
rect 59146 -79900 59226 -79830
rect 59276 -79900 59356 -79830
rect 59396 -79900 59476 -79830
rect 59966 -79340 60326 -79320
rect 59966 -79374 60326 -79340
rect 59966 -79380 60326 -79374
rect 59856 -79394 59916 -79380
rect 59856 -79428 59874 -79394
rect 59874 -79428 59908 -79394
rect 59908 -79428 59916 -79394
rect 59856 -79440 59916 -79428
rect 60376 -79394 60436 -79380
rect 60376 -79428 60384 -79394
rect 60384 -79428 60418 -79394
rect 60418 -79428 60436 -79394
rect 60376 -79440 60436 -79428
rect 61056 -79440 61126 -79340
rect 59806 -79720 59916 -79610
rect 60446 -79750 60526 -79630
rect 59646 -79900 59706 -79840
rect 58986 -80360 59126 -80220
rect 59996 -80300 60106 -80190
rect 55500 -81300 56200 -80900
rect 55440 -82160 55720 -81880
rect 53480 -82740 53780 -82540
rect 54150 -82508 54860 -82338
rect 54150 -82578 54850 -82508
rect 54850 -82578 54860 -82508
rect 53520 -82968 53640 -82858
rect 54750 -82908 54850 -82838
rect 54750 -82918 54840 -82908
rect 55430 -82888 55520 -82818
rect 55290 -82998 55390 -82928
rect 53050 -84908 53250 -83158
rect 53950 -83128 53998 -83098
rect 53998 -83128 54020 -83098
rect 53950 -83198 54020 -83128
rect 54920 -83090 54990 -83078
rect 54920 -83128 54926 -83090
rect 54926 -83128 54960 -83090
rect 54960 -83128 54990 -83090
rect 54920 -83168 54990 -83128
rect 53860 -83638 53920 -83528
rect 55230 -83428 55290 -83258
rect 55290 -83428 55320 -83258
rect 55430 -83418 55510 -83248
rect 55960 -82888 56040 -82738
rect 56190 -82968 56390 -82758
rect 56506 -82830 57016 -82580
rect 58966 -82630 59126 -82470
rect 59956 -82660 60166 -82500
rect 55880 -83056 55970 -83018
rect 55880 -83090 55882 -83056
rect 55882 -83090 55970 -83056
rect 55880 -83098 55970 -83090
rect 55000 -83638 55090 -83538
rect 54770 -83840 54840 -83838
rect 54770 -83928 54802 -83840
rect 54802 -83928 54840 -83840
rect 55540 -83638 55630 -83538
rect 56590 -83398 56660 -83268
rect 58906 -83020 58966 -82970
rect 58906 -83030 58926 -83020
rect 58926 -83030 58966 -83020
rect 59216 -83030 59276 -82970
rect 59326 -83030 59386 -82970
rect 59436 -83030 59496 -82970
rect 59636 -83030 59696 -82970
rect 59546 -83101 59606 -83090
rect 59286 -83155 59346 -83130
rect 59546 -83135 59560 -83101
rect 59560 -83135 59594 -83101
rect 59594 -83135 59606 -83101
rect 59286 -83189 59346 -83155
rect 59546 -83150 59606 -83135
rect 59286 -83190 59346 -83189
rect 59016 -83209 59076 -83200
rect 59016 -83243 59032 -83209
rect 59032 -83243 59066 -83209
rect 59066 -83243 59076 -83209
rect 59016 -83260 59076 -83243
rect 59546 -83270 59606 -83210
rect 58906 -83390 58966 -83330
rect 59216 -83380 59276 -83320
rect 59336 -83380 59396 -83320
rect 59436 -83380 59496 -83320
rect 55140 -84008 55200 -83938
rect 55030 -84128 55110 -84048
rect 55740 -84128 55810 -84048
rect 55880 -84128 55970 -84038
rect 56480 -83606 56550 -83588
rect 56480 -83640 56492 -83606
rect 56492 -83640 56530 -83606
rect 56530 -83640 56550 -83606
rect 56480 -83648 56550 -83640
rect 59866 -83230 59966 -83140
rect 60446 -83220 60526 -83120
rect 59636 -83390 59696 -83330
rect 59076 -83478 59166 -83440
rect 59076 -83510 59103 -83478
rect 59103 -83510 59137 -83478
rect 59137 -83510 59166 -83478
rect 60046 -83374 60126 -83340
rect 59856 -83428 59916 -83410
rect 60046 -83400 60126 -83374
rect 59856 -83462 59874 -83428
rect 59874 -83462 59908 -83428
rect 59908 -83462 59916 -83428
rect 59856 -83480 59916 -83462
rect 60376 -83428 60446 -83420
rect 60376 -83462 60384 -83428
rect 60384 -83462 60418 -83428
rect 60418 -83462 60446 -83428
rect 59976 -83516 60316 -83500
rect 60376 -83480 60446 -83462
rect 57098 -83589 57368 -83564
rect 57098 -83623 57125 -83589
rect 57125 -83623 57159 -83589
rect 57159 -83623 57217 -83589
rect 57217 -83623 57251 -83589
rect 57251 -83623 57309 -83589
rect 57309 -83623 57343 -83589
rect 57343 -83623 57368 -83589
rect 54770 -84328 54802 -84248
rect 54802 -84328 54840 -84248
rect 53850 -84648 53920 -84538
rect 54920 -84468 54980 -84398
rect 55000 -84638 55090 -84538
rect 55540 -84638 55630 -84538
rect 55220 -84918 55280 -84748
rect 55280 -84918 55310 -84748
rect 55410 -84928 55500 -84758
rect 53950 -85050 54010 -85008
rect 53950 -85088 53988 -85050
rect 53988 -85088 54010 -85050
rect 54910 -85050 54980 -84998
rect 54910 -85088 54916 -85050
rect 54916 -85088 54950 -85050
rect 54950 -85088 54980 -85050
rect 54910 -85098 54980 -85088
rect 53510 -85248 53630 -85128
rect 54740 -85344 54850 -85268
rect 54740 -85358 54850 -85344
rect 55240 -85218 55370 -85158
rect 55410 -85338 55510 -85248
rect 57098 -83680 57368 -83623
rect 57098 -83704 57368 -83680
rect 56900 -84148 57020 -84018
rect 58576 -84240 58736 -84080
rect 57098 -84480 57368 -84474
rect 56480 -84534 56550 -84528
rect 56480 -84568 56492 -84534
rect 56492 -84568 56530 -84534
rect 56530 -84568 56550 -84534
rect 56480 -84588 56550 -84568
rect 57098 -84565 57368 -84480
rect 57098 -84599 57125 -84565
rect 57125 -84599 57159 -84565
rect 57159 -84599 57217 -84565
rect 57217 -84599 57251 -84565
rect 57251 -84599 57309 -84565
rect 57309 -84599 57343 -84565
rect 57343 -84599 57368 -84565
rect 57098 -84614 57368 -84599
rect 59976 -83552 60316 -83516
rect 59176 -83720 59196 -83640
rect 59196 -83720 59236 -83640
rect 59176 -83920 59196 -83840
rect 59196 -83920 59236 -83840
rect 59076 -84040 59103 -84010
rect 59103 -84040 59137 -84010
rect 59137 -84040 59166 -84010
rect 59076 -84080 59166 -84040
rect 59576 -83698 59636 -83670
rect 59576 -83730 59580 -83698
rect 59580 -83730 59636 -83698
rect 59476 -83920 59502 -83850
rect 59502 -83920 59536 -83850
rect 59576 -83958 59590 -83790
rect 59590 -83958 59624 -83790
rect 59624 -83958 59636 -83790
rect 59576 -83960 59636 -83958
rect 59076 -84208 59166 -84170
rect 59076 -84240 59103 -84208
rect 59103 -84240 59137 -84208
rect 59137 -84240 59166 -84208
rect 59206 -84240 59266 -84170
rect 61206 -83700 61346 -83520
rect 59806 -83940 59818 -83800
rect 59818 -83940 59852 -83800
rect 59852 -83940 59866 -83800
rect 59916 -83782 60006 -83780
rect 59916 -83958 59940 -83782
rect 59940 -83958 60006 -83782
rect 59916 -83960 60006 -83958
rect 60306 -83890 60456 -83750
rect 59826 -84042 59862 -84010
rect 59862 -84042 59896 -84010
rect 59896 -84042 59916 -84010
rect 59826 -84080 59916 -84042
rect 59166 -84410 59196 -84330
rect 59196 -84410 59226 -84330
rect 59166 -84640 59196 -84560
rect 59196 -84640 59226 -84560
rect 59466 -84410 59501 -84330
rect 59501 -84410 59526 -84330
rect 59586 -84450 59589 -84310
rect 59589 -84450 59623 -84310
rect 59623 -84450 59646 -84310
rect 59516 -84521 59596 -84520
rect 59516 -84555 59545 -84521
rect 59545 -84555 59579 -84521
rect 59579 -84555 59596 -84521
rect 59516 -84580 59596 -84555
rect 59826 -84211 59926 -84170
rect 59826 -84240 59861 -84211
rect 59861 -84240 59895 -84211
rect 59895 -84240 59926 -84211
rect 60096 -84083 60127 -84080
rect 60127 -84083 60161 -84080
rect 60161 -84083 60176 -84080
rect 60096 -84141 60176 -84083
rect 60096 -84175 60127 -84141
rect 60127 -84175 60161 -84141
rect 60161 -84175 60176 -84141
rect 60096 -84233 60176 -84175
rect 60096 -84240 60127 -84233
rect 60127 -84240 60161 -84233
rect 60161 -84240 60176 -84233
rect 59796 -84295 59856 -84290
rect 59796 -84470 59817 -84295
rect 59817 -84470 59851 -84295
rect 59851 -84470 59856 -84295
rect 59916 -84295 60006 -84290
rect 59916 -84471 59939 -84295
rect 59939 -84471 60006 -84295
rect 59916 -84480 60006 -84471
rect 60476 -84325 60536 -84310
rect 60476 -84359 60484 -84325
rect 60484 -84359 60536 -84325
rect 60476 -84370 60536 -84359
rect 61036 -83930 61126 -83820
rect 61276 -84083 61291 -84050
rect 61291 -84083 61325 -84050
rect 61325 -84083 61356 -84050
rect 61276 -84141 61356 -84083
rect 61276 -84175 61291 -84141
rect 61291 -84175 61325 -84141
rect 61325 -84175 61356 -84141
rect 61276 -84233 61356 -84175
rect 61276 -84260 61291 -84233
rect 61291 -84260 61325 -84233
rect 61325 -84260 61356 -84233
rect 60476 -84460 60536 -84450
rect 60476 -84500 60486 -84460
rect 60486 -84500 60526 -84460
rect 60526 -84500 60536 -84460
rect 60476 -84510 60536 -84500
rect 60616 -84460 60736 -84450
rect 60616 -84500 60626 -84460
rect 60626 -84500 60666 -84460
rect 60666 -84500 60736 -84460
rect 60616 -84510 60736 -84500
rect 60756 -84460 60816 -84450
rect 60756 -84500 60766 -84460
rect 60766 -84500 60806 -84460
rect 60806 -84500 60816 -84460
rect 60756 -84510 60816 -84500
rect 60896 -84460 60956 -84450
rect 60896 -84500 60906 -84460
rect 60906 -84500 60946 -84460
rect 60946 -84500 60956 -84460
rect 60896 -84510 60956 -84500
rect 56380 -84888 56440 -84768
rect 55880 -85080 55970 -85078
rect 55880 -85114 55882 -85080
rect 55882 -85114 55970 -85080
rect 55880 -85158 55970 -85114
rect 55220 -85528 55330 -85418
rect 55530 -85602 55610 -85578
rect 55530 -85636 55560 -85602
rect 55560 -85636 55610 -85602
rect 55530 -85668 55610 -85636
rect 54140 -85708 54150 -85688
rect 54150 -85708 54840 -85688
rect 54840 -85708 54850 -85688
rect 54140 -85948 54850 -85708
rect 55320 -85748 55470 -85728
rect 55320 -85808 55470 -85748
rect 55320 -85868 55470 -85808
rect 56020 -85408 56080 -85258
rect 56170 -85408 56390 -85208
rect 56654 -85486 56998 -85268
rect 59076 -84770 59103 -84740
rect 59103 -84770 59137 -84740
rect 59137 -84770 59166 -84740
rect 59076 -84800 59166 -84770
rect 58926 -84910 58986 -84860
rect 58926 -84930 58966 -84910
rect 58966 -84930 58986 -84910
rect 59146 -84930 59226 -84860
rect 59276 -84930 59356 -84860
rect 59396 -84930 59476 -84860
rect 59646 -84920 59706 -84860
rect 59546 -85008 59606 -85000
rect 59256 -85062 59366 -85030
rect 59546 -85042 59560 -85008
rect 59560 -85042 59594 -85008
rect 59594 -85042 59606 -85008
rect 59016 -85116 59076 -85100
rect 59256 -85090 59366 -85062
rect 59546 -85060 59606 -85042
rect 59016 -85150 59032 -85116
rect 59032 -85150 59066 -85116
rect 59066 -85150 59076 -85116
rect 59016 -85160 59076 -85150
rect 58906 -85300 58926 -85230
rect 58926 -85300 58966 -85230
rect 58966 -85300 58986 -85230
rect 59146 -85300 59226 -85230
rect 59276 -85300 59356 -85230
rect 59396 -85300 59476 -85230
rect 59966 -84740 60326 -84720
rect 59966 -84774 60326 -84740
rect 59966 -84780 60326 -84774
rect 59856 -84794 59916 -84780
rect 59856 -84828 59874 -84794
rect 59874 -84828 59908 -84794
rect 59908 -84828 59916 -84794
rect 59856 -84840 59916 -84828
rect 60376 -84794 60436 -84780
rect 60376 -84828 60384 -84794
rect 60384 -84828 60418 -84794
rect 60418 -84828 60436 -84794
rect 60376 -84840 60436 -84828
rect 61056 -84840 61126 -84740
rect 59806 -85120 59916 -85010
rect 60446 -85150 60526 -85030
rect 59646 -85300 59706 -85240
rect 58986 -85760 59126 -85620
rect 59996 -85700 60106 -85590
rect 55500 -86600 56100 -86300
<< metal2 >>
rect 37800 2800 41600 3000
rect 37800 1400 38000 2800
rect 41400 1400 41600 2800
rect 37800 1200 41600 1400
rect 42800 2400 46600 2600
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 800 46600 1000
rect 56880 1020 59080 1030
rect 50800 820 53200 900
rect 42800 0 46600 200
rect 37800 -400 41600 -300
rect 37800 -3600 37900 -400
rect 41500 -3600 41600 -400
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 50800 -20 50900 820
rect 53100 -20 53200 820
rect 50800 -100 53200 -20
rect 56880 -50 59080 -40
rect 51400 -800 52600 -100
rect 51400 -1000 51500 -800
rect 52500 -1000 52600 -800
rect 42800 -1600 46600 -1400
rect 47000 -1300 48100 -1100
rect 37800 -3700 41600 -3600
rect 47000 -1700 47700 -1300
rect 48000 -1700 48100 -1300
rect 36200 -5000 37200 -4800
rect 36200 -5800 36400 -5000
rect 37000 -5800 37200 -5000
rect 47000 -5300 48100 -1700
rect 20800 -6600 22200 -6400
rect 20800 -7400 21000 -6600
rect 22000 -7400 22200 -6600
rect 20800 -7482 22200 -7400
rect 20800 -7600 21390 -7482
rect 21156 -7612 21390 -7600
rect 21620 -7600 22200 -7482
rect 21620 -7612 21856 -7600
rect 21156 -7679 21856 -7612
rect 20804 -7875 20878 -7865
rect 21156 -7969 21306 -7679
rect 21156 -8029 21186 -7969
rect 21276 -8029 21306 -7969
rect 21716 -7969 21856 -7679
rect 21716 -8029 21726 -7969
rect 21186 -11489 21276 -11479
rect 21816 -8029 21856 -7969
rect 22070 -7872 22140 -7862
rect 21726 -11489 21816 -11479
rect 20804 -11639 20878 -11629
rect 24600 -8700 25800 -8600
rect 24600 -9400 24700 -8700
rect 25700 -9400 25800 -8700
rect 24600 -11422 25800 -9400
rect 22140 -11432 25800 -11422
rect 22140 -11632 24730 -11432
rect 25190 -11632 25800 -11432
rect 22070 -11642 25800 -11632
rect 21070 -11702 21910 -11692
rect 20800 -12002 20880 -11992
rect 20250 -12082 20260 -12022
rect 20340 -12082 20800 -12022
rect 20260 -12092 20800 -12082
rect 20800 -12102 20880 -12092
rect 21070 -12182 21910 -11772
rect 24600 -11800 25800 -11642
rect 27000 -10600 34600 -10400
rect 16730 -12222 24910 -12182
rect 25090 -12222 25210 -11800
rect 16730 -12262 24909 -12222
rect 16527 -12329 16586 -12319
rect 16527 -13107 16586 -13106
rect 16526 -13116 16586 -13107
rect 16730 -12330 16789 -12262
rect 16933 -12329 16992 -12319
rect 16933 -13107 16992 -13106
rect 16526 -13162 16585 -13116
rect 16730 -13117 16789 -13107
rect 16932 -13116 16992 -13107
rect 17136 -12330 17195 -12262
rect 17339 -12329 17398 -12319
rect 17339 -13107 17398 -13106
rect 16932 -13162 16991 -13116
rect 17136 -13117 17195 -13107
rect 17338 -13116 17398 -13107
rect 17542 -12330 17601 -12262
rect 17745 -12329 17804 -12319
rect 17745 -13107 17804 -13106
rect 17338 -13162 17397 -13116
rect 17542 -13117 17601 -13107
rect 17744 -13116 17804 -13107
rect 17948 -12330 18007 -12262
rect 18151 -12329 18210 -12319
rect 18151 -13107 18210 -13106
rect 17744 -13162 17803 -13116
rect 17948 -13117 18007 -13107
rect 18150 -13116 18210 -13107
rect 18354 -12330 18413 -12262
rect 18557 -12329 18616 -12319
rect 18557 -13107 18616 -13106
rect 18150 -13162 18209 -13116
rect 18354 -13117 18413 -13107
rect 18556 -13116 18616 -13107
rect 18760 -12330 18819 -12262
rect 18963 -12329 19022 -12319
rect 18963 -13107 19022 -13106
rect 18556 -13162 18615 -13116
rect 18760 -13117 18819 -13107
rect 18962 -13116 19022 -13107
rect 19166 -12330 19225 -12262
rect 19369 -12329 19428 -12319
rect 19369 -13107 19428 -13106
rect 18962 -13162 19021 -13116
rect 19166 -13117 19225 -13107
rect 19368 -13116 19428 -13107
rect 19572 -12330 19631 -12262
rect 19775 -12329 19834 -12319
rect 19775 -13107 19834 -13106
rect 19368 -13162 19427 -13116
rect 19572 -13117 19631 -13107
rect 19774 -13116 19834 -13107
rect 19978 -12330 20037 -12262
rect 20181 -12329 20240 -12319
rect 20181 -13107 20240 -13106
rect 19774 -13162 19833 -13116
rect 19978 -13117 20037 -13107
rect 20180 -13116 20240 -13107
rect 20384 -12330 20443 -12262
rect 20993 -12329 21052 -12319
rect 20580 -12352 20640 -12342
rect 20580 -13052 20640 -13042
rect 20801 -12351 20861 -12341
rect 20801 -13051 20861 -13041
rect 20993 -13107 21052 -13106
rect 20180 -13162 20239 -13116
rect 20384 -13117 20443 -13107
rect 20992 -13116 21052 -13107
rect 21196 -12330 21255 -12262
rect 21399 -12329 21458 -12319
rect 21399 -13107 21458 -13106
rect 20992 -13162 21051 -13116
rect 21196 -13117 21255 -13107
rect 21398 -13116 21458 -13107
rect 21602 -12330 21661 -12262
rect 21805 -12329 21864 -12319
rect 21805 -13107 21864 -13106
rect 21398 -13162 21457 -13116
rect 21602 -13117 21661 -13107
rect 21804 -13116 21864 -13107
rect 22008 -12330 22067 -12262
rect 22211 -12329 22270 -12319
rect 22211 -13107 22270 -13106
rect 21804 -13162 21863 -13116
rect 22008 -13117 22067 -13107
rect 22210 -13116 22270 -13107
rect 22414 -12330 22473 -12262
rect 22617 -12329 22676 -12319
rect 22617 -13107 22676 -13106
rect 22210 -13162 22269 -13116
rect 22414 -13117 22473 -13107
rect 22616 -13116 22676 -13107
rect 22820 -12330 22879 -12262
rect 23023 -12329 23082 -12319
rect 23023 -13107 23082 -13106
rect 22616 -13162 22675 -13116
rect 22820 -13117 22879 -13107
rect 23022 -13116 23082 -13107
rect 23226 -12330 23285 -12262
rect 23429 -12329 23488 -12319
rect 23429 -13107 23488 -13106
rect 23022 -13162 23081 -13116
rect 23226 -13117 23285 -13107
rect 23428 -13116 23488 -13107
rect 23632 -12330 23691 -12262
rect 23835 -12329 23894 -12319
rect 23835 -13107 23894 -13106
rect 23428 -13162 23487 -13116
rect 23632 -13117 23691 -13107
rect 23834 -13116 23894 -13107
rect 24038 -12330 24097 -12262
rect 24241 -12329 24300 -12319
rect 24241 -13107 24300 -13106
rect 23834 -13162 23893 -13116
rect 24038 -13117 24097 -13107
rect 24240 -13116 24300 -13107
rect 24444 -12330 24503 -12262
rect 24647 -12329 24706 -12319
rect 24647 -13107 24706 -13106
rect 24240 -13162 24299 -13116
rect 24444 -13117 24503 -13107
rect 24646 -13116 24706 -13107
rect 24850 -12330 24909 -12262
rect 25090 -12302 25210 -12292
rect 24646 -13162 24705 -13116
rect 24850 -13117 24909 -13107
rect 27000 -13000 27200 -10600
rect 34400 -13000 34600 -10600
rect 16526 -13214 24705 -13162
rect 27000 -13200 34600 -13000
rect 16526 -13254 24706 -13214
rect 16526 -13255 17000 -13254
rect 17338 -13255 17397 -13254
rect 17744 -13255 17803 -13254
rect 18150 -13255 18209 -13254
rect 18556 -13255 18615 -13254
rect 18962 -13255 19021 -13254
rect 19368 -13255 19427 -13254
rect 19774 -13255 19833 -13254
rect 20180 -13255 20239 -13254
rect 20586 -13255 20645 -13254
rect 20992 -13255 21051 -13254
rect 21398 -13255 21457 -13254
rect 21804 -13255 21863 -13254
rect 22210 -13255 22269 -13254
rect 22616 -13255 22675 -13254
rect 23022 -13255 23081 -13254
rect 23428 -13255 23487 -13254
rect 23834 -13255 23893 -13254
rect 24240 -13255 24299 -13254
rect 24646 -13255 24705 -13254
rect 16530 -13312 17000 -13255
rect 16590 -13522 17000 -13312
rect 20570 -13312 20670 -13302
rect 20570 -13402 20670 -13392
rect 16580 -13532 17000 -13522
rect 16990 -14642 17000 -13532
rect 16580 -14652 17000 -14642
rect 16590 -14902 17000 -14652
rect 16580 -14912 17000 -14902
rect 16990 -16022 17000 -14912
rect 16580 -16032 16990 -16022
rect 14400 -26400 20000 -25800
rect 14400 -31200 15000 -26400
rect 19400 -31200 20000 -26400
rect 26000 -26400 35600 -25800
rect 26000 -30400 26600 -26400
rect 35200 -30400 35600 -26400
rect 26000 -31000 35600 -30400
rect 14400 -31800 20000 -31200
rect 36200 -32000 37200 -5800
rect 46400 -6780 48100 -5300
rect 46400 -7200 47640 -6780
rect 48080 -7200 48100 -6780
rect 46400 -8700 48100 -7200
rect 46400 -9400 46700 -8700
rect 47800 -9400 48100 -8700
rect 36000 -32200 37200 -32000
rect 36000 -33000 36200 -32200
rect 36800 -33000 37200 -32200
rect 36000 -33200 37200 -33000
rect 37500 -10700 38200 -10600
rect 37500 -11100 37600 -10700
rect 38100 -11100 38200 -10700
rect 37500 -33600 38200 -11100
rect 46400 -12220 48100 -9400
rect 46400 -12640 47700 -12220
rect 48080 -12640 48100 -12220
rect 35900 -33700 38200 -33600
rect 35900 -34700 36000 -33700
rect 38100 -34700 38200 -33700
rect 35900 -34800 38200 -34700
rect 38400 -16000 39100 -15900
rect 38400 -16600 38500 -16000
rect 39000 -16600 39100 -16000
rect 38400 -35200 39100 -16600
rect 46400 -17620 48100 -12640
rect 46400 -18100 47640 -17620
rect 48080 -18100 48100 -17620
rect 35900 -35300 39100 -35200
rect 35900 -36300 36000 -35300
rect 39000 -36300 39100 -35300
rect 35900 -36400 39100 -36300
rect 39400 -21400 40100 -21300
rect 39400 -22000 39500 -21400
rect 40000 -22000 40100 -21400
rect 39400 -36800 40100 -22000
rect 46400 -23020 48100 -18100
rect 46400 -23440 47680 -23020
rect 48080 -23440 48100 -23020
rect 35900 -36900 40100 -36800
rect 14000 -38000 25000 -37000
rect 35900 -37900 36000 -36900
rect 40000 -37900 40100 -36900
rect 35900 -38000 40100 -37900
rect 40300 -26800 41100 -26700
rect 40300 -27400 40400 -26800
rect 41000 -27400 41100 -26800
rect 14000 -49000 15000 -38000
rect 24000 -49000 25000 -38000
rect 40300 -38400 41100 -27400
rect 46400 -28460 48100 -23440
rect 46400 -28840 47800 -28460
rect 48080 -28840 48100 -28460
rect 35900 -38500 41100 -38400
rect 35900 -39500 36000 -38500
rect 41000 -39500 41100 -38500
rect 35900 -39600 41100 -39500
rect 41400 -32200 42200 -32100
rect 41400 -32800 41500 -32200
rect 42100 -32800 42200 -32200
rect 41400 -40000 42200 -32800
rect 46400 -33860 48100 -28840
rect 46400 -34200 47760 -33860
rect 48080 -34200 48100 -33860
rect 35900 -40100 42200 -40000
rect 35900 -41100 36000 -40100
rect 42100 -41100 42200 -40100
rect 35900 -41200 42200 -41100
rect 42400 -37600 43200 -37500
rect 42400 -38200 42500 -37600
rect 43100 -38200 43200 -37600
rect 42400 -41600 43200 -38200
rect 35900 -41700 43200 -41600
rect 35900 -42700 36000 -41700
rect 43100 -42700 43200 -41700
rect 35900 -42800 43200 -42700
rect 46400 -39220 48100 -34200
rect 46400 -39640 47760 -39220
rect 48080 -39640 48100 -39220
rect 43100 -43100 44400 -43000
rect 43100 -43200 43200 -43100
rect 35900 -43300 43200 -43200
rect 35900 -44300 36000 -43300
rect 44300 -44300 44400 -43100
rect 35900 -44400 44400 -44300
rect 46400 -44640 48100 -39640
rect 35900 -44900 44400 -44800
rect 35900 -45900 36000 -44900
rect 44300 -45900 44400 -44900
rect 35900 -46000 44400 -45900
rect 35900 -46500 43500 -46400
rect 35900 -47500 36000 -46500
rect 43400 -47500 43500 -46500
rect 35900 -47600 43500 -47500
rect 14000 -50000 25000 -49000
rect 35900 -48100 42600 -48000
rect 35900 -49100 36000 -48100
rect 42500 -49100 42600 -48100
rect 35900 -49200 42600 -49100
rect 35900 -49700 41700 -49600
rect 35900 -50700 36000 -49700
rect 41600 -50700 41700 -49700
rect 35900 -50800 41700 -50700
rect 35900 -51300 40800 -51200
rect 35900 -52300 36000 -51300
rect 40700 -52300 40800 -51300
rect 35900 -52400 40800 -52300
rect 35900 -52900 39900 -52800
rect 35900 -53900 36000 -52900
rect 39800 -53900 39900 -52900
rect 35900 -54000 39900 -53900
rect 35900 -54500 38900 -54400
rect 35900 -55500 36000 -54500
rect 38800 -55500 38900 -54500
rect 35900 -55600 38900 -55500
rect 35900 -56100 37800 -56000
rect 35900 -57100 36000 -56100
rect 37700 -57100 37800 -56100
rect 35900 -57200 37800 -57100
rect 24400 -58800 36000 -58200
rect 14600 -60000 20200 -59400
rect 14600 -64800 15200 -60000
rect 19600 -64800 20200 -60000
rect 14600 -65400 20200 -64800
rect 24400 -64800 25000 -58800
rect 35400 -64800 36000 -58800
rect 24400 -65400 36000 -64800
rect 37100 -86200 37800 -57200
rect 38200 -80800 38900 -55600
rect 39200 -75400 39900 -54000
rect 40100 -70000 40800 -52400
rect 41000 -64600 41700 -50800
rect 41900 -59200 42600 -49200
rect 42800 -53800 43500 -47600
rect 43700 -48400 44400 -46000
rect 43700 -49000 43800 -48400
rect 44300 -49000 44400 -48400
rect 43700 -49100 44400 -49000
rect 46400 -45060 47820 -44640
rect 48080 -45060 48100 -44640
rect 42800 -54400 42900 -53800
rect 43400 -54400 43500 -53800
rect 42800 -54500 43500 -54400
rect 46400 -49980 48100 -45060
rect 46400 -50480 47740 -49980
rect 48080 -50480 48100 -49980
rect 41900 -59800 42000 -59200
rect 42500 -59800 42600 -59200
rect 41900 -59900 42600 -59800
rect 46400 -55460 48100 -50480
rect 46400 -55820 47820 -55460
rect 48080 -55820 48100 -55460
rect 41000 -65200 41100 -64600
rect 41600 -65200 41700 -64600
rect 41000 -65300 41700 -65200
rect 46400 -60760 48100 -55820
rect 46400 -61300 47680 -60760
rect 48080 -61300 48100 -60760
rect 40100 -70600 40200 -70000
rect 40700 -70600 40800 -70000
rect 40100 -70700 40800 -70600
rect 46400 -66220 48100 -61300
rect 46400 -66660 47860 -66220
rect 48080 -66660 48100 -66220
rect 39200 -76000 39300 -75400
rect 39800 -76000 39900 -75400
rect 39200 -76100 39900 -76000
rect 46400 -71600 48100 -66660
rect 46400 -72060 47720 -71600
rect 48080 -72060 48100 -71600
rect 38200 -81400 38300 -80800
rect 38800 -81400 38900 -80800
rect 38200 -81500 38900 -81400
rect 46400 -76940 48100 -72060
rect 46400 -77500 47780 -76940
rect 48080 -77500 48100 -76940
rect 46400 -82380 48100 -77500
rect 46400 -82860 47800 -82380
rect 48080 -82860 48100 -82380
rect 46400 -82960 48100 -82860
rect 51400 -6300 52600 -1000
rect 55300 -600 55800 -500
rect 55300 -1000 55400 -600
rect 55700 -1000 55800 -600
rect 55300 -1100 55800 -1000
rect 53300 -1400 53800 -1300
rect 53300 -1600 53400 -1400
rect 53700 -1600 53800 -1400
rect 54140 -1338 56390 -1328
rect 54140 -1578 54150 -1338
rect 54860 -1578 56390 -1338
rect 58946 -1470 59146 -1450
rect 54140 -1588 56390 -1578
rect 53300 -1700 53800 -1600
rect 54850 -1818 55530 -1808
rect 53510 -1968 53520 -1858
rect 53640 -1968 53650 -1858
rect 54740 -1918 54750 -1838
rect 54850 -1888 55430 -1818
rect 55520 -1888 55530 -1818
rect 55950 -1888 55960 -1738
rect 56040 -1888 56050 -1738
rect 56170 -1758 56390 -1588
rect 56506 -1580 57016 -1570
rect 54840 -1918 54850 -1908
rect 55270 -2008 55280 -1918
rect 55400 -2008 55410 -1918
rect 56170 -1968 56190 -1758
rect 56390 -1968 56400 -1758
rect 58946 -1630 58966 -1470
rect 59126 -1630 59146 -1470
rect 58946 -1650 59146 -1630
rect 59316 -1500 60176 -1490
rect 59316 -1510 59956 -1500
rect 59316 -1650 59336 -1510
rect 59416 -1650 59956 -1510
rect 59316 -1660 59956 -1650
rect 60166 -1660 60176 -1500
rect 59316 -1670 60176 -1660
rect 56506 -1840 57016 -1830
rect 58956 -1720 61136 -1710
rect 58956 -1730 61056 -1720
rect 58956 -1840 58996 -1730
rect 59106 -1740 61056 -1730
rect 59106 -1840 59516 -1740
rect 59616 -1840 61056 -1740
rect 58396 -1930 58896 -1840
rect 58956 -1850 61056 -1840
rect 61126 -1850 61136 -1720
rect 58956 -1860 61136 -1850
rect 55850 -2048 55880 -2018
rect 53940 -2078 55880 -2048
rect 53940 -2098 54920 -2078
rect 53040 -3908 53050 -2158
rect 53250 -3908 53260 -2158
rect 53940 -2198 53950 -2098
rect 54020 -2148 54920 -2098
rect 54020 -2198 54030 -2148
rect 54910 -2168 54920 -2148
rect 54990 -2098 55880 -2078
rect 55970 -2048 55980 -2018
rect 54990 -2148 55970 -2098
rect 54990 -2168 55000 -2148
rect 55220 -2428 55230 -2258
rect 55320 -2428 55330 -2258
rect 55420 -2418 55430 -2248
rect 55510 -2258 55520 -2248
rect 55510 -2268 56670 -2258
rect 55510 -2398 55600 -2268
rect 55710 -2398 56590 -2268
rect 56660 -2398 56670 -2268
rect 55510 -2408 56670 -2398
rect 58396 -2290 58486 -1930
rect 58816 -1950 58896 -1930
rect 59646 -1950 59706 -1930
rect 58816 -1970 59706 -1950
rect 58816 -2030 58906 -1970
rect 58966 -2030 59216 -1970
rect 59276 -2030 59326 -1970
rect 59386 -2030 59436 -1970
rect 59496 -2030 59636 -1970
rect 59696 -2030 59706 -1970
rect 58816 -2040 59706 -2030
rect 58816 -2290 58896 -2040
rect 59536 -2090 59616 -2080
rect 59276 -2130 59356 -2120
rect 59276 -2190 59286 -2130
rect 59346 -2190 59356 -2130
rect 59536 -2150 59546 -2090
rect 59606 -2150 59616 -2090
rect 59536 -2170 59616 -2150
rect 58996 -2200 59076 -2190
rect 58996 -2260 59006 -2200
rect 59076 -2220 59086 -2200
rect 59536 -2210 59616 -2200
rect 59536 -2220 59546 -2210
rect 59076 -2260 59546 -2220
rect 58996 -2270 59076 -2260
rect 59536 -2270 59546 -2260
rect 59606 -2270 59616 -2210
rect 59536 -2280 59616 -2270
rect 58396 -2310 58896 -2290
rect 59646 -2310 59706 -2040
rect 60436 -2120 60536 -2110
rect 59856 -2140 59976 -2130
rect 59856 -2230 59866 -2140
rect 59966 -2230 59976 -2140
rect 60436 -2220 60446 -2120
rect 60526 -2220 60536 -2120
rect 60436 -2230 60536 -2220
rect 59856 -2240 59976 -2230
rect 58396 -2320 59706 -2310
rect 58396 -2330 59216 -2320
rect 58396 -2390 58906 -2330
rect 58966 -2380 59216 -2330
rect 59276 -2380 59336 -2320
rect 59396 -2380 59436 -2320
rect 59496 -2330 59706 -2320
rect 59496 -2380 59636 -2330
rect 58966 -2390 59636 -2380
rect 59696 -2390 59706 -2330
rect 58396 -2400 59706 -2390
rect 60036 -2320 60136 -2310
rect 60036 -2400 60046 -2320
rect 60126 -2400 60136 -2320
rect 55510 -2418 55520 -2408
rect 59646 -2410 59706 -2400
rect 60546 -2410 60636 -2400
rect 59066 -2440 59176 -2430
rect 59066 -2510 59076 -2440
rect 59166 -2510 59176 -2440
rect 59846 -2480 59856 -2410
rect 59916 -2430 59926 -2410
rect 60356 -2420 60556 -2410
rect 60356 -2430 60376 -2420
rect 59916 -2460 60376 -2430
rect 59916 -2480 59926 -2460
rect 60356 -2480 60376 -2460
rect 60446 -2480 60556 -2420
rect 60356 -2490 60556 -2480
rect 60626 -2490 60636 -2410
rect 59066 -2520 59176 -2510
rect 59966 -2500 60326 -2490
rect 53850 -2638 53860 -2528
rect 53920 -2538 55600 -2528
rect 53920 -2638 55000 -2538
rect 55090 -2638 55540 -2538
rect 55630 -2638 55640 -2538
rect 59966 -2560 59976 -2500
rect 60316 -2560 60326 -2500
rect 60546 -2510 60636 -2490
rect 61186 -2520 61366 -2510
rect 54770 -2838 54850 -2638
rect 56470 -2648 56480 -2588
rect 56550 -2648 56560 -2588
rect 57088 -2704 57098 -2564
rect 57368 -2704 57378 -2564
rect 59166 -2630 59376 -2620
rect 59166 -2640 59286 -2630
rect 59166 -2720 59176 -2640
rect 59236 -2720 59286 -2640
rect 59366 -2720 59376 -2630
rect 59166 -2730 59376 -2720
rect 59526 -2670 59646 -2650
rect 59526 -2730 59576 -2670
rect 59636 -2730 59646 -2670
rect 61186 -2700 61206 -2520
rect 61346 -2700 61366 -2520
rect 61186 -2710 61366 -2700
rect 59526 -2760 59646 -2730
rect 60286 -2750 60476 -2740
rect 59906 -2780 60016 -2770
rect 59806 -2790 59866 -2780
rect 54760 -2928 54770 -2838
rect 54840 -2928 54850 -2838
rect 59166 -2840 59536 -2830
rect 59166 -2920 59176 -2840
rect 59236 -2920 59286 -2840
rect 54920 -2938 55210 -2928
rect 54920 -3008 55140 -2938
rect 55200 -3008 55210 -2938
rect 59166 -2930 59286 -2920
rect 59356 -2850 59536 -2840
rect 59356 -2920 59476 -2850
rect 59356 -2930 59536 -2920
rect 59166 -2940 59536 -2930
rect 59566 -2960 59576 -2790
rect 59636 -2800 59866 -2790
rect 59636 -2940 59806 -2800
rect 59636 -2960 59866 -2940
rect 59906 -2960 59916 -2780
rect 60006 -2960 60016 -2780
rect 60286 -2890 60306 -2750
rect 60456 -2890 60476 -2750
rect 60286 -2900 60476 -2890
rect 61026 -2820 61136 -2810
rect 61026 -2930 61036 -2820
rect 61126 -2930 61136 -2820
rect 61026 -2940 61136 -2930
rect 59566 -2970 59636 -2960
rect 59906 -2970 60016 -2960
rect 54760 -3328 54770 -3248
rect 54840 -3328 54850 -3248
rect 54770 -3538 54850 -3328
rect 54920 -3398 54980 -3008
rect 55880 -3038 56900 -3018
rect 55010 -3128 55020 -3048
rect 55120 -3128 55740 -3048
rect 55810 -3128 55820 -3048
rect 55870 -3128 55880 -3038
rect 55970 -3128 56480 -3038
rect 56550 -3128 56900 -3038
rect 55880 -3148 56900 -3128
rect 57020 -3020 57040 -3018
rect 57800 -3020 58240 -3010
rect 57020 -3140 57800 -3020
rect 57020 -3148 57040 -3140
rect 57800 -3150 58240 -3140
rect 58516 -3060 58796 -2990
rect 58516 -3260 58556 -3060
rect 58756 -3260 58796 -3060
rect 59066 -3010 59936 -3000
rect 59066 -3080 59076 -3010
rect 59166 -3030 59826 -3010
rect 59166 -3080 59316 -3030
rect 59066 -3090 59316 -3080
rect 59376 -3080 59826 -3030
rect 59916 -3080 59936 -3010
rect 59376 -3090 59936 -3080
rect 60076 -3080 60196 -3040
rect 59066 -3170 59936 -3160
rect 59066 -3240 59076 -3170
rect 59166 -3240 59206 -3170
rect 59266 -3240 59826 -3170
rect 59926 -3240 59936 -3170
rect 59066 -3250 59936 -3240
rect 60076 -3240 60096 -3080
rect 60176 -3240 60196 -3080
rect 58516 -3340 58796 -3260
rect 60076 -3280 60196 -3240
rect 61266 -3050 61366 -3040
rect 61266 -3260 61276 -3050
rect 61356 -3260 61366 -3050
rect 61266 -3270 61366 -3260
rect 59586 -3290 59656 -3280
rect 59796 -3290 59866 -3280
rect 59586 -3310 59796 -3290
rect 59156 -3320 59536 -3310
rect 59156 -3330 59266 -3320
rect 54910 -3468 54920 -3398
rect 54980 -3468 54990 -3398
rect 59156 -3410 59166 -3330
rect 59226 -3410 59266 -3330
rect 59366 -3330 59536 -3320
rect 59366 -3410 59466 -3330
rect 59526 -3410 59536 -3330
rect 59156 -3430 59536 -3410
rect 59646 -3450 59796 -3310
rect 59586 -3470 59796 -3450
rect 59856 -3470 59866 -3290
rect 53840 -3648 53850 -3538
rect 53920 -3638 55000 -3538
rect 55090 -3638 55540 -3538
rect 55630 -3638 55640 -3538
rect 56470 -3588 56480 -3528
rect 56550 -3588 56560 -3528
rect 57088 -3614 57098 -3474
rect 57368 -3614 57378 -3474
rect 59796 -3480 59866 -3470
rect 59906 -3290 60016 -3280
rect 59906 -3480 59916 -3290
rect 60006 -3480 60016 -3290
rect 60476 -3310 60546 -3300
rect 60536 -3370 60546 -3310
rect 60476 -3380 60546 -3370
rect 60966 -3430 61486 -3420
rect 60966 -3440 61336 -3430
rect 59906 -3490 60016 -3480
rect 60466 -3450 61336 -3440
rect 59506 -3510 59606 -3500
rect 59156 -3560 59376 -3540
rect 53920 -3648 55640 -3638
rect 59156 -3640 59166 -3560
rect 59226 -3640 59266 -3560
rect 59156 -3650 59266 -3640
rect 59366 -3650 59376 -3560
rect 59506 -3580 59516 -3510
rect 59596 -3580 59606 -3510
rect 60466 -3510 60476 -3450
rect 60536 -3510 60616 -3450
rect 60736 -3510 60756 -3450
rect 60816 -3510 60896 -3450
rect 60956 -3510 61336 -3450
rect 60466 -3520 61336 -3510
rect 60966 -3560 61336 -3520
rect 61456 -3560 61486 -3430
rect 60966 -3570 61486 -3560
rect 59506 -3590 59606 -3580
rect 59156 -3660 59376 -3650
rect 59306 -3720 60336 -3700
rect 59066 -3740 59176 -3730
rect 55210 -3918 55220 -3748
rect 55310 -3918 55320 -3748
rect 55400 -3928 55410 -3758
rect 55500 -3768 55510 -3758
rect 55500 -3888 56380 -3768
rect 56440 -3888 56450 -3768
rect 59066 -3800 59076 -3740
rect 59166 -3800 59176 -3740
rect 59306 -3780 59316 -3720
rect 59376 -3740 59966 -3720
rect 59376 -3780 59816 -3740
rect 59306 -3790 59816 -3780
rect 59846 -3780 59916 -3770
rect 59066 -3810 59176 -3800
rect 59846 -3840 59856 -3780
rect 59946 -3780 59966 -3740
rect 60326 -3780 60336 -3720
rect 59946 -3790 60336 -3780
rect 60366 -3740 61146 -3730
rect 60366 -3780 61056 -3740
rect 59646 -3850 59716 -3840
rect 59846 -3850 59916 -3840
rect 60366 -3840 60376 -3780
rect 60436 -3840 61056 -3780
rect 61126 -3840 61146 -3740
rect 55500 -3908 56450 -3888
rect 58396 -3860 59716 -3850
rect 55500 -3928 55510 -3908
rect 58396 -3930 58926 -3860
rect 58986 -3930 59146 -3860
rect 59226 -3930 59276 -3860
rect 59356 -3930 59396 -3860
rect 59476 -3920 59646 -3860
rect 59706 -3920 59716 -3860
rect 60366 -3870 61146 -3840
rect 59476 -3930 59716 -3920
rect 58396 -3940 59716 -3930
rect 54900 -4008 54910 -3998
rect 53940 -4088 53950 -4008
rect 54010 -4088 54910 -4008
rect 53940 -4098 54910 -4088
rect 54980 -4018 54990 -3998
rect 54980 -4078 55980 -4018
rect 54980 -4098 55880 -4078
rect 53940 -4118 55880 -4098
rect 53500 -4248 53510 -4128
rect 53630 -4248 53640 -4128
rect 55850 -4158 55880 -4118
rect 55970 -4158 55980 -4078
rect 55230 -4218 55240 -4158
rect 55370 -4178 55710 -4158
rect 55370 -4188 55720 -4178
rect 55370 -4208 55620 -4188
rect 55370 -4218 55380 -4208
rect 55400 -4268 55410 -4248
rect 54730 -4358 54740 -4268
rect 54850 -4338 55410 -4268
rect 55510 -4338 55520 -4248
rect 55600 -4278 55620 -4208
rect 55710 -4278 55720 -4188
rect 54850 -4358 55520 -4338
rect 55210 -4528 55220 -4418
rect 55330 -4528 55340 -4418
rect 55850 -4578 55980 -4158
rect 56010 -4408 56020 -4258
rect 56080 -4408 56090 -4258
rect 56160 -4408 56170 -4208
rect 56390 -4408 56400 -4208
rect 58396 -4220 58896 -3940
rect 59006 -4100 59076 -4080
rect 59246 -4090 59256 -4030
rect 59366 -4090 59376 -4030
rect 59536 -4060 59546 -3990
rect 59606 -4060 59616 -3990
rect 59536 -4070 59616 -4060
rect 59006 -4160 59016 -4100
rect 59536 -4110 59616 -4100
rect 59076 -4120 59086 -4110
rect 59536 -4120 59546 -4110
rect 59076 -4160 59546 -4120
rect 59006 -4170 59546 -4160
rect 59606 -4170 59616 -4110
rect 59006 -4190 59076 -4170
rect 59536 -4190 59616 -4170
rect 59646 -4220 59716 -3940
rect 59796 -4010 59926 -4000
rect 59796 -4120 59806 -4010
rect 59916 -4120 59926 -4010
rect 59796 -4130 59926 -4120
rect 60436 -4030 60536 -4010
rect 60436 -4150 60446 -4030
rect 60526 -4150 60536 -4030
rect 60436 -4160 60536 -4150
rect 58396 -4230 59716 -4220
rect 56654 -4268 56998 -4258
rect 55520 -4668 55530 -4578
rect 55610 -4668 55980 -4578
rect 54130 -4948 54140 -4688
rect 54850 -4948 54860 -4688
rect 55310 -4868 55320 -4728
rect 55470 -4868 55480 -4728
rect 56170 -4938 56390 -4408
rect 58396 -4300 58906 -4230
rect 58986 -4300 59146 -4230
rect 59226 -4300 59276 -4230
rect 59356 -4300 59396 -4230
rect 59476 -4240 59716 -4230
rect 59476 -4300 59646 -4240
rect 59706 -4300 59716 -4240
rect 58396 -4310 59716 -4300
rect 58396 -4350 58896 -4310
rect 59646 -4320 59716 -4310
rect 56654 -4496 56998 -4486
rect 59006 -4400 60416 -4390
rect 59006 -4440 60266 -4400
rect 59006 -4510 59016 -4440
rect 59076 -4510 59546 -4440
rect 59606 -4510 60266 -4440
rect 59006 -4530 60266 -4510
rect 60406 -4530 60416 -4400
rect 59006 -4540 60416 -4530
rect 59986 -4590 60116 -4580
rect 58956 -4600 59156 -4590
rect 58956 -4780 58966 -4600
rect 59146 -4780 59156 -4600
rect 59986 -4700 59996 -4590
rect 60106 -4700 60116 -4590
rect 59986 -4710 60116 -4700
rect 58956 -4790 59156 -4780
rect 55680 -4948 56390 -4938
rect 54130 -5108 56390 -4948
rect 55680 -5118 56390 -5108
rect 59600 -4900 60500 -4800
rect 59600 -5200 59700 -4900
rect 60400 -5200 60500 -4900
rect 55500 -5300 56000 -5200
rect 59600 -5300 60500 -5200
rect 68000 -4900 68700 -4800
rect 68000 -5200 68100 -4900
rect 68600 -5200 68700 -4900
rect 55500 -5600 55600 -5300
rect 55900 -5600 56000 -5300
rect 55500 -5700 56000 -5600
rect 51400 -6500 51500 -6300
rect 52500 -6500 52600 -6300
rect 51400 -11700 52600 -6500
rect 55300 -6200 55800 -6100
rect 55300 -6500 55400 -6200
rect 55700 -6500 55800 -6200
rect 55300 -6600 55800 -6500
rect 54140 -6738 56390 -6728
rect 53500 -6860 53800 -6840
rect 53500 -7120 53520 -6860
rect 53780 -7120 53800 -6860
rect 54140 -6978 54150 -6738
rect 54860 -6978 56390 -6738
rect 58946 -6870 59146 -6850
rect 54140 -6988 56390 -6978
rect 53500 -7140 53800 -7120
rect 54850 -7218 55530 -7208
rect 53510 -7368 53520 -7258
rect 53640 -7368 53650 -7258
rect 54740 -7318 54750 -7238
rect 54850 -7288 55430 -7218
rect 55520 -7288 55530 -7218
rect 55950 -7288 55960 -7138
rect 56040 -7288 56050 -7138
rect 56170 -7158 56390 -6988
rect 56506 -6980 57016 -6970
rect 54840 -7318 54850 -7308
rect 55270 -7408 55280 -7318
rect 55400 -7408 55410 -7318
rect 56170 -7368 56190 -7158
rect 56390 -7368 56400 -7158
rect 58946 -7030 58966 -6870
rect 59126 -7030 59146 -6870
rect 58946 -7050 59146 -7030
rect 59316 -6900 60176 -6890
rect 59316 -6910 59956 -6900
rect 59316 -7050 59336 -6910
rect 59416 -7050 59956 -6910
rect 59316 -7060 59956 -7050
rect 60166 -7060 60176 -6900
rect 59316 -7070 60176 -7060
rect 56506 -7240 57016 -7230
rect 58956 -7120 61136 -7110
rect 58956 -7130 61056 -7120
rect 58956 -7240 58996 -7130
rect 59106 -7140 61056 -7130
rect 59106 -7240 59516 -7140
rect 59616 -7240 61056 -7140
rect 58396 -7330 58896 -7240
rect 58956 -7250 61056 -7240
rect 61126 -7250 61136 -7120
rect 58956 -7260 61136 -7250
rect 55850 -7448 55880 -7418
rect 53940 -7478 55880 -7448
rect 53940 -7498 54920 -7478
rect 53040 -9308 53050 -7558
rect 53250 -9308 53260 -7558
rect 53940 -7598 53950 -7498
rect 54020 -7548 54920 -7498
rect 54020 -7598 54030 -7548
rect 54910 -7568 54920 -7548
rect 54990 -7498 55880 -7478
rect 55970 -7448 55980 -7418
rect 54990 -7548 55970 -7498
rect 54990 -7568 55000 -7548
rect 55220 -7828 55230 -7658
rect 55320 -7828 55330 -7658
rect 55420 -7818 55430 -7648
rect 55510 -7658 55520 -7648
rect 55510 -7668 56670 -7658
rect 55510 -7798 55600 -7668
rect 55710 -7798 56590 -7668
rect 56660 -7798 56670 -7668
rect 55510 -7808 56670 -7798
rect 58396 -7690 58486 -7330
rect 58816 -7350 58896 -7330
rect 59646 -7350 59706 -7330
rect 58816 -7370 59706 -7350
rect 58816 -7430 58906 -7370
rect 58966 -7430 59216 -7370
rect 59276 -7430 59326 -7370
rect 59386 -7430 59436 -7370
rect 59496 -7430 59636 -7370
rect 59696 -7430 59706 -7370
rect 58816 -7440 59706 -7430
rect 58816 -7690 58896 -7440
rect 59536 -7490 59616 -7480
rect 59276 -7530 59356 -7520
rect 59276 -7590 59286 -7530
rect 59346 -7590 59356 -7530
rect 59536 -7550 59546 -7490
rect 59606 -7550 59616 -7490
rect 59536 -7570 59616 -7550
rect 58996 -7600 59076 -7590
rect 58996 -7660 59006 -7600
rect 59076 -7620 59086 -7600
rect 59536 -7610 59616 -7600
rect 59536 -7620 59546 -7610
rect 59076 -7660 59546 -7620
rect 58996 -7670 59076 -7660
rect 59536 -7670 59546 -7660
rect 59606 -7670 59616 -7610
rect 59536 -7680 59616 -7670
rect 58396 -7710 58896 -7690
rect 59646 -7710 59706 -7440
rect 60436 -7520 60536 -7510
rect 59856 -7540 59976 -7530
rect 59856 -7630 59866 -7540
rect 59966 -7630 59976 -7540
rect 60436 -7620 60446 -7520
rect 60526 -7620 60536 -7520
rect 60436 -7630 60536 -7620
rect 59856 -7640 59976 -7630
rect 58396 -7720 59706 -7710
rect 58396 -7730 59216 -7720
rect 58396 -7790 58906 -7730
rect 58966 -7780 59216 -7730
rect 59276 -7780 59336 -7720
rect 59396 -7780 59436 -7720
rect 59496 -7730 59706 -7720
rect 59496 -7780 59636 -7730
rect 58966 -7790 59636 -7780
rect 59696 -7790 59706 -7730
rect 58396 -7800 59706 -7790
rect 60036 -7720 60136 -7710
rect 60036 -7800 60046 -7720
rect 60126 -7800 60136 -7720
rect 55510 -7818 55520 -7808
rect 59646 -7810 59706 -7800
rect 60546 -7810 60636 -7800
rect 59066 -7840 59176 -7830
rect 59066 -7910 59076 -7840
rect 59166 -7910 59176 -7840
rect 59846 -7880 59856 -7810
rect 59916 -7830 59926 -7810
rect 60356 -7820 60556 -7810
rect 60356 -7830 60376 -7820
rect 59916 -7860 60376 -7830
rect 59916 -7880 59926 -7860
rect 60356 -7880 60376 -7860
rect 60446 -7880 60556 -7820
rect 60356 -7890 60556 -7880
rect 60626 -7890 60636 -7810
rect 59066 -7920 59176 -7910
rect 59966 -7900 60326 -7890
rect 53850 -8038 53860 -7928
rect 53920 -7938 55600 -7928
rect 53920 -8038 55000 -7938
rect 55090 -8038 55540 -7938
rect 55630 -8038 55640 -7938
rect 59966 -7960 59976 -7900
rect 60316 -7960 60326 -7900
rect 60546 -7910 60636 -7890
rect 61186 -7920 61366 -7910
rect 54770 -8238 54850 -8038
rect 56470 -8048 56480 -7988
rect 56550 -8048 56560 -7988
rect 57088 -8104 57098 -7964
rect 57368 -8104 57378 -7964
rect 59166 -8030 59376 -8020
rect 59166 -8040 59286 -8030
rect 59166 -8120 59176 -8040
rect 59236 -8120 59286 -8040
rect 59366 -8120 59376 -8030
rect 59166 -8130 59376 -8120
rect 59526 -8070 59646 -8050
rect 59526 -8130 59576 -8070
rect 59636 -8130 59646 -8070
rect 61186 -8100 61206 -7920
rect 61346 -8100 61366 -7920
rect 61186 -8110 61366 -8100
rect 59526 -8160 59646 -8130
rect 60286 -8150 60476 -8140
rect 59906 -8180 60016 -8170
rect 59806 -8190 59866 -8180
rect 54760 -8328 54770 -8238
rect 54840 -8328 54850 -8238
rect 59166 -8240 59536 -8230
rect 59166 -8320 59176 -8240
rect 59236 -8320 59286 -8240
rect 54920 -8338 55210 -8328
rect 54920 -8408 55140 -8338
rect 55200 -8408 55210 -8338
rect 59166 -8330 59286 -8320
rect 59356 -8250 59536 -8240
rect 59356 -8320 59476 -8250
rect 59356 -8330 59536 -8320
rect 59166 -8340 59536 -8330
rect 59566 -8360 59576 -8190
rect 59636 -8200 59866 -8190
rect 59636 -8340 59806 -8200
rect 59636 -8360 59866 -8340
rect 59906 -8360 59916 -8180
rect 60006 -8360 60016 -8180
rect 60286 -8290 60306 -8150
rect 60456 -8290 60476 -8150
rect 60286 -8300 60476 -8290
rect 61026 -8220 61136 -8210
rect 61026 -8330 61036 -8220
rect 61126 -8330 61136 -8220
rect 61026 -8340 61136 -8330
rect 59566 -8370 59636 -8360
rect 59906 -8370 60016 -8360
rect 54760 -8728 54770 -8648
rect 54840 -8728 54850 -8648
rect 54770 -8938 54850 -8728
rect 54920 -8798 54980 -8408
rect 55880 -8438 56900 -8418
rect 55010 -8528 55020 -8448
rect 55120 -8528 55740 -8448
rect 55810 -8528 55820 -8448
rect 55870 -8528 55880 -8438
rect 55970 -8528 56480 -8438
rect 56550 -8528 56900 -8438
rect 55880 -8548 56900 -8528
rect 57020 -8420 57040 -8418
rect 57800 -8420 58240 -8410
rect 57020 -8540 57800 -8420
rect 57020 -8548 57040 -8540
rect 57800 -8550 58240 -8540
rect 58516 -8460 58796 -8390
rect 58516 -8660 58556 -8460
rect 58756 -8660 58796 -8460
rect 59066 -8410 59936 -8400
rect 59066 -8480 59076 -8410
rect 59166 -8430 59826 -8410
rect 59166 -8480 59316 -8430
rect 59066 -8490 59316 -8480
rect 59376 -8480 59826 -8430
rect 59916 -8480 59936 -8410
rect 59376 -8490 59936 -8480
rect 60076 -8480 60196 -8440
rect 59066 -8570 59936 -8560
rect 59066 -8640 59076 -8570
rect 59166 -8640 59206 -8570
rect 59266 -8640 59826 -8570
rect 59926 -8640 59936 -8570
rect 59066 -8650 59936 -8640
rect 60076 -8640 60096 -8480
rect 60176 -8640 60196 -8480
rect 58516 -8740 58796 -8660
rect 60076 -8680 60196 -8640
rect 61266 -8450 61366 -8440
rect 61266 -8660 61276 -8450
rect 61356 -8660 61366 -8450
rect 61266 -8670 61366 -8660
rect 59586 -8690 59656 -8680
rect 59796 -8690 59866 -8680
rect 59586 -8710 59796 -8690
rect 59156 -8720 59536 -8710
rect 59156 -8730 59266 -8720
rect 54910 -8868 54920 -8798
rect 54980 -8868 54990 -8798
rect 59156 -8810 59166 -8730
rect 59226 -8810 59266 -8730
rect 59366 -8730 59536 -8720
rect 59366 -8810 59466 -8730
rect 59526 -8810 59536 -8730
rect 59156 -8830 59536 -8810
rect 59646 -8850 59796 -8710
rect 59586 -8870 59796 -8850
rect 59856 -8870 59866 -8690
rect 53840 -9048 53850 -8938
rect 53920 -9038 55000 -8938
rect 55090 -9038 55540 -8938
rect 55630 -9038 55640 -8938
rect 56470 -8988 56480 -8928
rect 56550 -8988 56560 -8928
rect 57088 -9014 57098 -8874
rect 57368 -9014 57378 -8874
rect 59796 -8880 59866 -8870
rect 59906 -8690 60016 -8680
rect 59906 -8880 59916 -8690
rect 60006 -8880 60016 -8690
rect 60476 -8710 60546 -8700
rect 60536 -8770 60546 -8710
rect 60476 -8780 60546 -8770
rect 60966 -8830 61486 -8820
rect 60966 -8840 61336 -8830
rect 59906 -8890 60016 -8880
rect 60466 -8850 61336 -8840
rect 59506 -8910 59606 -8900
rect 59156 -8960 59376 -8940
rect 53920 -9048 55640 -9038
rect 59156 -9040 59166 -8960
rect 59226 -9040 59266 -8960
rect 59156 -9050 59266 -9040
rect 59366 -9050 59376 -8960
rect 59506 -8980 59516 -8910
rect 59596 -8980 59606 -8910
rect 60466 -8910 60476 -8850
rect 60536 -8910 60616 -8850
rect 60736 -8910 60756 -8850
rect 60816 -8910 60896 -8850
rect 60956 -8910 61336 -8850
rect 60466 -8920 61336 -8910
rect 60966 -8960 61336 -8920
rect 61456 -8960 61486 -8830
rect 60966 -8970 61486 -8960
rect 59506 -8990 59606 -8980
rect 59156 -9060 59376 -9050
rect 59306 -9120 60336 -9100
rect 59066 -9140 59176 -9130
rect 55210 -9318 55220 -9148
rect 55310 -9318 55320 -9148
rect 55400 -9328 55410 -9158
rect 55500 -9168 55510 -9158
rect 55500 -9288 56380 -9168
rect 56440 -9288 56450 -9168
rect 59066 -9200 59076 -9140
rect 59166 -9200 59176 -9140
rect 59306 -9180 59316 -9120
rect 59376 -9140 59966 -9120
rect 59376 -9180 59816 -9140
rect 59306 -9190 59816 -9180
rect 59846 -9180 59916 -9170
rect 59066 -9210 59176 -9200
rect 59846 -9240 59856 -9180
rect 59946 -9180 59966 -9140
rect 60326 -9180 60336 -9120
rect 59946 -9190 60336 -9180
rect 60366 -9140 61146 -9130
rect 60366 -9180 61056 -9140
rect 59646 -9250 59716 -9240
rect 59846 -9250 59916 -9240
rect 60366 -9240 60376 -9180
rect 60436 -9240 61056 -9180
rect 61126 -9240 61146 -9140
rect 55500 -9308 56450 -9288
rect 58396 -9260 59716 -9250
rect 55500 -9328 55510 -9308
rect 58396 -9330 58926 -9260
rect 58986 -9330 59146 -9260
rect 59226 -9330 59276 -9260
rect 59356 -9330 59396 -9260
rect 59476 -9320 59646 -9260
rect 59706 -9320 59716 -9260
rect 60366 -9270 61146 -9240
rect 59476 -9330 59716 -9320
rect 58396 -9340 59716 -9330
rect 54900 -9408 54910 -9398
rect 53940 -9488 53950 -9408
rect 54010 -9488 54910 -9408
rect 53940 -9498 54910 -9488
rect 54980 -9418 54990 -9398
rect 54980 -9478 55980 -9418
rect 54980 -9498 55880 -9478
rect 53940 -9518 55880 -9498
rect 53500 -9648 53510 -9528
rect 53630 -9648 53640 -9528
rect 55850 -9558 55880 -9518
rect 55970 -9558 55980 -9478
rect 55230 -9618 55240 -9558
rect 55370 -9578 55710 -9558
rect 55370 -9588 55720 -9578
rect 55370 -9608 55620 -9588
rect 55370 -9618 55380 -9608
rect 55400 -9668 55410 -9648
rect 54730 -9758 54740 -9668
rect 54850 -9738 55410 -9668
rect 55510 -9738 55520 -9648
rect 55600 -9678 55620 -9608
rect 55710 -9678 55720 -9588
rect 54850 -9758 55520 -9738
rect 55210 -9928 55220 -9818
rect 55330 -9928 55340 -9818
rect 55850 -9978 55980 -9558
rect 56010 -9808 56020 -9658
rect 56080 -9808 56090 -9658
rect 56160 -9808 56170 -9608
rect 56390 -9808 56400 -9608
rect 58396 -9620 58896 -9340
rect 59006 -9500 59076 -9480
rect 59246 -9490 59256 -9430
rect 59366 -9490 59376 -9430
rect 59536 -9460 59546 -9390
rect 59606 -9460 59616 -9390
rect 59536 -9470 59616 -9460
rect 59006 -9560 59016 -9500
rect 59536 -9510 59616 -9500
rect 59076 -9520 59086 -9510
rect 59536 -9520 59546 -9510
rect 59076 -9560 59546 -9520
rect 59006 -9570 59546 -9560
rect 59606 -9570 59616 -9510
rect 59006 -9590 59076 -9570
rect 59536 -9590 59616 -9570
rect 59646 -9620 59716 -9340
rect 59796 -9410 59926 -9400
rect 59796 -9520 59806 -9410
rect 59916 -9520 59926 -9410
rect 59796 -9530 59926 -9520
rect 60436 -9430 60536 -9410
rect 60436 -9550 60446 -9430
rect 60526 -9550 60536 -9430
rect 60436 -9560 60536 -9550
rect 58396 -9630 59716 -9620
rect 56654 -9668 56998 -9658
rect 55520 -10068 55530 -9978
rect 55610 -10068 55980 -9978
rect 54130 -10348 54140 -10088
rect 54850 -10348 54860 -10088
rect 55310 -10268 55320 -10128
rect 55470 -10268 55480 -10128
rect 56170 -10338 56390 -9808
rect 58396 -9700 58906 -9630
rect 58986 -9700 59146 -9630
rect 59226 -9700 59276 -9630
rect 59356 -9700 59396 -9630
rect 59476 -9640 59716 -9630
rect 59476 -9700 59646 -9640
rect 59706 -9700 59716 -9640
rect 58396 -9710 59716 -9700
rect 58396 -9750 58896 -9710
rect 59646 -9720 59716 -9710
rect 56654 -9896 56998 -9886
rect 59006 -9800 60416 -9790
rect 59006 -9840 60266 -9800
rect 59006 -9910 59016 -9840
rect 59076 -9910 59546 -9840
rect 59606 -9910 60266 -9840
rect 59006 -9930 60266 -9910
rect 60406 -9930 60416 -9800
rect 59006 -9940 60416 -9930
rect 59986 -9990 60116 -9980
rect 58956 -10000 59156 -9990
rect 58956 -10180 58966 -10000
rect 59146 -10180 59156 -10000
rect 59986 -10100 59996 -9990
rect 60106 -10100 60116 -9990
rect 59986 -10110 60116 -10100
rect 58956 -10190 59156 -10180
rect 55680 -10348 56390 -10338
rect 54130 -10508 56390 -10348
rect 55680 -10518 56390 -10508
rect 59600 -10300 60500 -10200
rect 55400 -10700 56100 -10600
rect 55400 -11100 55500 -10700
rect 56000 -11100 56100 -10700
rect 59600 -10700 59700 -10300
rect 60400 -10700 60500 -10300
rect 59600 -10800 60500 -10700
rect 66800 -10300 67500 -10200
rect 66800 -10700 66900 -10300
rect 67400 -10700 67500 -10300
rect 55400 -11200 56100 -11100
rect 51400 -11900 51500 -11700
rect 52500 -11900 52600 -11700
rect 51400 -17100 52600 -11900
rect 55320 -11660 55800 -11600
rect 55320 -11980 55380 -11660
rect 55740 -11980 55800 -11660
rect 55320 -12040 55800 -11980
rect 54140 -12138 56390 -12128
rect 53460 -12340 53800 -12320
rect 53460 -12540 53480 -12340
rect 53780 -12540 53800 -12340
rect 54140 -12378 54150 -12138
rect 54860 -12378 56390 -12138
rect 58946 -12270 59146 -12250
rect 54140 -12388 56390 -12378
rect 53460 -12560 53800 -12540
rect 54850 -12618 55530 -12608
rect 53510 -12768 53520 -12658
rect 53640 -12768 53650 -12658
rect 54740 -12718 54750 -12638
rect 54850 -12688 55430 -12618
rect 55520 -12688 55530 -12618
rect 55950 -12688 55960 -12538
rect 56040 -12688 56050 -12538
rect 56170 -12558 56390 -12388
rect 56506 -12380 57016 -12370
rect 54840 -12718 54850 -12708
rect 55270 -12808 55280 -12718
rect 55400 -12808 55410 -12718
rect 56170 -12768 56190 -12558
rect 56390 -12768 56400 -12558
rect 58946 -12430 58966 -12270
rect 59126 -12430 59146 -12270
rect 58946 -12450 59146 -12430
rect 59316 -12300 60176 -12290
rect 59316 -12310 59956 -12300
rect 59316 -12450 59336 -12310
rect 59416 -12450 59956 -12310
rect 59316 -12460 59956 -12450
rect 60166 -12460 60176 -12300
rect 59316 -12470 60176 -12460
rect 56506 -12640 57016 -12630
rect 58956 -12520 61136 -12510
rect 58956 -12530 61056 -12520
rect 58956 -12640 58996 -12530
rect 59106 -12540 61056 -12530
rect 59106 -12640 59516 -12540
rect 59616 -12640 61056 -12540
rect 58396 -12730 58896 -12640
rect 58956 -12650 61056 -12640
rect 61126 -12650 61136 -12520
rect 58956 -12660 61136 -12650
rect 55850 -12848 55880 -12818
rect 53940 -12878 55880 -12848
rect 53940 -12898 54920 -12878
rect 53040 -14708 53050 -12958
rect 53250 -14708 53260 -12958
rect 53940 -12998 53950 -12898
rect 54020 -12948 54920 -12898
rect 54020 -12998 54030 -12948
rect 54910 -12968 54920 -12948
rect 54990 -12898 55880 -12878
rect 55970 -12848 55980 -12818
rect 54990 -12948 55970 -12898
rect 54990 -12968 55000 -12948
rect 55220 -13228 55230 -13058
rect 55320 -13228 55330 -13058
rect 55420 -13218 55430 -13048
rect 55510 -13058 55520 -13048
rect 55510 -13068 56670 -13058
rect 55510 -13198 55600 -13068
rect 55710 -13198 56590 -13068
rect 56660 -13198 56670 -13068
rect 55510 -13208 56670 -13198
rect 58396 -13090 58486 -12730
rect 58816 -12750 58896 -12730
rect 59646 -12750 59706 -12730
rect 58816 -12770 59706 -12750
rect 58816 -12830 58906 -12770
rect 58966 -12830 59216 -12770
rect 59276 -12830 59326 -12770
rect 59386 -12830 59436 -12770
rect 59496 -12830 59636 -12770
rect 59696 -12830 59706 -12770
rect 58816 -12840 59706 -12830
rect 58816 -13090 58896 -12840
rect 59536 -12890 59616 -12880
rect 59276 -12930 59356 -12920
rect 59276 -12990 59286 -12930
rect 59346 -12990 59356 -12930
rect 59536 -12950 59546 -12890
rect 59606 -12950 59616 -12890
rect 59536 -12970 59616 -12950
rect 58996 -13000 59076 -12990
rect 58996 -13060 59006 -13000
rect 59076 -13020 59086 -13000
rect 59536 -13010 59616 -13000
rect 59536 -13020 59546 -13010
rect 59076 -13060 59546 -13020
rect 58996 -13070 59076 -13060
rect 59536 -13070 59546 -13060
rect 59606 -13070 59616 -13010
rect 59536 -13080 59616 -13070
rect 58396 -13110 58896 -13090
rect 59646 -13110 59706 -12840
rect 60436 -12920 60536 -12910
rect 59856 -12940 59976 -12930
rect 59856 -13030 59866 -12940
rect 59966 -13030 59976 -12940
rect 60436 -13020 60446 -12920
rect 60526 -13020 60536 -12920
rect 60436 -13030 60536 -13020
rect 59856 -13040 59976 -13030
rect 58396 -13120 59706 -13110
rect 58396 -13130 59216 -13120
rect 58396 -13190 58906 -13130
rect 58966 -13180 59216 -13130
rect 59276 -13180 59336 -13120
rect 59396 -13180 59436 -13120
rect 59496 -13130 59706 -13120
rect 59496 -13180 59636 -13130
rect 58966 -13190 59636 -13180
rect 59696 -13190 59706 -13130
rect 58396 -13200 59706 -13190
rect 60036 -13120 60136 -13110
rect 60036 -13200 60046 -13120
rect 60126 -13200 60136 -13120
rect 55510 -13218 55520 -13208
rect 59646 -13210 59706 -13200
rect 60546 -13210 60636 -13200
rect 59066 -13240 59176 -13230
rect 59066 -13310 59076 -13240
rect 59166 -13310 59176 -13240
rect 59846 -13280 59856 -13210
rect 59916 -13230 59926 -13210
rect 60356 -13220 60556 -13210
rect 60356 -13230 60376 -13220
rect 59916 -13260 60376 -13230
rect 59916 -13280 59926 -13260
rect 60356 -13280 60376 -13260
rect 60446 -13280 60556 -13220
rect 60356 -13290 60556 -13280
rect 60626 -13290 60636 -13210
rect 59066 -13320 59176 -13310
rect 59966 -13300 60326 -13290
rect 53850 -13438 53860 -13328
rect 53920 -13338 55600 -13328
rect 53920 -13438 55000 -13338
rect 55090 -13438 55540 -13338
rect 55630 -13438 55640 -13338
rect 59966 -13360 59976 -13300
rect 60316 -13360 60326 -13300
rect 60546 -13310 60636 -13290
rect 61186 -13320 61366 -13310
rect 54770 -13638 54850 -13438
rect 56470 -13448 56480 -13388
rect 56550 -13448 56560 -13388
rect 57088 -13504 57098 -13364
rect 57368 -13504 57378 -13364
rect 59166 -13430 59376 -13420
rect 59166 -13440 59286 -13430
rect 59166 -13520 59176 -13440
rect 59236 -13520 59286 -13440
rect 59366 -13520 59376 -13430
rect 59166 -13530 59376 -13520
rect 59526 -13470 59646 -13450
rect 59526 -13530 59576 -13470
rect 59636 -13530 59646 -13470
rect 61186 -13500 61206 -13320
rect 61346 -13500 61366 -13320
rect 61186 -13510 61366 -13500
rect 59526 -13560 59646 -13530
rect 60286 -13550 60476 -13540
rect 59906 -13580 60016 -13570
rect 59806 -13590 59866 -13580
rect 54760 -13728 54770 -13638
rect 54840 -13728 54850 -13638
rect 59166 -13640 59536 -13630
rect 59166 -13720 59176 -13640
rect 59236 -13720 59286 -13640
rect 54920 -13738 55210 -13728
rect 54920 -13808 55140 -13738
rect 55200 -13808 55210 -13738
rect 59166 -13730 59286 -13720
rect 59356 -13650 59536 -13640
rect 59356 -13720 59476 -13650
rect 59356 -13730 59536 -13720
rect 59166 -13740 59536 -13730
rect 59566 -13760 59576 -13590
rect 59636 -13600 59866 -13590
rect 59636 -13740 59806 -13600
rect 59636 -13760 59866 -13740
rect 59906 -13760 59916 -13580
rect 60006 -13760 60016 -13580
rect 60286 -13690 60306 -13550
rect 60456 -13690 60476 -13550
rect 60286 -13700 60476 -13690
rect 61026 -13620 61136 -13610
rect 61026 -13730 61036 -13620
rect 61126 -13730 61136 -13620
rect 61026 -13740 61136 -13730
rect 59566 -13770 59636 -13760
rect 59906 -13770 60016 -13760
rect 54760 -14128 54770 -14048
rect 54840 -14128 54850 -14048
rect 54770 -14338 54850 -14128
rect 54920 -14198 54980 -13808
rect 55880 -13838 56900 -13818
rect 55010 -13928 55020 -13848
rect 55120 -13928 55740 -13848
rect 55810 -13928 55820 -13848
rect 55870 -13928 55880 -13838
rect 55970 -13928 56480 -13838
rect 56550 -13928 56900 -13838
rect 55880 -13948 56900 -13928
rect 57020 -13820 57040 -13818
rect 57800 -13820 58240 -13810
rect 57020 -13940 57800 -13820
rect 57020 -13948 57040 -13940
rect 57800 -13950 58240 -13940
rect 58516 -13860 58796 -13790
rect 58516 -14060 58556 -13860
rect 58756 -14060 58796 -13860
rect 59066 -13810 59936 -13800
rect 59066 -13880 59076 -13810
rect 59166 -13830 59826 -13810
rect 59166 -13880 59316 -13830
rect 59066 -13890 59316 -13880
rect 59376 -13880 59826 -13830
rect 59916 -13880 59936 -13810
rect 59376 -13890 59936 -13880
rect 60076 -13880 60196 -13840
rect 59066 -13970 59936 -13960
rect 59066 -14040 59076 -13970
rect 59166 -14040 59206 -13970
rect 59266 -14040 59826 -13970
rect 59926 -14040 59936 -13970
rect 59066 -14050 59936 -14040
rect 60076 -14040 60096 -13880
rect 60176 -14040 60196 -13880
rect 58516 -14140 58796 -14060
rect 60076 -14080 60196 -14040
rect 61266 -13850 61366 -13840
rect 61266 -14060 61276 -13850
rect 61356 -14060 61366 -13850
rect 61266 -14070 61366 -14060
rect 59586 -14090 59656 -14080
rect 59796 -14090 59866 -14080
rect 59586 -14110 59796 -14090
rect 59156 -14120 59536 -14110
rect 59156 -14130 59266 -14120
rect 54910 -14268 54920 -14198
rect 54980 -14268 54990 -14198
rect 59156 -14210 59166 -14130
rect 59226 -14210 59266 -14130
rect 59366 -14130 59536 -14120
rect 59366 -14210 59466 -14130
rect 59526 -14210 59536 -14130
rect 59156 -14230 59536 -14210
rect 59646 -14250 59796 -14110
rect 59586 -14270 59796 -14250
rect 59856 -14270 59866 -14090
rect 53840 -14448 53850 -14338
rect 53920 -14438 55000 -14338
rect 55090 -14438 55540 -14338
rect 55630 -14438 55640 -14338
rect 56470 -14388 56480 -14328
rect 56550 -14388 56560 -14328
rect 57088 -14414 57098 -14274
rect 57368 -14414 57378 -14274
rect 59796 -14280 59866 -14270
rect 59906 -14090 60016 -14080
rect 59906 -14280 59916 -14090
rect 60006 -14280 60016 -14090
rect 60476 -14110 60546 -14100
rect 60536 -14170 60546 -14110
rect 60476 -14180 60546 -14170
rect 60966 -14230 61486 -14220
rect 60966 -14240 61336 -14230
rect 59906 -14290 60016 -14280
rect 60466 -14250 61336 -14240
rect 59506 -14310 59606 -14300
rect 59156 -14360 59376 -14340
rect 53920 -14448 55640 -14438
rect 59156 -14440 59166 -14360
rect 59226 -14440 59266 -14360
rect 59156 -14450 59266 -14440
rect 59366 -14450 59376 -14360
rect 59506 -14380 59516 -14310
rect 59596 -14380 59606 -14310
rect 60466 -14310 60476 -14250
rect 60536 -14310 60616 -14250
rect 60736 -14310 60756 -14250
rect 60816 -14310 60896 -14250
rect 60956 -14310 61336 -14250
rect 60466 -14320 61336 -14310
rect 60966 -14360 61336 -14320
rect 61456 -14360 61486 -14230
rect 60966 -14370 61486 -14360
rect 59506 -14390 59606 -14380
rect 59156 -14460 59376 -14450
rect 59306 -14520 60336 -14500
rect 59066 -14540 59176 -14530
rect 55210 -14718 55220 -14548
rect 55310 -14718 55320 -14548
rect 55400 -14728 55410 -14558
rect 55500 -14568 55510 -14558
rect 55500 -14688 56380 -14568
rect 56440 -14688 56450 -14568
rect 59066 -14600 59076 -14540
rect 59166 -14600 59176 -14540
rect 59306 -14580 59316 -14520
rect 59376 -14540 59966 -14520
rect 59376 -14580 59816 -14540
rect 59306 -14590 59816 -14580
rect 59846 -14580 59916 -14570
rect 59066 -14610 59176 -14600
rect 59846 -14640 59856 -14580
rect 59946 -14580 59966 -14540
rect 60326 -14580 60336 -14520
rect 59946 -14590 60336 -14580
rect 60366 -14540 61146 -14530
rect 60366 -14580 61056 -14540
rect 59646 -14650 59716 -14640
rect 59846 -14650 59916 -14640
rect 60366 -14640 60376 -14580
rect 60436 -14640 61056 -14580
rect 61126 -14640 61146 -14540
rect 55500 -14708 56450 -14688
rect 58396 -14660 59716 -14650
rect 55500 -14728 55510 -14708
rect 58396 -14730 58926 -14660
rect 58986 -14730 59146 -14660
rect 59226 -14730 59276 -14660
rect 59356 -14730 59396 -14660
rect 59476 -14720 59646 -14660
rect 59706 -14720 59716 -14660
rect 60366 -14670 61146 -14640
rect 59476 -14730 59716 -14720
rect 58396 -14740 59716 -14730
rect 54900 -14808 54910 -14798
rect 53940 -14888 53950 -14808
rect 54010 -14888 54910 -14808
rect 53940 -14898 54910 -14888
rect 54980 -14818 54990 -14798
rect 54980 -14878 55980 -14818
rect 54980 -14898 55880 -14878
rect 53940 -14918 55880 -14898
rect 53500 -15048 53510 -14928
rect 53630 -15048 53640 -14928
rect 55850 -14958 55880 -14918
rect 55970 -14958 55980 -14878
rect 55230 -15018 55240 -14958
rect 55370 -14978 55710 -14958
rect 55370 -14988 55720 -14978
rect 55370 -15008 55620 -14988
rect 55370 -15018 55380 -15008
rect 55400 -15068 55410 -15048
rect 54730 -15158 54740 -15068
rect 54850 -15138 55410 -15068
rect 55510 -15138 55520 -15048
rect 55600 -15078 55620 -15008
rect 55710 -15078 55720 -14988
rect 54850 -15158 55520 -15138
rect 55210 -15328 55220 -15218
rect 55330 -15328 55340 -15218
rect 55850 -15378 55980 -14958
rect 56010 -15208 56020 -15058
rect 56080 -15208 56090 -15058
rect 56160 -15208 56170 -15008
rect 56390 -15208 56400 -15008
rect 58396 -15020 58896 -14740
rect 59006 -14900 59076 -14880
rect 59246 -14890 59256 -14830
rect 59366 -14890 59376 -14830
rect 59536 -14860 59546 -14790
rect 59606 -14860 59616 -14790
rect 59536 -14870 59616 -14860
rect 59006 -14960 59016 -14900
rect 59536 -14910 59616 -14900
rect 59076 -14920 59086 -14910
rect 59536 -14920 59546 -14910
rect 59076 -14960 59546 -14920
rect 59006 -14970 59546 -14960
rect 59606 -14970 59616 -14910
rect 59006 -14990 59076 -14970
rect 59536 -14990 59616 -14970
rect 59646 -15020 59716 -14740
rect 59796 -14810 59926 -14800
rect 59796 -14920 59806 -14810
rect 59916 -14920 59926 -14810
rect 59796 -14930 59926 -14920
rect 60436 -14830 60536 -14810
rect 60436 -14950 60446 -14830
rect 60526 -14950 60536 -14830
rect 60436 -14960 60536 -14950
rect 58396 -15030 59716 -15020
rect 56654 -15068 56998 -15058
rect 55520 -15468 55530 -15378
rect 55610 -15468 55980 -15378
rect 54130 -15748 54140 -15488
rect 54850 -15748 54860 -15488
rect 55310 -15668 55320 -15528
rect 55470 -15668 55480 -15528
rect 56170 -15738 56390 -15208
rect 58396 -15100 58906 -15030
rect 58986 -15100 59146 -15030
rect 59226 -15100 59276 -15030
rect 59356 -15100 59396 -15030
rect 59476 -15040 59716 -15030
rect 59476 -15100 59646 -15040
rect 59706 -15100 59716 -15040
rect 58396 -15110 59716 -15100
rect 58396 -15150 58896 -15110
rect 59646 -15120 59716 -15110
rect 56654 -15296 56998 -15286
rect 59006 -15200 60416 -15190
rect 59006 -15240 60266 -15200
rect 59006 -15310 59016 -15240
rect 59076 -15310 59546 -15240
rect 59606 -15310 60266 -15240
rect 59006 -15330 60266 -15310
rect 60406 -15330 60416 -15200
rect 59006 -15340 60416 -15330
rect 59986 -15390 60116 -15380
rect 58956 -15400 59156 -15390
rect 58956 -15580 58966 -15400
rect 59146 -15580 59156 -15400
rect 59986 -15500 59996 -15390
rect 60106 -15500 60116 -15390
rect 58956 -15590 59156 -15580
rect 55680 -15748 56390 -15738
rect 54130 -15908 56390 -15748
rect 55680 -15918 56390 -15908
rect 59700 -15600 60400 -15500
rect 59700 -15900 59800 -15600
rect 60300 -15900 60400 -15600
rect 59700 -16000 60400 -15900
rect 65800 -15600 66500 -15500
rect 65800 -15900 65900 -15600
rect 66400 -15900 66500 -15600
rect 55400 -16100 56100 -16000
rect 55400 -16500 55500 -16100
rect 56000 -16500 56100 -16100
rect 55400 -16600 56100 -16500
rect 51400 -17300 51500 -17100
rect 52500 -17300 52600 -17100
rect 51400 -22500 52600 -17300
rect 55360 -17100 55740 -17060
rect 55360 -17400 55400 -17100
rect 55700 -17400 55740 -17100
rect 55360 -17420 55740 -17400
rect 54140 -17538 56390 -17528
rect 53480 -17740 53800 -17720
rect 53480 -17940 53500 -17740
rect 53780 -17940 53800 -17740
rect 54140 -17778 54150 -17538
rect 54860 -17778 56390 -17538
rect 58946 -17670 59146 -17650
rect 54140 -17788 56390 -17778
rect 53480 -17960 53800 -17940
rect 54850 -18018 55530 -18008
rect 53510 -18168 53520 -18058
rect 53640 -18168 53650 -18058
rect 54740 -18118 54750 -18038
rect 54850 -18088 55430 -18018
rect 55520 -18088 55530 -18018
rect 55950 -18088 55960 -17938
rect 56040 -18088 56050 -17938
rect 56170 -17958 56390 -17788
rect 56506 -17780 57016 -17770
rect 54840 -18118 54850 -18108
rect 55270 -18208 55280 -18118
rect 55400 -18208 55410 -18118
rect 56170 -18168 56190 -17958
rect 56390 -18168 56400 -17958
rect 58946 -17830 58966 -17670
rect 59126 -17830 59146 -17670
rect 58946 -17850 59146 -17830
rect 59316 -17700 60176 -17690
rect 59316 -17710 59956 -17700
rect 59316 -17850 59336 -17710
rect 59416 -17850 59956 -17710
rect 59316 -17860 59956 -17850
rect 60166 -17860 60176 -17700
rect 59316 -17870 60176 -17860
rect 56506 -18040 57016 -18030
rect 58956 -17920 61136 -17910
rect 58956 -17930 61056 -17920
rect 58956 -18040 58996 -17930
rect 59106 -17940 61056 -17930
rect 59106 -18040 59516 -17940
rect 59616 -18040 61056 -17940
rect 58396 -18130 58896 -18040
rect 58956 -18050 61056 -18040
rect 61126 -18050 61136 -17920
rect 58956 -18060 61136 -18050
rect 55850 -18248 55880 -18218
rect 53940 -18278 55880 -18248
rect 53940 -18298 54920 -18278
rect 53040 -20108 53050 -18358
rect 53250 -20108 53260 -18358
rect 53940 -18398 53950 -18298
rect 54020 -18348 54920 -18298
rect 54020 -18398 54030 -18348
rect 54910 -18368 54920 -18348
rect 54990 -18298 55880 -18278
rect 55970 -18248 55980 -18218
rect 54990 -18348 55970 -18298
rect 54990 -18368 55000 -18348
rect 55220 -18628 55230 -18458
rect 55320 -18628 55330 -18458
rect 55420 -18618 55430 -18448
rect 55510 -18458 55520 -18448
rect 55510 -18468 56670 -18458
rect 55510 -18598 55600 -18468
rect 55710 -18598 56590 -18468
rect 56660 -18598 56670 -18468
rect 55510 -18608 56670 -18598
rect 58396 -18490 58486 -18130
rect 58816 -18150 58896 -18130
rect 59646 -18150 59706 -18130
rect 58816 -18170 59706 -18150
rect 58816 -18230 58906 -18170
rect 58966 -18230 59216 -18170
rect 59276 -18230 59326 -18170
rect 59386 -18230 59436 -18170
rect 59496 -18230 59636 -18170
rect 59696 -18230 59706 -18170
rect 58816 -18240 59706 -18230
rect 58816 -18490 58896 -18240
rect 59536 -18290 59616 -18280
rect 59276 -18330 59356 -18320
rect 59276 -18390 59286 -18330
rect 59346 -18390 59356 -18330
rect 59536 -18350 59546 -18290
rect 59606 -18350 59616 -18290
rect 59536 -18370 59616 -18350
rect 58996 -18400 59076 -18390
rect 58996 -18460 59006 -18400
rect 59076 -18420 59086 -18400
rect 59536 -18410 59616 -18400
rect 59536 -18420 59546 -18410
rect 59076 -18460 59546 -18420
rect 58996 -18470 59076 -18460
rect 59536 -18470 59546 -18460
rect 59606 -18470 59616 -18410
rect 59536 -18480 59616 -18470
rect 58396 -18510 58896 -18490
rect 59646 -18510 59706 -18240
rect 60436 -18320 60536 -18310
rect 59856 -18340 59976 -18330
rect 59856 -18430 59866 -18340
rect 59966 -18430 59976 -18340
rect 60436 -18420 60446 -18320
rect 60526 -18420 60536 -18320
rect 60436 -18430 60536 -18420
rect 59856 -18440 59976 -18430
rect 58396 -18520 59706 -18510
rect 58396 -18530 59216 -18520
rect 58396 -18590 58906 -18530
rect 58966 -18580 59216 -18530
rect 59276 -18580 59336 -18520
rect 59396 -18580 59436 -18520
rect 59496 -18530 59706 -18520
rect 59496 -18580 59636 -18530
rect 58966 -18590 59636 -18580
rect 59696 -18590 59706 -18530
rect 58396 -18600 59706 -18590
rect 60036 -18520 60136 -18510
rect 60036 -18600 60046 -18520
rect 60126 -18600 60136 -18520
rect 55510 -18618 55520 -18608
rect 59646 -18610 59706 -18600
rect 60546 -18610 60636 -18600
rect 59066 -18640 59176 -18630
rect 59066 -18710 59076 -18640
rect 59166 -18710 59176 -18640
rect 59846 -18680 59856 -18610
rect 59916 -18630 59926 -18610
rect 60356 -18620 60556 -18610
rect 60356 -18630 60376 -18620
rect 59916 -18660 60376 -18630
rect 59916 -18680 59926 -18660
rect 60356 -18680 60376 -18660
rect 60446 -18680 60556 -18620
rect 60356 -18690 60556 -18680
rect 60626 -18690 60636 -18610
rect 59066 -18720 59176 -18710
rect 59966 -18700 60326 -18690
rect 53850 -18838 53860 -18728
rect 53920 -18738 55600 -18728
rect 53920 -18838 55000 -18738
rect 55090 -18838 55540 -18738
rect 55630 -18838 55640 -18738
rect 59966 -18760 59976 -18700
rect 60316 -18760 60326 -18700
rect 60546 -18710 60636 -18690
rect 61186 -18720 61366 -18710
rect 54770 -19038 54850 -18838
rect 56470 -18848 56480 -18788
rect 56550 -18848 56560 -18788
rect 57088 -18904 57098 -18764
rect 57368 -18904 57378 -18764
rect 59166 -18830 59376 -18820
rect 59166 -18840 59286 -18830
rect 59166 -18920 59176 -18840
rect 59236 -18920 59286 -18840
rect 59366 -18920 59376 -18830
rect 59166 -18930 59376 -18920
rect 59526 -18870 59646 -18850
rect 59526 -18930 59576 -18870
rect 59636 -18930 59646 -18870
rect 61186 -18900 61206 -18720
rect 61346 -18900 61366 -18720
rect 61186 -18910 61366 -18900
rect 59526 -18960 59646 -18930
rect 60286 -18950 60476 -18940
rect 59906 -18980 60016 -18970
rect 59806 -18990 59866 -18980
rect 54760 -19128 54770 -19038
rect 54840 -19128 54850 -19038
rect 59166 -19040 59536 -19030
rect 59166 -19120 59176 -19040
rect 59236 -19120 59286 -19040
rect 54920 -19138 55210 -19128
rect 54920 -19208 55140 -19138
rect 55200 -19208 55210 -19138
rect 59166 -19130 59286 -19120
rect 59356 -19050 59536 -19040
rect 59356 -19120 59476 -19050
rect 59356 -19130 59536 -19120
rect 59166 -19140 59536 -19130
rect 59566 -19160 59576 -18990
rect 59636 -19000 59866 -18990
rect 59636 -19140 59806 -19000
rect 59636 -19160 59866 -19140
rect 59906 -19160 59916 -18980
rect 60006 -19160 60016 -18980
rect 60286 -19090 60306 -18950
rect 60456 -19090 60476 -18950
rect 60286 -19100 60476 -19090
rect 61026 -19020 61136 -19010
rect 61026 -19130 61036 -19020
rect 61126 -19130 61136 -19020
rect 61026 -19140 61136 -19130
rect 59566 -19170 59636 -19160
rect 59906 -19170 60016 -19160
rect 54760 -19528 54770 -19448
rect 54840 -19528 54850 -19448
rect 54770 -19738 54850 -19528
rect 54920 -19598 54980 -19208
rect 55880 -19238 56900 -19218
rect 55010 -19328 55020 -19248
rect 55120 -19328 55740 -19248
rect 55810 -19328 55820 -19248
rect 55870 -19328 55880 -19238
rect 55970 -19328 56480 -19238
rect 56550 -19328 56900 -19238
rect 55880 -19348 56900 -19328
rect 57020 -19220 57040 -19218
rect 57800 -19220 58240 -19210
rect 57020 -19340 57800 -19220
rect 57020 -19348 57040 -19340
rect 57800 -19350 58240 -19340
rect 58516 -19260 58796 -19190
rect 58516 -19460 58556 -19260
rect 58756 -19460 58796 -19260
rect 59066 -19210 59936 -19200
rect 59066 -19280 59076 -19210
rect 59166 -19230 59826 -19210
rect 59166 -19280 59316 -19230
rect 59066 -19290 59316 -19280
rect 59376 -19280 59826 -19230
rect 59916 -19280 59936 -19210
rect 59376 -19290 59936 -19280
rect 60076 -19280 60196 -19240
rect 59066 -19370 59936 -19360
rect 59066 -19440 59076 -19370
rect 59166 -19440 59206 -19370
rect 59266 -19440 59826 -19370
rect 59926 -19440 59936 -19370
rect 59066 -19450 59936 -19440
rect 60076 -19440 60096 -19280
rect 60176 -19440 60196 -19280
rect 58516 -19540 58796 -19460
rect 60076 -19480 60196 -19440
rect 61266 -19250 61366 -19240
rect 61266 -19460 61276 -19250
rect 61356 -19460 61366 -19250
rect 61266 -19470 61366 -19460
rect 59586 -19490 59656 -19480
rect 59796 -19490 59866 -19480
rect 59586 -19510 59796 -19490
rect 59156 -19520 59536 -19510
rect 59156 -19530 59266 -19520
rect 54910 -19668 54920 -19598
rect 54980 -19668 54990 -19598
rect 59156 -19610 59166 -19530
rect 59226 -19610 59266 -19530
rect 59366 -19530 59536 -19520
rect 59366 -19610 59466 -19530
rect 59526 -19610 59536 -19530
rect 59156 -19630 59536 -19610
rect 59646 -19650 59796 -19510
rect 59586 -19670 59796 -19650
rect 59856 -19670 59866 -19490
rect 53840 -19848 53850 -19738
rect 53920 -19838 55000 -19738
rect 55090 -19838 55540 -19738
rect 55630 -19838 55640 -19738
rect 56470 -19788 56480 -19728
rect 56550 -19788 56560 -19728
rect 57088 -19814 57098 -19674
rect 57368 -19814 57378 -19674
rect 59796 -19680 59866 -19670
rect 59906 -19490 60016 -19480
rect 59906 -19680 59916 -19490
rect 60006 -19680 60016 -19490
rect 60476 -19510 60546 -19500
rect 60536 -19570 60546 -19510
rect 60476 -19580 60546 -19570
rect 60966 -19630 61486 -19620
rect 60966 -19640 61336 -19630
rect 59906 -19690 60016 -19680
rect 60466 -19650 61336 -19640
rect 59506 -19710 59606 -19700
rect 59156 -19760 59376 -19740
rect 53920 -19848 55640 -19838
rect 59156 -19840 59166 -19760
rect 59226 -19840 59266 -19760
rect 59156 -19850 59266 -19840
rect 59366 -19850 59376 -19760
rect 59506 -19780 59516 -19710
rect 59596 -19780 59606 -19710
rect 60466 -19710 60476 -19650
rect 60536 -19710 60616 -19650
rect 60736 -19710 60756 -19650
rect 60816 -19710 60896 -19650
rect 60956 -19710 61336 -19650
rect 60466 -19720 61336 -19710
rect 60966 -19760 61336 -19720
rect 61456 -19760 61486 -19630
rect 60966 -19770 61486 -19760
rect 59506 -19790 59606 -19780
rect 59156 -19860 59376 -19850
rect 59306 -19920 60336 -19900
rect 59066 -19940 59176 -19930
rect 55210 -20118 55220 -19948
rect 55310 -20118 55320 -19948
rect 55400 -20128 55410 -19958
rect 55500 -19968 55510 -19958
rect 55500 -20088 56380 -19968
rect 56440 -20088 56450 -19968
rect 59066 -20000 59076 -19940
rect 59166 -20000 59176 -19940
rect 59306 -19980 59316 -19920
rect 59376 -19940 59966 -19920
rect 59376 -19980 59816 -19940
rect 59306 -19990 59816 -19980
rect 59846 -19980 59916 -19970
rect 59066 -20010 59176 -20000
rect 59846 -20040 59856 -19980
rect 59946 -19980 59966 -19940
rect 60326 -19980 60336 -19920
rect 59946 -19990 60336 -19980
rect 60366 -19940 61146 -19930
rect 60366 -19980 61056 -19940
rect 59646 -20050 59716 -20040
rect 59846 -20050 59916 -20040
rect 60366 -20040 60376 -19980
rect 60436 -20040 61056 -19980
rect 61126 -20040 61146 -19940
rect 55500 -20108 56450 -20088
rect 58396 -20060 59716 -20050
rect 55500 -20128 55510 -20108
rect 58396 -20130 58926 -20060
rect 58986 -20130 59146 -20060
rect 59226 -20130 59276 -20060
rect 59356 -20130 59396 -20060
rect 59476 -20120 59646 -20060
rect 59706 -20120 59716 -20060
rect 60366 -20070 61146 -20040
rect 59476 -20130 59716 -20120
rect 58396 -20140 59716 -20130
rect 54900 -20208 54910 -20198
rect 53940 -20288 53950 -20208
rect 54010 -20288 54910 -20208
rect 53940 -20298 54910 -20288
rect 54980 -20218 54990 -20198
rect 54980 -20278 55980 -20218
rect 54980 -20298 55880 -20278
rect 53940 -20318 55880 -20298
rect 53500 -20448 53510 -20328
rect 53630 -20448 53640 -20328
rect 55850 -20358 55880 -20318
rect 55970 -20358 55980 -20278
rect 55230 -20418 55240 -20358
rect 55370 -20378 55710 -20358
rect 55370 -20388 55720 -20378
rect 55370 -20408 55620 -20388
rect 55370 -20418 55380 -20408
rect 55400 -20468 55410 -20448
rect 54730 -20558 54740 -20468
rect 54850 -20538 55410 -20468
rect 55510 -20538 55520 -20448
rect 55600 -20478 55620 -20408
rect 55710 -20478 55720 -20388
rect 54850 -20558 55520 -20538
rect 55210 -20728 55220 -20618
rect 55330 -20728 55340 -20618
rect 55850 -20778 55980 -20358
rect 56010 -20608 56020 -20458
rect 56080 -20608 56090 -20458
rect 56160 -20608 56170 -20408
rect 56390 -20608 56400 -20408
rect 58396 -20420 58896 -20140
rect 59006 -20300 59076 -20280
rect 59246 -20290 59256 -20230
rect 59366 -20290 59376 -20230
rect 59536 -20260 59546 -20190
rect 59606 -20260 59616 -20190
rect 59536 -20270 59616 -20260
rect 59006 -20360 59016 -20300
rect 59536 -20310 59616 -20300
rect 59076 -20320 59086 -20310
rect 59536 -20320 59546 -20310
rect 59076 -20360 59546 -20320
rect 59006 -20370 59546 -20360
rect 59606 -20370 59616 -20310
rect 59006 -20390 59076 -20370
rect 59536 -20390 59616 -20370
rect 59646 -20420 59716 -20140
rect 59796 -20210 59926 -20200
rect 59796 -20320 59806 -20210
rect 59916 -20320 59926 -20210
rect 59796 -20330 59926 -20320
rect 60436 -20230 60536 -20210
rect 60436 -20350 60446 -20230
rect 60526 -20350 60536 -20230
rect 60436 -20360 60536 -20350
rect 58396 -20430 59716 -20420
rect 56654 -20468 56998 -20458
rect 55520 -20868 55530 -20778
rect 55610 -20868 55980 -20778
rect 54130 -21148 54140 -20888
rect 54850 -21148 54860 -20888
rect 55310 -21068 55320 -20928
rect 55470 -21068 55480 -20928
rect 56170 -21138 56390 -20608
rect 58396 -20500 58906 -20430
rect 58986 -20500 59146 -20430
rect 59226 -20500 59276 -20430
rect 59356 -20500 59396 -20430
rect 59476 -20440 59716 -20430
rect 59476 -20500 59646 -20440
rect 59706 -20500 59716 -20440
rect 58396 -20510 59716 -20500
rect 58396 -20550 58896 -20510
rect 59646 -20520 59716 -20510
rect 56654 -20696 56998 -20686
rect 59006 -20600 60416 -20590
rect 59006 -20640 60266 -20600
rect 59006 -20710 59016 -20640
rect 59076 -20710 59546 -20640
rect 59606 -20710 60266 -20640
rect 59006 -20730 60266 -20710
rect 60406 -20730 60416 -20600
rect 59006 -20740 60416 -20730
rect 59986 -20790 60116 -20780
rect 58956 -20800 59156 -20790
rect 58956 -20980 58966 -20800
rect 59146 -20980 59156 -20800
rect 59986 -20900 59996 -20790
rect 60106 -20900 60116 -20790
rect 58956 -20990 59156 -20980
rect 55680 -21148 56390 -21138
rect 54130 -21308 56390 -21148
rect 55680 -21318 56390 -21308
rect 59700 -21000 60400 -20900
rect 59700 -21300 59800 -21000
rect 60300 -21300 60400 -21000
rect 59700 -21400 60400 -21300
rect 64800 -21000 65500 -20900
rect 64800 -21300 64900 -21000
rect 65400 -21300 65500 -21000
rect 55400 -21500 56200 -21400
rect 55400 -21900 55500 -21500
rect 56100 -21900 56200 -21500
rect 55400 -22000 56200 -21900
rect 51400 -22700 51500 -22500
rect 52500 -22700 52600 -22500
rect 51400 -27900 52600 -22700
rect 55420 -22480 55740 -22460
rect 55420 -22760 55440 -22480
rect 55720 -22760 55740 -22480
rect 55420 -22780 55740 -22760
rect 54140 -22938 56390 -22928
rect 53460 -23140 53800 -23120
rect 53460 -23340 53480 -23140
rect 53780 -23340 53800 -23140
rect 54140 -23178 54150 -22938
rect 54860 -23178 56390 -22938
rect 58946 -23070 59146 -23050
rect 54140 -23188 56390 -23178
rect 53460 -23360 53800 -23340
rect 54850 -23418 55530 -23408
rect 53510 -23568 53520 -23458
rect 53640 -23568 53650 -23458
rect 54740 -23518 54750 -23438
rect 54850 -23488 55430 -23418
rect 55520 -23488 55530 -23418
rect 55950 -23488 55960 -23338
rect 56040 -23488 56050 -23338
rect 56170 -23358 56390 -23188
rect 56506 -23180 57016 -23170
rect 54840 -23518 54850 -23508
rect 55270 -23608 55280 -23518
rect 55400 -23608 55410 -23518
rect 56170 -23568 56190 -23358
rect 56390 -23568 56400 -23358
rect 58946 -23230 58966 -23070
rect 59126 -23230 59146 -23070
rect 58946 -23250 59146 -23230
rect 59316 -23100 60176 -23090
rect 59316 -23110 59956 -23100
rect 59316 -23250 59336 -23110
rect 59416 -23250 59956 -23110
rect 59316 -23260 59956 -23250
rect 60166 -23260 60176 -23100
rect 59316 -23270 60176 -23260
rect 56506 -23440 57016 -23430
rect 58956 -23320 61136 -23310
rect 58956 -23330 61056 -23320
rect 58956 -23440 58996 -23330
rect 59106 -23340 61056 -23330
rect 59106 -23440 59516 -23340
rect 59616 -23440 61056 -23340
rect 58396 -23530 58896 -23440
rect 58956 -23450 61056 -23440
rect 61126 -23450 61136 -23320
rect 58956 -23460 61136 -23450
rect 55850 -23648 55880 -23618
rect 53940 -23678 55880 -23648
rect 53940 -23698 54920 -23678
rect 53040 -25508 53050 -23758
rect 53250 -25508 53260 -23758
rect 53940 -23798 53950 -23698
rect 54020 -23748 54920 -23698
rect 54020 -23798 54030 -23748
rect 54910 -23768 54920 -23748
rect 54990 -23698 55880 -23678
rect 55970 -23648 55980 -23618
rect 54990 -23748 55970 -23698
rect 54990 -23768 55000 -23748
rect 55220 -24028 55230 -23858
rect 55320 -24028 55330 -23858
rect 55420 -24018 55430 -23848
rect 55510 -23858 55520 -23848
rect 55510 -23868 56670 -23858
rect 55510 -23998 55600 -23868
rect 55710 -23998 56590 -23868
rect 56660 -23998 56670 -23868
rect 55510 -24008 56670 -23998
rect 58396 -23890 58486 -23530
rect 58816 -23550 58896 -23530
rect 59646 -23550 59706 -23530
rect 58816 -23570 59706 -23550
rect 58816 -23630 58906 -23570
rect 58966 -23630 59216 -23570
rect 59276 -23630 59326 -23570
rect 59386 -23630 59436 -23570
rect 59496 -23630 59636 -23570
rect 59696 -23630 59706 -23570
rect 58816 -23640 59706 -23630
rect 58816 -23890 58896 -23640
rect 59536 -23690 59616 -23680
rect 59276 -23730 59356 -23720
rect 59276 -23790 59286 -23730
rect 59346 -23790 59356 -23730
rect 59536 -23750 59546 -23690
rect 59606 -23750 59616 -23690
rect 59536 -23770 59616 -23750
rect 58996 -23800 59076 -23790
rect 58996 -23860 59006 -23800
rect 59076 -23820 59086 -23800
rect 59536 -23810 59616 -23800
rect 59536 -23820 59546 -23810
rect 59076 -23860 59546 -23820
rect 58996 -23870 59076 -23860
rect 59536 -23870 59546 -23860
rect 59606 -23870 59616 -23810
rect 59536 -23880 59616 -23870
rect 58396 -23910 58896 -23890
rect 59646 -23910 59706 -23640
rect 60436 -23720 60536 -23710
rect 59856 -23740 59976 -23730
rect 59856 -23830 59866 -23740
rect 59966 -23830 59976 -23740
rect 60436 -23820 60446 -23720
rect 60526 -23820 60536 -23720
rect 60436 -23830 60536 -23820
rect 59856 -23840 59976 -23830
rect 58396 -23920 59706 -23910
rect 58396 -23930 59216 -23920
rect 58396 -23990 58906 -23930
rect 58966 -23980 59216 -23930
rect 59276 -23980 59336 -23920
rect 59396 -23980 59436 -23920
rect 59496 -23930 59706 -23920
rect 59496 -23980 59636 -23930
rect 58966 -23990 59636 -23980
rect 59696 -23990 59706 -23930
rect 58396 -24000 59706 -23990
rect 60036 -23920 60136 -23910
rect 60036 -24000 60046 -23920
rect 60126 -24000 60136 -23920
rect 55510 -24018 55520 -24008
rect 59646 -24010 59706 -24000
rect 60546 -24010 60636 -24000
rect 59066 -24040 59176 -24030
rect 59066 -24110 59076 -24040
rect 59166 -24110 59176 -24040
rect 59846 -24080 59856 -24010
rect 59916 -24030 59926 -24010
rect 60356 -24020 60556 -24010
rect 60356 -24030 60376 -24020
rect 59916 -24060 60376 -24030
rect 59916 -24080 59926 -24060
rect 60356 -24080 60376 -24060
rect 60446 -24080 60556 -24020
rect 60356 -24090 60556 -24080
rect 60626 -24090 60636 -24010
rect 59066 -24120 59176 -24110
rect 59966 -24100 60326 -24090
rect 53850 -24238 53860 -24128
rect 53920 -24138 55600 -24128
rect 53920 -24238 55000 -24138
rect 55090 -24238 55540 -24138
rect 55630 -24238 55640 -24138
rect 59966 -24160 59976 -24100
rect 60316 -24160 60326 -24100
rect 60546 -24110 60636 -24090
rect 61186 -24120 61366 -24110
rect 54770 -24438 54850 -24238
rect 56470 -24248 56480 -24188
rect 56550 -24248 56560 -24188
rect 57088 -24304 57098 -24164
rect 57368 -24304 57378 -24164
rect 59166 -24230 59376 -24220
rect 59166 -24240 59286 -24230
rect 59166 -24320 59176 -24240
rect 59236 -24320 59286 -24240
rect 59366 -24320 59376 -24230
rect 59166 -24330 59376 -24320
rect 59526 -24270 59646 -24250
rect 59526 -24330 59576 -24270
rect 59636 -24330 59646 -24270
rect 61186 -24300 61206 -24120
rect 61346 -24300 61366 -24120
rect 61186 -24310 61366 -24300
rect 59526 -24360 59646 -24330
rect 60286 -24350 60476 -24340
rect 59906 -24380 60016 -24370
rect 59806 -24390 59866 -24380
rect 54760 -24528 54770 -24438
rect 54840 -24528 54850 -24438
rect 59166 -24440 59536 -24430
rect 59166 -24520 59176 -24440
rect 59236 -24520 59286 -24440
rect 54920 -24538 55210 -24528
rect 54920 -24608 55140 -24538
rect 55200 -24608 55210 -24538
rect 59166 -24530 59286 -24520
rect 59356 -24450 59536 -24440
rect 59356 -24520 59476 -24450
rect 59356 -24530 59536 -24520
rect 59166 -24540 59536 -24530
rect 59566 -24560 59576 -24390
rect 59636 -24400 59866 -24390
rect 59636 -24540 59806 -24400
rect 59636 -24560 59866 -24540
rect 59906 -24560 59916 -24380
rect 60006 -24560 60016 -24380
rect 60286 -24490 60306 -24350
rect 60456 -24490 60476 -24350
rect 60286 -24500 60476 -24490
rect 61026 -24420 61136 -24410
rect 61026 -24530 61036 -24420
rect 61126 -24530 61136 -24420
rect 61026 -24540 61136 -24530
rect 59566 -24570 59636 -24560
rect 59906 -24570 60016 -24560
rect 54760 -24928 54770 -24848
rect 54840 -24928 54850 -24848
rect 54770 -25138 54850 -24928
rect 54920 -24998 54980 -24608
rect 55880 -24638 56900 -24618
rect 55010 -24728 55020 -24648
rect 55120 -24728 55740 -24648
rect 55810 -24728 55820 -24648
rect 55870 -24728 55880 -24638
rect 55970 -24728 56480 -24638
rect 56550 -24728 56900 -24638
rect 55880 -24748 56900 -24728
rect 57020 -24620 57040 -24618
rect 57800 -24620 58240 -24610
rect 57020 -24740 57800 -24620
rect 57020 -24748 57040 -24740
rect 57800 -24750 58240 -24740
rect 58516 -24660 58796 -24590
rect 58516 -24860 58556 -24660
rect 58756 -24860 58796 -24660
rect 59066 -24610 59936 -24600
rect 59066 -24680 59076 -24610
rect 59166 -24630 59826 -24610
rect 59166 -24680 59316 -24630
rect 59066 -24690 59316 -24680
rect 59376 -24680 59826 -24630
rect 59916 -24680 59936 -24610
rect 59376 -24690 59936 -24680
rect 60076 -24680 60196 -24640
rect 59066 -24770 59936 -24760
rect 59066 -24840 59076 -24770
rect 59166 -24840 59206 -24770
rect 59266 -24840 59826 -24770
rect 59926 -24840 59936 -24770
rect 59066 -24850 59936 -24840
rect 60076 -24840 60096 -24680
rect 60176 -24840 60196 -24680
rect 58516 -24940 58796 -24860
rect 60076 -24880 60196 -24840
rect 61266 -24650 61366 -24640
rect 61266 -24860 61276 -24650
rect 61356 -24860 61366 -24650
rect 61266 -24870 61366 -24860
rect 59586 -24890 59656 -24880
rect 59796 -24890 59866 -24880
rect 59586 -24910 59796 -24890
rect 59156 -24920 59536 -24910
rect 59156 -24930 59266 -24920
rect 54910 -25068 54920 -24998
rect 54980 -25068 54990 -24998
rect 59156 -25010 59166 -24930
rect 59226 -25010 59266 -24930
rect 59366 -24930 59536 -24920
rect 59366 -25010 59466 -24930
rect 59526 -25010 59536 -24930
rect 59156 -25030 59536 -25010
rect 59646 -25050 59796 -24910
rect 59586 -25070 59796 -25050
rect 59856 -25070 59866 -24890
rect 53840 -25248 53850 -25138
rect 53920 -25238 55000 -25138
rect 55090 -25238 55540 -25138
rect 55630 -25238 55640 -25138
rect 56470 -25188 56480 -25128
rect 56550 -25188 56560 -25128
rect 57088 -25214 57098 -25074
rect 57368 -25214 57378 -25074
rect 59796 -25080 59866 -25070
rect 59906 -24890 60016 -24880
rect 59906 -25080 59916 -24890
rect 60006 -25080 60016 -24890
rect 60476 -24910 60546 -24900
rect 60536 -24970 60546 -24910
rect 60476 -24980 60546 -24970
rect 60966 -25030 61486 -25020
rect 60966 -25040 61336 -25030
rect 59906 -25090 60016 -25080
rect 60466 -25050 61336 -25040
rect 59506 -25110 59606 -25100
rect 59156 -25160 59376 -25140
rect 53920 -25248 55640 -25238
rect 59156 -25240 59166 -25160
rect 59226 -25240 59266 -25160
rect 59156 -25250 59266 -25240
rect 59366 -25250 59376 -25160
rect 59506 -25180 59516 -25110
rect 59596 -25180 59606 -25110
rect 60466 -25110 60476 -25050
rect 60536 -25110 60616 -25050
rect 60736 -25110 60756 -25050
rect 60816 -25110 60896 -25050
rect 60956 -25110 61336 -25050
rect 60466 -25120 61336 -25110
rect 60966 -25160 61336 -25120
rect 61456 -25160 61486 -25030
rect 60966 -25170 61486 -25160
rect 59506 -25190 59606 -25180
rect 59156 -25260 59376 -25250
rect 59306 -25320 60336 -25300
rect 59066 -25340 59176 -25330
rect 55210 -25518 55220 -25348
rect 55310 -25518 55320 -25348
rect 55400 -25528 55410 -25358
rect 55500 -25368 55510 -25358
rect 55500 -25488 56380 -25368
rect 56440 -25488 56450 -25368
rect 59066 -25400 59076 -25340
rect 59166 -25400 59176 -25340
rect 59306 -25380 59316 -25320
rect 59376 -25340 59966 -25320
rect 59376 -25380 59816 -25340
rect 59306 -25390 59816 -25380
rect 59846 -25380 59916 -25370
rect 59066 -25410 59176 -25400
rect 59846 -25440 59856 -25380
rect 59946 -25380 59966 -25340
rect 60326 -25380 60336 -25320
rect 59946 -25390 60336 -25380
rect 60366 -25340 61146 -25330
rect 60366 -25380 61056 -25340
rect 59646 -25450 59716 -25440
rect 59846 -25450 59916 -25440
rect 60366 -25440 60376 -25380
rect 60436 -25440 61056 -25380
rect 61126 -25440 61146 -25340
rect 55500 -25508 56450 -25488
rect 58396 -25460 59716 -25450
rect 55500 -25528 55510 -25508
rect 58396 -25530 58926 -25460
rect 58986 -25530 59146 -25460
rect 59226 -25530 59276 -25460
rect 59356 -25530 59396 -25460
rect 59476 -25520 59646 -25460
rect 59706 -25520 59716 -25460
rect 60366 -25470 61146 -25440
rect 59476 -25530 59716 -25520
rect 58396 -25540 59716 -25530
rect 54900 -25608 54910 -25598
rect 53940 -25688 53950 -25608
rect 54010 -25688 54910 -25608
rect 53940 -25698 54910 -25688
rect 54980 -25618 54990 -25598
rect 54980 -25678 55980 -25618
rect 54980 -25698 55880 -25678
rect 53940 -25718 55880 -25698
rect 53500 -25848 53510 -25728
rect 53630 -25848 53640 -25728
rect 55850 -25758 55880 -25718
rect 55970 -25758 55980 -25678
rect 55230 -25818 55240 -25758
rect 55370 -25778 55710 -25758
rect 55370 -25788 55720 -25778
rect 55370 -25808 55620 -25788
rect 55370 -25818 55380 -25808
rect 55400 -25868 55410 -25848
rect 54730 -25958 54740 -25868
rect 54850 -25938 55410 -25868
rect 55510 -25938 55520 -25848
rect 55600 -25878 55620 -25808
rect 55710 -25878 55720 -25788
rect 54850 -25958 55520 -25938
rect 55210 -26128 55220 -26018
rect 55330 -26128 55340 -26018
rect 55850 -26178 55980 -25758
rect 56010 -26008 56020 -25858
rect 56080 -26008 56090 -25858
rect 56160 -26008 56170 -25808
rect 56390 -26008 56400 -25808
rect 58396 -25820 58896 -25540
rect 59006 -25700 59076 -25680
rect 59246 -25690 59256 -25630
rect 59366 -25690 59376 -25630
rect 59536 -25660 59546 -25590
rect 59606 -25660 59616 -25590
rect 59536 -25670 59616 -25660
rect 59006 -25760 59016 -25700
rect 59536 -25710 59616 -25700
rect 59076 -25720 59086 -25710
rect 59536 -25720 59546 -25710
rect 59076 -25760 59546 -25720
rect 59006 -25770 59546 -25760
rect 59606 -25770 59616 -25710
rect 59006 -25790 59076 -25770
rect 59536 -25790 59616 -25770
rect 59646 -25820 59716 -25540
rect 59796 -25610 59926 -25600
rect 59796 -25720 59806 -25610
rect 59916 -25720 59926 -25610
rect 59796 -25730 59926 -25720
rect 60436 -25630 60536 -25610
rect 60436 -25750 60446 -25630
rect 60526 -25750 60536 -25630
rect 60436 -25760 60536 -25750
rect 58396 -25830 59716 -25820
rect 56654 -25868 56998 -25858
rect 55520 -26268 55530 -26178
rect 55610 -26268 55980 -26178
rect 54130 -26548 54140 -26288
rect 54850 -26548 54860 -26288
rect 55310 -26468 55320 -26328
rect 55470 -26468 55480 -26328
rect 56170 -26538 56390 -26008
rect 58396 -25900 58906 -25830
rect 58986 -25900 59146 -25830
rect 59226 -25900 59276 -25830
rect 59356 -25900 59396 -25830
rect 59476 -25840 59716 -25830
rect 59476 -25900 59646 -25840
rect 59706 -25900 59716 -25840
rect 58396 -25910 59716 -25900
rect 58396 -25950 58896 -25910
rect 59646 -25920 59716 -25910
rect 56654 -26096 56998 -26086
rect 59006 -26000 60416 -25990
rect 59006 -26040 60266 -26000
rect 59006 -26110 59016 -26040
rect 59076 -26110 59546 -26040
rect 59606 -26110 60266 -26040
rect 59006 -26130 60266 -26110
rect 60406 -26130 60416 -26000
rect 59006 -26140 60416 -26130
rect 59986 -26190 60116 -26180
rect 58956 -26200 59156 -26190
rect 58956 -26380 58966 -26200
rect 59146 -26380 59156 -26200
rect 59986 -26300 59996 -26190
rect 60106 -26300 60116 -26190
rect 58956 -26390 59156 -26380
rect 55680 -26548 56390 -26538
rect 54130 -26708 56390 -26548
rect 55680 -26718 56390 -26708
rect 59600 -26400 60500 -26300
rect 59600 -26800 59700 -26400
rect 60400 -26800 60500 -26400
rect 55400 -26900 56200 -26800
rect 59600 -26900 60500 -26800
rect 63600 -26400 64200 -26300
rect 63600 -26800 63700 -26400
rect 64100 -26800 64200 -26400
rect 55400 -27300 55500 -26900
rect 56100 -27300 56200 -26900
rect 55400 -27400 56200 -27300
rect 51400 -28100 51500 -27900
rect 52500 -28100 52600 -27900
rect 51400 -33300 52600 -28100
rect 55440 -27880 55740 -27860
rect 55440 -28160 55460 -27880
rect 55720 -28160 55740 -27880
rect 55440 -28180 55740 -28160
rect 54140 -28338 56390 -28328
rect 53460 -28540 53800 -28520
rect 53460 -28740 53480 -28540
rect 53780 -28740 53800 -28540
rect 54140 -28578 54150 -28338
rect 54860 -28578 56390 -28338
rect 58946 -28470 59146 -28450
rect 54140 -28588 56390 -28578
rect 53460 -28760 53800 -28740
rect 54850 -28818 55530 -28808
rect 53510 -28968 53520 -28858
rect 53640 -28968 53650 -28858
rect 54740 -28918 54750 -28838
rect 54850 -28888 55430 -28818
rect 55520 -28888 55530 -28818
rect 55950 -28888 55960 -28738
rect 56040 -28888 56050 -28738
rect 56170 -28758 56390 -28588
rect 56506 -28580 57016 -28570
rect 54840 -28918 54850 -28908
rect 55270 -29008 55280 -28918
rect 55400 -29008 55410 -28918
rect 56170 -28968 56190 -28758
rect 56390 -28968 56400 -28758
rect 58946 -28630 58966 -28470
rect 59126 -28630 59146 -28470
rect 58946 -28650 59146 -28630
rect 59316 -28500 60176 -28490
rect 59316 -28510 59956 -28500
rect 59316 -28650 59336 -28510
rect 59416 -28650 59956 -28510
rect 59316 -28660 59956 -28650
rect 60166 -28660 60176 -28500
rect 59316 -28670 60176 -28660
rect 56506 -28840 57016 -28830
rect 58956 -28720 61136 -28710
rect 58956 -28730 61056 -28720
rect 58956 -28840 58996 -28730
rect 59106 -28740 61056 -28730
rect 59106 -28840 59516 -28740
rect 59616 -28840 61056 -28740
rect 58396 -28930 58896 -28840
rect 58956 -28850 61056 -28840
rect 61126 -28850 61136 -28720
rect 58956 -28860 61136 -28850
rect 55850 -29048 55880 -29018
rect 53940 -29078 55880 -29048
rect 53940 -29098 54920 -29078
rect 53040 -30908 53050 -29158
rect 53250 -30908 53260 -29158
rect 53940 -29198 53950 -29098
rect 54020 -29148 54920 -29098
rect 54020 -29198 54030 -29148
rect 54910 -29168 54920 -29148
rect 54990 -29098 55880 -29078
rect 55970 -29048 55980 -29018
rect 54990 -29148 55970 -29098
rect 54990 -29168 55000 -29148
rect 55220 -29428 55230 -29258
rect 55320 -29428 55330 -29258
rect 55420 -29418 55430 -29248
rect 55510 -29258 55520 -29248
rect 55510 -29268 56670 -29258
rect 55510 -29398 55600 -29268
rect 55710 -29398 56590 -29268
rect 56660 -29398 56670 -29268
rect 55510 -29408 56670 -29398
rect 58396 -29290 58486 -28930
rect 58816 -28950 58896 -28930
rect 59646 -28950 59706 -28930
rect 58816 -28970 59706 -28950
rect 58816 -29030 58906 -28970
rect 58966 -29030 59216 -28970
rect 59276 -29030 59326 -28970
rect 59386 -29030 59436 -28970
rect 59496 -29030 59636 -28970
rect 59696 -29030 59706 -28970
rect 58816 -29040 59706 -29030
rect 58816 -29290 58896 -29040
rect 59536 -29090 59616 -29080
rect 59276 -29130 59356 -29120
rect 59276 -29190 59286 -29130
rect 59346 -29190 59356 -29130
rect 59536 -29150 59546 -29090
rect 59606 -29150 59616 -29090
rect 59536 -29170 59616 -29150
rect 58996 -29200 59076 -29190
rect 58996 -29260 59006 -29200
rect 59076 -29220 59086 -29200
rect 59536 -29210 59616 -29200
rect 59536 -29220 59546 -29210
rect 59076 -29260 59546 -29220
rect 58996 -29270 59076 -29260
rect 59536 -29270 59546 -29260
rect 59606 -29270 59616 -29210
rect 59536 -29280 59616 -29270
rect 58396 -29310 58896 -29290
rect 59646 -29310 59706 -29040
rect 60436 -29120 60536 -29110
rect 59856 -29140 59976 -29130
rect 59856 -29230 59866 -29140
rect 59966 -29230 59976 -29140
rect 60436 -29220 60446 -29120
rect 60526 -29220 60536 -29120
rect 60436 -29230 60536 -29220
rect 59856 -29240 59976 -29230
rect 58396 -29320 59706 -29310
rect 58396 -29330 59216 -29320
rect 58396 -29390 58906 -29330
rect 58966 -29380 59216 -29330
rect 59276 -29380 59336 -29320
rect 59396 -29380 59436 -29320
rect 59496 -29330 59706 -29320
rect 59496 -29380 59636 -29330
rect 58966 -29390 59636 -29380
rect 59696 -29390 59706 -29330
rect 58396 -29400 59706 -29390
rect 60036 -29320 60136 -29310
rect 60036 -29400 60046 -29320
rect 60126 -29400 60136 -29320
rect 55510 -29418 55520 -29408
rect 59646 -29410 59706 -29400
rect 60546 -29410 60636 -29400
rect 59066 -29440 59176 -29430
rect 59066 -29510 59076 -29440
rect 59166 -29510 59176 -29440
rect 59846 -29480 59856 -29410
rect 59916 -29430 59926 -29410
rect 60356 -29420 60556 -29410
rect 60356 -29430 60376 -29420
rect 59916 -29460 60376 -29430
rect 59916 -29480 59926 -29460
rect 60356 -29480 60376 -29460
rect 60446 -29480 60556 -29420
rect 60356 -29490 60556 -29480
rect 60626 -29490 60636 -29410
rect 59066 -29520 59176 -29510
rect 59966 -29500 60326 -29490
rect 53850 -29638 53860 -29528
rect 53920 -29538 55600 -29528
rect 53920 -29638 55000 -29538
rect 55090 -29638 55540 -29538
rect 55630 -29638 55640 -29538
rect 59966 -29560 59976 -29500
rect 60316 -29560 60326 -29500
rect 60546 -29510 60636 -29490
rect 61186 -29520 61366 -29510
rect 54770 -29838 54850 -29638
rect 56470 -29648 56480 -29588
rect 56550 -29648 56560 -29588
rect 57088 -29704 57098 -29564
rect 57368 -29704 57378 -29564
rect 59166 -29630 59376 -29620
rect 59166 -29640 59286 -29630
rect 59166 -29720 59176 -29640
rect 59236 -29720 59286 -29640
rect 59366 -29720 59376 -29630
rect 59166 -29730 59376 -29720
rect 59526 -29670 59646 -29650
rect 59526 -29730 59576 -29670
rect 59636 -29730 59646 -29670
rect 61186 -29700 61206 -29520
rect 61346 -29700 61366 -29520
rect 61186 -29710 61366 -29700
rect 59526 -29760 59646 -29730
rect 60286 -29750 60476 -29740
rect 59906 -29780 60016 -29770
rect 59806 -29790 59866 -29780
rect 54760 -29928 54770 -29838
rect 54840 -29928 54850 -29838
rect 59166 -29840 59536 -29830
rect 59166 -29920 59176 -29840
rect 59236 -29920 59286 -29840
rect 54920 -29938 55210 -29928
rect 54920 -30008 55140 -29938
rect 55200 -30008 55210 -29938
rect 59166 -29930 59286 -29920
rect 59356 -29850 59536 -29840
rect 59356 -29920 59476 -29850
rect 59356 -29930 59536 -29920
rect 59166 -29940 59536 -29930
rect 59566 -29960 59576 -29790
rect 59636 -29800 59866 -29790
rect 59636 -29940 59806 -29800
rect 59636 -29960 59866 -29940
rect 59906 -29960 59916 -29780
rect 60006 -29960 60016 -29780
rect 60286 -29890 60306 -29750
rect 60456 -29890 60476 -29750
rect 60286 -29900 60476 -29890
rect 61026 -29820 61136 -29810
rect 61026 -29930 61036 -29820
rect 61126 -29930 61136 -29820
rect 61026 -29940 61136 -29930
rect 59566 -29970 59636 -29960
rect 59906 -29970 60016 -29960
rect 54760 -30328 54770 -30248
rect 54840 -30328 54850 -30248
rect 54770 -30538 54850 -30328
rect 54920 -30398 54980 -30008
rect 55880 -30038 56900 -30018
rect 55010 -30128 55020 -30048
rect 55120 -30128 55740 -30048
rect 55810 -30128 55820 -30048
rect 55870 -30128 55880 -30038
rect 55970 -30128 56480 -30038
rect 56550 -30128 56900 -30038
rect 55880 -30148 56900 -30128
rect 57020 -30020 57040 -30018
rect 57800 -30020 58240 -30010
rect 57020 -30140 57800 -30020
rect 57020 -30148 57040 -30140
rect 57800 -30150 58240 -30140
rect 58516 -30060 58796 -29990
rect 58516 -30260 58556 -30060
rect 58756 -30260 58796 -30060
rect 59066 -30010 59936 -30000
rect 59066 -30080 59076 -30010
rect 59166 -30030 59826 -30010
rect 59166 -30080 59316 -30030
rect 59066 -30090 59316 -30080
rect 59376 -30080 59826 -30030
rect 59916 -30080 59936 -30010
rect 59376 -30090 59936 -30080
rect 60076 -30080 60196 -30040
rect 59066 -30170 59936 -30160
rect 59066 -30240 59076 -30170
rect 59166 -30240 59206 -30170
rect 59266 -30240 59826 -30170
rect 59926 -30240 59936 -30170
rect 59066 -30250 59936 -30240
rect 60076 -30240 60096 -30080
rect 60176 -30240 60196 -30080
rect 58516 -30340 58796 -30260
rect 60076 -30280 60196 -30240
rect 61266 -30050 61366 -30040
rect 61266 -30260 61276 -30050
rect 61356 -30260 61366 -30050
rect 61266 -30270 61366 -30260
rect 59586 -30290 59656 -30280
rect 59796 -30290 59866 -30280
rect 59586 -30310 59796 -30290
rect 59156 -30320 59536 -30310
rect 59156 -30330 59266 -30320
rect 54910 -30468 54920 -30398
rect 54980 -30468 54990 -30398
rect 59156 -30410 59166 -30330
rect 59226 -30410 59266 -30330
rect 59366 -30330 59536 -30320
rect 59366 -30410 59466 -30330
rect 59526 -30410 59536 -30330
rect 59156 -30430 59536 -30410
rect 59646 -30450 59796 -30310
rect 59586 -30470 59796 -30450
rect 59856 -30470 59866 -30290
rect 53840 -30648 53850 -30538
rect 53920 -30638 55000 -30538
rect 55090 -30638 55540 -30538
rect 55630 -30638 55640 -30538
rect 56470 -30588 56480 -30528
rect 56550 -30588 56560 -30528
rect 57088 -30614 57098 -30474
rect 57368 -30614 57378 -30474
rect 59796 -30480 59866 -30470
rect 59906 -30290 60016 -30280
rect 59906 -30480 59916 -30290
rect 60006 -30480 60016 -30290
rect 60476 -30310 60546 -30300
rect 60536 -30370 60546 -30310
rect 60476 -30380 60546 -30370
rect 60966 -30430 61486 -30420
rect 60966 -30440 61336 -30430
rect 59906 -30490 60016 -30480
rect 60466 -30450 61336 -30440
rect 59506 -30510 59606 -30500
rect 59156 -30560 59376 -30540
rect 53920 -30648 55640 -30638
rect 59156 -30640 59166 -30560
rect 59226 -30640 59266 -30560
rect 59156 -30650 59266 -30640
rect 59366 -30650 59376 -30560
rect 59506 -30580 59516 -30510
rect 59596 -30580 59606 -30510
rect 60466 -30510 60476 -30450
rect 60536 -30510 60616 -30450
rect 60736 -30510 60756 -30450
rect 60816 -30510 60896 -30450
rect 60956 -30510 61336 -30450
rect 60466 -30520 61336 -30510
rect 60966 -30560 61336 -30520
rect 61456 -30560 61486 -30430
rect 60966 -30570 61486 -30560
rect 59506 -30590 59606 -30580
rect 59156 -30660 59376 -30650
rect 59306 -30720 60336 -30700
rect 59066 -30740 59176 -30730
rect 55210 -30918 55220 -30748
rect 55310 -30918 55320 -30748
rect 55400 -30928 55410 -30758
rect 55500 -30768 55510 -30758
rect 55500 -30888 56380 -30768
rect 56440 -30888 56450 -30768
rect 59066 -30800 59076 -30740
rect 59166 -30800 59176 -30740
rect 59306 -30780 59316 -30720
rect 59376 -30740 59966 -30720
rect 59376 -30780 59816 -30740
rect 59306 -30790 59816 -30780
rect 59846 -30780 59916 -30770
rect 59066 -30810 59176 -30800
rect 59846 -30840 59856 -30780
rect 59946 -30780 59966 -30740
rect 60326 -30780 60336 -30720
rect 59946 -30790 60336 -30780
rect 60366 -30740 61146 -30730
rect 60366 -30780 61056 -30740
rect 59646 -30850 59716 -30840
rect 59846 -30850 59916 -30840
rect 60366 -30840 60376 -30780
rect 60436 -30840 61056 -30780
rect 61126 -30840 61146 -30740
rect 55500 -30908 56450 -30888
rect 58396 -30860 59716 -30850
rect 55500 -30928 55510 -30908
rect 58396 -30930 58926 -30860
rect 58986 -30930 59146 -30860
rect 59226 -30930 59276 -30860
rect 59356 -30930 59396 -30860
rect 59476 -30920 59646 -30860
rect 59706 -30920 59716 -30860
rect 60366 -30870 61146 -30840
rect 59476 -30930 59716 -30920
rect 58396 -30940 59716 -30930
rect 54900 -31008 54910 -30998
rect 53940 -31088 53950 -31008
rect 54010 -31088 54910 -31008
rect 53940 -31098 54910 -31088
rect 54980 -31018 54990 -30998
rect 54980 -31078 55980 -31018
rect 54980 -31098 55880 -31078
rect 53940 -31118 55880 -31098
rect 53500 -31248 53510 -31128
rect 53630 -31248 53640 -31128
rect 55850 -31158 55880 -31118
rect 55970 -31158 55980 -31078
rect 55230 -31218 55240 -31158
rect 55370 -31178 55710 -31158
rect 55370 -31188 55720 -31178
rect 55370 -31208 55620 -31188
rect 55370 -31218 55380 -31208
rect 55400 -31268 55410 -31248
rect 54730 -31358 54740 -31268
rect 54850 -31338 55410 -31268
rect 55510 -31338 55520 -31248
rect 55600 -31278 55620 -31208
rect 55710 -31278 55720 -31188
rect 54850 -31358 55520 -31338
rect 55210 -31528 55220 -31418
rect 55330 -31528 55340 -31418
rect 55850 -31578 55980 -31158
rect 56010 -31408 56020 -31258
rect 56080 -31408 56090 -31258
rect 56160 -31408 56170 -31208
rect 56390 -31408 56400 -31208
rect 58396 -31220 58896 -30940
rect 59006 -31100 59076 -31080
rect 59246 -31090 59256 -31030
rect 59366 -31090 59376 -31030
rect 59536 -31060 59546 -30990
rect 59606 -31060 59616 -30990
rect 59536 -31070 59616 -31060
rect 59006 -31160 59016 -31100
rect 59536 -31110 59616 -31100
rect 59076 -31120 59086 -31110
rect 59536 -31120 59546 -31110
rect 59076 -31160 59546 -31120
rect 59006 -31170 59546 -31160
rect 59606 -31170 59616 -31110
rect 59006 -31190 59076 -31170
rect 59536 -31190 59616 -31170
rect 59646 -31220 59716 -30940
rect 59796 -31010 59926 -31000
rect 59796 -31120 59806 -31010
rect 59916 -31120 59926 -31010
rect 59796 -31130 59926 -31120
rect 60436 -31030 60536 -31010
rect 60436 -31150 60446 -31030
rect 60526 -31150 60536 -31030
rect 60436 -31160 60536 -31150
rect 58396 -31230 59716 -31220
rect 56654 -31268 56998 -31258
rect 55520 -31668 55530 -31578
rect 55610 -31668 55980 -31578
rect 54130 -31948 54140 -31688
rect 54850 -31948 54860 -31688
rect 55310 -31868 55320 -31728
rect 55470 -31868 55480 -31728
rect 56170 -31938 56390 -31408
rect 58396 -31300 58906 -31230
rect 58986 -31300 59146 -31230
rect 59226 -31300 59276 -31230
rect 59356 -31300 59396 -31230
rect 59476 -31240 59716 -31230
rect 59476 -31300 59646 -31240
rect 59706 -31300 59716 -31240
rect 58396 -31310 59716 -31300
rect 58396 -31350 58896 -31310
rect 59646 -31320 59716 -31310
rect 56654 -31496 56998 -31486
rect 59006 -31400 60416 -31390
rect 59006 -31440 60266 -31400
rect 59006 -31510 59016 -31440
rect 59076 -31510 59546 -31440
rect 59606 -31510 60266 -31440
rect 59006 -31530 60266 -31510
rect 60406 -31530 60416 -31400
rect 59006 -31540 60416 -31530
rect 59986 -31590 60116 -31580
rect 58956 -31600 59156 -31590
rect 58956 -31780 58966 -31600
rect 59146 -31780 59156 -31600
rect 59986 -31700 59996 -31590
rect 60106 -31700 60116 -31590
rect 58956 -31790 59156 -31780
rect 55680 -31948 56390 -31938
rect 54130 -32108 56390 -31948
rect 55680 -32118 56390 -32108
rect 59700 -31800 60400 -31700
rect 59700 -32100 59800 -31800
rect 60300 -32100 60400 -31800
rect 59700 -32200 60400 -32100
rect 62800 -31800 63400 -31700
rect 62800 -32100 62900 -31800
rect 63300 -32100 63400 -31800
rect 55400 -32300 56200 -32200
rect 55400 -32700 55500 -32300
rect 56100 -32700 56200 -32300
rect 55400 -32800 56200 -32700
rect 51400 -33500 51500 -33300
rect 52500 -33500 52600 -33300
rect 51400 -38700 52600 -33500
rect 55440 -33280 55740 -33260
rect 55440 -33560 55460 -33280
rect 55720 -33560 55740 -33280
rect 55440 -33580 55740 -33560
rect 54140 -33738 56390 -33728
rect 53460 -33940 53800 -33920
rect 53460 -34140 53480 -33940
rect 53780 -34140 53800 -33940
rect 54140 -33978 54150 -33738
rect 54860 -33978 56390 -33738
rect 58946 -33870 59146 -33850
rect 54140 -33988 56390 -33978
rect 53460 -34160 53800 -34140
rect 54850 -34218 55530 -34208
rect 53510 -34368 53520 -34258
rect 53640 -34368 53650 -34258
rect 54740 -34318 54750 -34238
rect 54850 -34288 55430 -34218
rect 55520 -34288 55530 -34218
rect 55950 -34288 55960 -34138
rect 56040 -34288 56050 -34138
rect 56170 -34158 56390 -33988
rect 56506 -33980 57016 -33970
rect 54840 -34318 54850 -34308
rect 55270 -34408 55280 -34318
rect 55400 -34408 55410 -34318
rect 56170 -34368 56190 -34158
rect 56390 -34368 56400 -34158
rect 58946 -34030 58966 -33870
rect 59126 -34030 59146 -33870
rect 58946 -34050 59146 -34030
rect 59316 -33900 60176 -33890
rect 59316 -33910 59956 -33900
rect 59316 -34050 59336 -33910
rect 59416 -34050 59956 -33910
rect 59316 -34060 59956 -34050
rect 60166 -34060 60176 -33900
rect 59316 -34070 60176 -34060
rect 56506 -34240 57016 -34230
rect 58956 -34120 61136 -34110
rect 58956 -34130 61056 -34120
rect 58956 -34240 58996 -34130
rect 59106 -34140 61056 -34130
rect 59106 -34240 59516 -34140
rect 59616 -34240 61056 -34140
rect 58396 -34330 58896 -34240
rect 58956 -34250 61056 -34240
rect 61126 -34250 61136 -34120
rect 58956 -34260 61136 -34250
rect 55850 -34448 55880 -34418
rect 53940 -34478 55880 -34448
rect 53940 -34498 54920 -34478
rect 53040 -36308 53050 -34558
rect 53250 -36308 53260 -34558
rect 53940 -34598 53950 -34498
rect 54020 -34548 54920 -34498
rect 54020 -34598 54030 -34548
rect 54910 -34568 54920 -34548
rect 54990 -34498 55880 -34478
rect 55970 -34448 55980 -34418
rect 54990 -34548 55970 -34498
rect 54990 -34568 55000 -34548
rect 55220 -34828 55230 -34658
rect 55320 -34828 55330 -34658
rect 55420 -34818 55430 -34648
rect 55510 -34658 55520 -34648
rect 55510 -34668 56670 -34658
rect 55510 -34798 55600 -34668
rect 55710 -34798 56590 -34668
rect 56660 -34798 56670 -34668
rect 55510 -34808 56670 -34798
rect 58396 -34690 58486 -34330
rect 58816 -34350 58896 -34330
rect 59646 -34350 59706 -34330
rect 58816 -34370 59706 -34350
rect 58816 -34430 58906 -34370
rect 58966 -34430 59216 -34370
rect 59276 -34430 59326 -34370
rect 59386 -34430 59436 -34370
rect 59496 -34430 59636 -34370
rect 59696 -34430 59706 -34370
rect 58816 -34440 59706 -34430
rect 58816 -34690 58896 -34440
rect 59536 -34490 59616 -34480
rect 59276 -34530 59356 -34520
rect 59276 -34590 59286 -34530
rect 59346 -34590 59356 -34530
rect 59536 -34550 59546 -34490
rect 59606 -34550 59616 -34490
rect 59536 -34570 59616 -34550
rect 58996 -34600 59076 -34590
rect 58996 -34660 59006 -34600
rect 59076 -34620 59086 -34600
rect 59536 -34610 59616 -34600
rect 59536 -34620 59546 -34610
rect 59076 -34660 59546 -34620
rect 58996 -34670 59076 -34660
rect 59536 -34670 59546 -34660
rect 59606 -34670 59616 -34610
rect 59536 -34680 59616 -34670
rect 58396 -34710 58896 -34690
rect 59646 -34710 59706 -34440
rect 60436 -34520 60536 -34510
rect 59856 -34540 59976 -34530
rect 59856 -34630 59866 -34540
rect 59966 -34630 59976 -34540
rect 60436 -34620 60446 -34520
rect 60526 -34620 60536 -34520
rect 60436 -34630 60536 -34620
rect 59856 -34640 59976 -34630
rect 58396 -34720 59706 -34710
rect 58396 -34730 59216 -34720
rect 58396 -34790 58906 -34730
rect 58966 -34780 59216 -34730
rect 59276 -34780 59336 -34720
rect 59396 -34780 59436 -34720
rect 59496 -34730 59706 -34720
rect 59496 -34780 59636 -34730
rect 58966 -34790 59636 -34780
rect 59696 -34790 59706 -34730
rect 58396 -34800 59706 -34790
rect 60036 -34720 60136 -34710
rect 60036 -34800 60046 -34720
rect 60126 -34800 60136 -34720
rect 55510 -34818 55520 -34808
rect 59646 -34810 59706 -34800
rect 60546 -34810 60636 -34800
rect 59066 -34840 59176 -34830
rect 59066 -34910 59076 -34840
rect 59166 -34910 59176 -34840
rect 59846 -34880 59856 -34810
rect 59916 -34830 59926 -34810
rect 60356 -34820 60556 -34810
rect 60356 -34830 60376 -34820
rect 59916 -34860 60376 -34830
rect 59916 -34880 59926 -34860
rect 60356 -34880 60376 -34860
rect 60446 -34880 60556 -34820
rect 60356 -34890 60556 -34880
rect 60626 -34890 60636 -34810
rect 59066 -34920 59176 -34910
rect 59966 -34900 60326 -34890
rect 53850 -35038 53860 -34928
rect 53920 -34938 55600 -34928
rect 53920 -35038 55000 -34938
rect 55090 -35038 55540 -34938
rect 55630 -35038 55640 -34938
rect 59966 -34960 59976 -34900
rect 60316 -34960 60326 -34900
rect 60546 -34910 60636 -34890
rect 61186 -34920 61366 -34910
rect 54770 -35238 54850 -35038
rect 56470 -35048 56480 -34988
rect 56550 -35048 56560 -34988
rect 57088 -35104 57098 -34964
rect 57368 -35104 57378 -34964
rect 59166 -35030 59376 -35020
rect 59166 -35040 59286 -35030
rect 59166 -35120 59176 -35040
rect 59236 -35120 59286 -35040
rect 59366 -35120 59376 -35030
rect 59166 -35130 59376 -35120
rect 59526 -35070 59646 -35050
rect 59526 -35130 59576 -35070
rect 59636 -35130 59646 -35070
rect 61186 -35100 61206 -34920
rect 61346 -35100 61366 -34920
rect 61186 -35110 61366 -35100
rect 59526 -35160 59646 -35130
rect 60286 -35150 60476 -35140
rect 59906 -35180 60016 -35170
rect 59806 -35190 59866 -35180
rect 54760 -35328 54770 -35238
rect 54840 -35328 54850 -35238
rect 59166 -35240 59536 -35230
rect 59166 -35320 59176 -35240
rect 59236 -35320 59286 -35240
rect 54920 -35338 55210 -35328
rect 54920 -35408 55140 -35338
rect 55200 -35408 55210 -35338
rect 59166 -35330 59286 -35320
rect 59356 -35250 59536 -35240
rect 59356 -35320 59476 -35250
rect 59356 -35330 59536 -35320
rect 59166 -35340 59536 -35330
rect 59566 -35360 59576 -35190
rect 59636 -35200 59866 -35190
rect 59636 -35340 59806 -35200
rect 59636 -35360 59866 -35340
rect 59906 -35360 59916 -35180
rect 60006 -35360 60016 -35180
rect 60286 -35290 60306 -35150
rect 60456 -35290 60476 -35150
rect 60286 -35300 60476 -35290
rect 61026 -35220 61136 -35210
rect 61026 -35330 61036 -35220
rect 61126 -35330 61136 -35220
rect 61026 -35340 61136 -35330
rect 59566 -35370 59636 -35360
rect 59906 -35370 60016 -35360
rect 54760 -35728 54770 -35648
rect 54840 -35728 54850 -35648
rect 54770 -35938 54850 -35728
rect 54920 -35798 54980 -35408
rect 55880 -35438 56900 -35418
rect 55010 -35528 55020 -35448
rect 55120 -35528 55740 -35448
rect 55810 -35528 55820 -35448
rect 55870 -35528 55880 -35438
rect 55970 -35528 56480 -35438
rect 56550 -35528 56900 -35438
rect 55880 -35548 56900 -35528
rect 57020 -35420 57040 -35418
rect 57800 -35420 58240 -35410
rect 57020 -35540 57800 -35420
rect 57020 -35548 57040 -35540
rect 57800 -35550 58240 -35540
rect 58516 -35460 58796 -35390
rect 58516 -35660 58556 -35460
rect 58756 -35660 58796 -35460
rect 59066 -35410 59936 -35400
rect 59066 -35480 59076 -35410
rect 59166 -35430 59826 -35410
rect 59166 -35480 59316 -35430
rect 59066 -35490 59316 -35480
rect 59376 -35480 59826 -35430
rect 59916 -35480 59936 -35410
rect 59376 -35490 59936 -35480
rect 60076 -35480 60196 -35440
rect 59066 -35570 59936 -35560
rect 59066 -35640 59076 -35570
rect 59166 -35640 59206 -35570
rect 59266 -35640 59826 -35570
rect 59926 -35640 59936 -35570
rect 59066 -35650 59936 -35640
rect 60076 -35640 60096 -35480
rect 60176 -35640 60196 -35480
rect 58516 -35740 58796 -35660
rect 60076 -35680 60196 -35640
rect 61266 -35450 61366 -35440
rect 61266 -35660 61276 -35450
rect 61356 -35660 61366 -35450
rect 61266 -35670 61366 -35660
rect 59586 -35690 59656 -35680
rect 59796 -35690 59866 -35680
rect 59586 -35710 59796 -35690
rect 59156 -35720 59536 -35710
rect 59156 -35730 59266 -35720
rect 54910 -35868 54920 -35798
rect 54980 -35868 54990 -35798
rect 59156 -35810 59166 -35730
rect 59226 -35810 59266 -35730
rect 59366 -35730 59536 -35720
rect 59366 -35810 59466 -35730
rect 59526 -35810 59536 -35730
rect 59156 -35830 59536 -35810
rect 59646 -35850 59796 -35710
rect 59586 -35870 59796 -35850
rect 59856 -35870 59866 -35690
rect 53840 -36048 53850 -35938
rect 53920 -36038 55000 -35938
rect 55090 -36038 55540 -35938
rect 55630 -36038 55640 -35938
rect 56470 -35988 56480 -35928
rect 56550 -35988 56560 -35928
rect 57088 -36014 57098 -35874
rect 57368 -36014 57378 -35874
rect 59796 -35880 59866 -35870
rect 59906 -35690 60016 -35680
rect 59906 -35880 59916 -35690
rect 60006 -35880 60016 -35690
rect 60476 -35710 60546 -35700
rect 60536 -35770 60546 -35710
rect 60476 -35780 60546 -35770
rect 60966 -35830 61486 -35820
rect 60966 -35840 61336 -35830
rect 59906 -35890 60016 -35880
rect 60466 -35850 61336 -35840
rect 59506 -35910 59606 -35900
rect 59156 -35960 59376 -35940
rect 53920 -36048 55640 -36038
rect 59156 -36040 59166 -35960
rect 59226 -36040 59266 -35960
rect 59156 -36050 59266 -36040
rect 59366 -36050 59376 -35960
rect 59506 -35980 59516 -35910
rect 59596 -35980 59606 -35910
rect 60466 -35910 60476 -35850
rect 60536 -35910 60616 -35850
rect 60736 -35910 60756 -35850
rect 60816 -35910 60896 -35850
rect 60956 -35910 61336 -35850
rect 60466 -35920 61336 -35910
rect 60966 -35960 61336 -35920
rect 61456 -35960 61486 -35830
rect 60966 -35970 61486 -35960
rect 59506 -35990 59606 -35980
rect 59156 -36060 59376 -36050
rect 59306 -36120 60336 -36100
rect 59066 -36140 59176 -36130
rect 55210 -36318 55220 -36148
rect 55310 -36318 55320 -36148
rect 55400 -36328 55410 -36158
rect 55500 -36168 55510 -36158
rect 55500 -36288 56380 -36168
rect 56440 -36288 56450 -36168
rect 59066 -36200 59076 -36140
rect 59166 -36200 59176 -36140
rect 59306 -36180 59316 -36120
rect 59376 -36140 59966 -36120
rect 59376 -36180 59816 -36140
rect 59306 -36190 59816 -36180
rect 59846 -36180 59916 -36170
rect 59066 -36210 59176 -36200
rect 59846 -36240 59856 -36180
rect 59946 -36180 59966 -36140
rect 60326 -36180 60336 -36120
rect 59946 -36190 60336 -36180
rect 60366 -36140 61146 -36130
rect 60366 -36180 61056 -36140
rect 59646 -36250 59716 -36240
rect 59846 -36250 59916 -36240
rect 60366 -36240 60376 -36180
rect 60436 -36240 61056 -36180
rect 61126 -36240 61146 -36140
rect 55500 -36308 56450 -36288
rect 58396 -36260 59716 -36250
rect 55500 -36328 55510 -36308
rect 58396 -36330 58926 -36260
rect 58986 -36330 59146 -36260
rect 59226 -36330 59276 -36260
rect 59356 -36330 59396 -36260
rect 59476 -36320 59646 -36260
rect 59706 -36320 59716 -36260
rect 60366 -36270 61146 -36240
rect 59476 -36330 59716 -36320
rect 58396 -36340 59716 -36330
rect 54900 -36408 54910 -36398
rect 53940 -36488 53950 -36408
rect 54010 -36488 54910 -36408
rect 53940 -36498 54910 -36488
rect 54980 -36418 54990 -36398
rect 54980 -36478 55980 -36418
rect 54980 -36498 55880 -36478
rect 53940 -36518 55880 -36498
rect 53500 -36648 53510 -36528
rect 53630 -36648 53640 -36528
rect 55850 -36558 55880 -36518
rect 55970 -36558 55980 -36478
rect 55230 -36618 55240 -36558
rect 55370 -36578 55710 -36558
rect 55370 -36588 55720 -36578
rect 55370 -36608 55620 -36588
rect 55370 -36618 55380 -36608
rect 55400 -36668 55410 -36648
rect 54730 -36758 54740 -36668
rect 54850 -36738 55410 -36668
rect 55510 -36738 55520 -36648
rect 55600 -36678 55620 -36608
rect 55710 -36678 55720 -36588
rect 54850 -36758 55520 -36738
rect 55210 -36928 55220 -36818
rect 55330 -36928 55340 -36818
rect 55850 -36978 55980 -36558
rect 56010 -36808 56020 -36658
rect 56080 -36808 56090 -36658
rect 56160 -36808 56170 -36608
rect 56390 -36808 56400 -36608
rect 58396 -36620 58896 -36340
rect 59006 -36500 59076 -36480
rect 59246 -36490 59256 -36430
rect 59366 -36490 59376 -36430
rect 59536 -36460 59546 -36390
rect 59606 -36460 59616 -36390
rect 59536 -36470 59616 -36460
rect 59006 -36560 59016 -36500
rect 59536 -36510 59616 -36500
rect 59076 -36520 59086 -36510
rect 59536 -36520 59546 -36510
rect 59076 -36560 59546 -36520
rect 59006 -36570 59546 -36560
rect 59606 -36570 59616 -36510
rect 59006 -36590 59076 -36570
rect 59536 -36590 59616 -36570
rect 59646 -36620 59716 -36340
rect 59796 -36410 59926 -36400
rect 59796 -36520 59806 -36410
rect 59916 -36520 59926 -36410
rect 59796 -36530 59926 -36520
rect 60436 -36430 60536 -36410
rect 60436 -36550 60446 -36430
rect 60526 -36550 60536 -36430
rect 60436 -36560 60536 -36550
rect 58396 -36630 59716 -36620
rect 56654 -36668 56998 -36658
rect 55520 -37068 55530 -36978
rect 55610 -37068 55980 -36978
rect 54130 -37348 54140 -37088
rect 54850 -37348 54860 -37088
rect 55310 -37268 55320 -37128
rect 55470 -37268 55480 -37128
rect 56170 -37338 56390 -36808
rect 58396 -36700 58906 -36630
rect 58986 -36700 59146 -36630
rect 59226 -36700 59276 -36630
rect 59356 -36700 59396 -36630
rect 59476 -36640 59716 -36630
rect 59476 -36700 59646 -36640
rect 59706 -36700 59716 -36640
rect 58396 -36710 59716 -36700
rect 58396 -36750 58896 -36710
rect 59646 -36720 59716 -36710
rect 56654 -36896 56998 -36886
rect 59006 -36800 60416 -36790
rect 59006 -36840 60266 -36800
rect 59006 -36910 59016 -36840
rect 59076 -36910 59546 -36840
rect 59606 -36910 60266 -36840
rect 59006 -36930 60266 -36910
rect 60406 -36930 60416 -36800
rect 59006 -36940 60416 -36930
rect 59986 -36990 60116 -36980
rect 58956 -37000 59156 -36990
rect 58956 -37180 58966 -37000
rect 59146 -37180 59156 -37000
rect 59986 -37100 59996 -36990
rect 60106 -37100 60116 -36990
rect 61900 -37100 62600 -37000
rect 58956 -37190 59156 -37180
rect 55680 -37348 56390 -37338
rect 54130 -37508 56390 -37348
rect 59800 -37200 60300 -37100
rect 59800 -37400 59900 -37200
rect 60200 -37400 60300 -37200
rect 59800 -37500 60300 -37400
rect 55680 -37518 56390 -37508
rect 55300 -37700 56200 -37600
rect 55300 -38100 55400 -37700
rect 56100 -38100 56200 -37700
rect 55300 -38200 56200 -38100
rect 61900 -37700 62000 -37100
rect 62500 -37700 62600 -37100
rect 51400 -38900 51500 -38700
rect 52500 -38900 52600 -38700
rect 51400 -44100 52600 -38900
rect 55440 -38680 55740 -38660
rect 55440 -38960 55460 -38680
rect 55720 -38960 55740 -38680
rect 55440 -38980 55740 -38960
rect 54140 -39138 56390 -39128
rect 53460 -39340 53800 -39320
rect 53460 -39540 53480 -39340
rect 53780 -39540 53800 -39340
rect 54140 -39378 54150 -39138
rect 54860 -39378 56390 -39138
rect 58946 -39270 59146 -39250
rect 54140 -39388 56390 -39378
rect 53460 -39560 53800 -39540
rect 54850 -39618 55530 -39608
rect 53510 -39768 53520 -39658
rect 53640 -39768 53650 -39658
rect 54740 -39718 54750 -39638
rect 54850 -39688 55430 -39618
rect 55520 -39688 55530 -39618
rect 55950 -39688 55960 -39538
rect 56040 -39688 56050 -39538
rect 56170 -39558 56390 -39388
rect 56506 -39380 57016 -39370
rect 54840 -39718 54850 -39708
rect 55270 -39808 55280 -39718
rect 55400 -39808 55410 -39718
rect 56170 -39768 56190 -39558
rect 56390 -39768 56400 -39558
rect 58946 -39430 58966 -39270
rect 59126 -39430 59146 -39270
rect 58946 -39450 59146 -39430
rect 59316 -39300 60176 -39290
rect 59316 -39310 59956 -39300
rect 59316 -39450 59336 -39310
rect 59416 -39450 59956 -39310
rect 59316 -39460 59956 -39450
rect 60166 -39460 60176 -39300
rect 59316 -39470 60176 -39460
rect 56506 -39640 57016 -39630
rect 58956 -39520 61136 -39510
rect 58956 -39530 61056 -39520
rect 58956 -39640 58996 -39530
rect 59106 -39540 61056 -39530
rect 59106 -39640 59516 -39540
rect 59616 -39640 61056 -39540
rect 58396 -39730 58896 -39640
rect 58956 -39650 61056 -39640
rect 61126 -39650 61136 -39520
rect 58956 -39660 61136 -39650
rect 55850 -39848 55880 -39818
rect 53940 -39878 55880 -39848
rect 53940 -39898 54920 -39878
rect 53040 -41708 53050 -39958
rect 53250 -41708 53260 -39958
rect 53940 -39998 53950 -39898
rect 54020 -39948 54920 -39898
rect 54020 -39998 54030 -39948
rect 54910 -39968 54920 -39948
rect 54990 -39898 55880 -39878
rect 55970 -39848 55980 -39818
rect 54990 -39948 55970 -39898
rect 54990 -39968 55000 -39948
rect 55220 -40228 55230 -40058
rect 55320 -40228 55330 -40058
rect 55420 -40218 55430 -40048
rect 55510 -40058 55520 -40048
rect 55510 -40068 56670 -40058
rect 55510 -40198 55600 -40068
rect 55710 -40198 56590 -40068
rect 56660 -40198 56670 -40068
rect 55510 -40208 56670 -40198
rect 58396 -40090 58486 -39730
rect 58816 -39750 58896 -39730
rect 59646 -39750 59706 -39730
rect 58816 -39770 59706 -39750
rect 58816 -39830 58906 -39770
rect 58966 -39830 59216 -39770
rect 59276 -39830 59326 -39770
rect 59386 -39830 59436 -39770
rect 59496 -39830 59636 -39770
rect 59696 -39830 59706 -39770
rect 58816 -39840 59706 -39830
rect 58816 -40090 58896 -39840
rect 59536 -39890 59616 -39880
rect 59276 -39930 59356 -39920
rect 59276 -39990 59286 -39930
rect 59346 -39990 59356 -39930
rect 59536 -39950 59546 -39890
rect 59606 -39950 59616 -39890
rect 59536 -39970 59616 -39950
rect 58996 -40000 59076 -39990
rect 58996 -40060 59006 -40000
rect 59076 -40020 59086 -40000
rect 59536 -40010 59616 -40000
rect 59536 -40020 59546 -40010
rect 59076 -40060 59546 -40020
rect 58996 -40070 59076 -40060
rect 59536 -40070 59546 -40060
rect 59606 -40070 59616 -40010
rect 59536 -40080 59616 -40070
rect 58396 -40110 58896 -40090
rect 59646 -40110 59706 -39840
rect 60436 -39920 60536 -39910
rect 59856 -39940 59976 -39930
rect 59856 -40030 59866 -39940
rect 59966 -40030 59976 -39940
rect 60436 -40020 60446 -39920
rect 60526 -40020 60536 -39920
rect 60436 -40030 60536 -40020
rect 59856 -40040 59976 -40030
rect 58396 -40120 59706 -40110
rect 58396 -40130 59216 -40120
rect 58396 -40190 58906 -40130
rect 58966 -40180 59216 -40130
rect 59276 -40180 59336 -40120
rect 59396 -40180 59436 -40120
rect 59496 -40130 59706 -40120
rect 59496 -40180 59636 -40130
rect 58966 -40190 59636 -40180
rect 59696 -40190 59706 -40130
rect 58396 -40200 59706 -40190
rect 60036 -40120 60136 -40110
rect 60036 -40200 60046 -40120
rect 60126 -40200 60136 -40120
rect 55510 -40218 55520 -40208
rect 59646 -40210 59706 -40200
rect 60546 -40210 60636 -40200
rect 59066 -40240 59176 -40230
rect 59066 -40310 59076 -40240
rect 59166 -40310 59176 -40240
rect 59846 -40280 59856 -40210
rect 59916 -40230 59926 -40210
rect 60356 -40220 60556 -40210
rect 60356 -40230 60376 -40220
rect 59916 -40260 60376 -40230
rect 59916 -40280 59926 -40260
rect 60356 -40280 60376 -40260
rect 60446 -40280 60556 -40220
rect 60356 -40290 60556 -40280
rect 60626 -40290 60636 -40210
rect 59066 -40320 59176 -40310
rect 59966 -40300 60326 -40290
rect 53850 -40438 53860 -40328
rect 53920 -40338 55600 -40328
rect 53920 -40438 55000 -40338
rect 55090 -40438 55540 -40338
rect 55630 -40438 55640 -40338
rect 59966 -40360 59976 -40300
rect 60316 -40360 60326 -40300
rect 60546 -40310 60636 -40290
rect 61186 -40320 61366 -40310
rect 54770 -40638 54850 -40438
rect 56470 -40448 56480 -40388
rect 56550 -40448 56560 -40388
rect 57088 -40504 57098 -40364
rect 57368 -40504 57378 -40364
rect 59166 -40430 59376 -40420
rect 59166 -40440 59286 -40430
rect 59166 -40520 59176 -40440
rect 59236 -40520 59286 -40440
rect 59366 -40520 59376 -40430
rect 59166 -40530 59376 -40520
rect 59526 -40470 59646 -40450
rect 59526 -40530 59576 -40470
rect 59636 -40530 59646 -40470
rect 61186 -40500 61206 -40320
rect 61346 -40500 61366 -40320
rect 61186 -40510 61366 -40500
rect 59526 -40560 59646 -40530
rect 60286 -40550 60476 -40540
rect 59906 -40580 60016 -40570
rect 59806 -40590 59866 -40580
rect 54760 -40728 54770 -40638
rect 54840 -40728 54850 -40638
rect 59166 -40640 59536 -40630
rect 59166 -40720 59176 -40640
rect 59236 -40720 59286 -40640
rect 54920 -40738 55210 -40728
rect 54920 -40808 55140 -40738
rect 55200 -40808 55210 -40738
rect 59166 -40730 59286 -40720
rect 59356 -40650 59536 -40640
rect 59356 -40720 59476 -40650
rect 59356 -40730 59536 -40720
rect 59166 -40740 59536 -40730
rect 59566 -40760 59576 -40590
rect 59636 -40600 59866 -40590
rect 59636 -40740 59806 -40600
rect 59636 -40760 59866 -40740
rect 59906 -40760 59916 -40580
rect 60006 -40760 60016 -40580
rect 60286 -40690 60306 -40550
rect 60456 -40690 60476 -40550
rect 60286 -40700 60476 -40690
rect 61026 -40620 61136 -40610
rect 61026 -40730 61036 -40620
rect 61126 -40730 61136 -40620
rect 61026 -40740 61136 -40730
rect 59566 -40770 59636 -40760
rect 59906 -40770 60016 -40760
rect 54760 -41128 54770 -41048
rect 54840 -41128 54850 -41048
rect 54770 -41338 54850 -41128
rect 54920 -41198 54980 -40808
rect 55880 -40838 56900 -40818
rect 55010 -40928 55020 -40848
rect 55120 -40928 55740 -40848
rect 55810 -40928 55820 -40848
rect 55870 -40928 55880 -40838
rect 55970 -40928 56480 -40838
rect 56550 -40928 56900 -40838
rect 55880 -40948 56900 -40928
rect 57020 -40820 57040 -40818
rect 57800 -40820 58240 -40810
rect 57020 -40940 57800 -40820
rect 57020 -40948 57040 -40940
rect 57800 -40950 58240 -40940
rect 58516 -40860 58796 -40790
rect 58516 -41060 58556 -40860
rect 58756 -41060 58796 -40860
rect 59066 -40810 59936 -40800
rect 59066 -40880 59076 -40810
rect 59166 -40830 59826 -40810
rect 59166 -40880 59316 -40830
rect 59066 -40890 59316 -40880
rect 59376 -40880 59826 -40830
rect 59916 -40880 59936 -40810
rect 59376 -40890 59936 -40880
rect 60076 -40880 60196 -40840
rect 59066 -40970 59936 -40960
rect 59066 -41040 59076 -40970
rect 59166 -41040 59206 -40970
rect 59266 -41040 59826 -40970
rect 59926 -41040 59936 -40970
rect 59066 -41050 59936 -41040
rect 60076 -41040 60096 -40880
rect 60176 -41040 60196 -40880
rect 58516 -41140 58796 -41060
rect 60076 -41080 60196 -41040
rect 61266 -40850 61366 -40840
rect 61266 -41060 61276 -40850
rect 61356 -41060 61366 -40850
rect 61266 -41070 61366 -41060
rect 59586 -41090 59656 -41080
rect 59796 -41090 59866 -41080
rect 59586 -41110 59796 -41090
rect 59156 -41120 59536 -41110
rect 59156 -41130 59266 -41120
rect 54910 -41268 54920 -41198
rect 54980 -41268 54990 -41198
rect 59156 -41210 59166 -41130
rect 59226 -41210 59266 -41130
rect 59366 -41130 59536 -41120
rect 59366 -41210 59466 -41130
rect 59526 -41210 59536 -41130
rect 59156 -41230 59536 -41210
rect 59646 -41250 59796 -41110
rect 59586 -41270 59796 -41250
rect 59856 -41270 59866 -41090
rect 53840 -41448 53850 -41338
rect 53920 -41438 55000 -41338
rect 55090 -41438 55540 -41338
rect 55630 -41438 55640 -41338
rect 56470 -41388 56480 -41328
rect 56550 -41388 56560 -41328
rect 57088 -41414 57098 -41274
rect 57368 -41414 57378 -41274
rect 59796 -41280 59866 -41270
rect 59906 -41090 60016 -41080
rect 59906 -41280 59916 -41090
rect 60006 -41280 60016 -41090
rect 60476 -41110 60546 -41100
rect 60536 -41170 60546 -41110
rect 60476 -41180 60546 -41170
rect 60966 -41230 61486 -41220
rect 60966 -41240 61336 -41230
rect 59906 -41290 60016 -41280
rect 60466 -41250 61336 -41240
rect 59506 -41310 59606 -41300
rect 59156 -41360 59376 -41340
rect 53920 -41448 55640 -41438
rect 59156 -41440 59166 -41360
rect 59226 -41440 59266 -41360
rect 59156 -41450 59266 -41440
rect 59366 -41450 59376 -41360
rect 59506 -41380 59516 -41310
rect 59596 -41380 59606 -41310
rect 60466 -41310 60476 -41250
rect 60536 -41310 60616 -41250
rect 60736 -41310 60756 -41250
rect 60816 -41310 60896 -41250
rect 60956 -41310 61336 -41250
rect 60466 -41320 61336 -41310
rect 60966 -41360 61336 -41320
rect 61456 -41360 61486 -41230
rect 60966 -41370 61486 -41360
rect 59506 -41390 59606 -41380
rect 59156 -41460 59376 -41450
rect 61900 -41500 62600 -37700
rect 62800 -41000 63400 -32100
rect 63600 -40660 64200 -26800
rect 64800 -40200 65500 -21300
rect 65800 -39800 66500 -15900
rect 66800 -39400 67500 -10700
rect 68000 -39000 68700 -5200
rect 71900 -34100 74100 -34000
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 72800 -38740 73100 -35600
rect 84700 -38050 85660 -37780
rect 75380 -38150 75560 -38140
rect 75380 -38270 75390 -38150
rect 75550 -38270 75560 -38150
rect 75380 -38280 75560 -38270
rect 78760 -38150 78900 -38140
rect 78760 -38270 78770 -38150
rect 78890 -38270 78900 -38150
rect 78760 -38280 78900 -38270
rect 72800 -38900 72820 -38740
rect 72810 -38920 72820 -38900
rect 73040 -38900 73100 -38740
rect 73210 -38360 73350 -38350
rect 73210 -38550 73220 -38360
rect 73340 -38550 73350 -38360
rect 73040 -38920 73050 -38900
rect 72810 -38930 73050 -38920
rect 68000 -39200 68100 -39000
rect 68600 -39200 68700 -39000
rect 68000 -39300 68700 -39200
rect 72810 -39070 73050 -39060
rect 72810 -39250 72820 -39070
rect 73040 -39250 73050 -39070
rect 72810 -39260 73050 -39250
rect 66800 -39600 66900 -39400
rect 67400 -39600 67500 -39400
rect 73210 -39340 73350 -38550
rect 73210 -39400 73230 -39340
rect 73330 -39400 73350 -39340
rect 66800 -39800 67500 -39600
rect 72810 -39560 73050 -39550
rect 72810 -39740 72820 -39560
rect 73040 -39740 73050 -39560
rect 72810 -39750 73050 -39740
rect 65800 -40000 65900 -39800
rect 66400 -40000 66500 -39800
rect 65800 -40100 66500 -40000
rect 72810 -39840 73050 -39830
rect 72810 -40020 72820 -39840
rect 73040 -40020 73050 -39840
rect 72810 -40030 73050 -40020
rect 64800 -40400 64900 -40200
rect 65400 -40400 65500 -40200
rect 64800 -40500 65500 -40400
rect 72810 -40300 73050 -40290
rect 72810 -40480 72820 -40300
rect 73040 -40480 73050 -40300
rect 72810 -40490 73050 -40480
rect 63600 -40800 63640 -40660
rect 64160 -40800 64200 -40660
rect 63600 -40840 64200 -40800
rect 72810 -40660 73050 -40650
rect 72810 -40840 72820 -40660
rect 73040 -40840 73050 -40660
rect 72810 -40850 73050 -40840
rect 62800 -41300 62900 -41000
rect 63300 -41300 63400 -41000
rect 72810 -41060 73050 -41050
rect 72810 -41240 72820 -41060
rect 73040 -41240 73050 -41060
rect 72810 -41250 73050 -41240
rect 62800 -41400 63400 -41300
rect 59306 -41520 60336 -41500
rect 59066 -41540 59176 -41530
rect 55210 -41718 55220 -41548
rect 55310 -41718 55320 -41548
rect 55400 -41728 55410 -41558
rect 55500 -41568 55510 -41558
rect 55500 -41688 56380 -41568
rect 56440 -41688 56450 -41568
rect 59066 -41600 59076 -41540
rect 59166 -41600 59176 -41540
rect 59306 -41580 59316 -41520
rect 59376 -41540 59966 -41520
rect 59376 -41580 59816 -41540
rect 59306 -41590 59816 -41580
rect 59846 -41580 59916 -41570
rect 59066 -41610 59176 -41600
rect 59846 -41640 59856 -41580
rect 59946 -41580 59966 -41540
rect 60326 -41580 60336 -41520
rect 59946 -41590 60336 -41580
rect 60366 -41540 61146 -41530
rect 60366 -41580 61056 -41540
rect 59646 -41650 59716 -41640
rect 59846 -41650 59916 -41640
rect 60366 -41640 60376 -41580
rect 60436 -41640 61056 -41580
rect 61126 -41640 61146 -41540
rect 55500 -41708 56450 -41688
rect 58396 -41660 59716 -41650
rect 55500 -41728 55510 -41708
rect 58396 -41730 58926 -41660
rect 58986 -41730 59146 -41660
rect 59226 -41730 59276 -41660
rect 59356 -41730 59396 -41660
rect 59476 -41720 59646 -41660
rect 59706 -41720 59716 -41660
rect 60366 -41670 61146 -41640
rect 59476 -41730 59716 -41720
rect 58396 -41740 59716 -41730
rect 54900 -41808 54910 -41798
rect 53940 -41888 53950 -41808
rect 54010 -41888 54910 -41808
rect 53940 -41898 54910 -41888
rect 54980 -41818 54990 -41798
rect 54980 -41878 55980 -41818
rect 54980 -41898 55880 -41878
rect 53940 -41918 55880 -41898
rect 53500 -42048 53510 -41928
rect 53630 -42048 53640 -41928
rect 55850 -41958 55880 -41918
rect 55970 -41958 55980 -41878
rect 55230 -42018 55240 -41958
rect 55370 -41978 55710 -41958
rect 55370 -41988 55720 -41978
rect 55370 -42008 55620 -41988
rect 55370 -42018 55380 -42008
rect 55400 -42068 55410 -42048
rect 54730 -42158 54740 -42068
rect 54850 -42138 55410 -42068
rect 55510 -42138 55520 -42048
rect 55600 -42078 55620 -42008
rect 55710 -42078 55720 -41988
rect 54850 -42158 55520 -42138
rect 55210 -42328 55220 -42218
rect 55330 -42328 55340 -42218
rect 55850 -42378 55980 -41958
rect 56010 -42208 56020 -42058
rect 56080 -42208 56090 -42058
rect 56160 -42208 56170 -42008
rect 56390 -42208 56400 -42008
rect 58396 -42020 58896 -41740
rect 59006 -41900 59076 -41880
rect 59246 -41890 59256 -41830
rect 59366 -41890 59376 -41830
rect 59536 -41860 59546 -41790
rect 59606 -41860 59616 -41790
rect 59536 -41870 59616 -41860
rect 59006 -41960 59016 -41900
rect 59536 -41910 59616 -41900
rect 59076 -41920 59086 -41910
rect 59536 -41920 59546 -41910
rect 59076 -41960 59546 -41920
rect 59006 -41970 59546 -41960
rect 59606 -41970 59616 -41910
rect 59006 -41990 59076 -41970
rect 59536 -41990 59616 -41970
rect 59646 -42020 59716 -41740
rect 61900 -41700 62000 -41500
rect 62500 -41700 62600 -41500
rect 72810 -41510 73050 -41500
rect 72810 -41690 72820 -41510
rect 73040 -41690 73050 -41510
rect 72810 -41700 73050 -41690
rect 61900 -41800 62600 -41700
rect 59796 -41810 59926 -41800
rect 59796 -41920 59806 -41810
rect 59916 -41920 59926 -41810
rect 59796 -41930 59926 -41920
rect 60436 -41830 60536 -41810
rect 60436 -41950 60446 -41830
rect 60526 -41950 60536 -41830
rect 60436 -41960 60536 -41950
rect 72810 -41880 73050 -41870
rect 58396 -42030 59716 -42020
rect 56654 -42068 56998 -42058
rect 55520 -42468 55530 -42378
rect 55610 -42468 55980 -42378
rect 54130 -42748 54140 -42488
rect 54850 -42748 54860 -42488
rect 55310 -42668 55320 -42528
rect 55470 -42668 55480 -42528
rect 56170 -42738 56390 -42208
rect 58396 -42100 58906 -42030
rect 58986 -42100 59146 -42030
rect 59226 -42100 59276 -42030
rect 59356 -42100 59396 -42030
rect 59476 -42040 59716 -42030
rect 59476 -42100 59646 -42040
rect 59706 -42100 59716 -42040
rect 72810 -42060 72820 -41880
rect 73040 -42060 73050 -41880
rect 72810 -42070 73050 -42060
rect 73210 -41900 73350 -39400
rect 73210 -42040 73220 -41900
rect 73340 -42040 73350 -41900
rect 73210 -42070 73350 -42040
rect 73460 -38360 73600 -38350
rect 73460 -38550 73470 -38360
rect 73590 -38550 73600 -38360
rect 73460 -39120 73600 -38550
rect 73460 -39180 73480 -39120
rect 73580 -39180 73600 -39120
rect 73460 -41530 73600 -39180
rect 73460 -41670 73470 -41530
rect 73590 -41670 73600 -41530
rect 58396 -42110 59716 -42100
rect 58396 -42150 58896 -42110
rect 59646 -42120 59716 -42110
rect 56654 -42296 56998 -42286
rect 59006 -42200 60416 -42190
rect 59006 -42240 60266 -42200
rect 59006 -42310 59016 -42240
rect 59076 -42310 59546 -42240
rect 59606 -42310 60266 -42240
rect 59006 -42330 60266 -42310
rect 60406 -42330 60416 -42200
rect 59006 -42340 60416 -42330
rect 59986 -42390 60116 -42380
rect 58956 -42400 59156 -42390
rect 58956 -42580 58966 -42400
rect 59146 -42580 59156 -42400
rect 59986 -42500 59996 -42390
rect 60106 -42500 60116 -42390
rect 59986 -42510 60116 -42500
rect 58956 -42590 59156 -42580
rect 55680 -42748 56390 -42738
rect 54130 -42908 56390 -42748
rect 55680 -42918 56390 -42908
rect 59600 -42800 60600 -42600
rect 55400 -43100 56200 -43000
rect 55400 -43500 55500 -43100
rect 56100 -43500 56200 -43100
rect 55400 -43600 56200 -43500
rect 59600 -43400 59800 -42800
rect 60400 -43400 60600 -42800
rect 59600 -43600 60600 -43400
rect 51400 -44300 51500 -44100
rect 52500 -44300 52600 -44100
rect 51400 -49500 52600 -44300
rect 55480 -44080 55740 -44060
rect 55480 -44360 55500 -44080
rect 55720 -44360 55740 -44080
rect 55480 -44380 55740 -44360
rect 73460 -44380 73600 -41670
rect 73710 -38360 73850 -38350
rect 73710 -38550 73720 -38360
rect 73840 -38550 73850 -38360
rect 73710 -38596 73850 -38550
rect 73710 -38648 73723 -38596
rect 73840 -38648 73850 -38596
rect 73710 -39230 73850 -38648
rect 73710 -39290 73730 -39230
rect 73830 -39290 73850 -39230
rect 73710 -41090 73850 -39290
rect 73710 -41220 73720 -41090
rect 73840 -41220 73850 -41090
rect 73710 -42930 73850 -41220
rect 73710 -43000 73720 -42930
rect 73840 -43000 73850 -42930
rect 73710 -43010 73850 -43000
rect 73960 -38360 74100 -38350
rect 73960 -38550 73970 -38360
rect 74090 -38550 74100 -38360
rect 73960 -39430 74100 -38550
rect 73960 -39490 73970 -39430
rect 74090 -39490 74100 -39430
rect 73960 -40680 74100 -39490
rect 74210 -38360 74350 -38350
rect 74210 -38550 74220 -38360
rect 74340 -38550 74350 -38360
rect 74210 -38760 74350 -38550
rect 74210 -38840 74220 -38760
rect 74340 -38840 74350 -38760
rect 74210 -39890 74350 -38840
rect 74210 -39950 74230 -39890
rect 74330 -39950 74350 -39890
rect 74210 -40390 74350 -39950
rect 74210 -40450 74220 -40390
rect 74340 -40450 74350 -40390
rect 74210 -40460 74350 -40450
rect 74460 -38360 74600 -38350
rect 74460 -38550 74470 -38360
rect 74590 -38550 74600 -38360
rect 74460 -38570 74600 -38550
rect 74460 -38674 74477 -38570
rect 74594 -38674 74600 -38570
rect 74460 -39860 74600 -38674
rect 74460 -40000 74470 -39860
rect 74590 -40000 74600 -39860
rect 74460 -40110 74600 -40000
rect 74460 -40180 74470 -40110
rect 74590 -40180 74600 -40110
rect 73960 -40820 73970 -40680
rect 74090 -40820 74100 -40680
rect 73460 -44440 73470 -44380
rect 73590 -44440 73600 -44380
rect 73460 -44460 73600 -44440
rect 73960 -43760 74100 -40820
rect 73960 -43830 73970 -43760
rect 74090 -43830 74100 -43760
rect 54140 -44538 56390 -44528
rect 53460 -44740 53800 -44720
rect 53460 -44940 53480 -44740
rect 53780 -44940 53800 -44740
rect 54140 -44778 54150 -44538
rect 54860 -44778 56390 -44538
rect 58946 -44670 59146 -44650
rect 54140 -44788 56390 -44778
rect 53460 -44960 53800 -44940
rect 54850 -45018 55530 -45008
rect 53510 -45168 53520 -45058
rect 53640 -45168 53650 -45058
rect 54740 -45118 54750 -45038
rect 54850 -45088 55430 -45018
rect 55520 -45088 55530 -45018
rect 55950 -45088 55960 -44938
rect 56040 -45088 56050 -44938
rect 56170 -44958 56390 -44788
rect 56506 -44780 57016 -44770
rect 54840 -45118 54850 -45108
rect 55270 -45208 55280 -45118
rect 55400 -45208 55410 -45118
rect 56170 -45168 56190 -44958
rect 56390 -45168 56400 -44958
rect 58946 -44830 58966 -44670
rect 59126 -44830 59146 -44670
rect 58946 -44850 59146 -44830
rect 59316 -44700 60176 -44690
rect 59316 -44710 59956 -44700
rect 59316 -44850 59336 -44710
rect 59416 -44850 59956 -44710
rect 59316 -44860 59956 -44850
rect 60166 -44860 60176 -44700
rect 73960 -44740 74100 -43830
rect 73960 -44800 73970 -44740
rect 74090 -44800 74100 -44740
rect 73960 -44810 74100 -44800
rect 74460 -41320 74600 -40180
rect 74460 -41380 74470 -41320
rect 74590 -41380 74600 -41320
rect 59316 -44870 60176 -44860
rect 56506 -45040 57016 -45030
rect 58956 -44920 61136 -44910
rect 58956 -44930 61056 -44920
rect 58956 -45040 58996 -44930
rect 59106 -44940 61056 -44930
rect 59106 -45040 59516 -44940
rect 59616 -45040 61056 -44940
rect 58396 -45130 58896 -45040
rect 58956 -45050 61056 -45040
rect 61126 -45050 61136 -44920
rect 58956 -45060 61136 -45050
rect 55850 -45248 55880 -45218
rect 53940 -45278 55880 -45248
rect 53940 -45298 54920 -45278
rect 53040 -47108 53050 -45358
rect 53250 -47108 53260 -45358
rect 53940 -45398 53950 -45298
rect 54020 -45348 54920 -45298
rect 54020 -45398 54030 -45348
rect 54910 -45368 54920 -45348
rect 54990 -45298 55880 -45278
rect 55970 -45248 55980 -45218
rect 54990 -45348 55970 -45298
rect 54990 -45368 55000 -45348
rect 55220 -45628 55230 -45458
rect 55320 -45628 55330 -45458
rect 55420 -45618 55430 -45448
rect 55510 -45458 55520 -45448
rect 55510 -45468 56670 -45458
rect 55510 -45598 55600 -45468
rect 55710 -45598 56590 -45468
rect 56660 -45598 56670 -45468
rect 55510 -45608 56670 -45598
rect 58396 -45490 58486 -45130
rect 58816 -45150 58896 -45130
rect 59646 -45150 59706 -45130
rect 58816 -45170 59706 -45150
rect 58816 -45230 58906 -45170
rect 58966 -45230 59216 -45170
rect 59276 -45230 59326 -45170
rect 59386 -45230 59436 -45170
rect 59496 -45230 59636 -45170
rect 59696 -45230 59706 -45170
rect 58816 -45240 59706 -45230
rect 58816 -45490 58896 -45240
rect 59536 -45290 59616 -45280
rect 59276 -45330 59356 -45320
rect 59276 -45390 59286 -45330
rect 59346 -45390 59356 -45330
rect 59536 -45350 59546 -45290
rect 59606 -45350 59616 -45290
rect 59536 -45370 59616 -45350
rect 58996 -45400 59076 -45390
rect 58996 -45460 59006 -45400
rect 59076 -45420 59086 -45400
rect 59536 -45410 59616 -45400
rect 59536 -45420 59546 -45410
rect 59076 -45460 59546 -45420
rect 58996 -45470 59076 -45460
rect 59536 -45470 59546 -45460
rect 59606 -45470 59616 -45410
rect 59536 -45480 59616 -45470
rect 58396 -45510 58896 -45490
rect 59646 -45510 59706 -45240
rect 60436 -45320 60536 -45310
rect 59856 -45340 59976 -45330
rect 59856 -45430 59866 -45340
rect 59966 -45430 59976 -45340
rect 60436 -45420 60446 -45320
rect 60526 -45420 60536 -45320
rect 60436 -45430 60536 -45420
rect 59856 -45440 59976 -45430
rect 74460 -45480 74600 -41380
rect 74710 -38360 74850 -38350
rect 74710 -38550 74720 -38360
rect 74840 -38550 74850 -38360
rect 74710 -38752 74850 -38550
rect 74710 -38830 74724 -38752
rect 74841 -38830 74850 -38752
rect 74710 -39580 74850 -38830
rect 74710 -39720 74720 -39580
rect 74840 -39720 74850 -39580
rect 74710 -39980 74850 -39720
rect 74710 -40040 74730 -39980
rect 74830 -40040 74850 -39980
rect 74710 -41630 74850 -40040
rect 74710 -41690 74720 -41630
rect 74840 -41690 74850 -41630
rect 74710 -41700 74850 -41690
rect 74960 -38360 75100 -38350
rect 74960 -38550 74970 -38360
rect 75090 -38550 75100 -38360
rect 74960 -39100 75100 -38550
rect 74960 -39220 74970 -39100
rect 75090 -39220 75100 -39100
rect 74960 -39780 75100 -39220
rect 74960 -39850 74980 -39780
rect 75080 -39850 75100 -39780
rect 74960 -42270 75100 -39850
rect 74960 -42330 74970 -42270
rect 75090 -42330 75100 -42270
rect 74960 -42340 75100 -42330
rect 75210 -38360 75350 -38350
rect 75210 -38550 75220 -38360
rect 75340 -38550 75350 -38360
rect 76910 -38410 77070 -38400
rect 75210 -38920 75350 -38550
rect 76635 -38440 76739 -38427
rect 76635 -38505 76648 -38440
rect 76726 -38505 76739 -38440
rect 75400 -38590 75480 -38580
rect 75400 -38650 75410 -38590
rect 75470 -38650 75480 -38590
rect 75400 -38660 75480 -38650
rect 75647 -38583 75777 -38570
rect 75400 -38661 75478 -38660
rect 75647 -38661 75673 -38583
rect 75751 -38661 75777 -38583
rect 75210 -39020 75220 -38920
rect 75340 -39020 75350 -38920
rect 75210 -40540 75350 -39020
rect 75647 -39090 75777 -38661
rect 75933 -38583 76063 -38570
rect 75933 -38661 75946 -38583
rect 76024 -38661 76063 -38583
rect 75933 -38940 76063 -38661
rect 76102 -38583 76193 -38570
rect 76180 -38661 76193 -38583
rect 76102 -38674 76193 -38661
rect 76230 -38583 76323 -38570
rect 76230 -38661 76232 -38583
rect 76310 -38661 76323 -38583
rect 76230 -38670 76323 -38661
rect 76232 -38882 76323 -38670
rect 76360 -38600 76460 -38580
rect 76360 -38660 76380 -38600
rect 76440 -38660 76460 -38600
rect 76360 -38680 76460 -38660
rect 76492 -38596 76596 -38583
rect 76492 -38661 76505 -38596
rect 76583 -38661 76596 -38596
rect 76492 -38674 76596 -38661
rect 76362 -38726 76453 -38680
rect 76362 -38804 76375 -38726
rect 76440 -38804 76453 -38726
rect 76362 -38817 76453 -38804
rect 75210 -40610 75220 -40540
rect 75340 -40610 75350 -40540
rect 75210 -41160 75350 -40610
rect 75210 -41240 75220 -41160
rect 75340 -41240 75350 -41160
rect 75210 -41770 75350 -41240
rect 75210 -41860 75220 -41770
rect 75340 -41860 75350 -41770
rect 58396 -45520 59706 -45510
rect 58396 -45530 59216 -45520
rect 58396 -45590 58906 -45530
rect 58966 -45580 59216 -45530
rect 59276 -45580 59336 -45520
rect 59396 -45580 59436 -45520
rect 59496 -45530 59706 -45520
rect 59496 -45580 59636 -45530
rect 58966 -45590 59636 -45580
rect 59696 -45590 59706 -45530
rect 58396 -45600 59706 -45590
rect 60036 -45520 60136 -45510
rect 60036 -45600 60046 -45520
rect 60126 -45600 60136 -45520
rect 74460 -45560 74470 -45480
rect 74590 -45560 74600 -45480
rect 74460 -45570 74600 -45560
rect 75210 -42410 75350 -41860
rect 75210 -42500 75220 -42410
rect 75340 -42500 75350 -42410
rect 75210 -43190 75350 -42500
rect 75210 -43250 75220 -43190
rect 75340 -43250 75350 -43190
rect 75210 -43620 75350 -43250
rect 75210 -43680 75220 -43620
rect 75340 -43680 75350 -43620
rect 75210 -44970 75350 -43680
rect 75640 -44270 75780 -39090
rect 75640 -44330 75660 -44270
rect 75760 -44330 75780 -44270
rect 75920 -43080 76070 -38940
rect 76219 -39080 76323 -38882
rect 76505 -39010 76596 -38674
rect 76635 -38596 76739 -38505
rect 76910 -38530 76920 -38410
rect 77060 -38530 77070 -38410
rect 76910 -38540 77070 -38530
rect 76635 -38674 76648 -38596
rect 76726 -38674 76739 -38596
rect 76635 -38687 76739 -38674
rect 76770 -38596 76870 -38580
rect 76770 -38630 76791 -38596
rect 76843 -38630 76870 -38596
rect 76770 -38700 76780 -38630
rect 76860 -38700 76870 -38630
rect 76770 -38720 76870 -38700
rect 78270 -38630 78360 -38620
rect 78270 -38700 78280 -38630
rect 78350 -38700 78360 -38630
rect 77160 -38790 77440 -38780
rect 75920 -43140 75940 -43080
rect 76050 -43140 76070 -43080
rect 76200 -43070 76350 -39080
rect 76200 -43130 76210 -43070
rect 76340 -43130 76350 -43070
rect 76200 -43140 76350 -43130
rect 75920 -44150 76070 -43140
rect 75920 -44240 75940 -44150
rect 76050 -44240 76070 -44150
rect 75920 -44840 76070 -44240
rect 75920 -44900 75940 -44840
rect 76050 -44900 76070 -44840
rect 76480 -44250 76620 -39010
rect 77160 -39040 77170 -38790
rect 77430 -39040 77440 -38790
rect 77160 -39050 77440 -39040
rect 78140 -39340 78220 -39330
rect 78140 -39400 78150 -39340
rect 78210 -39400 78220 -39340
rect 77220 -39440 77320 -39430
rect 77220 -39500 77230 -39440
rect 77310 -39500 77320 -39440
rect 77220 -39510 77320 -39500
rect 76910 -39570 77070 -39560
rect 76910 -39720 76920 -39570
rect 77060 -39720 77070 -39570
rect 76910 -39730 77070 -39720
rect 77160 -39780 77270 -39770
rect 77160 -39850 77170 -39780
rect 77260 -39850 77270 -39780
rect 77160 -39860 77270 -39850
rect 78140 -39790 78220 -39400
rect 78270 -39340 78360 -38700
rect 78270 -39400 78280 -39340
rect 78340 -39400 78360 -39340
rect 78270 -39410 78360 -39400
rect 78570 -39320 78650 -39310
rect 78570 -39380 78580 -39320
rect 78640 -39380 78650 -39320
rect 78140 -40080 78150 -39790
rect 78210 -40080 78220 -39790
rect 78570 -39840 78650 -39380
rect 78790 -39330 78870 -38280
rect 84700 -38480 84960 -38050
rect 85400 -38480 85660 -38050
rect 84700 -38690 85660 -38480
rect 87880 -38390 88840 -38140
rect 87880 -38820 88150 -38390
rect 88590 -38820 88840 -38390
rect 82760 -39010 82910 -38990
rect 82760 -39100 82780 -39010
rect 82890 -39100 82910 -39010
rect 80050 -39270 80460 -39240
rect 78790 -39390 78800 -39330
rect 78860 -39390 78870 -39330
rect 78790 -39400 78870 -39390
rect 79060 -39350 79270 -39330
rect 79060 -39510 79080 -39350
rect 79250 -39510 79270 -39350
rect 79060 -39520 79270 -39510
rect 80050 -39580 80080 -39270
rect 80430 -39580 80460 -39270
rect 82760 -39270 82910 -39100
rect 82760 -39520 82780 -39270
rect 82890 -39520 82910 -39270
rect 83350 -39010 83760 -38990
rect 83350 -39080 83370 -39010
rect 83740 -39080 83760 -39010
rect 83350 -39370 83760 -39080
rect 84850 -39000 85260 -38990
rect 84850 -39070 84870 -39000
rect 85240 -39070 85260 -39000
rect 84220 -39250 84320 -39240
rect 83350 -39380 83790 -39370
rect 83350 -39450 83370 -39380
rect 83770 -39450 83790 -39380
rect 83350 -39460 83790 -39450
rect 82760 -39560 82910 -39520
rect 84220 -39540 84230 -39250
rect 84310 -39540 84320 -39250
rect 84850 -39380 85260 -39070
rect 86310 -39000 86720 -38990
rect 86310 -39070 86330 -39000
rect 86700 -39070 86720 -39000
rect 84850 -39450 84870 -39380
rect 85240 -39450 85260 -39380
rect 84850 -39460 85260 -39450
rect 85700 -39260 85800 -39240
rect 80050 -39610 80460 -39580
rect 78570 -39900 78580 -39840
rect 78640 -39900 78650 -39840
rect 78570 -39920 78650 -39900
rect 80050 -39680 80460 -39650
rect 78140 -40100 78220 -40080
rect 80050 -40060 80080 -39680
rect 80430 -40060 80460 -39680
rect 84220 -39700 84320 -39540
rect 80050 -40090 80460 -40060
rect 83000 -39830 83640 -39700
rect 84220 -39810 84230 -39700
rect 84310 -39810 84320 -39700
rect 84220 -39820 84320 -39810
rect 85700 -39550 85710 -39260
rect 85790 -39550 85800 -39260
rect 86310 -39380 86720 -39070
rect 87440 -39000 87770 -38990
rect 87440 -39070 87460 -39000
rect 87750 -39070 87770 -39000
rect 87880 -39050 88840 -38820
rect 86310 -39450 86320 -39380
rect 86710 -39450 86720 -39380
rect 86310 -39460 86720 -39450
rect 87170 -39240 87270 -39230
rect 85700 -39700 85800 -39550
rect 85700 -39810 85710 -39700
rect 85790 -39810 85800 -39700
rect 85700 -39820 85800 -39810
rect 87170 -39510 87180 -39240
rect 87260 -39510 87270 -39240
rect 87440 -39380 87770 -39070
rect 87440 -39450 87450 -39380
rect 87760 -39450 87770 -39380
rect 87440 -39460 87770 -39450
rect 88640 -39250 88740 -39240
rect 87170 -39700 87270 -39510
rect 87170 -39810 87180 -39700
rect 87260 -39810 87270 -39700
rect 87170 -39820 87270 -39810
rect 88640 -39540 88650 -39250
rect 88730 -39540 88740 -39250
rect 88640 -39700 88740 -39540
rect 88640 -39810 88650 -39700
rect 88730 -39810 88740 -39700
rect 88640 -39820 88740 -39810
rect 91750 -39580 92160 -39550
rect 77400 -40110 77490 -40100
rect 77400 -40180 77410 -40110
rect 77480 -40180 77490 -40110
rect 79730 -40130 79920 -40120
rect 77400 -40190 77490 -40180
rect 79400 -40150 79690 -40140
rect 77770 -40390 77850 -40380
rect 77770 -40450 77780 -40390
rect 77840 -40450 77850 -40390
rect 79400 -40390 79410 -40150
rect 79680 -40390 79690 -40150
rect 79400 -40400 79690 -40390
rect 79730 -40370 79780 -40130
rect 79910 -40370 79920 -40130
rect 83000 -40180 83150 -39830
rect 83510 -40180 83640 -39830
rect 91750 -39960 91780 -39580
rect 92130 -39960 92160 -39580
rect 77440 -40540 77530 -40530
rect 77440 -40610 77450 -40540
rect 77520 -40610 77530 -40540
rect 77440 -40620 77530 -40610
rect 77770 -40570 77850 -40450
rect 77770 -40630 77780 -40570
rect 77840 -40630 77850 -40570
rect 77770 -40640 77850 -40630
rect 78300 -40650 78420 -40640
rect 78300 -40760 78310 -40650
rect 78410 -40760 78420 -40650
rect 78300 -40770 78420 -40760
rect 76910 -40820 77070 -40810
rect 76910 -40960 76920 -40820
rect 77060 -40960 77070 -40820
rect 76910 -40970 77070 -40960
rect 78050 -41090 78130 -41080
rect 77770 -41140 77850 -41130
rect 77440 -41160 77540 -41150
rect 77440 -41240 77450 -41160
rect 77530 -41240 77540 -41160
rect 77440 -41250 77540 -41240
rect 77770 -41200 77780 -41140
rect 77840 -41200 77850 -41140
rect 77770 -41320 77850 -41200
rect 77770 -41380 77780 -41320
rect 77840 -41380 77850 -41320
rect 77770 -41390 77850 -41380
rect 78050 -41180 78060 -41090
rect 78120 -41180 78130 -41090
rect 78340 -41130 78420 -40770
rect 77770 -41630 77850 -41620
rect 77770 -41690 77780 -41630
rect 77840 -41690 77850 -41630
rect 77480 -41770 77590 -41760
rect 77480 -41860 77490 -41770
rect 77580 -41860 77590 -41770
rect 77480 -41870 77590 -41860
rect 77770 -41810 77850 -41690
rect 77770 -41870 77780 -41810
rect 77840 -41870 77850 -41810
rect 77770 -41880 77850 -41870
rect 76910 -42060 77070 -42050
rect 76910 -42220 76920 -42060
rect 77060 -42220 77070 -42060
rect 76910 -42230 77070 -42220
rect 77770 -42270 77850 -42260
rect 77770 -42330 77780 -42270
rect 77840 -42330 77850 -42270
rect 77770 -42380 77850 -42330
rect 77460 -42410 77570 -42400
rect 77460 -42500 77470 -42410
rect 77560 -42500 77570 -42410
rect 77770 -42440 77780 -42380
rect 77840 -42440 77850 -42380
rect 77770 -42450 77850 -42440
rect 78050 -42330 78130 -41180
rect 78160 -41140 78300 -41130
rect 78160 -41240 78180 -41140
rect 78290 -41240 78300 -41140
rect 78340 -41190 78350 -41130
rect 78410 -41190 78420 -41130
rect 78340 -41200 78420 -41190
rect 78660 -41030 78790 -41020
rect 78160 -41260 78300 -41240
rect 78200 -41720 78300 -41260
rect 78660 -41380 78670 -41030
rect 78780 -41380 78790 -41030
rect 78660 -41390 78790 -41380
rect 79400 -41380 79690 -41370
rect 79400 -41620 79410 -41380
rect 79680 -41620 79690 -41380
rect 79400 -41630 79690 -41620
rect 78160 -41730 78300 -41720
rect 78160 -42000 78170 -41730
rect 78290 -42000 78300 -41730
rect 78160 -42010 78300 -42000
rect 78520 -41730 78600 -41720
rect 78520 -42000 78530 -41730
rect 78590 -42000 78600 -41730
rect 78050 -42340 78310 -42330
rect 77460 -42510 77570 -42500
rect 78050 -42640 78060 -42340
rect 78120 -42370 78310 -42340
rect 78120 -42470 78160 -42370
rect 78260 -42470 78310 -42370
rect 78120 -42640 78310 -42470
rect 78050 -42650 78310 -42640
rect 78520 -42530 78600 -42000
rect 79040 -42360 79170 -42340
rect 79040 -42470 79050 -42360
rect 79150 -42470 79170 -42360
rect 78520 -42650 78710 -42530
rect 78230 -42880 78310 -42650
rect 77460 -42930 77550 -42920
rect 77460 -43000 77470 -42930
rect 77540 -43000 77550 -42930
rect 78230 -42940 78240 -42880
rect 78300 -42940 78310 -42880
rect 78230 -42950 78310 -42940
rect 77460 -43010 77550 -43000
rect 77850 -43050 77930 -43040
rect 77190 -43080 77270 -43070
rect 77190 -43140 77200 -43080
rect 77260 -43140 77270 -43080
rect 77850 -43110 77860 -43050
rect 77920 -43110 77930 -43050
rect 78620 -43080 78710 -42650
rect 77850 -43120 77930 -43110
rect 76910 -43310 77070 -43300
rect 76910 -43450 76920 -43310
rect 77060 -43450 77070 -43310
rect 76910 -43460 77070 -43450
rect 77190 -43530 77270 -43140
rect 77190 -43590 77200 -43530
rect 77260 -43590 77270 -43530
rect 77190 -43600 77270 -43590
rect 77860 -43500 77920 -43120
rect 78340 -43140 78410 -43080
rect 77950 -43190 78030 -43180
rect 77950 -43250 77960 -43190
rect 78020 -43250 78030 -43190
rect 78620 -43140 78630 -43080
rect 78700 -43140 78710 -43080
rect 78620 -43150 78710 -43140
rect 78850 -42920 78990 -42910
rect 78340 -43210 78410 -43200
rect 78850 -43210 78860 -42920
rect 78980 -43210 78990 -42920
rect 77950 -43260 78030 -43250
rect 78350 -43480 78400 -43210
rect 78850 -43220 78990 -43210
rect 78240 -43500 78420 -43480
rect 77860 -43680 77920 -43670
rect 77960 -43620 78040 -43610
rect 77960 -43680 77970 -43620
rect 78030 -43680 78040 -43620
rect 77960 -43690 78040 -43680
rect 77420 -43760 77510 -43750
rect 77420 -43830 77430 -43760
rect 77500 -43830 77510 -43760
rect 77420 -43840 77510 -43830
rect 78300 -43870 78420 -43500
rect 78240 -43880 78420 -43870
rect 76480 -44310 76490 -44250
rect 76610 -44310 76620 -44250
rect 76480 -44880 76620 -44310
rect 78170 -44130 78310 -44120
rect 77960 -44350 78040 -44340
rect 77750 -44420 77830 -44410
rect 77750 -44480 77760 -44420
rect 77820 -44480 77830 -44420
rect 77960 -44470 77970 -44350
rect 78030 -44470 78040 -44350
rect 77960 -44480 78040 -44470
rect 78170 -44470 78180 -44130
rect 78300 -44470 78310 -44130
rect 77750 -44490 77830 -44480
rect 78170 -44510 78310 -44470
rect 76910 -44520 77070 -44510
rect 76910 -44610 76920 -44520
rect 77060 -44610 77070 -44520
rect 76910 -44620 77070 -44610
rect 77750 -44740 77830 -44730
rect 77750 -44800 77760 -44740
rect 77820 -44800 77830 -44740
rect 77750 -44810 77830 -44800
rect 75210 -45060 75230 -44970
rect 75330 -45060 75350 -44970
rect 75210 -45500 75350 -45060
rect 76480 -44950 76490 -44880
rect 76610 -44950 76620 -44880
rect 77950 -44850 78030 -44840
rect 77950 -44920 77960 -44850
rect 78020 -44920 78030 -44850
rect 77950 -44930 78030 -44920
rect 76480 -45350 76620 -44950
rect 76480 -45420 76500 -45350
rect 76600 -45420 76620 -45350
rect 75210 -45570 75230 -45500
rect 75330 -45570 75350 -45500
rect 55510 -45618 55520 -45608
rect 59646 -45610 59706 -45600
rect 60546 -45610 60636 -45600
rect 59066 -45640 59176 -45630
rect 59066 -45710 59076 -45640
rect 59166 -45710 59176 -45640
rect 59846 -45680 59856 -45610
rect 59916 -45630 59926 -45610
rect 60356 -45620 60556 -45610
rect 60356 -45630 60376 -45620
rect 59916 -45660 60376 -45630
rect 59916 -45680 59926 -45660
rect 60356 -45680 60376 -45660
rect 60446 -45680 60556 -45620
rect 60356 -45690 60556 -45680
rect 60626 -45690 60636 -45610
rect 59066 -45720 59176 -45710
rect 59966 -45700 60326 -45690
rect 53850 -45838 53860 -45728
rect 53920 -45738 55600 -45728
rect 53920 -45838 55000 -45738
rect 55090 -45838 55540 -45738
rect 55630 -45838 55640 -45738
rect 59966 -45760 59976 -45700
rect 60316 -45760 60326 -45700
rect 60546 -45710 60636 -45690
rect 61186 -45720 61366 -45710
rect 54770 -46038 54850 -45838
rect 56470 -45848 56480 -45788
rect 56550 -45848 56560 -45788
rect 57088 -45904 57098 -45764
rect 57368 -45904 57378 -45764
rect 59166 -45830 59376 -45820
rect 59166 -45840 59286 -45830
rect 59166 -45920 59176 -45840
rect 59236 -45920 59286 -45840
rect 59366 -45920 59376 -45830
rect 59166 -45930 59376 -45920
rect 59526 -45870 59646 -45850
rect 59526 -45930 59576 -45870
rect 59636 -45930 59646 -45870
rect 61186 -45900 61206 -45720
rect 61346 -45900 61366 -45720
rect 61186 -45910 61366 -45900
rect 75210 -45890 75350 -45570
rect 78060 -45480 78150 -45470
rect 78060 -45590 78070 -45480
rect 78140 -45590 78150 -45480
rect 77590 -45610 77720 -45600
rect 76910 -45640 77070 -45630
rect 76910 -45740 76920 -45640
rect 77060 -45740 77070 -45640
rect 77590 -45680 77600 -45610
rect 77710 -45680 77720 -45610
rect 77590 -45690 77720 -45680
rect 76910 -45750 77070 -45740
rect 59526 -45960 59646 -45930
rect 60286 -45950 60476 -45940
rect 59906 -45980 60016 -45970
rect 59806 -45990 59866 -45980
rect 54760 -46128 54770 -46038
rect 54840 -46128 54850 -46038
rect 59166 -46040 59536 -46030
rect 59166 -46120 59176 -46040
rect 59236 -46120 59286 -46040
rect 54920 -46138 55210 -46128
rect 54920 -46208 55140 -46138
rect 55200 -46208 55210 -46138
rect 59166 -46130 59286 -46120
rect 59356 -46050 59536 -46040
rect 59356 -46120 59476 -46050
rect 59356 -46130 59536 -46120
rect 59166 -46140 59536 -46130
rect 59566 -46160 59576 -45990
rect 59636 -46000 59866 -45990
rect 59636 -46140 59806 -46000
rect 59636 -46160 59866 -46140
rect 59906 -46160 59916 -45980
rect 60006 -46160 60016 -45980
rect 60286 -46090 60306 -45950
rect 60456 -46090 60476 -45950
rect 75210 -45950 75220 -45890
rect 75340 -45950 75350 -45890
rect 75210 -45960 75350 -45950
rect 78060 -45890 78150 -45590
rect 78230 -45530 78310 -44510
rect 78770 -44770 78930 -44760
rect 78770 -44890 78780 -44770
rect 78920 -44890 78930 -44770
rect 79040 -44800 79170 -42470
rect 79400 -42640 79690 -42630
rect 79400 -42880 79410 -42640
rect 79680 -42880 79690 -42640
rect 79400 -42890 79690 -42880
rect 79400 -43860 79690 -43850
rect 79400 -44100 79410 -43860
rect 79680 -44100 79690 -43860
rect 79400 -44110 79690 -44100
rect 79040 -44870 79070 -44800
rect 79140 -44870 79170 -44800
rect 79040 -44890 79170 -44870
rect 78770 -44900 78930 -44890
rect 78230 -45590 78240 -45530
rect 78300 -45590 78310 -45530
rect 78230 -45600 78310 -45590
rect 78630 -44950 78760 -44940
rect 78630 -45090 78640 -44950
rect 78750 -45090 78760 -44950
rect 78630 -45510 78760 -45090
rect 78630 -45600 78640 -45510
rect 78740 -45600 78760 -45510
rect 78630 -45610 78760 -45600
rect 78800 -45550 78880 -44900
rect 79400 -45120 79690 -45110
rect 79400 -45360 79410 -45120
rect 79680 -45360 79690 -45120
rect 78800 -45610 78810 -45550
rect 78870 -45610 78880 -45550
rect 78800 -45620 78880 -45610
rect 79060 -45380 79210 -45360
rect 79400 -45370 79690 -45360
rect 79060 -45680 79080 -45380
rect 79190 -45680 79210 -45380
rect 79060 -45700 79210 -45680
rect 78060 -45950 78070 -45890
rect 78140 -45950 78150 -45890
rect 78060 -45960 78150 -45950
rect 60286 -46100 60476 -46090
rect 61026 -46020 61136 -46010
rect 61026 -46130 61036 -46020
rect 61126 -46130 61136 -46020
rect 61026 -46140 61136 -46130
rect 59566 -46170 59636 -46160
rect 59906 -46170 60016 -46160
rect 75380 -46190 75560 -46180
rect 54760 -46528 54770 -46448
rect 54840 -46528 54850 -46448
rect 54770 -46738 54850 -46528
rect 54920 -46598 54980 -46208
rect 55880 -46238 56900 -46218
rect 55010 -46328 55020 -46248
rect 55120 -46328 55740 -46248
rect 55810 -46328 55820 -46248
rect 55870 -46328 55880 -46238
rect 55970 -46328 56480 -46238
rect 56550 -46328 56900 -46238
rect 55880 -46348 56900 -46328
rect 57020 -46220 57040 -46218
rect 57800 -46220 58240 -46210
rect 57020 -46340 57800 -46220
rect 57020 -46348 57040 -46340
rect 57800 -46350 58240 -46340
rect 58516 -46260 58796 -46190
rect 58516 -46460 58556 -46260
rect 58756 -46460 58796 -46260
rect 59066 -46210 59936 -46200
rect 59066 -46280 59076 -46210
rect 59166 -46230 59826 -46210
rect 59166 -46280 59316 -46230
rect 59066 -46290 59316 -46280
rect 59376 -46280 59826 -46230
rect 59916 -46280 59936 -46210
rect 59376 -46290 59936 -46280
rect 60076 -46280 60196 -46240
rect 59066 -46370 59936 -46360
rect 59066 -46440 59076 -46370
rect 59166 -46440 59206 -46370
rect 59266 -46440 59826 -46370
rect 59926 -46440 59936 -46370
rect 59066 -46450 59936 -46440
rect 60076 -46440 60096 -46280
rect 60176 -46440 60196 -46280
rect 58516 -46540 58796 -46460
rect 60076 -46480 60196 -46440
rect 61266 -46250 61366 -46240
rect 61266 -46460 61276 -46250
rect 61356 -46460 61366 -46250
rect 75380 -46310 75390 -46190
rect 75550 -46310 75560 -46190
rect 75380 -46320 75560 -46310
rect 78760 -46190 78900 -46180
rect 78760 -46310 78770 -46190
rect 78890 -46310 78900 -46190
rect 78760 -46320 78900 -46310
rect 79730 -46190 79920 -40370
rect 81110 -40250 81600 -40220
rect 81110 -40510 81140 -40250
rect 81570 -40510 81600 -40250
rect 83000 -40290 83640 -40180
rect 87520 -40240 88480 -39980
rect 91750 -39990 92160 -39960
rect 81110 -40540 81600 -40510
rect 87520 -40590 87830 -40240
rect 88190 -40590 88480 -40240
rect 80050 -40910 80460 -40880
rect 80050 -41290 80080 -40910
rect 80430 -41290 80460 -40910
rect 80050 -41320 80460 -41290
rect 82430 -40910 82980 -40880
rect 87520 -40890 88480 -40590
rect 82430 -41290 82460 -40910
rect 82950 -41290 82980 -40910
rect 82430 -41320 82980 -41290
rect 79980 -42910 80390 -42880
rect 79980 -43290 80010 -42910
rect 80360 -43290 80390 -42910
rect 79980 -43320 80390 -43290
rect 82090 -42910 82520 -42880
rect 82090 -43290 82120 -42910
rect 82490 -43290 82520 -42910
rect 82090 -43320 82520 -43290
rect 79980 -45430 80390 -45400
rect 79980 -45810 80010 -45430
rect 80360 -45810 80390 -45430
rect 79980 -45840 80390 -45810
rect 81480 -45430 81960 -45400
rect 81480 -45810 81510 -45430
rect 81930 -45810 81960 -45430
rect 81480 -45840 81960 -45810
rect 79730 -46310 79740 -46190
rect 79910 -46310 79920 -46190
rect 79730 -46320 79920 -46310
rect 61266 -46470 61366 -46460
rect 73210 -46400 73350 -46390
rect 59586 -46490 59656 -46480
rect 59796 -46490 59866 -46480
rect 59586 -46510 59796 -46490
rect 59156 -46520 59536 -46510
rect 59156 -46530 59266 -46520
rect 54910 -46668 54920 -46598
rect 54980 -46668 54990 -46598
rect 59156 -46610 59166 -46530
rect 59226 -46610 59266 -46530
rect 59366 -46530 59536 -46520
rect 59366 -46610 59466 -46530
rect 59526 -46610 59536 -46530
rect 59156 -46630 59536 -46610
rect 59646 -46650 59796 -46510
rect 59586 -46670 59796 -46650
rect 59856 -46670 59866 -46490
rect 53840 -46848 53850 -46738
rect 53920 -46838 55000 -46738
rect 55090 -46838 55540 -46738
rect 55630 -46838 55640 -46738
rect 56470 -46788 56480 -46728
rect 56550 -46788 56560 -46728
rect 57088 -46814 57098 -46674
rect 57368 -46814 57378 -46674
rect 59796 -46680 59866 -46670
rect 59906 -46490 60016 -46480
rect 59906 -46680 59916 -46490
rect 60006 -46680 60016 -46490
rect 60476 -46510 60546 -46500
rect 60536 -46570 60546 -46510
rect 60476 -46580 60546 -46570
rect 73210 -46590 73220 -46400
rect 73340 -46590 73350 -46400
rect 60966 -46630 61486 -46620
rect 60966 -46640 61336 -46630
rect 59906 -46690 60016 -46680
rect 60466 -46650 61336 -46640
rect 59506 -46710 59606 -46700
rect 59156 -46760 59376 -46740
rect 53920 -46848 55640 -46838
rect 59156 -46840 59166 -46760
rect 59226 -46840 59266 -46760
rect 59156 -46850 59266 -46840
rect 59366 -46850 59376 -46760
rect 59506 -46780 59516 -46710
rect 59596 -46780 59606 -46710
rect 60466 -46710 60476 -46650
rect 60536 -46710 60616 -46650
rect 60736 -46710 60756 -46650
rect 60816 -46710 60896 -46650
rect 60956 -46710 61336 -46650
rect 60466 -46720 61336 -46710
rect 60966 -46760 61336 -46720
rect 61456 -46760 61486 -46630
rect 60966 -46770 61486 -46760
rect 59506 -46790 59606 -46780
rect 59156 -46860 59376 -46850
rect 72810 -46900 73050 -46890
rect 59306 -46920 60336 -46900
rect 59066 -46940 59176 -46930
rect 55210 -47118 55220 -46948
rect 55310 -47118 55320 -46948
rect 55400 -47128 55410 -46958
rect 55500 -46968 55510 -46958
rect 55500 -47088 56380 -46968
rect 56440 -47088 56450 -46968
rect 59066 -47000 59076 -46940
rect 59166 -47000 59176 -46940
rect 59306 -46980 59316 -46920
rect 59376 -46940 59966 -46920
rect 59376 -46980 59816 -46940
rect 59306 -46990 59816 -46980
rect 59846 -46980 59916 -46970
rect 59066 -47010 59176 -47000
rect 59846 -47040 59856 -46980
rect 59946 -46980 59966 -46940
rect 60326 -46980 60336 -46920
rect 59946 -46990 60336 -46980
rect 60366 -46940 61146 -46930
rect 60366 -46980 61056 -46940
rect 59646 -47050 59716 -47040
rect 59846 -47050 59916 -47040
rect 60366 -47040 60376 -46980
rect 60436 -47040 61056 -46980
rect 61126 -47040 61146 -46940
rect 55500 -47108 56450 -47088
rect 58396 -47060 59716 -47050
rect 55500 -47128 55510 -47108
rect 58396 -47130 58926 -47060
rect 58986 -47130 59146 -47060
rect 59226 -47130 59276 -47060
rect 59356 -47130 59396 -47060
rect 59476 -47120 59646 -47060
rect 59706 -47120 59716 -47060
rect 60366 -47070 61146 -47040
rect 72810 -47080 72820 -46900
rect 73040 -47080 73050 -46900
rect 72810 -47090 73050 -47080
rect 59476 -47130 59716 -47120
rect 58396 -47140 59716 -47130
rect 54900 -47208 54910 -47198
rect 53940 -47288 53950 -47208
rect 54010 -47288 54910 -47208
rect 53940 -47298 54910 -47288
rect 54980 -47218 54990 -47198
rect 54980 -47278 55980 -47218
rect 54980 -47298 55880 -47278
rect 53940 -47318 55880 -47298
rect 53500 -47448 53510 -47328
rect 53630 -47448 53640 -47328
rect 55850 -47358 55880 -47318
rect 55970 -47358 55980 -47278
rect 55230 -47418 55240 -47358
rect 55370 -47378 55710 -47358
rect 55370 -47388 55720 -47378
rect 55370 -47408 55620 -47388
rect 55370 -47418 55380 -47408
rect 55400 -47468 55410 -47448
rect 54730 -47558 54740 -47468
rect 54850 -47538 55410 -47468
rect 55510 -47538 55520 -47448
rect 55600 -47478 55620 -47408
rect 55710 -47478 55720 -47388
rect 54850 -47558 55520 -47538
rect 55210 -47728 55220 -47618
rect 55330 -47728 55340 -47618
rect 55850 -47778 55980 -47358
rect 56010 -47608 56020 -47458
rect 56080 -47608 56090 -47458
rect 56160 -47608 56170 -47408
rect 56390 -47608 56400 -47408
rect 58396 -47420 58896 -47140
rect 59006 -47300 59076 -47280
rect 59246 -47290 59256 -47230
rect 59366 -47290 59376 -47230
rect 59536 -47260 59546 -47190
rect 59606 -47260 59616 -47190
rect 59536 -47270 59616 -47260
rect 59006 -47360 59016 -47300
rect 59536 -47310 59616 -47300
rect 59076 -47320 59086 -47310
rect 59536 -47320 59546 -47310
rect 59076 -47360 59546 -47320
rect 59006 -47370 59546 -47360
rect 59606 -47370 59616 -47310
rect 59006 -47390 59076 -47370
rect 59536 -47390 59616 -47370
rect 59646 -47420 59716 -47140
rect 62400 -47200 63000 -47100
rect 59796 -47210 59926 -47200
rect 59796 -47320 59806 -47210
rect 59916 -47320 59926 -47210
rect 59796 -47330 59926 -47320
rect 60436 -47230 60536 -47210
rect 60436 -47350 60446 -47230
rect 60526 -47350 60536 -47230
rect 60436 -47360 60536 -47350
rect 58396 -47430 59716 -47420
rect 56654 -47468 56998 -47458
rect 55520 -47868 55530 -47778
rect 55610 -47868 55980 -47778
rect 54130 -48148 54140 -47888
rect 54850 -48148 54860 -47888
rect 55310 -48068 55320 -47928
rect 55470 -48068 55480 -47928
rect 56170 -48138 56390 -47608
rect 58396 -47500 58906 -47430
rect 58986 -47500 59146 -47430
rect 59226 -47500 59276 -47430
rect 59356 -47500 59396 -47430
rect 59476 -47440 59716 -47430
rect 59476 -47500 59646 -47440
rect 59706 -47500 59716 -47440
rect 58396 -47510 59716 -47500
rect 58396 -47550 58896 -47510
rect 59646 -47520 59716 -47510
rect 62400 -47500 62500 -47200
rect 62900 -47500 63000 -47200
rect 72810 -47230 73050 -47220
rect 72810 -47410 72820 -47230
rect 73040 -47410 73050 -47230
rect 72810 -47420 73050 -47410
rect 73210 -47380 73350 -46590
rect 56654 -47696 56998 -47686
rect 59006 -47600 60416 -47590
rect 59006 -47640 60266 -47600
rect 59006 -47710 59016 -47640
rect 59076 -47710 59546 -47640
rect 59606 -47710 60266 -47640
rect 59006 -47730 60266 -47710
rect 60406 -47730 60416 -47600
rect 59006 -47740 60416 -47730
rect 59986 -47790 60116 -47780
rect 58956 -47800 59156 -47790
rect 58956 -47980 58966 -47800
rect 59146 -47980 59156 -47800
rect 59986 -47900 59996 -47790
rect 60106 -47900 60116 -47790
rect 58956 -47990 59156 -47980
rect 55680 -48148 56390 -48138
rect 54130 -48308 56390 -48148
rect 55680 -48318 56390 -48308
rect 59600 -48000 60500 -47900
rect 59600 -48400 59700 -48000
rect 60400 -48400 60500 -48000
rect 55400 -48500 56200 -48400
rect 59600 -48500 60500 -48400
rect 62400 -48000 63000 -47500
rect 73210 -47440 73230 -47380
rect 73330 -47440 73350 -47380
rect 62400 -48400 62500 -48000
rect 62900 -48400 63000 -48000
rect 62400 -48500 63000 -48400
rect 64100 -47700 64600 -47600
rect 64100 -47900 64200 -47700
rect 64500 -47900 64600 -47700
rect 55400 -48900 55500 -48500
rect 56100 -48900 56200 -48500
rect 55400 -49000 56200 -48900
rect 51400 -49700 51500 -49500
rect 52500 -49700 52600 -49500
rect 51400 -54900 52600 -49700
rect 55440 -49480 55740 -49460
rect 55440 -49760 55460 -49480
rect 55720 -49760 55740 -49480
rect 55440 -49780 55740 -49760
rect 54140 -49938 56390 -49928
rect 53440 -50140 53800 -50120
rect 53440 -50340 53460 -50140
rect 53780 -50340 53800 -50140
rect 54140 -50178 54150 -49938
rect 54860 -50178 56390 -49938
rect 58946 -50070 59146 -50050
rect 54140 -50188 56390 -50178
rect 53440 -50360 53800 -50340
rect 54850 -50418 55530 -50408
rect 53510 -50568 53520 -50458
rect 53640 -50568 53650 -50458
rect 54740 -50518 54750 -50438
rect 54850 -50488 55430 -50418
rect 55520 -50488 55530 -50418
rect 55950 -50488 55960 -50338
rect 56040 -50488 56050 -50338
rect 56170 -50358 56390 -50188
rect 56506 -50180 57016 -50170
rect 54840 -50518 54850 -50508
rect 55270 -50608 55280 -50518
rect 55400 -50608 55410 -50518
rect 56170 -50568 56190 -50358
rect 56390 -50568 56400 -50358
rect 58946 -50230 58966 -50070
rect 59126 -50230 59146 -50070
rect 58946 -50250 59146 -50230
rect 59316 -50100 60176 -50090
rect 59316 -50110 59956 -50100
rect 59316 -50250 59336 -50110
rect 59416 -50250 59956 -50110
rect 59316 -50260 59956 -50250
rect 60166 -50260 60176 -50100
rect 59316 -50270 60176 -50260
rect 56506 -50440 57016 -50430
rect 58956 -50320 61136 -50310
rect 58956 -50330 61056 -50320
rect 58956 -50440 58996 -50330
rect 59106 -50340 61056 -50330
rect 59106 -50440 59516 -50340
rect 59616 -50440 61056 -50340
rect 58396 -50530 58896 -50440
rect 58956 -50450 61056 -50440
rect 61126 -50450 61136 -50320
rect 58956 -50460 61136 -50450
rect 55850 -50648 55880 -50618
rect 53940 -50678 55880 -50648
rect 53940 -50698 54920 -50678
rect 53040 -52508 53050 -50758
rect 53250 -52508 53260 -50758
rect 53940 -50798 53950 -50698
rect 54020 -50748 54920 -50698
rect 54020 -50798 54030 -50748
rect 54910 -50768 54920 -50748
rect 54990 -50698 55880 -50678
rect 55970 -50648 55980 -50618
rect 54990 -50748 55970 -50698
rect 54990 -50768 55000 -50748
rect 55220 -51028 55230 -50858
rect 55320 -51028 55330 -50858
rect 55420 -51018 55430 -50848
rect 55510 -50858 55520 -50848
rect 55510 -50868 56670 -50858
rect 55510 -50998 55600 -50868
rect 55710 -50998 56590 -50868
rect 56660 -50998 56670 -50868
rect 55510 -51008 56670 -50998
rect 58396 -50890 58486 -50530
rect 58816 -50550 58896 -50530
rect 59646 -50550 59706 -50530
rect 58816 -50570 59706 -50550
rect 58816 -50630 58906 -50570
rect 58966 -50630 59216 -50570
rect 59276 -50630 59326 -50570
rect 59386 -50630 59436 -50570
rect 59496 -50630 59636 -50570
rect 59696 -50630 59706 -50570
rect 58816 -50640 59706 -50630
rect 58816 -50890 58896 -50640
rect 59536 -50690 59616 -50680
rect 59276 -50730 59356 -50720
rect 59276 -50790 59286 -50730
rect 59346 -50790 59356 -50730
rect 59536 -50750 59546 -50690
rect 59606 -50750 59616 -50690
rect 59536 -50770 59616 -50750
rect 58996 -50800 59076 -50790
rect 58996 -50860 59006 -50800
rect 59076 -50820 59086 -50800
rect 59536 -50810 59616 -50800
rect 59536 -50820 59546 -50810
rect 59076 -50860 59546 -50820
rect 58996 -50870 59076 -50860
rect 59536 -50870 59546 -50860
rect 59606 -50870 59616 -50810
rect 59536 -50880 59616 -50870
rect 58396 -50910 58896 -50890
rect 59646 -50910 59706 -50640
rect 60436 -50720 60536 -50710
rect 59856 -50740 59976 -50730
rect 59856 -50830 59866 -50740
rect 59966 -50830 59976 -50740
rect 60436 -50820 60446 -50720
rect 60526 -50820 60536 -50720
rect 60436 -50830 60536 -50820
rect 59856 -50840 59976 -50830
rect 58396 -50920 59706 -50910
rect 58396 -50930 59216 -50920
rect 58396 -50990 58906 -50930
rect 58966 -50980 59216 -50930
rect 59276 -50980 59336 -50920
rect 59396 -50980 59436 -50920
rect 59496 -50930 59706 -50920
rect 59496 -50980 59636 -50930
rect 58966 -50990 59636 -50980
rect 59696 -50990 59706 -50930
rect 58396 -51000 59706 -50990
rect 60036 -50920 60136 -50910
rect 60036 -51000 60046 -50920
rect 60126 -51000 60136 -50920
rect 55510 -51018 55520 -51008
rect 59646 -51010 59706 -51000
rect 60546 -51010 60636 -51000
rect 59066 -51040 59176 -51030
rect 59066 -51110 59076 -51040
rect 59166 -51110 59176 -51040
rect 59846 -51080 59856 -51010
rect 59916 -51030 59926 -51010
rect 60356 -51020 60556 -51010
rect 60356 -51030 60376 -51020
rect 59916 -51060 60376 -51030
rect 59916 -51080 59926 -51060
rect 60356 -51080 60376 -51060
rect 60446 -51080 60556 -51020
rect 60356 -51090 60556 -51080
rect 60626 -51090 60636 -51010
rect 59066 -51120 59176 -51110
rect 59966 -51100 60326 -51090
rect 53850 -51238 53860 -51128
rect 53920 -51138 55600 -51128
rect 53920 -51238 55000 -51138
rect 55090 -51238 55540 -51138
rect 55630 -51238 55640 -51138
rect 59966 -51160 59976 -51100
rect 60316 -51160 60326 -51100
rect 60546 -51110 60636 -51090
rect 61186 -51120 61366 -51110
rect 54770 -51438 54850 -51238
rect 56470 -51248 56480 -51188
rect 56550 -51248 56560 -51188
rect 57088 -51304 57098 -51164
rect 57368 -51304 57378 -51164
rect 59166 -51230 59376 -51220
rect 59166 -51240 59286 -51230
rect 59166 -51320 59176 -51240
rect 59236 -51320 59286 -51240
rect 59366 -51320 59376 -51230
rect 59166 -51330 59376 -51320
rect 59526 -51270 59646 -51250
rect 59526 -51330 59576 -51270
rect 59636 -51330 59646 -51270
rect 61186 -51300 61206 -51120
rect 61346 -51300 61366 -51120
rect 61186 -51310 61366 -51300
rect 59526 -51360 59646 -51330
rect 60286 -51350 60476 -51340
rect 59906 -51380 60016 -51370
rect 59806 -51390 59866 -51380
rect 54760 -51528 54770 -51438
rect 54840 -51528 54850 -51438
rect 59166 -51440 59536 -51430
rect 59166 -51520 59176 -51440
rect 59236 -51520 59286 -51440
rect 54920 -51538 55210 -51528
rect 54920 -51608 55140 -51538
rect 55200 -51608 55210 -51538
rect 59166 -51530 59286 -51520
rect 59356 -51450 59536 -51440
rect 59356 -51520 59476 -51450
rect 59356 -51530 59536 -51520
rect 59166 -51540 59536 -51530
rect 59566 -51560 59576 -51390
rect 59636 -51400 59866 -51390
rect 59636 -51540 59806 -51400
rect 59636 -51560 59866 -51540
rect 59906 -51560 59916 -51380
rect 60006 -51560 60016 -51380
rect 60286 -51490 60306 -51350
rect 60456 -51490 60476 -51350
rect 60286 -51500 60476 -51490
rect 61026 -51420 61136 -51410
rect 61026 -51530 61036 -51420
rect 61126 -51530 61136 -51420
rect 61026 -51540 61136 -51530
rect 59566 -51570 59636 -51560
rect 59906 -51570 60016 -51560
rect 54760 -51928 54770 -51848
rect 54840 -51928 54850 -51848
rect 54770 -52138 54850 -51928
rect 54920 -51998 54980 -51608
rect 55880 -51638 56900 -51618
rect 55010 -51728 55020 -51648
rect 55120 -51728 55740 -51648
rect 55810 -51728 55820 -51648
rect 55870 -51728 55880 -51638
rect 55970 -51728 56480 -51638
rect 56550 -51728 56900 -51638
rect 55880 -51748 56900 -51728
rect 57020 -51620 57040 -51618
rect 57800 -51620 58240 -51610
rect 57020 -51740 57800 -51620
rect 57020 -51748 57040 -51740
rect 57800 -51750 58240 -51740
rect 58516 -51660 58796 -51590
rect 58516 -51860 58556 -51660
rect 58756 -51860 58796 -51660
rect 59066 -51610 59936 -51600
rect 59066 -51680 59076 -51610
rect 59166 -51630 59826 -51610
rect 59166 -51680 59316 -51630
rect 59066 -51690 59316 -51680
rect 59376 -51680 59826 -51630
rect 59916 -51680 59936 -51610
rect 59376 -51690 59936 -51680
rect 60076 -51680 60196 -51640
rect 59066 -51770 59936 -51760
rect 59066 -51840 59076 -51770
rect 59166 -51840 59206 -51770
rect 59266 -51840 59826 -51770
rect 59926 -51840 59936 -51770
rect 59066 -51850 59936 -51840
rect 60076 -51840 60096 -51680
rect 60176 -51840 60196 -51680
rect 58516 -51940 58796 -51860
rect 60076 -51880 60196 -51840
rect 61266 -51650 61366 -51640
rect 61266 -51860 61276 -51650
rect 61356 -51860 61366 -51650
rect 61266 -51870 61366 -51860
rect 59586 -51890 59656 -51880
rect 59796 -51890 59866 -51880
rect 59586 -51910 59796 -51890
rect 59156 -51920 59536 -51910
rect 59156 -51930 59266 -51920
rect 54910 -52068 54920 -51998
rect 54980 -52068 54990 -51998
rect 59156 -52010 59166 -51930
rect 59226 -52010 59266 -51930
rect 59366 -51930 59536 -51920
rect 59366 -52010 59466 -51930
rect 59526 -52010 59536 -51930
rect 59156 -52030 59536 -52010
rect 59646 -52050 59796 -51910
rect 59586 -52070 59796 -52050
rect 59856 -52070 59866 -51890
rect 53840 -52248 53850 -52138
rect 53920 -52238 55000 -52138
rect 55090 -52238 55540 -52138
rect 55630 -52238 55640 -52138
rect 56470 -52188 56480 -52128
rect 56550 -52188 56560 -52128
rect 57088 -52214 57098 -52074
rect 57368 -52214 57378 -52074
rect 59796 -52080 59866 -52070
rect 59906 -51890 60016 -51880
rect 59906 -52080 59916 -51890
rect 60006 -52080 60016 -51890
rect 60476 -51910 60546 -51900
rect 60536 -51970 60546 -51910
rect 60476 -51980 60546 -51970
rect 60966 -52030 61486 -52020
rect 60966 -52040 61336 -52030
rect 59906 -52090 60016 -52080
rect 60466 -52050 61336 -52040
rect 59506 -52110 59606 -52100
rect 59156 -52160 59376 -52140
rect 53920 -52248 55640 -52238
rect 59156 -52240 59166 -52160
rect 59226 -52240 59266 -52160
rect 59156 -52250 59266 -52240
rect 59366 -52250 59376 -52160
rect 59506 -52180 59516 -52110
rect 59596 -52180 59606 -52110
rect 60466 -52110 60476 -52050
rect 60536 -52110 60616 -52050
rect 60736 -52110 60756 -52050
rect 60816 -52110 60896 -52050
rect 60956 -52110 61336 -52050
rect 60466 -52120 61336 -52110
rect 60966 -52160 61336 -52120
rect 61456 -52160 61486 -52030
rect 60966 -52170 61486 -52160
rect 59506 -52190 59606 -52180
rect 59156 -52260 59376 -52250
rect 59306 -52320 60336 -52300
rect 59066 -52340 59176 -52330
rect 55210 -52518 55220 -52348
rect 55310 -52518 55320 -52348
rect 55400 -52528 55410 -52358
rect 55500 -52368 55510 -52358
rect 55500 -52488 56380 -52368
rect 56440 -52488 56450 -52368
rect 59066 -52400 59076 -52340
rect 59166 -52400 59176 -52340
rect 59306 -52380 59316 -52320
rect 59376 -52340 59966 -52320
rect 59376 -52380 59816 -52340
rect 59306 -52390 59816 -52380
rect 59846 -52380 59916 -52370
rect 59066 -52410 59176 -52400
rect 59846 -52440 59856 -52380
rect 59946 -52380 59966 -52340
rect 60326 -52380 60336 -52320
rect 59946 -52390 60336 -52380
rect 60366 -52340 61146 -52330
rect 60366 -52380 61056 -52340
rect 59646 -52450 59716 -52440
rect 59846 -52450 59916 -52440
rect 60366 -52440 60376 -52380
rect 60436 -52440 61056 -52380
rect 61126 -52440 61146 -52340
rect 55500 -52508 56450 -52488
rect 58396 -52460 59716 -52450
rect 55500 -52528 55510 -52508
rect 58396 -52530 58926 -52460
rect 58986 -52530 59146 -52460
rect 59226 -52530 59276 -52460
rect 59356 -52530 59396 -52460
rect 59476 -52520 59646 -52460
rect 59706 -52520 59716 -52460
rect 60366 -52470 61146 -52440
rect 59476 -52530 59716 -52520
rect 58396 -52540 59716 -52530
rect 54900 -52608 54910 -52598
rect 53940 -52688 53950 -52608
rect 54010 -52688 54910 -52608
rect 53940 -52698 54910 -52688
rect 54980 -52618 54990 -52598
rect 54980 -52678 55980 -52618
rect 54980 -52698 55880 -52678
rect 53940 -52718 55880 -52698
rect 53500 -52848 53510 -52728
rect 53630 -52848 53640 -52728
rect 55850 -52758 55880 -52718
rect 55970 -52758 55980 -52678
rect 55230 -52818 55240 -52758
rect 55370 -52778 55710 -52758
rect 55370 -52788 55720 -52778
rect 55370 -52808 55620 -52788
rect 55370 -52818 55380 -52808
rect 55400 -52868 55410 -52848
rect 54730 -52958 54740 -52868
rect 54850 -52938 55410 -52868
rect 55510 -52938 55520 -52848
rect 55600 -52878 55620 -52808
rect 55710 -52878 55720 -52788
rect 54850 -52958 55520 -52938
rect 55210 -53128 55220 -53018
rect 55330 -53128 55340 -53018
rect 55850 -53178 55980 -52758
rect 56010 -53008 56020 -52858
rect 56080 -53008 56090 -52858
rect 56160 -53008 56170 -52808
rect 56390 -53008 56400 -52808
rect 58396 -52820 58896 -52540
rect 59006 -52700 59076 -52680
rect 59246 -52690 59256 -52630
rect 59366 -52690 59376 -52630
rect 59536 -52660 59546 -52590
rect 59606 -52660 59616 -52590
rect 59536 -52670 59616 -52660
rect 59006 -52760 59016 -52700
rect 59536 -52710 59616 -52700
rect 59076 -52720 59086 -52710
rect 59536 -52720 59546 -52710
rect 59076 -52760 59546 -52720
rect 59006 -52770 59546 -52760
rect 59606 -52770 59616 -52710
rect 59006 -52790 59076 -52770
rect 59536 -52790 59616 -52770
rect 59646 -52820 59716 -52540
rect 59796 -52610 59926 -52600
rect 59796 -52720 59806 -52610
rect 59916 -52720 59926 -52610
rect 59796 -52730 59926 -52720
rect 60436 -52630 60536 -52610
rect 60436 -52750 60446 -52630
rect 60526 -52750 60536 -52630
rect 60436 -52760 60536 -52750
rect 58396 -52830 59716 -52820
rect 56654 -52868 56998 -52858
rect 55520 -53268 55530 -53178
rect 55610 -53268 55980 -53178
rect 54130 -53548 54140 -53288
rect 54850 -53548 54860 -53288
rect 55310 -53468 55320 -53328
rect 55470 -53468 55480 -53328
rect 56170 -53538 56390 -53008
rect 58396 -52900 58906 -52830
rect 58986 -52900 59146 -52830
rect 59226 -52900 59276 -52830
rect 59356 -52900 59396 -52830
rect 59476 -52840 59716 -52830
rect 59476 -52900 59646 -52840
rect 59706 -52900 59716 -52840
rect 58396 -52910 59716 -52900
rect 58396 -52950 58896 -52910
rect 59646 -52920 59716 -52910
rect 56654 -53096 56998 -53086
rect 59006 -53000 60416 -52990
rect 59006 -53040 60266 -53000
rect 59006 -53110 59016 -53040
rect 59076 -53110 59546 -53040
rect 59606 -53110 60266 -53040
rect 59006 -53130 60266 -53110
rect 60406 -53130 60416 -53000
rect 59006 -53140 60416 -53130
rect 59986 -53190 60116 -53180
rect 58956 -53200 59156 -53190
rect 58956 -53380 58966 -53200
rect 59146 -53380 59156 -53200
rect 59986 -53300 59996 -53190
rect 60106 -53300 60116 -53190
rect 58956 -53390 59156 -53380
rect 55680 -53548 56390 -53538
rect 54130 -53708 56390 -53548
rect 55680 -53718 56390 -53708
rect 59600 -53400 60500 -53300
rect 59600 -53800 59700 -53400
rect 60400 -53800 60500 -53400
rect 55300 -53900 56200 -53800
rect 59600 -53900 60500 -53800
rect 64100 -53400 64600 -47900
rect 72810 -47720 73050 -47710
rect 72810 -47900 72820 -47720
rect 73040 -47900 73050 -47720
rect 72810 -47910 73050 -47900
rect 72810 -48000 73050 -47990
rect 64100 -53800 64200 -53400
rect 64500 -53800 64600 -53400
rect 64100 -53900 64600 -53800
rect 65000 -48100 65500 -48000
rect 65000 -48300 65100 -48100
rect 65400 -48300 65500 -48100
rect 72810 -48180 72820 -48000
rect 73040 -48180 73050 -48000
rect 72810 -48190 73050 -48180
rect 55300 -54300 55400 -53900
rect 56100 -54300 56200 -53900
rect 55300 -54400 56200 -54300
rect 51400 -55100 51500 -54900
rect 52500 -55100 52600 -54900
rect 51400 -60300 52600 -55100
rect 55440 -54880 55740 -54860
rect 55440 -55160 55460 -54880
rect 55720 -55160 55740 -54880
rect 55440 -55180 55740 -55160
rect 54140 -55338 56390 -55328
rect 53460 -55540 53800 -55520
rect 53460 -55740 53480 -55540
rect 53780 -55740 53800 -55540
rect 54140 -55578 54150 -55338
rect 54860 -55578 56390 -55338
rect 58946 -55470 59146 -55450
rect 54140 -55588 56390 -55578
rect 53460 -55760 53800 -55740
rect 54850 -55818 55530 -55808
rect 53510 -55968 53520 -55858
rect 53640 -55968 53650 -55858
rect 54740 -55918 54750 -55838
rect 54850 -55888 55430 -55818
rect 55520 -55888 55530 -55818
rect 55950 -55888 55960 -55738
rect 56040 -55888 56050 -55738
rect 56170 -55758 56390 -55588
rect 56506 -55580 57016 -55570
rect 54840 -55918 54850 -55908
rect 55270 -56008 55280 -55918
rect 55400 -56008 55410 -55918
rect 56170 -55968 56190 -55758
rect 56390 -55968 56400 -55758
rect 58946 -55630 58966 -55470
rect 59126 -55630 59146 -55470
rect 58946 -55650 59146 -55630
rect 59316 -55500 60176 -55490
rect 59316 -55510 59956 -55500
rect 59316 -55650 59336 -55510
rect 59416 -55650 59956 -55510
rect 59316 -55660 59956 -55650
rect 60166 -55660 60176 -55500
rect 59316 -55670 60176 -55660
rect 56506 -55840 57016 -55830
rect 58956 -55720 61136 -55710
rect 58956 -55730 61056 -55720
rect 58956 -55840 58996 -55730
rect 59106 -55740 61056 -55730
rect 59106 -55840 59516 -55740
rect 59616 -55840 61056 -55740
rect 58396 -55930 58896 -55840
rect 58956 -55850 61056 -55840
rect 61126 -55850 61136 -55720
rect 58956 -55860 61136 -55850
rect 55850 -56048 55880 -56018
rect 53940 -56078 55880 -56048
rect 53940 -56098 54920 -56078
rect 53040 -57908 53050 -56158
rect 53250 -57908 53260 -56158
rect 53940 -56198 53950 -56098
rect 54020 -56148 54920 -56098
rect 54020 -56198 54030 -56148
rect 54910 -56168 54920 -56148
rect 54990 -56098 55880 -56078
rect 55970 -56048 55980 -56018
rect 54990 -56148 55970 -56098
rect 54990 -56168 55000 -56148
rect 55220 -56428 55230 -56258
rect 55320 -56428 55330 -56258
rect 55420 -56418 55430 -56248
rect 55510 -56258 55520 -56248
rect 55510 -56268 56670 -56258
rect 55510 -56398 55600 -56268
rect 55710 -56398 56590 -56268
rect 56660 -56398 56670 -56268
rect 55510 -56408 56670 -56398
rect 58396 -56290 58486 -55930
rect 58816 -55950 58896 -55930
rect 59646 -55950 59706 -55930
rect 58816 -55970 59706 -55950
rect 58816 -56030 58906 -55970
rect 58966 -56030 59216 -55970
rect 59276 -56030 59326 -55970
rect 59386 -56030 59436 -55970
rect 59496 -56030 59636 -55970
rect 59696 -56030 59706 -55970
rect 58816 -56040 59706 -56030
rect 58816 -56290 58896 -56040
rect 59536 -56090 59616 -56080
rect 59276 -56130 59356 -56120
rect 59276 -56190 59286 -56130
rect 59346 -56190 59356 -56130
rect 59536 -56150 59546 -56090
rect 59606 -56150 59616 -56090
rect 59536 -56170 59616 -56150
rect 58996 -56200 59076 -56190
rect 58996 -56260 59006 -56200
rect 59076 -56220 59086 -56200
rect 59536 -56210 59616 -56200
rect 59536 -56220 59546 -56210
rect 59076 -56260 59546 -56220
rect 58996 -56270 59076 -56260
rect 59536 -56270 59546 -56260
rect 59606 -56270 59616 -56210
rect 59536 -56280 59616 -56270
rect 58396 -56310 58896 -56290
rect 59646 -56310 59706 -56040
rect 60436 -56120 60536 -56110
rect 59856 -56140 59976 -56130
rect 59856 -56230 59866 -56140
rect 59966 -56230 59976 -56140
rect 60436 -56220 60446 -56120
rect 60526 -56220 60536 -56120
rect 60436 -56230 60536 -56220
rect 59856 -56240 59976 -56230
rect 58396 -56320 59706 -56310
rect 58396 -56330 59216 -56320
rect 58396 -56390 58906 -56330
rect 58966 -56380 59216 -56330
rect 59276 -56380 59336 -56320
rect 59396 -56380 59436 -56320
rect 59496 -56330 59706 -56320
rect 59496 -56380 59636 -56330
rect 58966 -56390 59636 -56380
rect 59696 -56390 59706 -56330
rect 58396 -56400 59706 -56390
rect 60036 -56320 60136 -56310
rect 60036 -56400 60046 -56320
rect 60126 -56400 60136 -56320
rect 55510 -56418 55520 -56408
rect 59646 -56410 59706 -56400
rect 60546 -56410 60636 -56400
rect 59066 -56440 59176 -56430
rect 59066 -56510 59076 -56440
rect 59166 -56510 59176 -56440
rect 59846 -56480 59856 -56410
rect 59916 -56430 59926 -56410
rect 60356 -56420 60556 -56410
rect 60356 -56430 60376 -56420
rect 59916 -56460 60376 -56430
rect 59916 -56480 59926 -56460
rect 60356 -56480 60376 -56460
rect 60446 -56480 60556 -56420
rect 60356 -56490 60556 -56480
rect 60626 -56490 60636 -56410
rect 59066 -56520 59176 -56510
rect 59966 -56500 60326 -56490
rect 53850 -56638 53860 -56528
rect 53920 -56538 55600 -56528
rect 53920 -56638 55000 -56538
rect 55090 -56638 55540 -56538
rect 55630 -56638 55640 -56538
rect 59966 -56560 59976 -56500
rect 60316 -56560 60326 -56500
rect 60546 -56510 60636 -56490
rect 61186 -56520 61366 -56510
rect 54770 -56838 54850 -56638
rect 56470 -56648 56480 -56588
rect 56550 -56648 56560 -56588
rect 57088 -56704 57098 -56564
rect 57368 -56704 57378 -56564
rect 59166 -56630 59376 -56620
rect 59166 -56640 59286 -56630
rect 59166 -56720 59176 -56640
rect 59236 -56720 59286 -56640
rect 59366 -56720 59376 -56630
rect 59166 -56730 59376 -56720
rect 59526 -56670 59646 -56650
rect 59526 -56730 59576 -56670
rect 59636 -56730 59646 -56670
rect 61186 -56700 61206 -56520
rect 61346 -56700 61366 -56520
rect 61186 -56710 61366 -56700
rect 59526 -56760 59646 -56730
rect 60286 -56750 60476 -56740
rect 59906 -56780 60016 -56770
rect 59806 -56790 59866 -56780
rect 54760 -56928 54770 -56838
rect 54840 -56928 54850 -56838
rect 59166 -56840 59536 -56830
rect 59166 -56920 59176 -56840
rect 59236 -56920 59286 -56840
rect 54920 -56938 55210 -56928
rect 54920 -57008 55140 -56938
rect 55200 -57008 55210 -56938
rect 59166 -56930 59286 -56920
rect 59356 -56850 59536 -56840
rect 59356 -56920 59476 -56850
rect 59356 -56930 59536 -56920
rect 59166 -56940 59536 -56930
rect 59566 -56960 59576 -56790
rect 59636 -56800 59866 -56790
rect 59636 -56940 59806 -56800
rect 59636 -56960 59866 -56940
rect 59906 -56960 59916 -56780
rect 60006 -56960 60016 -56780
rect 60286 -56890 60306 -56750
rect 60456 -56890 60476 -56750
rect 60286 -56900 60476 -56890
rect 61026 -56820 61136 -56810
rect 61026 -56930 61036 -56820
rect 61126 -56930 61136 -56820
rect 61026 -56940 61136 -56930
rect 59566 -56970 59636 -56960
rect 59906 -56970 60016 -56960
rect 54760 -57328 54770 -57248
rect 54840 -57328 54850 -57248
rect 54770 -57538 54850 -57328
rect 54920 -57398 54980 -57008
rect 55880 -57038 56900 -57018
rect 55010 -57128 55020 -57048
rect 55120 -57128 55740 -57048
rect 55810 -57128 55820 -57048
rect 55870 -57128 55880 -57038
rect 55970 -57128 56480 -57038
rect 56550 -57128 56900 -57038
rect 55880 -57148 56900 -57128
rect 57020 -57020 57040 -57018
rect 57800 -57020 58240 -57010
rect 57020 -57140 57800 -57020
rect 57020 -57148 57040 -57140
rect 57800 -57150 58240 -57140
rect 58516 -57060 58796 -56990
rect 58516 -57260 58556 -57060
rect 58756 -57260 58796 -57060
rect 59066 -57010 59936 -57000
rect 59066 -57080 59076 -57010
rect 59166 -57030 59826 -57010
rect 59166 -57080 59316 -57030
rect 59066 -57090 59316 -57080
rect 59376 -57080 59826 -57030
rect 59916 -57080 59936 -57010
rect 59376 -57090 59936 -57080
rect 60076 -57080 60196 -57040
rect 59066 -57170 59936 -57160
rect 59066 -57240 59076 -57170
rect 59166 -57240 59206 -57170
rect 59266 -57240 59826 -57170
rect 59926 -57240 59936 -57170
rect 59066 -57250 59936 -57240
rect 60076 -57240 60096 -57080
rect 60176 -57240 60196 -57080
rect 58516 -57340 58796 -57260
rect 60076 -57280 60196 -57240
rect 61266 -57050 61366 -57040
rect 61266 -57260 61276 -57050
rect 61356 -57260 61366 -57050
rect 61266 -57270 61366 -57260
rect 59586 -57290 59656 -57280
rect 59796 -57290 59866 -57280
rect 59586 -57310 59796 -57290
rect 59156 -57320 59536 -57310
rect 59156 -57330 59266 -57320
rect 54910 -57468 54920 -57398
rect 54980 -57468 54990 -57398
rect 59156 -57410 59166 -57330
rect 59226 -57410 59266 -57330
rect 59366 -57330 59536 -57320
rect 59366 -57410 59466 -57330
rect 59526 -57410 59536 -57330
rect 59156 -57430 59536 -57410
rect 59646 -57450 59796 -57310
rect 59586 -57470 59796 -57450
rect 59856 -57470 59866 -57290
rect 53840 -57648 53850 -57538
rect 53920 -57638 55000 -57538
rect 55090 -57638 55540 -57538
rect 55630 -57638 55640 -57538
rect 56470 -57588 56480 -57528
rect 56550 -57588 56560 -57528
rect 57088 -57614 57098 -57474
rect 57368 -57614 57378 -57474
rect 59796 -57480 59866 -57470
rect 59906 -57290 60016 -57280
rect 59906 -57480 59916 -57290
rect 60006 -57480 60016 -57290
rect 60476 -57310 60546 -57300
rect 60536 -57370 60546 -57310
rect 60476 -57380 60546 -57370
rect 60966 -57430 61486 -57420
rect 60966 -57440 61336 -57430
rect 59906 -57490 60016 -57480
rect 60466 -57450 61336 -57440
rect 59506 -57510 59606 -57500
rect 59156 -57560 59376 -57540
rect 53920 -57648 55640 -57638
rect 59156 -57640 59166 -57560
rect 59226 -57640 59266 -57560
rect 59156 -57650 59266 -57640
rect 59366 -57650 59376 -57560
rect 59506 -57580 59516 -57510
rect 59596 -57580 59606 -57510
rect 60466 -57510 60476 -57450
rect 60536 -57510 60616 -57450
rect 60736 -57510 60756 -57450
rect 60816 -57510 60896 -57450
rect 60956 -57510 61336 -57450
rect 60466 -57520 61336 -57510
rect 60966 -57560 61336 -57520
rect 61456 -57560 61486 -57430
rect 60966 -57570 61486 -57560
rect 59506 -57590 59606 -57580
rect 59156 -57660 59376 -57650
rect 59306 -57720 60336 -57700
rect 59066 -57740 59176 -57730
rect 55210 -57918 55220 -57748
rect 55310 -57918 55320 -57748
rect 55400 -57928 55410 -57758
rect 55500 -57768 55510 -57758
rect 55500 -57888 56380 -57768
rect 56440 -57888 56450 -57768
rect 59066 -57800 59076 -57740
rect 59166 -57800 59176 -57740
rect 59306 -57780 59316 -57720
rect 59376 -57740 59966 -57720
rect 59376 -57780 59816 -57740
rect 59306 -57790 59816 -57780
rect 59846 -57780 59916 -57770
rect 59066 -57810 59176 -57800
rect 59846 -57840 59856 -57780
rect 59946 -57780 59966 -57740
rect 60326 -57780 60336 -57720
rect 59946 -57790 60336 -57780
rect 60366 -57740 61146 -57730
rect 60366 -57780 61056 -57740
rect 59646 -57850 59716 -57840
rect 59846 -57850 59916 -57840
rect 60366 -57840 60376 -57780
rect 60436 -57840 61056 -57780
rect 61126 -57840 61146 -57740
rect 55500 -57908 56450 -57888
rect 58396 -57860 59716 -57850
rect 55500 -57928 55510 -57908
rect 58396 -57930 58926 -57860
rect 58986 -57930 59146 -57860
rect 59226 -57930 59276 -57860
rect 59356 -57930 59396 -57860
rect 59476 -57920 59646 -57860
rect 59706 -57920 59716 -57860
rect 60366 -57870 61146 -57840
rect 59476 -57930 59716 -57920
rect 58396 -57940 59716 -57930
rect 54900 -58008 54910 -57998
rect 53940 -58088 53950 -58008
rect 54010 -58088 54910 -58008
rect 53940 -58098 54910 -58088
rect 54980 -58018 54990 -57998
rect 54980 -58078 55980 -58018
rect 54980 -58098 55880 -58078
rect 53940 -58118 55880 -58098
rect 53500 -58248 53510 -58128
rect 53630 -58248 53640 -58128
rect 55850 -58158 55880 -58118
rect 55970 -58158 55980 -58078
rect 55230 -58218 55240 -58158
rect 55370 -58178 55710 -58158
rect 55370 -58188 55720 -58178
rect 55370 -58208 55620 -58188
rect 55370 -58218 55380 -58208
rect 55400 -58268 55410 -58248
rect 54730 -58358 54740 -58268
rect 54850 -58338 55410 -58268
rect 55510 -58338 55520 -58248
rect 55600 -58278 55620 -58208
rect 55710 -58278 55720 -58188
rect 54850 -58358 55520 -58338
rect 55210 -58528 55220 -58418
rect 55330 -58528 55340 -58418
rect 55850 -58578 55980 -58158
rect 56010 -58408 56020 -58258
rect 56080 -58408 56090 -58258
rect 56160 -58408 56170 -58208
rect 56390 -58408 56400 -58208
rect 58396 -58220 58896 -57940
rect 59006 -58100 59076 -58080
rect 59246 -58090 59256 -58030
rect 59366 -58090 59376 -58030
rect 59536 -58060 59546 -57990
rect 59606 -58060 59616 -57990
rect 59536 -58070 59616 -58060
rect 59006 -58160 59016 -58100
rect 59536 -58110 59616 -58100
rect 59076 -58120 59086 -58110
rect 59536 -58120 59546 -58110
rect 59076 -58160 59546 -58120
rect 59006 -58170 59546 -58160
rect 59606 -58170 59616 -58110
rect 59006 -58190 59076 -58170
rect 59536 -58190 59616 -58170
rect 59646 -58220 59716 -57940
rect 59796 -58010 59926 -58000
rect 59796 -58120 59806 -58010
rect 59916 -58120 59926 -58010
rect 59796 -58130 59926 -58120
rect 60436 -58030 60536 -58010
rect 60436 -58150 60446 -58030
rect 60526 -58150 60536 -58030
rect 60436 -58160 60536 -58150
rect 58396 -58230 59716 -58220
rect 56654 -58268 56998 -58258
rect 55520 -58668 55530 -58578
rect 55610 -58668 55980 -58578
rect 54130 -58948 54140 -58688
rect 54850 -58948 54860 -58688
rect 55310 -58868 55320 -58728
rect 55470 -58868 55480 -58728
rect 56170 -58938 56390 -58408
rect 58396 -58300 58906 -58230
rect 58986 -58300 59146 -58230
rect 59226 -58300 59276 -58230
rect 59356 -58300 59396 -58230
rect 59476 -58240 59716 -58230
rect 59476 -58300 59646 -58240
rect 59706 -58300 59716 -58240
rect 58396 -58310 59716 -58300
rect 58396 -58350 58896 -58310
rect 59646 -58320 59716 -58310
rect 56654 -58496 56998 -58486
rect 59006 -58400 60416 -58390
rect 59006 -58440 60266 -58400
rect 59006 -58510 59016 -58440
rect 59076 -58510 59546 -58440
rect 59606 -58510 60266 -58440
rect 59006 -58530 60266 -58510
rect 60406 -58530 60416 -58400
rect 59006 -58540 60416 -58530
rect 59986 -58590 60116 -58580
rect 58956 -58600 59156 -58590
rect 58956 -58780 58966 -58600
rect 59146 -58780 59156 -58600
rect 59986 -58700 59996 -58590
rect 60106 -58700 60116 -58590
rect 58956 -58790 59156 -58780
rect 55680 -58948 56390 -58938
rect 54130 -59108 56390 -58948
rect 55680 -59118 56390 -59108
rect 59600 -58800 60500 -58700
rect 59600 -59200 59700 -58800
rect 60400 -59200 60500 -58800
rect 55400 -59300 56200 -59200
rect 59600 -59300 60500 -59200
rect 65000 -58800 65500 -48300
rect 65000 -59200 65100 -58800
rect 65400 -59200 65500 -58800
rect 65000 -59300 65500 -59200
rect 66000 -48500 66500 -48400
rect 66000 -48700 66100 -48500
rect 66400 -48700 66500 -48500
rect 72810 -48460 73050 -48450
rect 72810 -48640 72820 -48460
rect 73040 -48640 73050 -48460
rect 72810 -48650 73050 -48640
rect 55400 -59700 55500 -59300
rect 56100 -59700 56200 -59300
rect 55400 -59800 56200 -59700
rect 51400 -60500 51500 -60300
rect 52500 -60500 52600 -60300
rect 51400 -65700 52600 -60500
rect 55440 -60280 55740 -60260
rect 55440 -60560 55460 -60280
rect 55720 -60560 55740 -60280
rect 55440 -60580 55740 -60560
rect 54140 -60738 56390 -60728
rect 53460 -60940 53800 -60920
rect 53460 -61140 53480 -60940
rect 53780 -61140 53800 -60940
rect 54140 -60978 54150 -60738
rect 54860 -60978 56390 -60738
rect 58946 -60870 59146 -60850
rect 54140 -60988 56390 -60978
rect 53460 -61160 53800 -61140
rect 54850 -61218 55530 -61208
rect 53510 -61368 53520 -61258
rect 53640 -61368 53650 -61258
rect 54740 -61318 54750 -61238
rect 54850 -61288 55430 -61218
rect 55520 -61288 55530 -61218
rect 55950 -61288 55960 -61138
rect 56040 -61288 56050 -61138
rect 56170 -61158 56390 -60988
rect 56506 -60980 57016 -60970
rect 54840 -61318 54850 -61308
rect 55270 -61408 55280 -61318
rect 55400 -61408 55410 -61318
rect 56170 -61368 56190 -61158
rect 56390 -61368 56400 -61158
rect 58946 -61030 58966 -60870
rect 59126 -61030 59146 -60870
rect 58946 -61050 59146 -61030
rect 59316 -60900 60176 -60890
rect 59316 -60910 59956 -60900
rect 59316 -61050 59336 -60910
rect 59416 -61050 59956 -60910
rect 59316 -61060 59956 -61050
rect 60166 -61060 60176 -60900
rect 59316 -61070 60176 -61060
rect 56506 -61240 57016 -61230
rect 58956 -61120 61136 -61110
rect 58956 -61130 61056 -61120
rect 58956 -61240 58996 -61130
rect 59106 -61140 61056 -61130
rect 59106 -61240 59516 -61140
rect 59616 -61240 61056 -61140
rect 58396 -61330 58896 -61240
rect 58956 -61250 61056 -61240
rect 61126 -61250 61136 -61120
rect 58956 -61260 61136 -61250
rect 55850 -61448 55880 -61418
rect 53940 -61478 55880 -61448
rect 53940 -61498 54920 -61478
rect 53040 -63308 53050 -61558
rect 53250 -63308 53260 -61558
rect 53940 -61598 53950 -61498
rect 54020 -61548 54920 -61498
rect 54020 -61598 54030 -61548
rect 54910 -61568 54920 -61548
rect 54990 -61498 55880 -61478
rect 55970 -61448 55980 -61418
rect 54990 -61548 55970 -61498
rect 54990 -61568 55000 -61548
rect 55220 -61828 55230 -61658
rect 55320 -61828 55330 -61658
rect 55420 -61818 55430 -61648
rect 55510 -61658 55520 -61648
rect 55510 -61668 56670 -61658
rect 55510 -61798 55600 -61668
rect 55710 -61798 56590 -61668
rect 56660 -61798 56670 -61668
rect 55510 -61808 56670 -61798
rect 58396 -61690 58486 -61330
rect 58816 -61350 58896 -61330
rect 59646 -61350 59706 -61330
rect 58816 -61370 59706 -61350
rect 58816 -61430 58906 -61370
rect 58966 -61430 59216 -61370
rect 59276 -61430 59326 -61370
rect 59386 -61430 59436 -61370
rect 59496 -61430 59636 -61370
rect 59696 -61430 59706 -61370
rect 58816 -61440 59706 -61430
rect 58816 -61690 58896 -61440
rect 59536 -61490 59616 -61480
rect 59276 -61530 59356 -61520
rect 59276 -61590 59286 -61530
rect 59346 -61590 59356 -61530
rect 59536 -61550 59546 -61490
rect 59606 -61550 59616 -61490
rect 59536 -61570 59616 -61550
rect 58996 -61600 59076 -61590
rect 58996 -61660 59006 -61600
rect 59076 -61620 59086 -61600
rect 59536 -61610 59616 -61600
rect 59536 -61620 59546 -61610
rect 59076 -61660 59546 -61620
rect 58996 -61670 59076 -61660
rect 59536 -61670 59546 -61660
rect 59606 -61670 59616 -61610
rect 59536 -61680 59616 -61670
rect 58396 -61710 58896 -61690
rect 59646 -61710 59706 -61440
rect 60436 -61520 60536 -61510
rect 59856 -61540 59976 -61530
rect 59856 -61630 59866 -61540
rect 59966 -61630 59976 -61540
rect 60436 -61620 60446 -61520
rect 60526 -61620 60536 -61520
rect 60436 -61630 60536 -61620
rect 59856 -61640 59976 -61630
rect 58396 -61720 59706 -61710
rect 58396 -61730 59216 -61720
rect 58396 -61790 58906 -61730
rect 58966 -61780 59216 -61730
rect 59276 -61780 59336 -61720
rect 59396 -61780 59436 -61720
rect 59496 -61730 59706 -61720
rect 59496 -61780 59636 -61730
rect 58966 -61790 59636 -61780
rect 59696 -61790 59706 -61730
rect 58396 -61800 59706 -61790
rect 60036 -61720 60136 -61710
rect 60036 -61800 60046 -61720
rect 60126 -61800 60136 -61720
rect 55510 -61818 55520 -61808
rect 59646 -61810 59706 -61800
rect 60546 -61810 60636 -61800
rect 59066 -61840 59176 -61830
rect 59066 -61910 59076 -61840
rect 59166 -61910 59176 -61840
rect 59846 -61880 59856 -61810
rect 59916 -61830 59926 -61810
rect 60356 -61820 60556 -61810
rect 60356 -61830 60376 -61820
rect 59916 -61860 60376 -61830
rect 59916 -61880 59926 -61860
rect 60356 -61880 60376 -61860
rect 60446 -61880 60556 -61820
rect 60356 -61890 60556 -61880
rect 60626 -61890 60636 -61810
rect 59066 -61920 59176 -61910
rect 59966 -61900 60326 -61890
rect 53850 -62038 53860 -61928
rect 53920 -61938 55600 -61928
rect 53920 -62038 55000 -61938
rect 55090 -62038 55540 -61938
rect 55630 -62038 55640 -61938
rect 59966 -61960 59976 -61900
rect 60316 -61960 60326 -61900
rect 60546 -61910 60636 -61890
rect 61186 -61920 61366 -61910
rect 54770 -62238 54850 -62038
rect 56470 -62048 56480 -61988
rect 56550 -62048 56560 -61988
rect 57088 -62104 57098 -61964
rect 57368 -62104 57378 -61964
rect 59166 -62030 59376 -62020
rect 59166 -62040 59286 -62030
rect 59166 -62120 59176 -62040
rect 59236 -62120 59286 -62040
rect 59366 -62120 59376 -62030
rect 59166 -62130 59376 -62120
rect 59526 -62070 59646 -62050
rect 59526 -62130 59576 -62070
rect 59636 -62130 59646 -62070
rect 61186 -62100 61206 -61920
rect 61346 -62100 61366 -61920
rect 61186 -62110 61366 -62100
rect 59526 -62160 59646 -62130
rect 60286 -62150 60476 -62140
rect 59906 -62180 60016 -62170
rect 59806 -62190 59866 -62180
rect 54760 -62328 54770 -62238
rect 54840 -62328 54850 -62238
rect 59166 -62240 59536 -62230
rect 59166 -62320 59176 -62240
rect 59236 -62320 59286 -62240
rect 54920 -62338 55210 -62328
rect 54920 -62408 55140 -62338
rect 55200 -62408 55210 -62338
rect 59166 -62330 59286 -62320
rect 59356 -62250 59536 -62240
rect 59356 -62320 59476 -62250
rect 59356 -62330 59536 -62320
rect 59166 -62340 59536 -62330
rect 59566 -62360 59576 -62190
rect 59636 -62200 59866 -62190
rect 59636 -62340 59806 -62200
rect 59636 -62360 59866 -62340
rect 59906 -62360 59916 -62180
rect 60006 -62360 60016 -62180
rect 60286 -62290 60306 -62150
rect 60456 -62290 60476 -62150
rect 60286 -62300 60476 -62290
rect 61026 -62220 61136 -62210
rect 61026 -62330 61036 -62220
rect 61126 -62330 61136 -62220
rect 61026 -62340 61136 -62330
rect 59566 -62370 59636 -62360
rect 59906 -62370 60016 -62360
rect 54760 -62728 54770 -62648
rect 54840 -62728 54850 -62648
rect 54770 -62938 54850 -62728
rect 54920 -62798 54980 -62408
rect 55880 -62438 56900 -62418
rect 55010 -62528 55020 -62448
rect 55120 -62528 55740 -62448
rect 55810 -62528 55820 -62448
rect 55870 -62528 55880 -62438
rect 55970 -62528 56480 -62438
rect 56550 -62528 56900 -62438
rect 55880 -62548 56900 -62528
rect 57020 -62420 57040 -62418
rect 57800 -62420 58240 -62410
rect 57020 -62540 57800 -62420
rect 57020 -62548 57040 -62540
rect 57800 -62550 58240 -62540
rect 58516 -62460 58796 -62390
rect 58516 -62660 58556 -62460
rect 58756 -62660 58796 -62460
rect 59066 -62410 59936 -62400
rect 59066 -62480 59076 -62410
rect 59166 -62430 59826 -62410
rect 59166 -62480 59316 -62430
rect 59066 -62490 59316 -62480
rect 59376 -62480 59826 -62430
rect 59916 -62480 59936 -62410
rect 59376 -62490 59936 -62480
rect 60076 -62480 60196 -62440
rect 59066 -62570 59936 -62560
rect 59066 -62640 59076 -62570
rect 59166 -62640 59206 -62570
rect 59266 -62640 59826 -62570
rect 59926 -62640 59936 -62570
rect 59066 -62650 59936 -62640
rect 60076 -62640 60096 -62480
rect 60176 -62640 60196 -62480
rect 58516 -62740 58796 -62660
rect 60076 -62680 60196 -62640
rect 61266 -62450 61366 -62440
rect 61266 -62660 61276 -62450
rect 61356 -62660 61366 -62450
rect 61266 -62670 61366 -62660
rect 59586 -62690 59656 -62680
rect 59796 -62690 59866 -62680
rect 59586 -62710 59796 -62690
rect 59156 -62720 59536 -62710
rect 59156 -62730 59266 -62720
rect 54910 -62868 54920 -62798
rect 54980 -62868 54990 -62798
rect 59156 -62810 59166 -62730
rect 59226 -62810 59266 -62730
rect 59366 -62730 59536 -62720
rect 59366 -62810 59466 -62730
rect 59526 -62810 59536 -62730
rect 59156 -62830 59536 -62810
rect 59646 -62850 59796 -62710
rect 59586 -62870 59796 -62850
rect 59856 -62870 59866 -62690
rect 53840 -63048 53850 -62938
rect 53920 -63038 55000 -62938
rect 55090 -63038 55540 -62938
rect 55630 -63038 55640 -62938
rect 56470 -62988 56480 -62928
rect 56550 -62988 56560 -62928
rect 57088 -63014 57098 -62874
rect 57368 -63014 57378 -62874
rect 59796 -62880 59866 -62870
rect 59906 -62690 60016 -62680
rect 59906 -62880 59916 -62690
rect 60006 -62880 60016 -62690
rect 60476 -62710 60546 -62700
rect 60536 -62770 60546 -62710
rect 60476 -62780 60546 -62770
rect 60966 -62830 61486 -62820
rect 60966 -62840 61336 -62830
rect 59906 -62890 60016 -62880
rect 60466 -62850 61336 -62840
rect 59506 -62910 59606 -62900
rect 59156 -62960 59376 -62940
rect 53920 -63048 55640 -63038
rect 59156 -63040 59166 -62960
rect 59226 -63040 59266 -62960
rect 59156 -63050 59266 -63040
rect 59366 -63050 59376 -62960
rect 59506 -62980 59516 -62910
rect 59596 -62980 59606 -62910
rect 60466 -62910 60476 -62850
rect 60536 -62910 60616 -62850
rect 60736 -62910 60756 -62850
rect 60816 -62910 60896 -62850
rect 60956 -62910 61336 -62850
rect 60466 -62920 61336 -62910
rect 60966 -62960 61336 -62920
rect 61456 -62960 61486 -62830
rect 60966 -62970 61486 -62960
rect 59506 -62990 59606 -62980
rect 59156 -63060 59376 -63050
rect 59306 -63120 60336 -63100
rect 59066 -63140 59176 -63130
rect 55210 -63318 55220 -63148
rect 55310 -63318 55320 -63148
rect 55400 -63328 55410 -63158
rect 55500 -63168 55510 -63158
rect 55500 -63288 56380 -63168
rect 56440 -63288 56450 -63168
rect 59066 -63200 59076 -63140
rect 59166 -63200 59176 -63140
rect 59306 -63180 59316 -63120
rect 59376 -63140 59966 -63120
rect 59376 -63180 59816 -63140
rect 59306 -63190 59816 -63180
rect 59846 -63180 59916 -63170
rect 59066 -63210 59176 -63200
rect 59846 -63240 59856 -63180
rect 59946 -63180 59966 -63140
rect 60326 -63180 60336 -63120
rect 59946 -63190 60336 -63180
rect 60366 -63140 61146 -63130
rect 60366 -63180 61056 -63140
rect 59646 -63250 59716 -63240
rect 59846 -63250 59916 -63240
rect 60366 -63240 60376 -63180
rect 60436 -63240 61056 -63180
rect 61126 -63240 61146 -63140
rect 55500 -63308 56450 -63288
rect 58396 -63260 59716 -63250
rect 55500 -63328 55510 -63308
rect 58396 -63330 58926 -63260
rect 58986 -63330 59146 -63260
rect 59226 -63330 59276 -63260
rect 59356 -63330 59396 -63260
rect 59476 -63320 59646 -63260
rect 59706 -63320 59716 -63260
rect 60366 -63270 61146 -63240
rect 59476 -63330 59716 -63320
rect 58396 -63340 59716 -63330
rect 54900 -63408 54910 -63398
rect 53940 -63488 53950 -63408
rect 54010 -63488 54910 -63408
rect 53940 -63498 54910 -63488
rect 54980 -63418 54990 -63398
rect 54980 -63478 55980 -63418
rect 54980 -63498 55880 -63478
rect 53940 -63518 55880 -63498
rect 53500 -63648 53510 -63528
rect 53630 -63648 53640 -63528
rect 55850 -63558 55880 -63518
rect 55970 -63558 55980 -63478
rect 55230 -63618 55240 -63558
rect 55370 -63578 55710 -63558
rect 55370 -63588 55720 -63578
rect 55370 -63608 55620 -63588
rect 55370 -63618 55380 -63608
rect 55400 -63668 55410 -63648
rect 54730 -63758 54740 -63668
rect 54850 -63738 55410 -63668
rect 55510 -63738 55520 -63648
rect 55600 -63678 55620 -63608
rect 55710 -63678 55720 -63588
rect 54850 -63758 55520 -63738
rect 55210 -63928 55220 -63818
rect 55330 -63928 55340 -63818
rect 55850 -63978 55980 -63558
rect 56010 -63808 56020 -63658
rect 56080 -63808 56090 -63658
rect 56160 -63808 56170 -63608
rect 56390 -63808 56400 -63608
rect 58396 -63620 58896 -63340
rect 59006 -63500 59076 -63480
rect 59246 -63490 59256 -63430
rect 59366 -63490 59376 -63430
rect 59536 -63460 59546 -63390
rect 59606 -63460 59616 -63390
rect 59536 -63470 59616 -63460
rect 59006 -63560 59016 -63500
rect 59536 -63510 59616 -63500
rect 59076 -63520 59086 -63510
rect 59536 -63520 59546 -63510
rect 59076 -63560 59546 -63520
rect 59006 -63570 59546 -63560
rect 59606 -63570 59616 -63510
rect 59006 -63590 59076 -63570
rect 59536 -63590 59616 -63570
rect 59646 -63620 59716 -63340
rect 59796 -63410 59926 -63400
rect 59796 -63520 59806 -63410
rect 59916 -63520 59926 -63410
rect 59796 -63530 59926 -63520
rect 60436 -63430 60536 -63410
rect 60436 -63550 60446 -63430
rect 60526 -63550 60536 -63430
rect 60436 -63560 60536 -63550
rect 58396 -63630 59716 -63620
rect 56654 -63668 56998 -63658
rect 55520 -64068 55530 -63978
rect 55610 -64068 55980 -63978
rect 54130 -64348 54140 -64088
rect 54850 -64348 54860 -64088
rect 55310 -64268 55320 -64128
rect 55470 -64268 55480 -64128
rect 56170 -64338 56390 -63808
rect 58396 -63700 58906 -63630
rect 58986 -63700 59146 -63630
rect 59226 -63700 59276 -63630
rect 59356 -63700 59396 -63630
rect 59476 -63640 59716 -63630
rect 59476 -63700 59646 -63640
rect 59706 -63700 59716 -63640
rect 58396 -63710 59716 -63700
rect 58396 -63750 58896 -63710
rect 59646 -63720 59716 -63710
rect 56654 -63896 56998 -63886
rect 59006 -63800 60416 -63790
rect 59006 -63840 60266 -63800
rect 59006 -63910 59016 -63840
rect 59076 -63910 59546 -63840
rect 59606 -63910 60266 -63840
rect 59006 -63930 60266 -63910
rect 60406 -63930 60416 -63800
rect 59006 -63940 60416 -63930
rect 59986 -63990 60116 -63980
rect 58956 -64000 59156 -63990
rect 58956 -64180 58966 -64000
rect 59146 -64180 59156 -64000
rect 59986 -64100 59996 -63990
rect 60106 -64100 60116 -63990
rect 58956 -64190 59156 -64180
rect 55680 -64348 56390 -64338
rect 54130 -64508 56390 -64348
rect 55680 -64518 56390 -64508
rect 59600 -64200 60500 -64100
rect 59600 -64600 59700 -64200
rect 60400 -64600 60500 -64200
rect 55400 -64700 56200 -64600
rect 59600 -64700 60500 -64600
rect 66000 -64200 66500 -48700
rect 66000 -64600 66100 -64200
rect 66400 -64600 66500 -64200
rect 66000 -64700 66500 -64600
rect 67000 -48900 67500 -48800
rect 67000 -49100 67100 -48900
rect 67400 -49100 67500 -48900
rect 72810 -48820 73050 -48810
rect 72810 -49000 72820 -48820
rect 73040 -49000 73050 -48820
rect 72810 -49010 73050 -49000
rect 55400 -65100 55500 -64700
rect 56100 -65100 56200 -64700
rect 55400 -65200 56200 -65100
rect 51400 -65900 51500 -65700
rect 52500 -65900 52600 -65700
rect 51400 -71100 52600 -65900
rect 55420 -65680 55740 -65660
rect 55420 -65960 55440 -65680
rect 55720 -65960 55740 -65680
rect 55420 -65980 55740 -65960
rect 54140 -66138 56390 -66128
rect 53460 -66340 53800 -66320
rect 53460 -66540 53480 -66340
rect 53780 -66540 53800 -66340
rect 54140 -66378 54150 -66138
rect 54860 -66378 56390 -66138
rect 58946 -66270 59146 -66250
rect 54140 -66388 56390 -66378
rect 53460 -66560 53800 -66540
rect 54850 -66618 55530 -66608
rect 53510 -66768 53520 -66658
rect 53640 -66768 53650 -66658
rect 54740 -66718 54750 -66638
rect 54850 -66688 55430 -66618
rect 55520 -66688 55530 -66618
rect 55950 -66688 55960 -66538
rect 56040 -66688 56050 -66538
rect 56170 -66558 56390 -66388
rect 56506 -66380 57016 -66370
rect 54840 -66718 54850 -66708
rect 55270 -66808 55280 -66718
rect 55400 -66808 55410 -66718
rect 56170 -66768 56190 -66558
rect 56390 -66768 56400 -66558
rect 58946 -66430 58966 -66270
rect 59126 -66430 59146 -66270
rect 58946 -66450 59146 -66430
rect 59316 -66300 60176 -66290
rect 59316 -66310 59956 -66300
rect 59316 -66450 59336 -66310
rect 59416 -66450 59956 -66310
rect 59316 -66460 59956 -66450
rect 60166 -66460 60176 -66300
rect 59316 -66470 60176 -66460
rect 56506 -66640 57016 -66630
rect 58956 -66520 61136 -66510
rect 58956 -66530 61056 -66520
rect 58956 -66640 58996 -66530
rect 59106 -66540 61056 -66530
rect 59106 -66640 59516 -66540
rect 59616 -66640 61056 -66540
rect 58396 -66730 58896 -66640
rect 58956 -66650 61056 -66640
rect 61126 -66650 61136 -66520
rect 58956 -66660 61136 -66650
rect 55850 -66848 55880 -66818
rect 53940 -66878 55880 -66848
rect 53940 -66898 54920 -66878
rect 53040 -68708 53050 -66958
rect 53250 -68708 53260 -66958
rect 53940 -66998 53950 -66898
rect 54020 -66948 54920 -66898
rect 54020 -66998 54030 -66948
rect 54910 -66968 54920 -66948
rect 54990 -66898 55880 -66878
rect 55970 -66848 55980 -66818
rect 54990 -66948 55970 -66898
rect 54990 -66968 55000 -66948
rect 55220 -67228 55230 -67058
rect 55320 -67228 55330 -67058
rect 55420 -67218 55430 -67048
rect 55510 -67058 55520 -67048
rect 55510 -67068 56670 -67058
rect 55510 -67198 55600 -67068
rect 55710 -67198 56590 -67068
rect 56660 -67198 56670 -67068
rect 55510 -67208 56670 -67198
rect 58396 -67090 58486 -66730
rect 58816 -66750 58896 -66730
rect 59646 -66750 59706 -66730
rect 58816 -66770 59706 -66750
rect 58816 -66830 58906 -66770
rect 58966 -66830 59216 -66770
rect 59276 -66830 59326 -66770
rect 59386 -66830 59436 -66770
rect 59496 -66830 59636 -66770
rect 59696 -66830 59706 -66770
rect 58816 -66840 59706 -66830
rect 58816 -67090 58896 -66840
rect 59536 -66890 59616 -66880
rect 59276 -66930 59356 -66920
rect 59276 -66990 59286 -66930
rect 59346 -66990 59356 -66930
rect 59536 -66950 59546 -66890
rect 59606 -66950 59616 -66890
rect 59536 -66970 59616 -66950
rect 58996 -67000 59076 -66990
rect 58996 -67060 59006 -67000
rect 59076 -67020 59086 -67000
rect 59536 -67010 59616 -67000
rect 59536 -67020 59546 -67010
rect 59076 -67060 59546 -67020
rect 58996 -67070 59076 -67060
rect 59536 -67070 59546 -67060
rect 59606 -67070 59616 -67010
rect 59536 -67080 59616 -67070
rect 58396 -67110 58896 -67090
rect 59646 -67110 59706 -66840
rect 60436 -66920 60536 -66910
rect 59856 -66940 59976 -66930
rect 59856 -67030 59866 -66940
rect 59966 -67030 59976 -66940
rect 60436 -67020 60446 -66920
rect 60526 -67020 60536 -66920
rect 60436 -67030 60536 -67020
rect 59856 -67040 59976 -67030
rect 58396 -67120 59706 -67110
rect 58396 -67130 59216 -67120
rect 58396 -67190 58906 -67130
rect 58966 -67180 59216 -67130
rect 59276 -67180 59336 -67120
rect 59396 -67180 59436 -67120
rect 59496 -67130 59706 -67120
rect 59496 -67180 59636 -67130
rect 58966 -67190 59636 -67180
rect 59696 -67190 59706 -67130
rect 58396 -67200 59706 -67190
rect 60036 -67120 60136 -67110
rect 60036 -67200 60046 -67120
rect 60126 -67200 60136 -67120
rect 55510 -67218 55520 -67208
rect 59646 -67210 59706 -67200
rect 60546 -67210 60636 -67200
rect 59066 -67240 59176 -67230
rect 59066 -67310 59076 -67240
rect 59166 -67310 59176 -67240
rect 59846 -67280 59856 -67210
rect 59916 -67230 59926 -67210
rect 60356 -67220 60556 -67210
rect 60356 -67230 60376 -67220
rect 59916 -67260 60376 -67230
rect 59916 -67280 59926 -67260
rect 60356 -67280 60376 -67260
rect 60446 -67280 60556 -67220
rect 60356 -67290 60556 -67280
rect 60626 -67290 60636 -67210
rect 59066 -67320 59176 -67310
rect 59966 -67300 60326 -67290
rect 53850 -67438 53860 -67328
rect 53920 -67338 55600 -67328
rect 53920 -67438 55000 -67338
rect 55090 -67438 55540 -67338
rect 55630 -67438 55640 -67338
rect 59966 -67360 59976 -67300
rect 60316 -67360 60326 -67300
rect 60546 -67310 60636 -67290
rect 61186 -67320 61366 -67310
rect 54770 -67638 54850 -67438
rect 56470 -67448 56480 -67388
rect 56550 -67448 56560 -67388
rect 57088 -67504 57098 -67364
rect 57368 -67504 57378 -67364
rect 59166 -67430 59376 -67420
rect 59166 -67440 59286 -67430
rect 59166 -67520 59176 -67440
rect 59236 -67520 59286 -67440
rect 59366 -67520 59376 -67430
rect 59166 -67530 59376 -67520
rect 59526 -67470 59646 -67450
rect 59526 -67530 59576 -67470
rect 59636 -67530 59646 -67470
rect 61186 -67500 61206 -67320
rect 61346 -67500 61366 -67320
rect 61186 -67510 61366 -67500
rect 59526 -67560 59646 -67530
rect 60286 -67550 60476 -67540
rect 59906 -67580 60016 -67570
rect 59806 -67590 59866 -67580
rect 54760 -67728 54770 -67638
rect 54840 -67728 54850 -67638
rect 59166 -67640 59536 -67630
rect 59166 -67720 59176 -67640
rect 59236 -67720 59286 -67640
rect 54920 -67738 55210 -67728
rect 54920 -67808 55140 -67738
rect 55200 -67808 55210 -67738
rect 59166 -67730 59286 -67720
rect 59356 -67650 59536 -67640
rect 59356 -67720 59476 -67650
rect 59356 -67730 59536 -67720
rect 59166 -67740 59536 -67730
rect 59566 -67760 59576 -67590
rect 59636 -67600 59866 -67590
rect 59636 -67740 59806 -67600
rect 59636 -67760 59866 -67740
rect 59906 -67760 59916 -67580
rect 60006 -67760 60016 -67580
rect 60286 -67690 60306 -67550
rect 60456 -67690 60476 -67550
rect 60286 -67700 60476 -67690
rect 61026 -67620 61136 -67610
rect 61026 -67730 61036 -67620
rect 61126 -67730 61136 -67620
rect 61026 -67740 61136 -67730
rect 59566 -67770 59636 -67760
rect 59906 -67770 60016 -67760
rect 54760 -68128 54770 -68048
rect 54840 -68128 54850 -68048
rect 54770 -68338 54850 -68128
rect 54920 -68198 54980 -67808
rect 55880 -67838 56900 -67818
rect 55010 -67928 55020 -67848
rect 55120 -67928 55740 -67848
rect 55810 -67928 55820 -67848
rect 55870 -67928 55880 -67838
rect 55970 -67928 56480 -67838
rect 56550 -67928 56900 -67838
rect 55880 -67948 56900 -67928
rect 57020 -67820 57040 -67818
rect 57800 -67820 58240 -67810
rect 57020 -67940 57800 -67820
rect 57020 -67948 57040 -67940
rect 57800 -67950 58240 -67940
rect 58516 -67860 58796 -67790
rect 58516 -68060 58556 -67860
rect 58756 -68060 58796 -67860
rect 59066 -67810 59936 -67800
rect 59066 -67880 59076 -67810
rect 59166 -67830 59826 -67810
rect 59166 -67880 59316 -67830
rect 59066 -67890 59316 -67880
rect 59376 -67880 59826 -67830
rect 59916 -67880 59936 -67810
rect 59376 -67890 59936 -67880
rect 60076 -67880 60196 -67840
rect 59066 -67970 59936 -67960
rect 59066 -68040 59076 -67970
rect 59166 -68040 59206 -67970
rect 59266 -68040 59826 -67970
rect 59926 -68040 59936 -67970
rect 59066 -68050 59936 -68040
rect 60076 -68040 60096 -67880
rect 60176 -68040 60196 -67880
rect 58516 -68140 58796 -68060
rect 60076 -68080 60196 -68040
rect 61266 -67850 61366 -67840
rect 61266 -68060 61276 -67850
rect 61356 -68060 61366 -67850
rect 61266 -68070 61366 -68060
rect 59586 -68090 59656 -68080
rect 59796 -68090 59866 -68080
rect 59586 -68110 59796 -68090
rect 59156 -68120 59536 -68110
rect 59156 -68130 59266 -68120
rect 54910 -68268 54920 -68198
rect 54980 -68268 54990 -68198
rect 59156 -68210 59166 -68130
rect 59226 -68210 59266 -68130
rect 59366 -68130 59536 -68120
rect 59366 -68210 59466 -68130
rect 59526 -68210 59536 -68130
rect 59156 -68230 59536 -68210
rect 59646 -68250 59796 -68110
rect 59586 -68270 59796 -68250
rect 59856 -68270 59866 -68090
rect 53840 -68448 53850 -68338
rect 53920 -68438 55000 -68338
rect 55090 -68438 55540 -68338
rect 55630 -68438 55640 -68338
rect 56470 -68388 56480 -68328
rect 56550 -68388 56560 -68328
rect 57088 -68414 57098 -68274
rect 57368 -68414 57378 -68274
rect 59796 -68280 59866 -68270
rect 59906 -68090 60016 -68080
rect 59906 -68280 59916 -68090
rect 60006 -68280 60016 -68090
rect 60476 -68110 60546 -68100
rect 60536 -68170 60546 -68110
rect 60476 -68180 60546 -68170
rect 60966 -68230 61486 -68220
rect 60966 -68240 61336 -68230
rect 59906 -68290 60016 -68280
rect 60466 -68250 61336 -68240
rect 59506 -68310 59606 -68300
rect 59156 -68360 59376 -68340
rect 53920 -68448 55640 -68438
rect 59156 -68440 59166 -68360
rect 59226 -68440 59266 -68360
rect 59156 -68450 59266 -68440
rect 59366 -68450 59376 -68360
rect 59506 -68380 59516 -68310
rect 59596 -68380 59606 -68310
rect 60466 -68310 60476 -68250
rect 60536 -68310 60616 -68250
rect 60736 -68310 60756 -68250
rect 60816 -68310 60896 -68250
rect 60956 -68310 61336 -68250
rect 60466 -68320 61336 -68310
rect 60966 -68360 61336 -68320
rect 61456 -68360 61486 -68230
rect 60966 -68370 61486 -68360
rect 59506 -68390 59606 -68380
rect 59156 -68460 59376 -68450
rect 59306 -68520 60336 -68500
rect 59066 -68540 59176 -68530
rect 55210 -68718 55220 -68548
rect 55310 -68718 55320 -68548
rect 55400 -68728 55410 -68558
rect 55500 -68568 55510 -68558
rect 55500 -68688 56380 -68568
rect 56440 -68688 56450 -68568
rect 59066 -68600 59076 -68540
rect 59166 -68600 59176 -68540
rect 59306 -68580 59316 -68520
rect 59376 -68540 59966 -68520
rect 59376 -68580 59816 -68540
rect 59306 -68590 59816 -68580
rect 59846 -68580 59916 -68570
rect 59066 -68610 59176 -68600
rect 59846 -68640 59856 -68580
rect 59946 -68580 59966 -68540
rect 60326 -68580 60336 -68520
rect 59946 -68590 60336 -68580
rect 60366 -68540 61146 -68530
rect 60366 -68580 61056 -68540
rect 59646 -68650 59716 -68640
rect 59846 -68650 59916 -68640
rect 60366 -68640 60376 -68580
rect 60436 -68640 61056 -68580
rect 61126 -68640 61146 -68540
rect 55500 -68708 56450 -68688
rect 58396 -68660 59716 -68650
rect 55500 -68728 55510 -68708
rect 58396 -68730 58926 -68660
rect 58986 -68730 59146 -68660
rect 59226 -68730 59276 -68660
rect 59356 -68730 59396 -68660
rect 59476 -68720 59646 -68660
rect 59706 -68720 59716 -68660
rect 60366 -68670 61146 -68640
rect 59476 -68730 59716 -68720
rect 58396 -68740 59716 -68730
rect 54900 -68808 54910 -68798
rect 53940 -68888 53950 -68808
rect 54010 -68888 54910 -68808
rect 53940 -68898 54910 -68888
rect 54980 -68818 54990 -68798
rect 54980 -68878 55980 -68818
rect 54980 -68898 55880 -68878
rect 53940 -68918 55880 -68898
rect 53500 -69048 53510 -68928
rect 53630 -69048 53640 -68928
rect 55850 -68958 55880 -68918
rect 55970 -68958 55980 -68878
rect 55230 -69018 55240 -68958
rect 55370 -68978 55710 -68958
rect 55370 -68988 55720 -68978
rect 55370 -69008 55620 -68988
rect 55370 -69018 55380 -69008
rect 55400 -69068 55410 -69048
rect 54730 -69158 54740 -69068
rect 54850 -69138 55410 -69068
rect 55510 -69138 55520 -69048
rect 55600 -69078 55620 -69008
rect 55710 -69078 55720 -68988
rect 54850 -69158 55520 -69138
rect 55210 -69328 55220 -69218
rect 55330 -69328 55340 -69218
rect 55850 -69378 55980 -68958
rect 56010 -69208 56020 -69058
rect 56080 -69208 56090 -69058
rect 56160 -69208 56170 -69008
rect 56390 -69208 56400 -69008
rect 58396 -69020 58896 -68740
rect 59006 -68900 59076 -68880
rect 59246 -68890 59256 -68830
rect 59366 -68890 59376 -68830
rect 59536 -68860 59546 -68790
rect 59606 -68860 59616 -68790
rect 59536 -68870 59616 -68860
rect 59006 -68960 59016 -68900
rect 59536 -68910 59616 -68900
rect 59076 -68920 59086 -68910
rect 59536 -68920 59546 -68910
rect 59076 -68960 59546 -68920
rect 59006 -68970 59546 -68960
rect 59606 -68970 59616 -68910
rect 59006 -68990 59076 -68970
rect 59536 -68990 59616 -68970
rect 59646 -69020 59716 -68740
rect 59796 -68810 59926 -68800
rect 59796 -68920 59806 -68810
rect 59916 -68920 59926 -68810
rect 59796 -68930 59926 -68920
rect 60436 -68830 60536 -68810
rect 60436 -68950 60446 -68830
rect 60526 -68950 60536 -68830
rect 60436 -68960 60536 -68950
rect 58396 -69030 59716 -69020
rect 56654 -69068 56998 -69058
rect 55520 -69468 55530 -69378
rect 55610 -69468 55980 -69378
rect 54130 -69748 54140 -69488
rect 54850 -69748 54860 -69488
rect 55310 -69668 55320 -69528
rect 55470 -69668 55480 -69528
rect 56170 -69738 56390 -69208
rect 58396 -69100 58906 -69030
rect 58986 -69100 59146 -69030
rect 59226 -69100 59276 -69030
rect 59356 -69100 59396 -69030
rect 59476 -69040 59716 -69030
rect 59476 -69100 59646 -69040
rect 59706 -69100 59716 -69040
rect 58396 -69110 59716 -69100
rect 58396 -69150 58896 -69110
rect 59646 -69120 59716 -69110
rect 56654 -69296 56998 -69286
rect 59006 -69200 60416 -69190
rect 59006 -69240 60266 -69200
rect 59006 -69310 59016 -69240
rect 59076 -69310 59546 -69240
rect 59606 -69310 60266 -69240
rect 59006 -69330 60266 -69310
rect 60406 -69330 60416 -69200
rect 59006 -69340 60416 -69330
rect 59986 -69390 60116 -69380
rect 58956 -69400 59156 -69390
rect 58956 -69580 58966 -69400
rect 59146 -69580 59156 -69400
rect 59986 -69500 59996 -69390
rect 60106 -69500 60116 -69390
rect 58956 -69590 59156 -69580
rect 55680 -69748 56390 -69738
rect 54130 -69908 56390 -69748
rect 55680 -69918 56390 -69908
rect 59600 -69600 60500 -69500
rect 59600 -70000 59700 -69600
rect 60400 -70000 60500 -69600
rect 55400 -70100 56200 -70000
rect 59600 -70100 60500 -70000
rect 67000 -69600 67500 -49100
rect 67000 -70000 67100 -69600
rect 67400 -70000 67500 -69600
rect 67000 -70100 67500 -70000
rect 67900 -49300 68400 -49200
rect 67900 -49500 68000 -49300
rect 68300 -49500 68400 -49300
rect 72810 -49220 73050 -49210
rect 72810 -49400 72820 -49220
rect 73040 -49400 73050 -49220
rect 72810 -49410 73050 -49400
rect 55400 -70500 55500 -70100
rect 56100 -70500 56200 -70100
rect 55400 -70600 56200 -70500
rect 51400 -71300 51500 -71100
rect 52500 -71300 52600 -71100
rect 51400 -76500 52600 -71300
rect 55440 -71080 55740 -71060
rect 55440 -71360 55460 -71080
rect 55720 -71360 55740 -71080
rect 55440 -71380 55740 -71360
rect 54140 -71538 56390 -71528
rect 53460 -71740 53800 -71720
rect 53460 -71940 53480 -71740
rect 53780 -71940 53800 -71740
rect 54140 -71778 54150 -71538
rect 54860 -71778 56390 -71538
rect 58946 -71670 59146 -71650
rect 54140 -71788 56390 -71778
rect 53460 -71960 53800 -71940
rect 54850 -72018 55530 -72008
rect 53510 -72168 53520 -72058
rect 53640 -72168 53650 -72058
rect 54740 -72118 54750 -72038
rect 54850 -72088 55430 -72018
rect 55520 -72088 55530 -72018
rect 55950 -72088 55960 -71938
rect 56040 -72088 56050 -71938
rect 56170 -71958 56390 -71788
rect 56506 -71780 57016 -71770
rect 54840 -72118 54850 -72108
rect 55270 -72208 55280 -72118
rect 55400 -72208 55410 -72118
rect 56170 -72168 56190 -71958
rect 56390 -72168 56400 -71958
rect 58946 -71830 58966 -71670
rect 59126 -71830 59146 -71670
rect 58946 -71850 59146 -71830
rect 59316 -71700 60176 -71690
rect 59316 -71710 59956 -71700
rect 59316 -71850 59336 -71710
rect 59416 -71850 59956 -71710
rect 59316 -71860 59956 -71850
rect 60166 -71860 60176 -71700
rect 59316 -71870 60176 -71860
rect 56506 -72040 57016 -72030
rect 58956 -71920 61136 -71910
rect 58956 -71930 61056 -71920
rect 58956 -72040 58996 -71930
rect 59106 -71940 61056 -71930
rect 59106 -72040 59516 -71940
rect 59616 -72040 61056 -71940
rect 58396 -72130 58896 -72040
rect 58956 -72050 61056 -72040
rect 61126 -72050 61136 -71920
rect 58956 -72060 61136 -72050
rect 55850 -72248 55880 -72218
rect 53940 -72278 55880 -72248
rect 53940 -72298 54920 -72278
rect 53040 -74108 53050 -72358
rect 53250 -74108 53260 -72358
rect 53940 -72398 53950 -72298
rect 54020 -72348 54920 -72298
rect 54020 -72398 54030 -72348
rect 54910 -72368 54920 -72348
rect 54990 -72298 55880 -72278
rect 55970 -72248 55980 -72218
rect 54990 -72348 55970 -72298
rect 54990 -72368 55000 -72348
rect 55220 -72628 55230 -72458
rect 55320 -72628 55330 -72458
rect 55420 -72618 55430 -72448
rect 55510 -72458 55520 -72448
rect 55510 -72468 56670 -72458
rect 55510 -72598 55600 -72468
rect 55710 -72598 56590 -72468
rect 56660 -72598 56670 -72468
rect 55510 -72608 56670 -72598
rect 58396 -72490 58486 -72130
rect 58816 -72150 58896 -72130
rect 59646 -72150 59706 -72130
rect 58816 -72170 59706 -72150
rect 58816 -72230 58906 -72170
rect 58966 -72230 59216 -72170
rect 59276 -72230 59326 -72170
rect 59386 -72230 59436 -72170
rect 59496 -72230 59636 -72170
rect 59696 -72230 59706 -72170
rect 58816 -72240 59706 -72230
rect 58816 -72490 58896 -72240
rect 59536 -72290 59616 -72280
rect 59276 -72330 59356 -72320
rect 59276 -72390 59286 -72330
rect 59346 -72390 59356 -72330
rect 59536 -72350 59546 -72290
rect 59606 -72350 59616 -72290
rect 59536 -72370 59616 -72350
rect 58996 -72400 59076 -72390
rect 58996 -72460 59006 -72400
rect 59076 -72420 59086 -72400
rect 59536 -72410 59616 -72400
rect 59536 -72420 59546 -72410
rect 59076 -72460 59546 -72420
rect 58996 -72470 59076 -72460
rect 59536 -72470 59546 -72460
rect 59606 -72470 59616 -72410
rect 59536 -72480 59616 -72470
rect 58396 -72510 58896 -72490
rect 59646 -72510 59706 -72240
rect 60436 -72320 60536 -72310
rect 59856 -72340 59976 -72330
rect 59856 -72430 59866 -72340
rect 59966 -72430 59976 -72340
rect 60436 -72420 60446 -72320
rect 60526 -72420 60536 -72320
rect 60436 -72430 60536 -72420
rect 59856 -72440 59976 -72430
rect 58396 -72520 59706 -72510
rect 58396 -72530 59216 -72520
rect 58396 -72590 58906 -72530
rect 58966 -72580 59216 -72530
rect 59276 -72580 59336 -72520
rect 59396 -72580 59436 -72520
rect 59496 -72530 59706 -72520
rect 59496 -72580 59636 -72530
rect 58966 -72590 59636 -72580
rect 59696 -72590 59706 -72530
rect 58396 -72600 59706 -72590
rect 60036 -72520 60136 -72510
rect 60036 -72600 60046 -72520
rect 60126 -72600 60136 -72520
rect 55510 -72618 55520 -72608
rect 59646 -72610 59706 -72600
rect 60546 -72610 60636 -72600
rect 59066 -72640 59176 -72630
rect 59066 -72710 59076 -72640
rect 59166 -72710 59176 -72640
rect 59846 -72680 59856 -72610
rect 59916 -72630 59926 -72610
rect 60356 -72620 60556 -72610
rect 60356 -72630 60376 -72620
rect 59916 -72660 60376 -72630
rect 59916 -72680 59926 -72660
rect 60356 -72680 60376 -72660
rect 60446 -72680 60556 -72620
rect 60356 -72690 60556 -72680
rect 60626 -72690 60636 -72610
rect 59066 -72720 59176 -72710
rect 59966 -72700 60326 -72690
rect 53850 -72838 53860 -72728
rect 53920 -72738 55600 -72728
rect 53920 -72838 55000 -72738
rect 55090 -72838 55540 -72738
rect 55630 -72838 55640 -72738
rect 59966 -72760 59976 -72700
rect 60316 -72760 60326 -72700
rect 60546 -72710 60636 -72690
rect 61186 -72720 61366 -72710
rect 54770 -73038 54850 -72838
rect 56470 -72848 56480 -72788
rect 56550 -72848 56560 -72788
rect 57088 -72904 57098 -72764
rect 57368 -72904 57378 -72764
rect 59166 -72830 59376 -72820
rect 59166 -72840 59286 -72830
rect 59166 -72920 59176 -72840
rect 59236 -72920 59286 -72840
rect 59366 -72920 59376 -72830
rect 59166 -72930 59376 -72920
rect 59526 -72870 59646 -72850
rect 59526 -72930 59576 -72870
rect 59636 -72930 59646 -72870
rect 61186 -72900 61206 -72720
rect 61346 -72900 61366 -72720
rect 61186 -72910 61366 -72900
rect 59526 -72960 59646 -72930
rect 60286 -72950 60476 -72940
rect 59906 -72980 60016 -72970
rect 59806 -72990 59866 -72980
rect 54760 -73128 54770 -73038
rect 54840 -73128 54850 -73038
rect 59166 -73040 59536 -73030
rect 59166 -73120 59176 -73040
rect 59236 -73120 59286 -73040
rect 54920 -73138 55210 -73128
rect 54920 -73208 55140 -73138
rect 55200 -73208 55210 -73138
rect 59166 -73130 59286 -73120
rect 59356 -73050 59536 -73040
rect 59356 -73120 59476 -73050
rect 59356 -73130 59536 -73120
rect 59166 -73140 59536 -73130
rect 59566 -73160 59576 -72990
rect 59636 -73000 59866 -72990
rect 59636 -73140 59806 -73000
rect 59636 -73160 59866 -73140
rect 59906 -73160 59916 -72980
rect 60006 -73160 60016 -72980
rect 60286 -73090 60306 -72950
rect 60456 -73090 60476 -72950
rect 60286 -73100 60476 -73090
rect 61026 -73020 61136 -73010
rect 61026 -73130 61036 -73020
rect 61126 -73130 61136 -73020
rect 61026 -73140 61136 -73130
rect 59566 -73170 59636 -73160
rect 59906 -73170 60016 -73160
rect 54760 -73528 54770 -73448
rect 54840 -73528 54850 -73448
rect 54770 -73738 54850 -73528
rect 54920 -73598 54980 -73208
rect 55880 -73238 56900 -73218
rect 55010 -73328 55020 -73248
rect 55120 -73328 55740 -73248
rect 55810 -73328 55820 -73248
rect 55870 -73328 55880 -73238
rect 55970 -73328 56480 -73238
rect 56550 -73328 56900 -73238
rect 55880 -73348 56900 -73328
rect 57020 -73220 57040 -73218
rect 57800 -73220 58240 -73210
rect 57020 -73340 57800 -73220
rect 57020 -73348 57040 -73340
rect 57800 -73350 58240 -73340
rect 58516 -73260 58796 -73190
rect 58516 -73460 58556 -73260
rect 58756 -73460 58796 -73260
rect 59066 -73210 59936 -73200
rect 59066 -73280 59076 -73210
rect 59166 -73230 59826 -73210
rect 59166 -73280 59316 -73230
rect 59066 -73290 59316 -73280
rect 59376 -73280 59826 -73230
rect 59916 -73280 59936 -73210
rect 59376 -73290 59936 -73280
rect 60076 -73280 60196 -73240
rect 59066 -73370 59936 -73360
rect 59066 -73440 59076 -73370
rect 59166 -73440 59206 -73370
rect 59266 -73440 59826 -73370
rect 59926 -73440 59936 -73370
rect 59066 -73450 59936 -73440
rect 60076 -73440 60096 -73280
rect 60176 -73440 60196 -73280
rect 58516 -73540 58796 -73460
rect 60076 -73480 60196 -73440
rect 61266 -73250 61366 -73240
rect 61266 -73460 61276 -73250
rect 61356 -73460 61366 -73250
rect 61266 -73470 61366 -73460
rect 59586 -73490 59656 -73480
rect 59796 -73490 59866 -73480
rect 59586 -73510 59796 -73490
rect 59156 -73520 59536 -73510
rect 59156 -73530 59266 -73520
rect 54910 -73668 54920 -73598
rect 54980 -73668 54990 -73598
rect 59156 -73610 59166 -73530
rect 59226 -73610 59266 -73530
rect 59366 -73530 59536 -73520
rect 59366 -73610 59466 -73530
rect 59526 -73610 59536 -73530
rect 59156 -73630 59536 -73610
rect 59646 -73650 59796 -73510
rect 59586 -73670 59796 -73650
rect 59856 -73670 59866 -73490
rect 53840 -73848 53850 -73738
rect 53920 -73838 55000 -73738
rect 55090 -73838 55540 -73738
rect 55630 -73838 55640 -73738
rect 56470 -73788 56480 -73728
rect 56550 -73788 56560 -73728
rect 57088 -73814 57098 -73674
rect 57368 -73814 57378 -73674
rect 59796 -73680 59866 -73670
rect 59906 -73490 60016 -73480
rect 59906 -73680 59916 -73490
rect 60006 -73680 60016 -73490
rect 60476 -73510 60546 -73500
rect 60536 -73570 60546 -73510
rect 60476 -73580 60546 -73570
rect 60966 -73630 61486 -73620
rect 60966 -73640 61336 -73630
rect 59906 -73690 60016 -73680
rect 60466 -73650 61336 -73640
rect 59506 -73710 59606 -73700
rect 59156 -73760 59376 -73740
rect 53920 -73848 55640 -73838
rect 59156 -73840 59166 -73760
rect 59226 -73840 59266 -73760
rect 59156 -73850 59266 -73840
rect 59366 -73850 59376 -73760
rect 59506 -73780 59516 -73710
rect 59596 -73780 59606 -73710
rect 60466 -73710 60476 -73650
rect 60536 -73710 60616 -73650
rect 60736 -73710 60756 -73650
rect 60816 -73710 60896 -73650
rect 60956 -73710 61336 -73650
rect 60466 -73720 61336 -73710
rect 60966 -73760 61336 -73720
rect 61456 -73760 61486 -73630
rect 60966 -73770 61486 -73760
rect 59506 -73790 59606 -73780
rect 59156 -73860 59376 -73850
rect 59306 -73920 60336 -73900
rect 59066 -73940 59176 -73930
rect 55210 -74118 55220 -73948
rect 55310 -74118 55320 -73948
rect 55400 -74128 55410 -73958
rect 55500 -73968 55510 -73958
rect 55500 -74088 56380 -73968
rect 56440 -74088 56450 -73968
rect 59066 -74000 59076 -73940
rect 59166 -74000 59176 -73940
rect 59306 -73980 59316 -73920
rect 59376 -73940 59966 -73920
rect 59376 -73980 59816 -73940
rect 59306 -73990 59816 -73980
rect 59846 -73980 59916 -73970
rect 59066 -74010 59176 -74000
rect 59846 -74040 59856 -73980
rect 59946 -73980 59966 -73940
rect 60326 -73980 60336 -73920
rect 59946 -73990 60336 -73980
rect 60366 -73940 61146 -73930
rect 60366 -73980 61056 -73940
rect 59646 -74050 59716 -74040
rect 59846 -74050 59916 -74040
rect 60366 -74040 60376 -73980
rect 60436 -74040 61056 -73980
rect 61126 -74040 61146 -73940
rect 55500 -74108 56450 -74088
rect 58396 -74060 59716 -74050
rect 55500 -74128 55510 -74108
rect 58396 -74130 58926 -74060
rect 58986 -74130 59146 -74060
rect 59226 -74130 59276 -74060
rect 59356 -74130 59396 -74060
rect 59476 -74120 59646 -74060
rect 59706 -74120 59716 -74060
rect 60366 -74070 61146 -74040
rect 59476 -74130 59716 -74120
rect 58396 -74140 59716 -74130
rect 54900 -74208 54910 -74198
rect 53940 -74288 53950 -74208
rect 54010 -74288 54910 -74208
rect 53940 -74298 54910 -74288
rect 54980 -74218 54990 -74198
rect 54980 -74278 55980 -74218
rect 54980 -74298 55880 -74278
rect 53940 -74318 55880 -74298
rect 53500 -74448 53510 -74328
rect 53630 -74448 53640 -74328
rect 55850 -74358 55880 -74318
rect 55970 -74358 55980 -74278
rect 55230 -74418 55240 -74358
rect 55370 -74378 55710 -74358
rect 55370 -74388 55720 -74378
rect 55370 -74408 55620 -74388
rect 55370 -74418 55380 -74408
rect 55400 -74468 55410 -74448
rect 54730 -74558 54740 -74468
rect 54850 -74538 55410 -74468
rect 55510 -74538 55520 -74448
rect 55600 -74478 55620 -74408
rect 55710 -74478 55720 -74388
rect 54850 -74558 55520 -74538
rect 55210 -74728 55220 -74618
rect 55330 -74728 55340 -74618
rect 55850 -74778 55980 -74358
rect 56010 -74608 56020 -74458
rect 56080 -74608 56090 -74458
rect 56160 -74608 56170 -74408
rect 56390 -74608 56400 -74408
rect 58396 -74420 58896 -74140
rect 59006 -74300 59076 -74280
rect 59246 -74290 59256 -74230
rect 59366 -74290 59376 -74230
rect 59536 -74260 59546 -74190
rect 59606 -74260 59616 -74190
rect 59536 -74270 59616 -74260
rect 59006 -74360 59016 -74300
rect 59536 -74310 59616 -74300
rect 59076 -74320 59086 -74310
rect 59536 -74320 59546 -74310
rect 59076 -74360 59546 -74320
rect 59006 -74370 59546 -74360
rect 59606 -74370 59616 -74310
rect 59006 -74390 59076 -74370
rect 59536 -74390 59616 -74370
rect 59646 -74420 59716 -74140
rect 59796 -74210 59926 -74200
rect 59796 -74320 59806 -74210
rect 59916 -74320 59926 -74210
rect 59796 -74330 59926 -74320
rect 60436 -74230 60536 -74210
rect 60436 -74350 60446 -74230
rect 60526 -74350 60536 -74230
rect 60436 -74360 60536 -74350
rect 58396 -74430 59716 -74420
rect 56654 -74468 56998 -74458
rect 55520 -74868 55530 -74778
rect 55610 -74868 55980 -74778
rect 54130 -75148 54140 -74888
rect 54850 -75148 54860 -74888
rect 55310 -75068 55320 -74928
rect 55470 -75068 55480 -74928
rect 56170 -75138 56390 -74608
rect 58396 -74500 58906 -74430
rect 58986 -74500 59146 -74430
rect 59226 -74500 59276 -74430
rect 59356 -74500 59396 -74430
rect 59476 -74440 59716 -74430
rect 59476 -74500 59646 -74440
rect 59706 -74500 59716 -74440
rect 58396 -74510 59716 -74500
rect 58396 -74550 58896 -74510
rect 59646 -74520 59716 -74510
rect 56654 -74696 56998 -74686
rect 59006 -74600 60416 -74590
rect 59006 -74640 60266 -74600
rect 59006 -74710 59016 -74640
rect 59076 -74710 59546 -74640
rect 59606 -74710 60266 -74640
rect 59006 -74730 60266 -74710
rect 60406 -74730 60416 -74600
rect 59006 -74740 60416 -74730
rect 59986 -74790 60116 -74780
rect 58956 -74800 59156 -74790
rect 58956 -74980 58966 -74800
rect 59146 -74980 59156 -74800
rect 59986 -74900 59996 -74790
rect 60106 -74900 60116 -74790
rect 58956 -74990 59156 -74980
rect 55680 -75148 56390 -75138
rect 54130 -75308 56390 -75148
rect 55680 -75318 56390 -75308
rect 59600 -75000 60500 -74900
rect 59600 -75400 59700 -75000
rect 60400 -75400 60500 -75000
rect 55400 -75500 56200 -75400
rect 59600 -75500 60500 -75400
rect 67900 -75000 68400 -49500
rect 67900 -75400 68000 -75000
rect 68300 -75400 68400 -75000
rect 67900 -75500 68400 -75400
rect 68900 -49700 69400 -49600
rect 68900 -49900 69000 -49700
rect 69300 -49900 69400 -49700
rect 72810 -49670 73050 -49660
rect 72810 -49850 72820 -49670
rect 73040 -49850 73050 -49670
rect 72810 -49860 73050 -49850
rect 55400 -75900 55500 -75500
rect 56100 -75900 56200 -75500
rect 55400 -76000 56200 -75900
rect 51400 -76700 51500 -76500
rect 52500 -76700 52600 -76500
rect 51400 -81900 52600 -76700
rect 55380 -76480 55740 -76460
rect 55380 -76760 55400 -76480
rect 55720 -76760 55740 -76480
rect 55380 -76780 55740 -76760
rect 54140 -76938 56390 -76928
rect 53460 -77140 53800 -77120
rect 53460 -77340 53480 -77140
rect 53780 -77340 53800 -77140
rect 54140 -77178 54150 -76938
rect 54860 -77178 56390 -76938
rect 58946 -77070 59146 -77050
rect 54140 -77188 56390 -77178
rect 53460 -77360 53800 -77340
rect 54850 -77418 55530 -77408
rect 53510 -77568 53520 -77458
rect 53640 -77568 53650 -77458
rect 54740 -77518 54750 -77438
rect 54850 -77488 55430 -77418
rect 55520 -77488 55530 -77418
rect 55950 -77488 55960 -77338
rect 56040 -77488 56050 -77338
rect 56170 -77358 56390 -77188
rect 56506 -77180 57016 -77170
rect 54840 -77518 54850 -77508
rect 55270 -77608 55280 -77518
rect 55400 -77608 55410 -77518
rect 56170 -77568 56190 -77358
rect 56390 -77568 56400 -77358
rect 58946 -77230 58966 -77070
rect 59126 -77230 59146 -77070
rect 58946 -77250 59146 -77230
rect 59316 -77100 60176 -77090
rect 59316 -77110 59956 -77100
rect 59316 -77250 59336 -77110
rect 59416 -77250 59956 -77110
rect 59316 -77260 59956 -77250
rect 60166 -77260 60176 -77100
rect 59316 -77270 60176 -77260
rect 56506 -77440 57016 -77430
rect 58956 -77320 61136 -77310
rect 58956 -77330 61056 -77320
rect 58956 -77440 58996 -77330
rect 59106 -77340 61056 -77330
rect 59106 -77440 59516 -77340
rect 59616 -77440 61056 -77340
rect 58396 -77530 58896 -77440
rect 58956 -77450 61056 -77440
rect 61126 -77450 61136 -77320
rect 58956 -77460 61136 -77450
rect 55850 -77648 55880 -77618
rect 53940 -77678 55880 -77648
rect 53940 -77698 54920 -77678
rect 53040 -79508 53050 -77758
rect 53250 -79508 53260 -77758
rect 53940 -77798 53950 -77698
rect 54020 -77748 54920 -77698
rect 54020 -77798 54030 -77748
rect 54910 -77768 54920 -77748
rect 54990 -77698 55880 -77678
rect 55970 -77648 55980 -77618
rect 54990 -77748 55970 -77698
rect 54990 -77768 55000 -77748
rect 55220 -78028 55230 -77858
rect 55320 -78028 55330 -77858
rect 55420 -78018 55430 -77848
rect 55510 -77858 55520 -77848
rect 55510 -77868 56670 -77858
rect 55510 -77998 55600 -77868
rect 55710 -77998 56590 -77868
rect 56660 -77998 56670 -77868
rect 55510 -78008 56670 -77998
rect 58396 -77890 58486 -77530
rect 58816 -77550 58896 -77530
rect 59646 -77550 59706 -77530
rect 58816 -77570 59706 -77550
rect 58816 -77630 58906 -77570
rect 58966 -77630 59216 -77570
rect 59276 -77630 59326 -77570
rect 59386 -77630 59436 -77570
rect 59496 -77630 59636 -77570
rect 59696 -77630 59706 -77570
rect 58816 -77640 59706 -77630
rect 58816 -77890 58896 -77640
rect 59536 -77690 59616 -77680
rect 59276 -77730 59356 -77720
rect 59276 -77790 59286 -77730
rect 59346 -77790 59356 -77730
rect 59536 -77750 59546 -77690
rect 59606 -77750 59616 -77690
rect 59536 -77770 59616 -77750
rect 58996 -77800 59076 -77790
rect 58996 -77860 59006 -77800
rect 59076 -77820 59086 -77800
rect 59536 -77810 59616 -77800
rect 59536 -77820 59546 -77810
rect 59076 -77860 59546 -77820
rect 58996 -77870 59076 -77860
rect 59536 -77870 59546 -77860
rect 59606 -77870 59616 -77810
rect 59536 -77880 59616 -77870
rect 58396 -77910 58896 -77890
rect 59646 -77910 59706 -77640
rect 60436 -77720 60536 -77710
rect 59856 -77740 59976 -77730
rect 59856 -77830 59866 -77740
rect 59966 -77830 59976 -77740
rect 60436 -77820 60446 -77720
rect 60526 -77820 60536 -77720
rect 60436 -77830 60536 -77820
rect 59856 -77840 59976 -77830
rect 58396 -77920 59706 -77910
rect 58396 -77930 59216 -77920
rect 58396 -77990 58906 -77930
rect 58966 -77980 59216 -77930
rect 59276 -77980 59336 -77920
rect 59396 -77980 59436 -77920
rect 59496 -77930 59706 -77920
rect 59496 -77980 59636 -77930
rect 58966 -77990 59636 -77980
rect 59696 -77990 59706 -77930
rect 58396 -78000 59706 -77990
rect 60036 -77920 60136 -77910
rect 60036 -78000 60046 -77920
rect 60126 -78000 60136 -77920
rect 55510 -78018 55520 -78008
rect 59646 -78010 59706 -78000
rect 60546 -78010 60636 -78000
rect 59066 -78040 59176 -78030
rect 59066 -78110 59076 -78040
rect 59166 -78110 59176 -78040
rect 59846 -78080 59856 -78010
rect 59916 -78030 59926 -78010
rect 60356 -78020 60556 -78010
rect 60356 -78030 60376 -78020
rect 59916 -78060 60376 -78030
rect 59916 -78080 59926 -78060
rect 60356 -78080 60376 -78060
rect 60446 -78080 60556 -78020
rect 60356 -78090 60556 -78080
rect 60626 -78090 60636 -78010
rect 59066 -78120 59176 -78110
rect 59966 -78100 60326 -78090
rect 53850 -78238 53860 -78128
rect 53920 -78138 55600 -78128
rect 53920 -78238 55000 -78138
rect 55090 -78238 55540 -78138
rect 55630 -78238 55640 -78138
rect 59966 -78160 59976 -78100
rect 60316 -78160 60326 -78100
rect 60546 -78110 60636 -78090
rect 61186 -78120 61366 -78110
rect 54770 -78438 54850 -78238
rect 56470 -78248 56480 -78188
rect 56550 -78248 56560 -78188
rect 57088 -78304 57098 -78164
rect 57368 -78304 57378 -78164
rect 59166 -78230 59376 -78220
rect 59166 -78240 59286 -78230
rect 59166 -78320 59176 -78240
rect 59236 -78320 59286 -78240
rect 59366 -78320 59376 -78230
rect 59166 -78330 59376 -78320
rect 59526 -78270 59646 -78250
rect 59526 -78330 59576 -78270
rect 59636 -78330 59646 -78270
rect 61186 -78300 61206 -78120
rect 61346 -78300 61366 -78120
rect 61186 -78310 61366 -78300
rect 59526 -78360 59646 -78330
rect 60286 -78350 60476 -78340
rect 59906 -78380 60016 -78370
rect 59806 -78390 59866 -78380
rect 54760 -78528 54770 -78438
rect 54840 -78528 54850 -78438
rect 59166 -78440 59536 -78430
rect 59166 -78520 59176 -78440
rect 59236 -78520 59286 -78440
rect 54920 -78538 55210 -78528
rect 54920 -78608 55140 -78538
rect 55200 -78608 55210 -78538
rect 59166 -78530 59286 -78520
rect 59356 -78450 59536 -78440
rect 59356 -78520 59476 -78450
rect 59356 -78530 59536 -78520
rect 59166 -78540 59536 -78530
rect 59566 -78560 59576 -78390
rect 59636 -78400 59866 -78390
rect 59636 -78540 59806 -78400
rect 59636 -78560 59866 -78540
rect 59906 -78560 59916 -78380
rect 60006 -78560 60016 -78380
rect 60286 -78490 60306 -78350
rect 60456 -78490 60476 -78350
rect 60286 -78500 60476 -78490
rect 61026 -78420 61136 -78410
rect 61026 -78530 61036 -78420
rect 61126 -78530 61136 -78420
rect 61026 -78540 61136 -78530
rect 59566 -78570 59636 -78560
rect 59906 -78570 60016 -78560
rect 54760 -78928 54770 -78848
rect 54840 -78928 54850 -78848
rect 54770 -79138 54850 -78928
rect 54920 -78998 54980 -78608
rect 55880 -78638 56900 -78618
rect 55010 -78728 55020 -78648
rect 55120 -78728 55740 -78648
rect 55810 -78728 55820 -78648
rect 55870 -78728 55880 -78638
rect 55970 -78728 56480 -78638
rect 56550 -78728 56900 -78638
rect 55880 -78748 56900 -78728
rect 57020 -78620 57040 -78618
rect 57800 -78620 58240 -78610
rect 57020 -78740 57800 -78620
rect 57020 -78748 57040 -78740
rect 57800 -78750 58240 -78740
rect 58516 -78660 58796 -78590
rect 58516 -78860 58556 -78660
rect 58756 -78860 58796 -78660
rect 59066 -78610 59936 -78600
rect 59066 -78680 59076 -78610
rect 59166 -78630 59826 -78610
rect 59166 -78680 59316 -78630
rect 59066 -78690 59316 -78680
rect 59376 -78680 59826 -78630
rect 59916 -78680 59936 -78610
rect 59376 -78690 59936 -78680
rect 60076 -78680 60196 -78640
rect 59066 -78770 59936 -78760
rect 59066 -78840 59076 -78770
rect 59166 -78840 59206 -78770
rect 59266 -78840 59826 -78770
rect 59926 -78840 59936 -78770
rect 59066 -78850 59936 -78840
rect 60076 -78840 60096 -78680
rect 60176 -78840 60196 -78680
rect 58516 -78940 58796 -78860
rect 60076 -78880 60196 -78840
rect 61266 -78650 61366 -78640
rect 61266 -78860 61276 -78650
rect 61356 -78860 61366 -78650
rect 61266 -78870 61366 -78860
rect 59586 -78890 59656 -78880
rect 59796 -78890 59866 -78880
rect 59586 -78910 59796 -78890
rect 59156 -78920 59536 -78910
rect 59156 -78930 59266 -78920
rect 54910 -79068 54920 -78998
rect 54980 -79068 54990 -78998
rect 59156 -79010 59166 -78930
rect 59226 -79010 59266 -78930
rect 59366 -78930 59536 -78920
rect 59366 -79010 59466 -78930
rect 59526 -79010 59536 -78930
rect 59156 -79030 59536 -79010
rect 59646 -79050 59796 -78910
rect 59586 -79070 59796 -79050
rect 59856 -79070 59866 -78890
rect 53840 -79248 53850 -79138
rect 53920 -79238 55000 -79138
rect 55090 -79238 55540 -79138
rect 55630 -79238 55640 -79138
rect 56470 -79188 56480 -79128
rect 56550 -79188 56560 -79128
rect 57088 -79214 57098 -79074
rect 57368 -79214 57378 -79074
rect 59796 -79080 59866 -79070
rect 59906 -78890 60016 -78880
rect 59906 -79080 59916 -78890
rect 60006 -79080 60016 -78890
rect 60476 -78910 60546 -78900
rect 60536 -78970 60546 -78910
rect 60476 -78980 60546 -78970
rect 60966 -79030 61486 -79020
rect 60966 -79040 61336 -79030
rect 59906 -79090 60016 -79080
rect 60466 -79050 61336 -79040
rect 59506 -79110 59606 -79100
rect 59156 -79160 59376 -79140
rect 53920 -79248 55640 -79238
rect 59156 -79240 59166 -79160
rect 59226 -79240 59266 -79160
rect 59156 -79250 59266 -79240
rect 59366 -79250 59376 -79160
rect 59506 -79180 59516 -79110
rect 59596 -79180 59606 -79110
rect 60466 -79110 60476 -79050
rect 60536 -79110 60616 -79050
rect 60736 -79110 60756 -79050
rect 60816 -79110 60896 -79050
rect 60956 -79110 61336 -79050
rect 60466 -79120 61336 -79110
rect 60966 -79160 61336 -79120
rect 61456 -79160 61486 -79030
rect 60966 -79170 61486 -79160
rect 59506 -79190 59606 -79180
rect 59156 -79260 59376 -79250
rect 59306 -79320 60336 -79300
rect 59066 -79340 59176 -79330
rect 55210 -79518 55220 -79348
rect 55310 -79518 55320 -79348
rect 55400 -79528 55410 -79358
rect 55500 -79368 55510 -79358
rect 55500 -79488 56380 -79368
rect 56440 -79488 56450 -79368
rect 59066 -79400 59076 -79340
rect 59166 -79400 59176 -79340
rect 59306 -79380 59316 -79320
rect 59376 -79340 59966 -79320
rect 59376 -79380 59816 -79340
rect 59306 -79390 59816 -79380
rect 59846 -79380 59916 -79370
rect 59066 -79410 59176 -79400
rect 59846 -79440 59856 -79380
rect 59946 -79380 59966 -79340
rect 60326 -79380 60336 -79320
rect 59946 -79390 60336 -79380
rect 60366 -79340 61146 -79330
rect 60366 -79380 61056 -79340
rect 59646 -79450 59716 -79440
rect 59846 -79450 59916 -79440
rect 60366 -79440 60376 -79380
rect 60436 -79440 61056 -79380
rect 61126 -79440 61146 -79340
rect 55500 -79508 56450 -79488
rect 58396 -79460 59716 -79450
rect 55500 -79528 55510 -79508
rect 58396 -79530 58926 -79460
rect 58986 -79530 59146 -79460
rect 59226 -79530 59276 -79460
rect 59356 -79530 59396 -79460
rect 59476 -79520 59646 -79460
rect 59706 -79520 59716 -79460
rect 60366 -79470 61146 -79440
rect 59476 -79530 59716 -79520
rect 58396 -79540 59716 -79530
rect 54900 -79608 54910 -79598
rect 53940 -79688 53950 -79608
rect 54010 -79688 54910 -79608
rect 53940 -79698 54910 -79688
rect 54980 -79618 54990 -79598
rect 54980 -79678 55980 -79618
rect 54980 -79698 55880 -79678
rect 53940 -79718 55880 -79698
rect 53500 -79848 53510 -79728
rect 53630 -79848 53640 -79728
rect 55850 -79758 55880 -79718
rect 55970 -79758 55980 -79678
rect 55230 -79818 55240 -79758
rect 55370 -79778 55710 -79758
rect 55370 -79788 55720 -79778
rect 55370 -79808 55620 -79788
rect 55370 -79818 55380 -79808
rect 55400 -79868 55410 -79848
rect 54730 -79958 54740 -79868
rect 54850 -79938 55410 -79868
rect 55510 -79938 55520 -79848
rect 55600 -79878 55620 -79808
rect 55710 -79878 55720 -79788
rect 54850 -79958 55520 -79938
rect 55210 -80128 55220 -80018
rect 55330 -80128 55340 -80018
rect 55850 -80178 55980 -79758
rect 56010 -80008 56020 -79858
rect 56080 -80008 56090 -79858
rect 56160 -80008 56170 -79808
rect 56390 -80008 56400 -79808
rect 58396 -79820 58896 -79540
rect 59006 -79700 59076 -79680
rect 59246 -79690 59256 -79630
rect 59366 -79690 59376 -79630
rect 59536 -79660 59546 -79590
rect 59606 -79660 59616 -79590
rect 59536 -79670 59616 -79660
rect 59006 -79760 59016 -79700
rect 59536 -79710 59616 -79700
rect 59076 -79720 59086 -79710
rect 59536 -79720 59546 -79710
rect 59076 -79760 59546 -79720
rect 59006 -79770 59546 -79760
rect 59606 -79770 59616 -79710
rect 59006 -79790 59076 -79770
rect 59536 -79790 59616 -79770
rect 59646 -79820 59716 -79540
rect 59796 -79610 59926 -79600
rect 59796 -79720 59806 -79610
rect 59916 -79720 59926 -79610
rect 59796 -79730 59926 -79720
rect 60436 -79630 60536 -79610
rect 60436 -79750 60446 -79630
rect 60526 -79750 60536 -79630
rect 60436 -79760 60536 -79750
rect 58396 -79830 59716 -79820
rect 56654 -79868 56998 -79858
rect 55520 -80268 55530 -80178
rect 55610 -80268 55980 -80178
rect 54130 -80548 54140 -80288
rect 54850 -80548 54860 -80288
rect 55310 -80468 55320 -80328
rect 55470 -80468 55480 -80328
rect 56170 -80538 56390 -80008
rect 58396 -79900 58906 -79830
rect 58986 -79900 59146 -79830
rect 59226 -79900 59276 -79830
rect 59356 -79900 59396 -79830
rect 59476 -79840 59716 -79830
rect 59476 -79900 59646 -79840
rect 59706 -79900 59716 -79840
rect 58396 -79910 59716 -79900
rect 58396 -79950 58896 -79910
rect 59646 -79920 59716 -79910
rect 56654 -80096 56998 -80086
rect 59006 -80000 60416 -79990
rect 59006 -80040 60266 -80000
rect 59006 -80110 59016 -80040
rect 59076 -80110 59546 -80040
rect 59606 -80110 60266 -80040
rect 59006 -80130 60266 -80110
rect 60406 -80130 60416 -80000
rect 59006 -80140 60416 -80130
rect 59986 -80190 60116 -80180
rect 58956 -80200 59156 -80190
rect 58956 -80380 58966 -80200
rect 59146 -80380 59156 -80200
rect 59986 -80300 59996 -80190
rect 60106 -80300 60116 -80190
rect 58956 -80390 59156 -80380
rect 55680 -80548 56390 -80538
rect 54130 -80708 56390 -80548
rect 55680 -80718 56390 -80708
rect 59600 -80400 60500 -80300
rect 59600 -80800 59700 -80400
rect 60400 -80800 60500 -80400
rect 55400 -80900 56300 -80800
rect 59600 -80900 60500 -80800
rect 68900 -80400 69400 -49900
rect 68900 -80800 69000 -80400
rect 69300 -80800 69400 -80400
rect 68900 -80900 69400 -80800
rect 69900 -50100 70400 -50000
rect 69900 -50300 70000 -50100
rect 70300 -50300 70400 -50100
rect 72810 -50040 73050 -50030
rect 72810 -50220 72820 -50040
rect 73040 -50220 73050 -50040
rect 72810 -50230 73050 -50220
rect 73210 -50060 73350 -47440
rect 73210 -50200 73220 -50060
rect 73340 -50200 73350 -50060
rect 73210 -50230 73350 -50200
rect 73460 -46400 73600 -46390
rect 73460 -46590 73470 -46400
rect 73590 -46590 73600 -46400
rect 73460 -47160 73600 -46590
rect 73460 -47220 73480 -47160
rect 73580 -47220 73600 -47160
rect 73460 -49690 73600 -47220
rect 73460 -49830 73470 -49690
rect 73590 -49830 73600 -49690
rect 55400 -81300 55500 -80900
rect 56200 -81300 56300 -80900
rect 55400 -81400 56300 -81300
rect 51400 -82100 51500 -81900
rect 52500 -82100 52600 -81900
rect 37100 -86700 37200 -86200
rect 37700 -86700 37800 -86200
rect 51400 -86700 52600 -82100
rect 55420 -81880 55740 -81860
rect 55420 -82160 55440 -81880
rect 55720 -82160 55740 -81880
rect 55420 -82180 55740 -82160
rect 54140 -82338 56390 -82328
rect 53460 -82540 53800 -82520
rect 53460 -82740 53480 -82540
rect 53780 -82740 53800 -82540
rect 54140 -82578 54150 -82338
rect 54860 -82578 56390 -82338
rect 58946 -82470 59146 -82450
rect 54140 -82588 56390 -82578
rect 53460 -82760 53800 -82740
rect 54850 -82818 55530 -82808
rect 53510 -82968 53520 -82858
rect 53640 -82968 53650 -82858
rect 54740 -82918 54750 -82838
rect 54850 -82888 55430 -82818
rect 55520 -82888 55530 -82818
rect 55950 -82888 55960 -82738
rect 56040 -82888 56050 -82738
rect 56170 -82758 56390 -82588
rect 56506 -82580 57016 -82570
rect 54840 -82918 54850 -82908
rect 55270 -83008 55280 -82918
rect 55400 -83008 55410 -82918
rect 56170 -82968 56190 -82758
rect 56390 -82968 56400 -82758
rect 58946 -82630 58966 -82470
rect 59126 -82630 59146 -82470
rect 58946 -82650 59146 -82630
rect 59316 -82500 60176 -82490
rect 59316 -82510 59956 -82500
rect 59316 -82650 59336 -82510
rect 59416 -82650 59956 -82510
rect 59316 -82660 59956 -82650
rect 60166 -82660 60176 -82500
rect 59316 -82670 60176 -82660
rect 56506 -82840 57016 -82830
rect 58956 -82720 61136 -82710
rect 58956 -82730 61056 -82720
rect 58956 -82840 58996 -82730
rect 59106 -82740 61056 -82730
rect 59106 -82840 59516 -82740
rect 59616 -82840 61056 -82740
rect 58396 -82930 58896 -82840
rect 58956 -82850 61056 -82840
rect 61126 -82850 61136 -82720
rect 58956 -82860 61136 -82850
rect 55850 -83048 55880 -83018
rect 53940 -83078 55880 -83048
rect 53940 -83098 54920 -83078
rect 53040 -84908 53050 -83158
rect 53250 -84908 53260 -83158
rect 53940 -83198 53950 -83098
rect 54020 -83148 54920 -83098
rect 54020 -83198 54030 -83148
rect 54910 -83168 54920 -83148
rect 54990 -83098 55880 -83078
rect 55970 -83048 55980 -83018
rect 54990 -83148 55970 -83098
rect 54990 -83168 55000 -83148
rect 55220 -83428 55230 -83258
rect 55320 -83428 55330 -83258
rect 55420 -83418 55430 -83248
rect 55510 -83258 55520 -83248
rect 55510 -83268 56670 -83258
rect 55510 -83398 55600 -83268
rect 55710 -83398 56590 -83268
rect 56660 -83398 56670 -83268
rect 55510 -83408 56670 -83398
rect 58396 -83290 58486 -82930
rect 58816 -82950 58896 -82930
rect 59646 -82950 59706 -82930
rect 58816 -82970 59706 -82950
rect 58816 -83030 58906 -82970
rect 58966 -83030 59216 -82970
rect 59276 -83030 59326 -82970
rect 59386 -83030 59436 -82970
rect 59496 -83030 59636 -82970
rect 59696 -83030 59706 -82970
rect 58816 -83040 59706 -83030
rect 58816 -83290 58896 -83040
rect 59536 -83090 59616 -83080
rect 59276 -83130 59356 -83120
rect 59276 -83190 59286 -83130
rect 59346 -83190 59356 -83130
rect 59536 -83150 59546 -83090
rect 59606 -83150 59616 -83090
rect 59536 -83170 59616 -83150
rect 58996 -83200 59076 -83190
rect 58996 -83260 59006 -83200
rect 59076 -83220 59086 -83200
rect 59536 -83210 59616 -83200
rect 59536 -83220 59546 -83210
rect 59076 -83260 59546 -83220
rect 58996 -83270 59076 -83260
rect 59536 -83270 59546 -83260
rect 59606 -83270 59616 -83210
rect 59536 -83280 59616 -83270
rect 58396 -83310 58896 -83290
rect 59646 -83310 59706 -83040
rect 60436 -83120 60536 -83110
rect 59856 -83140 59976 -83130
rect 59856 -83230 59866 -83140
rect 59966 -83230 59976 -83140
rect 60436 -83220 60446 -83120
rect 60526 -83220 60536 -83120
rect 60436 -83230 60536 -83220
rect 59856 -83240 59976 -83230
rect 58396 -83320 59706 -83310
rect 58396 -83330 59216 -83320
rect 58396 -83390 58906 -83330
rect 58966 -83380 59216 -83330
rect 59276 -83380 59336 -83320
rect 59396 -83380 59436 -83320
rect 59496 -83330 59706 -83320
rect 59496 -83380 59636 -83330
rect 58966 -83390 59636 -83380
rect 59696 -83390 59706 -83330
rect 58396 -83400 59706 -83390
rect 60036 -83320 60136 -83310
rect 60036 -83400 60046 -83320
rect 60126 -83400 60136 -83320
rect 55510 -83418 55520 -83408
rect 59646 -83410 59706 -83400
rect 60546 -83410 60636 -83400
rect 59066 -83440 59176 -83430
rect 59066 -83510 59076 -83440
rect 59166 -83510 59176 -83440
rect 59846 -83480 59856 -83410
rect 59916 -83430 59926 -83410
rect 60356 -83420 60556 -83410
rect 60356 -83430 60376 -83420
rect 59916 -83460 60376 -83430
rect 59916 -83480 59926 -83460
rect 60356 -83480 60376 -83460
rect 60446 -83480 60556 -83420
rect 60356 -83490 60556 -83480
rect 60626 -83490 60636 -83410
rect 59066 -83520 59176 -83510
rect 59966 -83500 60326 -83490
rect 53850 -83638 53860 -83528
rect 53920 -83538 55600 -83528
rect 53920 -83638 55000 -83538
rect 55090 -83638 55540 -83538
rect 55630 -83638 55640 -83538
rect 59966 -83560 59976 -83500
rect 60316 -83560 60326 -83500
rect 60546 -83510 60636 -83490
rect 61186 -83520 61366 -83510
rect 54770 -83838 54850 -83638
rect 56470 -83648 56480 -83588
rect 56550 -83648 56560 -83588
rect 57088 -83704 57098 -83564
rect 57368 -83704 57378 -83564
rect 59166 -83630 59376 -83620
rect 59166 -83640 59286 -83630
rect 59166 -83720 59176 -83640
rect 59236 -83720 59286 -83640
rect 59366 -83720 59376 -83630
rect 59166 -83730 59376 -83720
rect 59526 -83670 59646 -83650
rect 59526 -83730 59576 -83670
rect 59636 -83730 59646 -83670
rect 61186 -83700 61206 -83520
rect 61346 -83700 61366 -83520
rect 61186 -83710 61366 -83700
rect 59526 -83760 59646 -83730
rect 60286 -83750 60476 -83740
rect 59906 -83780 60016 -83770
rect 59806 -83790 59866 -83780
rect 54760 -83928 54770 -83838
rect 54840 -83928 54850 -83838
rect 59166 -83840 59536 -83830
rect 59166 -83920 59176 -83840
rect 59236 -83920 59286 -83840
rect 54920 -83938 55210 -83928
rect 54920 -84008 55140 -83938
rect 55200 -84008 55210 -83938
rect 59166 -83930 59286 -83920
rect 59356 -83850 59536 -83840
rect 59356 -83920 59476 -83850
rect 59356 -83930 59536 -83920
rect 59166 -83940 59536 -83930
rect 59566 -83960 59576 -83790
rect 59636 -83800 59866 -83790
rect 59636 -83940 59806 -83800
rect 59636 -83960 59866 -83940
rect 59906 -83960 59916 -83780
rect 60006 -83960 60016 -83780
rect 60286 -83890 60306 -83750
rect 60456 -83890 60476 -83750
rect 60286 -83900 60476 -83890
rect 61026 -83820 61136 -83810
rect 61026 -83930 61036 -83820
rect 61126 -83930 61136 -83820
rect 61026 -83940 61136 -83930
rect 59566 -83970 59636 -83960
rect 59906 -83970 60016 -83960
rect 54760 -84328 54770 -84248
rect 54840 -84328 54850 -84248
rect 54770 -84538 54850 -84328
rect 54920 -84398 54980 -84008
rect 55880 -84038 56900 -84018
rect 55010 -84128 55020 -84048
rect 55120 -84128 55740 -84048
rect 55810 -84128 55820 -84048
rect 55870 -84128 55880 -84038
rect 55970 -84128 56480 -84038
rect 56550 -84128 56900 -84038
rect 55880 -84148 56900 -84128
rect 57020 -84020 57040 -84018
rect 57800 -84020 58240 -84010
rect 57020 -84140 57800 -84020
rect 57020 -84148 57040 -84140
rect 57800 -84150 58240 -84140
rect 58516 -84060 58796 -83990
rect 58516 -84260 58556 -84060
rect 58756 -84260 58796 -84060
rect 59066 -84010 59936 -84000
rect 59066 -84080 59076 -84010
rect 59166 -84030 59826 -84010
rect 59166 -84080 59316 -84030
rect 59066 -84090 59316 -84080
rect 59376 -84080 59826 -84030
rect 59916 -84080 59936 -84010
rect 59376 -84090 59936 -84080
rect 60076 -84080 60196 -84040
rect 59066 -84170 59936 -84160
rect 59066 -84240 59076 -84170
rect 59166 -84240 59206 -84170
rect 59266 -84240 59826 -84170
rect 59926 -84240 59936 -84170
rect 59066 -84250 59936 -84240
rect 60076 -84240 60096 -84080
rect 60176 -84240 60196 -84080
rect 58516 -84340 58796 -84260
rect 60076 -84280 60196 -84240
rect 61266 -84050 61366 -84040
rect 61266 -84260 61276 -84050
rect 61356 -84260 61366 -84050
rect 61266 -84270 61366 -84260
rect 59586 -84290 59656 -84280
rect 59796 -84290 59866 -84280
rect 59586 -84310 59796 -84290
rect 59156 -84320 59536 -84310
rect 59156 -84330 59266 -84320
rect 54910 -84468 54920 -84398
rect 54980 -84468 54990 -84398
rect 59156 -84410 59166 -84330
rect 59226 -84410 59266 -84330
rect 59366 -84330 59536 -84320
rect 59366 -84410 59466 -84330
rect 59526 -84410 59536 -84330
rect 59156 -84430 59536 -84410
rect 59646 -84450 59796 -84310
rect 59586 -84470 59796 -84450
rect 59856 -84470 59866 -84290
rect 53840 -84648 53850 -84538
rect 53920 -84638 55000 -84538
rect 55090 -84638 55540 -84538
rect 55630 -84638 55640 -84538
rect 56470 -84588 56480 -84528
rect 56550 -84588 56560 -84528
rect 57088 -84614 57098 -84474
rect 57368 -84614 57378 -84474
rect 59796 -84480 59866 -84470
rect 59906 -84290 60016 -84280
rect 59906 -84480 59916 -84290
rect 60006 -84480 60016 -84290
rect 60476 -84310 60546 -84300
rect 60536 -84370 60546 -84310
rect 60476 -84380 60546 -84370
rect 60966 -84430 61486 -84420
rect 60966 -84440 61336 -84430
rect 59906 -84490 60016 -84480
rect 60466 -84450 61336 -84440
rect 59506 -84510 59606 -84500
rect 59156 -84560 59376 -84540
rect 53920 -84648 55640 -84638
rect 59156 -84640 59166 -84560
rect 59226 -84640 59266 -84560
rect 59156 -84650 59266 -84640
rect 59366 -84650 59376 -84560
rect 59506 -84580 59516 -84510
rect 59596 -84580 59606 -84510
rect 60466 -84510 60476 -84450
rect 60536 -84510 60616 -84450
rect 60736 -84510 60756 -84450
rect 60816 -84510 60896 -84450
rect 60956 -84510 61336 -84450
rect 60466 -84520 61336 -84510
rect 60966 -84560 61336 -84520
rect 61456 -84560 61486 -84430
rect 60966 -84570 61486 -84560
rect 59506 -84590 59606 -84580
rect 59156 -84660 59376 -84650
rect 59306 -84720 60336 -84700
rect 59066 -84740 59176 -84730
rect 55210 -84918 55220 -84748
rect 55310 -84918 55320 -84748
rect 55400 -84928 55410 -84758
rect 55500 -84768 55510 -84758
rect 55500 -84888 56380 -84768
rect 56440 -84888 56450 -84768
rect 59066 -84800 59076 -84740
rect 59166 -84800 59176 -84740
rect 59306 -84780 59316 -84720
rect 59376 -84740 59966 -84720
rect 59376 -84780 59816 -84740
rect 59306 -84790 59816 -84780
rect 59846 -84780 59916 -84770
rect 59066 -84810 59176 -84800
rect 59846 -84840 59856 -84780
rect 59946 -84780 59966 -84740
rect 60326 -84780 60336 -84720
rect 59946 -84790 60336 -84780
rect 60366 -84740 61146 -84730
rect 60366 -84780 61056 -84740
rect 59646 -84850 59716 -84840
rect 59846 -84850 59916 -84840
rect 60366 -84840 60376 -84780
rect 60436 -84840 61056 -84780
rect 61126 -84840 61146 -84740
rect 55500 -84908 56450 -84888
rect 58396 -84860 59716 -84850
rect 55500 -84928 55510 -84908
rect 58396 -84930 58926 -84860
rect 58986 -84930 59146 -84860
rect 59226 -84930 59276 -84860
rect 59356 -84930 59396 -84860
rect 59476 -84920 59646 -84860
rect 59706 -84920 59716 -84860
rect 60366 -84870 61146 -84840
rect 59476 -84930 59716 -84920
rect 58396 -84940 59716 -84930
rect 54900 -85008 54910 -84998
rect 53940 -85088 53950 -85008
rect 54010 -85088 54910 -85008
rect 53940 -85098 54910 -85088
rect 54980 -85018 54990 -84998
rect 54980 -85078 55980 -85018
rect 54980 -85098 55880 -85078
rect 53940 -85118 55880 -85098
rect 53500 -85248 53510 -85128
rect 53630 -85248 53640 -85128
rect 55850 -85158 55880 -85118
rect 55970 -85158 55980 -85078
rect 55230 -85218 55240 -85158
rect 55370 -85178 55710 -85158
rect 55370 -85188 55720 -85178
rect 55370 -85208 55620 -85188
rect 55370 -85218 55380 -85208
rect 55400 -85268 55410 -85248
rect 54730 -85358 54740 -85268
rect 54850 -85338 55410 -85268
rect 55510 -85338 55520 -85248
rect 55600 -85278 55620 -85208
rect 55710 -85278 55720 -85188
rect 54850 -85358 55520 -85338
rect 55210 -85528 55220 -85418
rect 55330 -85528 55340 -85418
rect 55850 -85578 55980 -85158
rect 56010 -85408 56020 -85258
rect 56080 -85408 56090 -85258
rect 56160 -85408 56170 -85208
rect 56390 -85408 56400 -85208
rect 58396 -85220 58896 -84940
rect 59006 -85100 59076 -85080
rect 59246 -85090 59256 -85030
rect 59366 -85090 59376 -85030
rect 59536 -85060 59546 -84990
rect 59606 -85060 59616 -84990
rect 59536 -85070 59616 -85060
rect 59006 -85160 59016 -85100
rect 59536 -85110 59616 -85100
rect 59076 -85120 59086 -85110
rect 59536 -85120 59546 -85110
rect 59076 -85160 59546 -85120
rect 59006 -85170 59546 -85160
rect 59606 -85170 59616 -85110
rect 59006 -85190 59076 -85170
rect 59536 -85190 59616 -85170
rect 59646 -85220 59716 -84940
rect 59796 -85010 59926 -85000
rect 59796 -85120 59806 -85010
rect 59916 -85120 59926 -85010
rect 59796 -85130 59926 -85120
rect 60436 -85030 60536 -85010
rect 60436 -85150 60446 -85030
rect 60526 -85150 60536 -85030
rect 60436 -85160 60536 -85150
rect 58396 -85230 59716 -85220
rect 56654 -85268 56998 -85258
rect 55520 -85668 55530 -85578
rect 55610 -85668 55980 -85578
rect 54130 -85948 54140 -85688
rect 54850 -85948 54860 -85688
rect 55310 -85868 55320 -85728
rect 55470 -85868 55480 -85728
rect 56170 -85938 56390 -85408
rect 58396 -85300 58906 -85230
rect 58986 -85300 59146 -85230
rect 59226 -85300 59276 -85230
rect 59356 -85300 59396 -85230
rect 59476 -85240 59716 -85230
rect 59476 -85300 59646 -85240
rect 59706 -85300 59716 -85240
rect 58396 -85310 59716 -85300
rect 58396 -85350 58896 -85310
rect 59646 -85320 59716 -85310
rect 56654 -85496 56998 -85486
rect 59006 -85400 60416 -85390
rect 59006 -85440 60266 -85400
rect 59006 -85510 59016 -85440
rect 59076 -85510 59546 -85440
rect 59606 -85510 60266 -85440
rect 59006 -85530 60266 -85510
rect 60406 -85530 60416 -85400
rect 59006 -85540 60416 -85530
rect 59986 -85590 60116 -85580
rect 58956 -85600 59156 -85590
rect 58956 -85780 58966 -85600
rect 59146 -85780 59156 -85600
rect 59986 -85700 59996 -85590
rect 60106 -85700 60116 -85590
rect 58956 -85790 59156 -85780
rect 55680 -85948 56390 -85938
rect 54130 -86108 56390 -85948
rect 55680 -86118 56390 -86108
rect 59600 -85800 60500 -85700
rect 59600 -86200 59700 -85800
rect 60400 -86200 60500 -85800
rect 55400 -86300 56200 -86200
rect 59600 -86300 60500 -86200
rect 69900 -85800 70400 -50300
rect 73460 -52420 73600 -49830
rect 73710 -46400 73850 -46390
rect 73710 -46590 73720 -46400
rect 73840 -46590 73850 -46400
rect 73710 -46636 73850 -46590
rect 73710 -46688 73723 -46636
rect 73840 -46688 73850 -46636
rect 73710 -47270 73850 -46688
rect 73710 -47330 73730 -47270
rect 73830 -47330 73850 -47270
rect 73710 -49240 73850 -47330
rect 73710 -49380 73720 -49240
rect 73840 -49380 73850 -49240
rect 73710 -50970 73850 -49380
rect 73710 -51040 73720 -50970
rect 73840 -51040 73850 -50970
rect 73710 -51050 73850 -51040
rect 73960 -46400 74100 -46390
rect 73960 -46590 73970 -46400
rect 74090 -46590 74100 -46400
rect 73960 -47470 74100 -46590
rect 73960 -47530 73970 -47470
rect 74090 -47530 74100 -47470
rect 73960 -48840 74100 -47530
rect 74210 -46400 74350 -46390
rect 74210 -46590 74220 -46400
rect 74340 -46590 74350 -46400
rect 74210 -46800 74350 -46590
rect 74210 -46880 74220 -46800
rect 74340 -46880 74350 -46800
rect 74210 -47930 74350 -46880
rect 74210 -47990 74230 -47930
rect 74330 -47990 74350 -47930
rect 74210 -48430 74350 -47990
rect 74210 -48490 74220 -48430
rect 74340 -48490 74350 -48430
rect 74210 -48500 74350 -48490
rect 74460 -46400 74600 -46390
rect 74460 -46590 74470 -46400
rect 74590 -46590 74600 -46400
rect 74460 -46610 74600 -46590
rect 74460 -46714 74477 -46610
rect 74594 -46714 74600 -46610
rect 74460 -48150 74600 -46714
rect 74460 -48220 74470 -48150
rect 74590 -48220 74600 -48150
rect 73960 -48980 73970 -48840
rect 74090 -48980 74100 -48840
rect 73460 -52480 73470 -52420
rect 73590 -52480 73600 -52420
rect 73460 -52500 73600 -52480
rect 73960 -51800 74100 -48980
rect 73960 -51870 73970 -51800
rect 74090 -51870 74100 -51800
rect 73960 -52780 74100 -51870
rect 73960 -52840 73970 -52780
rect 74090 -52840 74100 -52780
rect 73960 -52850 74100 -52840
rect 74460 -49360 74600 -48220
rect 74460 -49420 74470 -49360
rect 74590 -49420 74600 -49360
rect 74460 -53520 74600 -49420
rect 74710 -46400 74850 -46390
rect 74710 -46590 74720 -46400
rect 74840 -46590 74850 -46400
rect 74710 -46792 74850 -46590
rect 74710 -46870 74724 -46792
rect 74841 -46870 74850 -46792
rect 74710 -47740 74850 -46870
rect 74710 -47880 74720 -47740
rect 74840 -47880 74850 -47740
rect 74710 -48020 74850 -47880
rect 74710 -48080 74730 -48020
rect 74830 -48080 74850 -48020
rect 74710 -49670 74850 -48080
rect 74710 -49730 74720 -49670
rect 74840 -49730 74850 -49670
rect 74710 -49740 74850 -49730
rect 74960 -46400 75100 -46390
rect 74960 -46590 74970 -46400
rect 75090 -46590 75100 -46400
rect 74960 -47260 75100 -46590
rect 74960 -47380 74970 -47260
rect 75090 -47380 75100 -47260
rect 74960 -47820 75100 -47380
rect 74960 -47890 74980 -47820
rect 75080 -47890 75100 -47820
rect 74960 -50310 75100 -47890
rect 74960 -50370 74970 -50310
rect 75090 -50370 75100 -50310
rect 74960 -50380 75100 -50370
rect 75210 -46400 75350 -46390
rect 75210 -46590 75220 -46400
rect 75340 -46590 75350 -46400
rect 76910 -46450 77070 -46440
rect 75210 -47080 75350 -46590
rect 76635 -46480 76739 -46467
rect 76635 -46545 76648 -46480
rect 76726 -46545 76739 -46480
rect 75400 -46630 75480 -46620
rect 75400 -46690 75410 -46630
rect 75470 -46690 75480 -46630
rect 75400 -46700 75480 -46690
rect 75647 -46623 75777 -46610
rect 75400 -46701 75478 -46700
rect 75647 -46701 75673 -46623
rect 75751 -46701 75777 -46623
rect 75210 -47180 75220 -47080
rect 75340 -47180 75350 -47080
rect 75647 -47130 75777 -46701
rect 75933 -46623 76063 -46610
rect 75933 -46701 75946 -46623
rect 76024 -46701 76063 -46623
rect 75933 -46980 76063 -46701
rect 76102 -46623 76193 -46610
rect 76180 -46701 76193 -46623
rect 76102 -46714 76193 -46701
rect 76230 -46623 76323 -46610
rect 76230 -46701 76232 -46623
rect 76310 -46701 76323 -46623
rect 76230 -46710 76323 -46701
rect 76232 -46922 76323 -46710
rect 76360 -46640 76460 -46620
rect 76360 -46700 76380 -46640
rect 76440 -46700 76460 -46640
rect 76360 -46720 76460 -46700
rect 76492 -46636 76596 -46623
rect 76492 -46701 76505 -46636
rect 76583 -46701 76596 -46636
rect 76492 -46714 76596 -46701
rect 76362 -46766 76453 -46720
rect 76362 -46844 76375 -46766
rect 76440 -46844 76453 -46766
rect 76362 -46857 76453 -46844
rect 75210 -48580 75350 -47180
rect 75210 -48650 75220 -48580
rect 75340 -48650 75350 -48580
rect 75210 -49200 75350 -48650
rect 75210 -49280 75220 -49200
rect 75340 -49280 75350 -49200
rect 75210 -49810 75350 -49280
rect 75210 -49900 75220 -49810
rect 75340 -49900 75350 -49810
rect 74460 -53600 74470 -53520
rect 74590 -53600 74600 -53520
rect 74460 -53610 74600 -53600
rect 75210 -50450 75350 -49900
rect 75210 -50540 75220 -50450
rect 75340 -50540 75350 -50450
rect 75210 -51230 75350 -50540
rect 75210 -51290 75220 -51230
rect 75340 -51290 75350 -51230
rect 75210 -51660 75350 -51290
rect 75210 -51720 75220 -51660
rect 75340 -51720 75350 -51660
rect 75210 -53010 75350 -51720
rect 75640 -52310 75780 -47130
rect 75640 -52370 75660 -52310
rect 75760 -52370 75780 -52310
rect 75920 -51120 76070 -46980
rect 76219 -47120 76323 -46922
rect 76505 -47050 76596 -46714
rect 76635 -46636 76739 -46545
rect 76910 -46570 76920 -46450
rect 77060 -46570 77070 -46450
rect 76910 -46580 77070 -46570
rect 76635 -46714 76648 -46636
rect 76726 -46714 76739 -46636
rect 76635 -46727 76739 -46714
rect 76770 -46636 76870 -46620
rect 76770 -46670 76791 -46636
rect 76843 -46670 76870 -46636
rect 76770 -46740 76780 -46670
rect 76860 -46740 76870 -46670
rect 76770 -46760 76870 -46740
rect 78270 -46670 78360 -46660
rect 78270 -46740 78280 -46670
rect 78350 -46740 78360 -46670
rect 77160 -46830 77440 -46820
rect 75920 -51180 75940 -51120
rect 76050 -51180 76070 -51120
rect 76200 -51110 76350 -47120
rect 76200 -51170 76210 -51110
rect 76340 -51170 76350 -51110
rect 76200 -51180 76350 -51170
rect 75920 -52190 76070 -51180
rect 75920 -52280 75940 -52190
rect 76050 -52280 76070 -52190
rect 75920 -52880 76070 -52280
rect 75920 -52940 75940 -52880
rect 76050 -52940 76070 -52880
rect 76480 -52290 76620 -47050
rect 77160 -47080 77170 -46830
rect 77430 -47080 77440 -46830
rect 77160 -47090 77440 -47080
rect 78140 -47380 78220 -47370
rect 78140 -47440 78150 -47380
rect 78210 -47440 78220 -47380
rect 77220 -47480 77320 -47470
rect 77220 -47540 77230 -47480
rect 77310 -47540 77320 -47480
rect 77220 -47550 77320 -47540
rect 76910 -47610 77070 -47600
rect 76910 -47760 76920 -47610
rect 77060 -47760 77070 -47610
rect 76910 -47770 77070 -47760
rect 77160 -47820 77270 -47810
rect 77160 -47890 77170 -47820
rect 77260 -47890 77270 -47820
rect 77160 -47900 77270 -47890
rect 78140 -47830 78220 -47440
rect 78270 -47380 78360 -46740
rect 78270 -47440 78280 -47380
rect 78340 -47440 78360 -47380
rect 78270 -47450 78360 -47440
rect 78570 -47360 78650 -47350
rect 78570 -47420 78580 -47360
rect 78640 -47420 78650 -47360
rect 78140 -48120 78150 -47830
rect 78210 -48120 78220 -47830
rect 78570 -47880 78650 -47420
rect 78790 -47370 78870 -46320
rect 80050 -47310 80460 -47280
rect 78790 -47430 78800 -47370
rect 78860 -47430 78870 -47370
rect 78790 -47440 78870 -47430
rect 79060 -47390 79270 -47370
rect 79060 -47550 79080 -47390
rect 79250 -47550 79270 -47390
rect 79060 -47560 79270 -47550
rect 80050 -47620 80080 -47310
rect 80430 -47620 80460 -47310
rect 80050 -47650 80460 -47620
rect 78570 -47940 78580 -47880
rect 78640 -47940 78650 -47880
rect 78570 -47960 78650 -47940
rect 80050 -47720 80460 -47690
rect 78140 -48140 78220 -48120
rect 80050 -48100 80080 -47720
rect 80430 -48100 80460 -47720
rect 80050 -48130 80460 -48100
rect 77400 -48150 77490 -48140
rect 77400 -48220 77410 -48150
rect 77480 -48220 77490 -48150
rect 77400 -48230 77490 -48220
rect 79400 -48190 79690 -48180
rect 77770 -48430 77850 -48420
rect 77770 -48490 77780 -48430
rect 77840 -48490 77850 -48430
rect 79400 -48430 79410 -48190
rect 79680 -48430 79690 -48190
rect 79400 -48440 79690 -48430
rect 77440 -48580 77530 -48570
rect 77440 -48650 77450 -48580
rect 77520 -48650 77530 -48580
rect 77440 -48660 77530 -48650
rect 77770 -48610 77850 -48490
rect 77770 -48670 77780 -48610
rect 77840 -48670 77850 -48610
rect 77770 -48680 77850 -48670
rect 78300 -48690 78420 -48680
rect 78300 -48800 78310 -48690
rect 78410 -48800 78420 -48690
rect 78300 -48810 78420 -48800
rect 76910 -48860 77070 -48850
rect 76910 -49000 76920 -48860
rect 77060 -49000 77070 -48860
rect 76910 -49010 77070 -49000
rect 78050 -49130 78130 -49120
rect 77770 -49180 77850 -49170
rect 77440 -49200 77540 -49190
rect 77440 -49280 77450 -49200
rect 77530 -49280 77540 -49200
rect 77440 -49290 77540 -49280
rect 77770 -49240 77780 -49180
rect 77840 -49240 77850 -49180
rect 77770 -49360 77850 -49240
rect 77770 -49420 77780 -49360
rect 77840 -49420 77850 -49360
rect 77770 -49430 77850 -49420
rect 78050 -49220 78060 -49130
rect 78120 -49220 78130 -49130
rect 78340 -49170 78420 -48810
rect 80050 -48950 80460 -48920
rect 77770 -49670 77850 -49660
rect 77770 -49730 77780 -49670
rect 77840 -49730 77850 -49670
rect 77480 -49810 77590 -49800
rect 77480 -49900 77490 -49810
rect 77580 -49900 77590 -49810
rect 77480 -49910 77590 -49900
rect 77770 -49850 77850 -49730
rect 77770 -49910 77780 -49850
rect 77840 -49910 77850 -49850
rect 77770 -49920 77850 -49910
rect 76910 -50100 77070 -50090
rect 76910 -50260 76920 -50100
rect 77060 -50260 77070 -50100
rect 76910 -50270 77070 -50260
rect 77770 -50310 77850 -50300
rect 77770 -50370 77780 -50310
rect 77840 -50370 77850 -50310
rect 77770 -50420 77850 -50370
rect 77460 -50450 77570 -50440
rect 77460 -50540 77470 -50450
rect 77560 -50540 77570 -50450
rect 77770 -50480 77780 -50420
rect 77840 -50480 77850 -50420
rect 77770 -50490 77850 -50480
rect 78050 -50370 78130 -49220
rect 78160 -49180 78300 -49170
rect 78160 -49280 78180 -49180
rect 78290 -49280 78300 -49180
rect 78340 -49230 78350 -49170
rect 78410 -49230 78420 -49170
rect 78340 -49240 78420 -49230
rect 78660 -49070 78790 -49060
rect 78160 -49300 78300 -49280
rect 78200 -49760 78300 -49300
rect 78660 -49420 78670 -49070
rect 78780 -49420 78790 -49070
rect 80050 -49330 80080 -48950
rect 80430 -49330 80460 -48950
rect 80050 -49360 80460 -49330
rect 78660 -49430 78790 -49420
rect 79400 -49420 79690 -49410
rect 79400 -49660 79410 -49420
rect 79680 -49660 79690 -49420
rect 79400 -49670 79690 -49660
rect 78160 -49770 78300 -49760
rect 78160 -50040 78170 -49770
rect 78290 -50040 78300 -49770
rect 78160 -50050 78300 -50040
rect 78520 -49770 78600 -49760
rect 78520 -50040 78530 -49770
rect 78590 -50040 78600 -49770
rect 78050 -50380 78310 -50370
rect 77460 -50550 77570 -50540
rect 78050 -50680 78060 -50380
rect 78120 -50410 78310 -50380
rect 78120 -50510 78160 -50410
rect 78260 -50510 78310 -50410
rect 78120 -50680 78310 -50510
rect 78050 -50690 78310 -50680
rect 78520 -50570 78600 -50040
rect 79040 -50400 79170 -50380
rect 79040 -50510 79050 -50400
rect 79150 -50510 79170 -50400
rect 78520 -50690 78710 -50570
rect 78230 -50920 78310 -50690
rect 77460 -50970 77550 -50960
rect 77460 -51040 77470 -50970
rect 77540 -51040 77550 -50970
rect 78230 -50980 78240 -50920
rect 78300 -50980 78310 -50920
rect 78230 -50990 78310 -50980
rect 77460 -51050 77550 -51040
rect 77850 -51090 77930 -51080
rect 77190 -51120 77270 -51110
rect 77190 -51180 77200 -51120
rect 77260 -51180 77270 -51120
rect 77850 -51150 77860 -51090
rect 77920 -51150 77930 -51090
rect 78620 -51120 78710 -50690
rect 77850 -51160 77930 -51150
rect 76910 -51350 77070 -51340
rect 76910 -51490 76920 -51350
rect 77060 -51490 77070 -51350
rect 76910 -51500 77070 -51490
rect 77190 -51570 77270 -51180
rect 77190 -51630 77200 -51570
rect 77260 -51630 77270 -51570
rect 77190 -51640 77270 -51630
rect 77860 -51540 77920 -51160
rect 78340 -51180 78410 -51120
rect 77950 -51230 78030 -51220
rect 77950 -51290 77960 -51230
rect 78020 -51290 78030 -51230
rect 78620 -51180 78630 -51120
rect 78700 -51180 78710 -51120
rect 78620 -51190 78710 -51180
rect 78850 -50960 78990 -50950
rect 78340 -51250 78410 -51240
rect 78850 -51250 78860 -50960
rect 78980 -51250 78990 -50960
rect 77950 -51300 78030 -51290
rect 78350 -51520 78400 -51250
rect 78850 -51260 78990 -51250
rect 78240 -51540 78420 -51520
rect 77860 -51720 77920 -51710
rect 77960 -51660 78040 -51650
rect 77960 -51720 77970 -51660
rect 78030 -51720 78040 -51660
rect 77960 -51730 78040 -51720
rect 77420 -51800 77510 -51790
rect 77420 -51870 77430 -51800
rect 77500 -51870 77510 -51800
rect 77420 -51880 77510 -51870
rect 78300 -51910 78420 -51540
rect 78240 -51920 78420 -51910
rect 76480 -52350 76490 -52290
rect 76610 -52350 76620 -52290
rect 76480 -52920 76620 -52350
rect 78170 -52170 78310 -52160
rect 77960 -52390 78040 -52380
rect 77750 -52460 77830 -52450
rect 77750 -52520 77760 -52460
rect 77820 -52520 77830 -52460
rect 77960 -52510 77970 -52390
rect 78030 -52510 78040 -52390
rect 77960 -52520 78040 -52510
rect 78170 -52510 78180 -52170
rect 78300 -52510 78310 -52170
rect 77750 -52530 77830 -52520
rect 78170 -52550 78310 -52510
rect 76910 -52560 77070 -52550
rect 76910 -52650 76920 -52560
rect 77060 -52650 77070 -52560
rect 76910 -52660 77070 -52650
rect 77750 -52780 77830 -52770
rect 77750 -52840 77760 -52780
rect 77820 -52840 77830 -52780
rect 77750 -52850 77830 -52840
rect 75210 -53100 75230 -53010
rect 75330 -53100 75350 -53010
rect 75210 -53540 75350 -53100
rect 76480 -52990 76490 -52920
rect 76610 -52990 76620 -52920
rect 77950 -52890 78030 -52880
rect 77950 -52960 77960 -52890
rect 78020 -52960 78030 -52890
rect 77950 -52970 78030 -52960
rect 76480 -53390 76620 -52990
rect 76480 -53460 76500 -53390
rect 76600 -53460 76620 -53390
rect 75210 -53610 75230 -53540
rect 75330 -53610 75350 -53540
rect 75210 -53930 75350 -53610
rect 78060 -53520 78150 -53510
rect 78060 -53630 78070 -53520
rect 78140 -53630 78150 -53520
rect 77590 -53650 77720 -53640
rect 76910 -53680 77070 -53670
rect 76910 -53780 76920 -53680
rect 77060 -53780 77070 -53680
rect 77590 -53720 77600 -53650
rect 77710 -53720 77720 -53650
rect 77590 -53730 77720 -53720
rect 76910 -53790 77070 -53780
rect 75210 -53990 75220 -53930
rect 75340 -53990 75350 -53930
rect 75210 -54000 75350 -53990
rect 78060 -53930 78150 -53630
rect 78230 -53570 78310 -52550
rect 78770 -52810 78930 -52800
rect 78770 -52930 78780 -52810
rect 78920 -52930 78930 -52810
rect 79040 -52840 79170 -50510
rect 79400 -50680 79690 -50670
rect 79400 -50920 79410 -50680
rect 79680 -50920 79690 -50680
rect 79400 -50930 79690 -50920
rect 79980 -50950 80390 -50920
rect 79980 -51330 80010 -50950
rect 80360 -51330 80390 -50950
rect 79980 -51360 80390 -51330
rect 81630 -51680 81770 -45840
rect 81940 -48020 82080 -48010
rect 81940 -48140 81950 -48020
rect 82070 -48140 82080 -48020
rect 81940 -51140 82080 -48140
rect 82210 -48020 82350 -43320
rect 82210 -48140 82220 -48020
rect 82340 -48140 82350 -48020
rect 82210 -48150 82350 -48140
rect 82460 -43890 82560 -43880
rect 82460 -44000 82470 -43890
rect 82550 -44000 82560 -43890
rect 82460 -48920 82560 -44000
rect 82630 -43890 82730 -41320
rect 82810 -42740 91440 -42710
rect 82810 -43310 82820 -42740
rect 91410 -43310 91440 -42740
rect 82810 -43340 91440 -43310
rect 85310 -43450 85400 -43440
rect 85310 -43540 85320 -43450
rect 85390 -43540 85400 -43450
rect 85310 -43810 85400 -43540
rect 82630 -44000 82640 -43890
rect 82720 -44000 82730 -43890
rect 82630 -44010 82730 -44000
rect 83030 -43890 83110 -43880
rect 83030 -44000 83040 -43890
rect 83100 -44000 83110 -43890
rect 83030 -44010 83110 -44000
rect 85310 -44000 85320 -43810
rect 85390 -44000 85400 -43810
rect 85580 -43450 86490 -43440
rect 85580 -43540 85590 -43450
rect 86480 -43540 86490 -43450
rect 85580 -43870 86490 -43540
rect 87030 -43450 87930 -43440
rect 87030 -43540 87040 -43450
rect 87920 -43540 87930 -43450
rect 85580 -43950 85590 -43870
rect 86480 -43950 86490 -43870
rect 85580 -43960 86490 -43950
rect 86790 -43790 86880 -43780
rect 85310 -44010 85400 -44000
rect 86790 -44000 86800 -43790
rect 86870 -44000 86880 -43790
rect 87030 -43870 87930 -43540
rect 88500 -43450 89400 -43440
rect 88500 -43540 88510 -43450
rect 89390 -43540 89400 -43450
rect 87030 -43950 87040 -43870
rect 87920 -43950 87930 -43870
rect 87030 -43960 87930 -43950
rect 88260 -43800 88350 -43790
rect 86790 -44230 86880 -44000
rect 86790 -44310 86800 -44230
rect 86870 -44310 86880 -44230
rect 86790 -44320 86880 -44310
rect 88260 -44000 88270 -43800
rect 88340 -44000 88350 -43800
rect 88500 -43880 89400 -43540
rect 89970 -43450 90770 -43440
rect 89970 -43540 89980 -43450
rect 90760 -43540 90770 -43450
rect 88500 -43950 88510 -43880
rect 89390 -43950 89400 -43880
rect 88500 -43960 89400 -43950
rect 89740 -43800 89820 -43790
rect 88260 -44230 88350 -44000
rect 88260 -44310 88270 -44230
rect 88340 -44310 88350 -44230
rect 88260 -44320 88350 -44310
rect 89810 -44010 89820 -43800
rect 89970 -43879 90770 -43540
rect 89970 -43951 89982 -43879
rect 90762 -43951 90770 -43879
rect 89970 -43961 90770 -43951
rect 91200 -43800 91290 -43790
rect 89740 -44230 89820 -44010
rect 89740 -44310 89750 -44230
rect 89810 -44310 89820 -44230
rect 89740 -44320 89820 -44310
rect 91200 -44010 91210 -43800
rect 91280 -44010 91290 -43800
rect 91200 -44230 91290 -44010
rect 91200 -44310 91210 -44230
rect 91280 -44310 91290 -44230
rect 91200 -44320 91290 -44310
rect 91750 -44080 92160 -44050
rect 82790 -44440 91440 -44410
rect 82790 -45010 82820 -44440
rect 91410 -45010 91440 -44440
rect 91750 -44460 91780 -44080
rect 92130 -44460 92160 -44080
rect 91750 -44490 92160 -44460
rect 82790 -45040 91440 -45010
rect 82794 -46878 91444 -46848
rect 82794 -47448 82824 -46878
rect 91414 -47448 91444 -46878
rect 82794 -47478 91444 -47448
rect 85314 -47588 85404 -47578
rect 85314 -47678 85324 -47588
rect 85394 -47678 85404 -47588
rect 85314 -47948 85404 -47678
rect 83030 -48020 83110 -48010
rect 83030 -48140 83040 -48020
rect 83100 -48140 83110 -48020
rect 83030 -48150 83110 -48140
rect 85314 -48138 85324 -47948
rect 85394 -48138 85404 -47948
rect 85584 -47588 86494 -47578
rect 85584 -47678 85594 -47588
rect 86484 -47678 86494 -47588
rect 85584 -48008 86494 -47678
rect 87034 -47588 87934 -47578
rect 87034 -47678 87044 -47588
rect 87924 -47678 87934 -47588
rect 85584 -48088 85594 -48008
rect 86484 -48088 86494 -48008
rect 85584 -48098 86494 -48088
rect 86794 -47928 86884 -47918
rect 85314 -48148 85404 -48138
rect 86794 -48138 86804 -47928
rect 86874 -48138 86884 -47928
rect 87034 -48008 87934 -47678
rect 88504 -47588 89404 -47578
rect 88504 -47678 88514 -47588
rect 89394 -47678 89404 -47588
rect 87034 -48088 87044 -48008
rect 87924 -48088 87934 -48008
rect 87034 -48098 87934 -48088
rect 88264 -47938 88354 -47928
rect 86794 -48368 86884 -48138
rect 86794 -48448 86804 -48368
rect 86874 -48448 86884 -48368
rect 86794 -48458 86884 -48448
rect 88264 -48138 88274 -47938
rect 88344 -48138 88354 -47938
rect 88504 -48018 89404 -47678
rect 89974 -47588 90774 -47578
rect 89974 -47678 89984 -47588
rect 90764 -47678 90774 -47588
rect 88504 -48088 88514 -48018
rect 89394 -48088 89404 -48018
rect 88504 -48098 89404 -48088
rect 89744 -47938 89824 -47928
rect 88264 -48368 88354 -48138
rect 88264 -48448 88274 -48368
rect 88344 -48448 88354 -48368
rect 88264 -48458 88354 -48448
rect 89814 -48148 89824 -47938
rect 89974 -48017 90774 -47678
rect 89974 -48089 89986 -48017
rect 90766 -48089 90774 -48017
rect 89974 -48099 90774 -48089
rect 91204 -47938 91294 -47928
rect 89744 -48368 89824 -48148
rect 89744 -48448 89754 -48368
rect 89814 -48448 89824 -48368
rect 89744 -48458 89824 -48448
rect 91204 -48148 91214 -47938
rect 91284 -48148 91294 -47938
rect 91204 -48368 91294 -48148
rect 91204 -48448 91214 -48368
rect 91284 -48448 91294 -48368
rect 91204 -48458 91294 -48448
rect 91750 -48240 92160 -48210
rect 82794 -48578 91444 -48548
rect 82420 -48950 82640 -48920
rect 82420 -49330 82450 -48950
rect 82610 -49330 82640 -48950
rect 82794 -49148 82824 -48578
rect 91414 -49148 91444 -48578
rect 91750 -48620 91780 -48240
rect 92130 -48620 92160 -48240
rect 91750 -48650 92160 -48620
rect 82794 -49178 91444 -49148
rect 82420 -49360 82640 -49330
rect 82790 -50530 91440 -50500
rect 82790 -51100 82820 -50530
rect 91410 -51100 91440 -50530
rect 82790 -51130 91440 -51100
rect 81940 -51350 81950 -51140
rect 82070 -51350 82080 -51140
rect 81940 -51360 82080 -51350
rect 85310 -51240 85400 -51230
rect 85310 -51330 85320 -51240
rect 85390 -51330 85400 -51240
rect 85310 -51600 85400 -51330
rect 81630 -51790 81640 -51680
rect 81760 -51790 81770 -51680
rect 81630 -51800 81770 -51790
rect 82280 -51680 82450 -51670
rect 82280 -51790 82290 -51680
rect 82440 -51790 82450 -51680
rect 79400 -51900 79690 -51890
rect 79400 -52140 79410 -51900
rect 79680 -52140 79690 -51900
rect 79400 -52150 79690 -52140
rect 79040 -52910 79070 -52840
rect 79140 -52910 79170 -52840
rect 79040 -52930 79170 -52910
rect 78770 -52940 78930 -52930
rect 78230 -53630 78240 -53570
rect 78300 -53630 78310 -53570
rect 78230 -53640 78310 -53630
rect 78630 -52990 78760 -52980
rect 78630 -53130 78640 -52990
rect 78750 -53130 78760 -52990
rect 78630 -53550 78760 -53130
rect 78630 -53640 78640 -53550
rect 78740 -53640 78760 -53550
rect 78630 -53650 78760 -53640
rect 78800 -53590 78880 -52940
rect 79400 -53160 79690 -53150
rect 79400 -53400 79410 -53160
rect 79680 -53400 79690 -53160
rect 78800 -53650 78810 -53590
rect 78870 -53650 78880 -53590
rect 78800 -53660 78880 -53650
rect 79060 -53420 79210 -53400
rect 79400 -53410 79690 -53400
rect 79060 -53720 79080 -53420
rect 79190 -53720 79210 -53420
rect 82280 -53440 82450 -51790
rect 83020 -51680 83110 -51670
rect 83020 -51790 83030 -51680
rect 83100 -51790 83110 -51680
rect 83020 -51800 83110 -51790
rect 85310 -51790 85320 -51600
rect 85390 -51790 85400 -51600
rect 85580 -51240 86490 -51230
rect 85580 -51330 85590 -51240
rect 86480 -51330 86490 -51240
rect 85580 -51660 86490 -51330
rect 87030 -51240 87930 -51230
rect 87030 -51330 87040 -51240
rect 87920 -51330 87930 -51240
rect 85580 -51740 85590 -51660
rect 86480 -51740 86490 -51660
rect 85580 -51750 86490 -51740
rect 86790 -51580 86880 -51570
rect 85310 -51800 85400 -51790
rect 86790 -51790 86800 -51580
rect 86870 -51790 86880 -51580
rect 87030 -51660 87930 -51330
rect 88500 -51240 89400 -51230
rect 88500 -51330 88510 -51240
rect 89390 -51330 89400 -51240
rect 87030 -51740 87040 -51660
rect 87920 -51740 87930 -51660
rect 87030 -51750 87930 -51740
rect 88260 -51590 88350 -51580
rect 86790 -52020 86880 -51790
rect 86790 -52100 86800 -52020
rect 86870 -52100 86880 -52020
rect 86790 -52110 86880 -52100
rect 88260 -51790 88270 -51590
rect 88340 -51790 88350 -51590
rect 88500 -51670 89400 -51330
rect 89970 -51240 90770 -51230
rect 89970 -51330 89980 -51240
rect 90760 -51330 90770 -51240
rect 88500 -51740 88510 -51670
rect 89390 -51740 89400 -51670
rect 88500 -51750 89400 -51740
rect 89740 -51590 89820 -51580
rect 88260 -52020 88350 -51790
rect 88260 -52100 88270 -52020
rect 88340 -52100 88350 -52020
rect 88260 -52110 88350 -52100
rect 89810 -51800 89820 -51590
rect 89970 -51669 90770 -51330
rect 89970 -51741 89982 -51669
rect 90762 -51741 90770 -51669
rect 89970 -51751 90770 -51741
rect 91200 -51590 91290 -51580
rect 89740 -52020 89820 -51800
rect 89740 -52100 89750 -52020
rect 89810 -52100 89820 -52020
rect 89740 -52110 89820 -52100
rect 91200 -51800 91210 -51590
rect 91280 -51800 91290 -51590
rect 91200 -52020 91290 -51800
rect 91200 -52100 91210 -52020
rect 91280 -52100 91290 -52020
rect 91200 -52110 91290 -52100
rect 91750 -51870 92160 -51840
rect 82790 -52230 91440 -52200
rect 82790 -52800 82820 -52230
rect 91410 -52800 91440 -52230
rect 91750 -52250 91780 -51870
rect 92130 -52250 92160 -51870
rect 91750 -52280 92160 -52250
rect 82790 -52830 91440 -52800
rect 79060 -53740 79210 -53720
rect 79980 -53470 80390 -53440
rect 79980 -53850 80010 -53470
rect 80360 -53850 80390 -53470
rect 79980 -53880 80390 -53850
rect 82110 -53470 82780 -53440
rect 82110 -53850 82140 -53470
rect 82750 -53850 82780 -53470
rect 82110 -53880 82780 -53850
rect 78060 -53990 78070 -53930
rect 78140 -53990 78150 -53930
rect 78060 -54000 78150 -53990
rect 69900 -86200 70000 -85800
rect 70300 -86200 70400 -85800
rect 69900 -86300 70400 -86200
rect 55400 -86600 55500 -86300
rect 56100 -86600 56200 -86300
rect 55400 -86700 56200 -86600
rect 37100 -86800 37800 -86700
<< via2 >>
rect 38000 1400 41400 2800
rect 43000 1000 46400 2400
rect 37900 -3600 41500 -400
rect 43000 -1400 46400 0
rect 56880 -40 59080 1020
rect 51500 -1000 52500 -800
rect 47700 -1700 48000 -1300
rect 36400 -5800 37000 -5000
rect 21000 -7400 22000 -6600
rect 20804 -11629 20878 -7875
rect 24700 -9400 25700 -8700
rect 20800 -12092 20880 -12002
rect 20580 -13042 20640 -12352
rect 20801 -13041 20861 -12351
rect 27200 -13000 34400 -10600
rect 20570 -13392 20670 -13312
rect 15000 -31200 19400 -26400
rect 26600 -30400 35200 -26400
rect 47640 -7200 48080 -6780
rect 46700 -9400 47800 -8700
rect 37600 -11100 38100 -10700
rect 47700 -12640 48080 -12220
rect 38500 -16600 39000 -16000
rect 47640 -18100 48080 -17620
rect 39500 -22000 40000 -21400
rect 47680 -23440 48080 -23020
rect 40400 -27400 41000 -26800
rect 15000 -49000 24000 -38000
rect 47800 -28840 48080 -28460
rect 41500 -32800 42100 -32200
rect 47760 -34200 48080 -33860
rect 42500 -38200 43100 -37600
rect 47760 -39640 48080 -39220
rect 43200 -43300 44300 -43100
rect 43200 -43800 44300 -43300
rect 15200 -64800 19600 -60000
rect 25000 -64800 35400 -58800
rect 43800 -49000 44300 -48400
rect 47820 -45060 48080 -44640
rect 42900 -54400 43400 -53800
rect 47740 -50480 48080 -49980
rect 42000 -59800 42500 -59200
rect 47820 -55820 48080 -55460
rect 41100 -65200 41600 -64600
rect 47680 -61300 48080 -60760
rect 40200 -70600 40700 -70000
rect 47860 -66660 48080 -66220
rect 39300 -76000 39800 -75400
rect 47720 -72060 48080 -71600
rect 38300 -81400 38800 -80800
rect 47780 -77500 48080 -76940
rect 47800 -82860 48080 -82380
rect 55400 -1000 55700 -600
rect 53400 -1600 53700 -1400
rect 53520 -1968 53640 -1858
rect 55960 -1888 56040 -1738
rect 55280 -1928 55400 -1918
rect 55280 -1998 55290 -1928
rect 55290 -1998 55390 -1928
rect 55390 -1998 55400 -1928
rect 55280 -2008 55400 -1998
rect 56506 -1830 57016 -1580
rect 58966 -1630 59126 -1470
rect 59336 -1650 59416 -1510
rect 60046 -1640 60126 -1520
rect 58996 -1840 59106 -1730
rect 59516 -1840 59616 -1740
rect 61056 -1850 61126 -1720
rect 53050 -3908 53250 -2158
rect 55880 -2098 55970 -2018
rect 55230 -2428 55320 -2258
rect 55600 -2398 55710 -2268
rect 58486 -2290 58816 -1930
rect 59286 -2190 59346 -2130
rect 59546 -2150 59606 -2090
rect 59006 -2260 59016 -2200
rect 59016 -2260 59066 -2200
rect 59546 -2270 59606 -2210
rect 59866 -2230 59966 -2140
rect 60446 -2220 60526 -2120
rect 60046 -2340 60126 -2320
rect 60046 -2400 60126 -2340
rect 59076 -2510 59166 -2440
rect 60556 -2490 60626 -2410
rect 59976 -2552 60316 -2500
rect 59976 -2560 60316 -2552
rect 56480 -2648 56550 -2588
rect 57098 -2704 57368 -2564
rect 59286 -2720 59366 -2630
rect 59576 -2730 59636 -2670
rect 61206 -2700 61346 -2520
rect 59286 -2930 59356 -2840
rect 59916 -2960 60006 -2780
rect 60306 -2890 60456 -2750
rect 61036 -2930 61126 -2820
rect 55020 -3128 55030 -3048
rect 55030 -3128 55110 -3048
rect 55110 -3128 55120 -3048
rect 55880 -3128 55970 -3038
rect 56480 -3128 56550 -3038
rect 57800 -3140 58240 -3020
rect 58556 -3080 58756 -3060
rect 58556 -3240 58576 -3080
rect 58576 -3240 58736 -3080
rect 58736 -3240 58756 -3080
rect 58556 -3260 58756 -3240
rect 59076 -3080 59166 -3010
rect 59316 -3090 59376 -3030
rect 59076 -3240 59166 -3170
rect 60096 -3240 60176 -3080
rect 61276 -3260 61356 -3050
rect 59266 -3410 59366 -3320
rect 56480 -3588 56550 -3528
rect 57098 -3614 57368 -3474
rect 59916 -3480 60006 -3290
rect 60476 -3370 60536 -3310
rect 59266 -3650 59366 -3560
rect 59516 -3520 59596 -3510
rect 59516 -3580 59596 -3520
rect 61336 -3560 61456 -3430
rect 55220 -3918 55310 -3748
rect 55410 -3928 55500 -3758
rect 59076 -3800 59166 -3740
rect 59316 -3780 59376 -3720
rect 59996 -3780 60106 -3720
rect 53510 -4248 53630 -4128
rect 55880 -4158 55970 -4078
rect 55620 -4278 55710 -4188
rect 55220 -4518 55320 -4418
rect 56020 -4408 56080 -4258
rect 59256 -4090 59366 -4030
rect 59546 -4000 59606 -3990
rect 59546 -4060 59606 -4000
rect 59016 -4160 59076 -4100
rect 59546 -4170 59606 -4110
rect 59806 -4120 59916 -4010
rect 60446 -4150 60526 -4030
rect 55320 -4868 55470 -4728
rect 56654 -4486 56998 -4268
rect 59016 -4510 59076 -4440
rect 59546 -4510 59606 -4440
rect 60266 -4530 60406 -4400
rect 58966 -4620 59146 -4600
rect 58966 -4760 58986 -4620
rect 58986 -4760 59126 -4620
rect 59126 -4760 59146 -4620
rect 58966 -4780 59146 -4760
rect 59996 -4700 60106 -4590
rect 59700 -5200 60400 -4900
rect 68100 -5200 68600 -4900
rect 55600 -5600 55900 -5300
rect 51500 -6500 52500 -6300
rect 55400 -6500 55700 -6200
rect 53520 -7120 53780 -6860
rect 53520 -7368 53640 -7258
rect 55960 -7288 56040 -7138
rect 55280 -7328 55400 -7318
rect 55280 -7398 55290 -7328
rect 55290 -7398 55390 -7328
rect 55390 -7398 55400 -7328
rect 55280 -7408 55400 -7398
rect 56506 -7230 57016 -6980
rect 58966 -7030 59126 -6870
rect 59336 -7050 59416 -6910
rect 60046 -7040 60126 -6920
rect 58996 -7240 59106 -7130
rect 59516 -7240 59616 -7140
rect 61056 -7250 61126 -7120
rect 53050 -9308 53250 -7558
rect 55880 -7498 55970 -7418
rect 55230 -7828 55320 -7658
rect 55600 -7798 55710 -7668
rect 58486 -7690 58816 -7330
rect 59286 -7590 59346 -7530
rect 59546 -7550 59606 -7490
rect 59006 -7660 59016 -7600
rect 59016 -7660 59066 -7600
rect 59546 -7670 59606 -7610
rect 59866 -7630 59966 -7540
rect 60446 -7620 60526 -7520
rect 60046 -7740 60126 -7720
rect 60046 -7800 60126 -7740
rect 59076 -7910 59166 -7840
rect 60556 -7890 60626 -7810
rect 59976 -7952 60316 -7900
rect 59976 -7960 60316 -7952
rect 56480 -8048 56550 -7988
rect 57098 -8104 57368 -7964
rect 59286 -8120 59366 -8030
rect 59576 -8130 59636 -8070
rect 61206 -8100 61346 -7920
rect 59286 -8330 59356 -8240
rect 59916 -8360 60006 -8180
rect 60306 -8290 60456 -8150
rect 61036 -8330 61126 -8220
rect 55020 -8528 55030 -8448
rect 55030 -8528 55110 -8448
rect 55110 -8528 55120 -8448
rect 55880 -8528 55970 -8438
rect 56480 -8528 56550 -8438
rect 57800 -8540 58240 -8420
rect 58556 -8480 58756 -8460
rect 58556 -8640 58576 -8480
rect 58576 -8640 58736 -8480
rect 58736 -8640 58756 -8480
rect 58556 -8660 58756 -8640
rect 59076 -8480 59166 -8410
rect 59316 -8490 59376 -8430
rect 59076 -8640 59166 -8570
rect 60096 -8640 60176 -8480
rect 61276 -8660 61356 -8450
rect 59266 -8810 59366 -8720
rect 56480 -8988 56550 -8928
rect 57098 -9014 57368 -8874
rect 59916 -8880 60006 -8690
rect 60476 -8770 60536 -8710
rect 59266 -9050 59366 -8960
rect 59516 -8920 59596 -8910
rect 59516 -8980 59596 -8920
rect 61336 -8960 61456 -8830
rect 55220 -9318 55310 -9148
rect 55410 -9328 55500 -9158
rect 59076 -9200 59166 -9140
rect 59316 -9180 59376 -9120
rect 59996 -9180 60106 -9120
rect 53510 -9648 53630 -9528
rect 55880 -9558 55970 -9478
rect 55620 -9678 55710 -9588
rect 55220 -9918 55320 -9818
rect 56020 -9808 56080 -9658
rect 59256 -9490 59366 -9430
rect 59546 -9400 59606 -9390
rect 59546 -9460 59606 -9400
rect 59016 -9560 59076 -9500
rect 59546 -9570 59606 -9510
rect 59806 -9520 59916 -9410
rect 60446 -9550 60526 -9430
rect 55320 -10268 55470 -10128
rect 56654 -9886 56998 -9668
rect 59016 -9910 59076 -9840
rect 59546 -9910 59606 -9840
rect 60266 -9930 60406 -9800
rect 58966 -10020 59146 -10000
rect 58966 -10160 58986 -10020
rect 58986 -10160 59126 -10020
rect 59126 -10160 59146 -10020
rect 58966 -10180 59146 -10160
rect 59996 -10100 60106 -9990
rect 55500 -11100 56000 -10700
rect 59700 -10700 60400 -10300
rect 66900 -10700 67400 -10300
rect 51500 -11900 52500 -11700
rect 55380 -11980 55740 -11660
rect 53480 -12540 53780 -12340
rect 53520 -12768 53640 -12658
rect 55960 -12688 56040 -12538
rect 55280 -12728 55400 -12718
rect 55280 -12798 55290 -12728
rect 55290 -12798 55390 -12728
rect 55390 -12798 55400 -12728
rect 55280 -12808 55400 -12798
rect 56506 -12630 57016 -12380
rect 58966 -12430 59126 -12270
rect 59336 -12450 59416 -12310
rect 60046 -12440 60126 -12320
rect 58996 -12640 59106 -12530
rect 59516 -12640 59616 -12540
rect 61056 -12650 61126 -12520
rect 53050 -14708 53250 -12958
rect 55880 -12898 55970 -12818
rect 55230 -13228 55320 -13058
rect 55600 -13198 55710 -13068
rect 58486 -13090 58816 -12730
rect 59286 -12990 59346 -12930
rect 59546 -12950 59606 -12890
rect 59006 -13060 59016 -13000
rect 59016 -13060 59066 -13000
rect 59546 -13070 59606 -13010
rect 59866 -13030 59966 -12940
rect 60446 -13020 60526 -12920
rect 60046 -13140 60126 -13120
rect 60046 -13200 60126 -13140
rect 59076 -13310 59166 -13240
rect 60556 -13290 60626 -13210
rect 59976 -13352 60316 -13300
rect 59976 -13360 60316 -13352
rect 56480 -13448 56550 -13388
rect 57098 -13504 57368 -13364
rect 59286 -13520 59366 -13430
rect 59576 -13530 59636 -13470
rect 61206 -13500 61346 -13320
rect 59286 -13730 59356 -13640
rect 59916 -13760 60006 -13580
rect 60306 -13690 60456 -13550
rect 61036 -13730 61126 -13620
rect 55020 -13928 55030 -13848
rect 55030 -13928 55110 -13848
rect 55110 -13928 55120 -13848
rect 55880 -13928 55970 -13838
rect 56480 -13928 56550 -13838
rect 57800 -13940 58240 -13820
rect 58556 -13880 58756 -13860
rect 58556 -14040 58576 -13880
rect 58576 -14040 58736 -13880
rect 58736 -14040 58756 -13880
rect 58556 -14060 58756 -14040
rect 59076 -13880 59166 -13810
rect 59316 -13890 59376 -13830
rect 59076 -14040 59166 -13970
rect 60096 -14040 60176 -13880
rect 61276 -14060 61356 -13850
rect 59266 -14210 59366 -14120
rect 56480 -14388 56550 -14328
rect 57098 -14414 57368 -14274
rect 59916 -14280 60006 -14090
rect 60476 -14170 60536 -14110
rect 59266 -14450 59366 -14360
rect 59516 -14320 59596 -14310
rect 59516 -14380 59596 -14320
rect 61336 -14360 61456 -14230
rect 55220 -14718 55310 -14548
rect 55410 -14728 55500 -14558
rect 59076 -14600 59166 -14540
rect 59316 -14580 59376 -14520
rect 59996 -14580 60106 -14520
rect 53510 -15048 53630 -14928
rect 55880 -14958 55970 -14878
rect 55620 -15078 55710 -14988
rect 55220 -15318 55320 -15218
rect 56020 -15208 56080 -15058
rect 59256 -14890 59366 -14830
rect 59546 -14800 59606 -14790
rect 59546 -14860 59606 -14800
rect 59016 -14960 59076 -14900
rect 59546 -14970 59606 -14910
rect 59806 -14920 59916 -14810
rect 60446 -14950 60526 -14830
rect 55320 -15668 55470 -15528
rect 56654 -15286 56998 -15068
rect 59016 -15310 59076 -15240
rect 59546 -15310 59606 -15240
rect 60266 -15330 60406 -15200
rect 58966 -15420 59146 -15400
rect 58966 -15560 58986 -15420
rect 58986 -15560 59126 -15420
rect 59126 -15560 59146 -15420
rect 58966 -15580 59146 -15560
rect 59996 -15500 60106 -15390
rect 59800 -15900 60300 -15600
rect 65900 -15900 66400 -15600
rect 55500 -16500 56000 -16100
rect 51500 -17300 52500 -17100
rect 55400 -17400 55700 -17100
rect 53500 -17940 53780 -17740
rect 53520 -18168 53640 -18058
rect 55960 -18088 56040 -17938
rect 55280 -18128 55400 -18118
rect 55280 -18198 55290 -18128
rect 55290 -18198 55390 -18128
rect 55390 -18198 55400 -18128
rect 55280 -18208 55400 -18198
rect 56506 -18030 57016 -17780
rect 58966 -17830 59126 -17670
rect 59336 -17850 59416 -17710
rect 60046 -17840 60126 -17720
rect 58996 -18040 59106 -17930
rect 59516 -18040 59616 -17940
rect 61056 -18050 61126 -17920
rect 53050 -20108 53250 -18358
rect 55880 -18298 55970 -18218
rect 55230 -18628 55320 -18458
rect 55600 -18598 55710 -18468
rect 58486 -18490 58816 -18130
rect 59286 -18390 59346 -18330
rect 59546 -18350 59606 -18290
rect 59006 -18460 59016 -18400
rect 59016 -18460 59066 -18400
rect 59546 -18470 59606 -18410
rect 59866 -18430 59966 -18340
rect 60446 -18420 60526 -18320
rect 60046 -18540 60126 -18520
rect 60046 -18600 60126 -18540
rect 59076 -18710 59166 -18640
rect 60556 -18690 60626 -18610
rect 59976 -18752 60316 -18700
rect 59976 -18760 60316 -18752
rect 56480 -18848 56550 -18788
rect 57098 -18904 57368 -18764
rect 59286 -18920 59366 -18830
rect 59576 -18930 59636 -18870
rect 61206 -18900 61346 -18720
rect 59286 -19130 59356 -19040
rect 59916 -19160 60006 -18980
rect 60306 -19090 60456 -18950
rect 61036 -19130 61126 -19020
rect 55020 -19328 55030 -19248
rect 55030 -19328 55110 -19248
rect 55110 -19328 55120 -19248
rect 55880 -19328 55970 -19238
rect 56480 -19328 56550 -19238
rect 57800 -19340 58240 -19220
rect 58556 -19280 58756 -19260
rect 58556 -19440 58576 -19280
rect 58576 -19440 58736 -19280
rect 58736 -19440 58756 -19280
rect 58556 -19460 58756 -19440
rect 59076 -19280 59166 -19210
rect 59316 -19290 59376 -19230
rect 59076 -19440 59166 -19370
rect 60096 -19440 60176 -19280
rect 61276 -19460 61356 -19250
rect 59266 -19610 59366 -19520
rect 56480 -19788 56550 -19728
rect 57098 -19814 57368 -19674
rect 59916 -19680 60006 -19490
rect 60476 -19570 60536 -19510
rect 59266 -19850 59366 -19760
rect 59516 -19720 59596 -19710
rect 59516 -19780 59596 -19720
rect 61336 -19760 61456 -19630
rect 55220 -20118 55310 -19948
rect 55410 -20128 55500 -19958
rect 59076 -20000 59166 -19940
rect 59316 -19980 59376 -19920
rect 59996 -19980 60106 -19920
rect 53510 -20448 53630 -20328
rect 55880 -20358 55970 -20278
rect 55620 -20478 55710 -20388
rect 55220 -20718 55320 -20618
rect 56020 -20608 56080 -20458
rect 59256 -20290 59366 -20230
rect 59546 -20200 59606 -20190
rect 59546 -20260 59606 -20200
rect 59016 -20360 59076 -20300
rect 59546 -20370 59606 -20310
rect 59806 -20320 59916 -20210
rect 60446 -20350 60526 -20230
rect 55320 -21068 55470 -20928
rect 56654 -20686 56998 -20468
rect 59016 -20710 59076 -20640
rect 59546 -20710 59606 -20640
rect 60266 -20730 60406 -20600
rect 58966 -20820 59146 -20800
rect 58966 -20960 58986 -20820
rect 58986 -20960 59126 -20820
rect 59126 -20960 59146 -20820
rect 58966 -20980 59146 -20960
rect 59996 -20900 60106 -20790
rect 59800 -21300 60300 -21000
rect 64900 -21300 65400 -21000
rect 55500 -21900 56100 -21500
rect 51500 -22700 52500 -22500
rect 55440 -22760 55720 -22480
rect 53480 -23340 53780 -23140
rect 53520 -23568 53640 -23458
rect 55960 -23488 56040 -23338
rect 55280 -23528 55400 -23518
rect 55280 -23598 55290 -23528
rect 55290 -23598 55390 -23528
rect 55390 -23598 55400 -23528
rect 55280 -23608 55400 -23598
rect 56506 -23430 57016 -23180
rect 58966 -23230 59126 -23070
rect 59336 -23250 59416 -23110
rect 60046 -23240 60126 -23120
rect 58996 -23440 59106 -23330
rect 59516 -23440 59616 -23340
rect 61056 -23450 61126 -23320
rect 53050 -25508 53250 -23758
rect 55880 -23698 55970 -23618
rect 55230 -24028 55320 -23858
rect 55600 -23998 55710 -23868
rect 58486 -23890 58816 -23530
rect 59286 -23790 59346 -23730
rect 59546 -23750 59606 -23690
rect 59006 -23860 59016 -23800
rect 59016 -23860 59066 -23800
rect 59546 -23870 59606 -23810
rect 59866 -23830 59966 -23740
rect 60446 -23820 60526 -23720
rect 60046 -23940 60126 -23920
rect 60046 -24000 60126 -23940
rect 59076 -24110 59166 -24040
rect 60556 -24090 60626 -24010
rect 59976 -24152 60316 -24100
rect 59976 -24160 60316 -24152
rect 56480 -24248 56550 -24188
rect 57098 -24304 57368 -24164
rect 59286 -24320 59366 -24230
rect 59576 -24330 59636 -24270
rect 61206 -24300 61346 -24120
rect 59286 -24530 59356 -24440
rect 59916 -24560 60006 -24380
rect 60306 -24490 60456 -24350
rect 61036 -24530 61126 -24420
rect 55020 -24728 55030 -24648
rect 55030 -24728 55110 -24648
rect 55110 -24728 55120 -24648
rect 55880 -24728 55970 -24638
rect 56480 -24728 56550 -24638
rect 57800 -24740 58240 -24620
rect 58556 -24680 58756 -24660
rect 58556 -24840 58576 -24680
rect 58576 -24840 58736 -24680
rect 58736 -24840 58756 -24680
rect 58556 -24860 58756 -24840
rect 59076 -24680 59166 -24610
rect 59316 -24690 59376 -24630
rect 59076 -24840 59166 -24770
rect 60096 -24840 60176 -24680
rect 61276 -24860 61356 -24650
rect 59266 -25010 59366 -24920
rect 56480 -25188 56550 -25128
rect 57098 -25214 57368 -25074
rect 59916 -25080 60006 -24890
rect 60476 -24970 60536 -24910
rect 59266 -25250 59366 -25160
rect 59516 -25120 59596 -25110
rect 59516 -25180 59596 -25120
rect 61336 -25160 61456 -25030
rect 55220 -25518 55310 -25348
rect 55410 -25528 55500 -25358
rect 59076 -25400 59166 -25340
rect 59316 -25380 59376 -25320
rect 59996 -25380 60106 -25320
rect 53510 -25848 53630 -25728
rect 55880 -25758 55970 -25678
rect 55620 -25878 55710 -25788
rect 55220 -26118 55320 -26018
rect 56020 -26008 56080 -25858
rect 59256 -25690 59366 -25630
rect 59546 -25600 59606 -25590
rect 59546 -25660 59606 -25600
rect 59016 -25760 59076 -25700
rect 59546 -25770 59606 -25710
rect 59806 -25720 59916 -25610
rect 60446 -25750 60526 -25630
rect 55320 -26468 55470 -26328
rect 56654 -26086 56998 -25868
rect 59016 -26110 59076 -26040
rect 59546 -26110 59606 -26040
rect 60266 -26130 60406 -26000
rect 58966 -26220 59146 -26200
rect 58966 -26360 58986 -26220
rect 58986 -26360 59126 -26220
rect 59126 -26360 59146 -26220
rect 58966 -26380 59146 -26360
rect 59996 -26300 60106 -26190
rect 59700 -26800 60400 -26400
rect 63700 -26800 64100 -26400
rect 55500 -27300 56100 -26900
rect 51500 -28100 52500 -27900
rect 55460 -28160 55720 -27880
rect 53480 -28740 53780 -28540
rect 53520 -28968 53640 -28858
rect 55960 -28888 56040 -28738
rect 55280 -28928 55400 -28918
rect 55280 -28998 55290 -28928
rect 55290 -28998 55390 -28928
rect 55390 -28998 55400 -28928
rect 55280 -29008 55400 -28998
rect 56506 -28830 57016 -28580
rect 58966 -28630 59126 -28470
rect 59336 -28650 59416 -28510
rect 60046 -28640 60126 -28520
rect 58996 -28840 59106 -28730
rect 59516 -28840 59616 -28740
rect 61056 -28850 61126 -28720
rect 53050 -30908 53250 -29158
rect 55880 -29098 55970 -29018
rect 55230 -29428 55320 -29258
rect 55600 -29398 55710 -29268
rect 58486 -29290 58816 -28930
rect 59286 -29190 59346 -29130
rect 59546 -29150 59606 -29090
rect 59006 -29260 59016 -29200
rect 59016 -29260 59066 -29200
rect 59546 -29270 59606 -29210
rect 59866 -29230 59966 -29140
rect 60446 -29220 60526 -29120
rect 60046 -29340 60126 -29320
rect 60046 -29400 60126 -29340
rect 59076 -29510 59166 -29440
rect 60556 -29490 60626 -29410
rect 59976 -29552 60316 -29500
rect 59976 -29560 60316 -29552
rect 56480 -29648 56550 -29588
rect 57098 -29704 57368 -29564
rect 59286 -29720 59366 -29630
rect 59576 -29730 59636 -29670
rect 61206 -29700 61346 -29520
rect 59286 -29930 59356 -29840
rect 59916 -29960 60006 -29780
rect 60306 -29890 60456 -29750
rect 61036 -29930 61126 -29820
rect 55020 -30128 55030 -30048
rect 55030 -30128 55110 -30048
rect 55110 -30128 55120 -30048
rect 55880 -30128 55970 -30038
rect 56480 -30128 56550 -30038
rect 57800 -30140 58240 -30020
rect 58556 -30080 58756 -30060
rect 58556 -30240 58576 -30080
rect 58576 -30240 58736 -30080
rect 58736 -30240 58756 -30080
rect 58556 -30260 58756 -30240
rect 59076 -30080 59166 -30010
rect 59316 -30090 59376 -30030
rect 59076 -30240 59166 -30170
rect 60096 -30240 60176 -30080
rect 61276 -30260 61356 -30050
rect 59266 -30410 59366 -30320
rect 56480 -30588 56550 -30528
rect 57098 -30614 57368 -30474
rect 59916 -30480 60006 -30290
rect 60476 -30370 60536 -30310
rect 59266 -30650 59366 -30560
rect 59516 -30520 59596 -30510
rect 59516 -30580 59596 -30520
rect 61336 -30560 61456 -30430
rect 55220 -30918 55310 -30748
rect 55410 -30928 55500 -30758
rect 59076 -30800 59166 -30740
rect 59316 -30780 59376 -30720
rect 59996 -30780 60106 -30720
rect 53510 -31248 53630 -31128
rect 55880 -31158 55970 -31078
rect 55620 -31278 55710 -31188
rect 55220 -31518 55320 -31418
rect 56020 -31408 56080 -31258
rect 59256 -31090 59366 -31030
rect 59546 -31000 59606 -30990
rect 59546 -31060 59606 -31000
rect 59016 -31160 59076 -31100
rect 59546 -31170 59606 -31110
rect 59806 -31120 59916 -31010
rect 60446 -31150 60526 -31030
rect 55320 -31868 55470 -31728
rect 56654 -31486 56998 -31268
rect 59016 -31510 59076 -31440
rect 59546 -31510 59606 -31440
rect 60266 -31530 60406 -31400
rect 58966 -31620 59146 -31600
rect 58966 -31760 58986 -31620
rect 58986 -31760 59126 -31620
rect 59126 -31760 59146 -31620
rect 58966 -31780 59146 -31760
rect 59996 -31700 60106 -31590
rect 59800 -32100 60300 -31800
rect 62900 -32100 63300 -31800
rect 55500 -32700 56100 -32300
rect 51500 -33500 52500 -33300
rect 55460 -33560 55720 -33280
rect 53480 -34140 53780 -33940
rect 53520 -34368 53640 -34258
rect 55960 -34288 56040 -34138
rect 55280 -34328 55400 -34318
rect 55280 -34398 55290 -34328
rect 55290 -34398 55390 -34328
rect 55390 -34398 55400 -34328
rect 55280 -34408 55400 -34398
rect 56506 -34230 57016 -33980
rect 58966 -34030 59126 -33870
rect 59336 -34050 59416 -33910
rect 60046 -34040 60126 -33920
rect 58996 -34240 59106 -34130
rect 59516 -34240 59616 -34140
rect 61056 -34250 61126 -34120
rect 53050 -36308 53250 -34558
rect 55880 -34498 55970 -34418
rect 55230 -34828 55320 -34658
rect 55600 -34798 55710 -34668
rect 58486 -34690 58816 -34330
rect 59286 -34590 59346 -34530
rect 59546 -34550 59606 -34490
rect 59006 -34660 59016 -34600
rect 59016 -34660 59066 -34600
rect 59546 -34670 59606 -34610
rect 59866 -34630 59966 -34540
rect 60446 -34620 60526 -34520
rect 60046 -34740 60126 -34720
rect 60046 -34800 60126 -34740
rect 59076 -34910 59166 -34840
rect 60556 -34890 60626 -34810
rect 59976 -34952 60316 -34900
rect 59976 -34960 60316 -34952
rect 56480 -35048 56550 -34988
rect 57098 -35104 57368 -34964
rect 59286 -35120 59366 -35030
rect 59576 -35130 59636 -35070
rect 61206 -35100 61346 -34920
rect 59286 -35330 59356 -35240
rect 59916 -35360 60006 -35180
rect 60306 -35290 60456 -35150
rect 61036 -35330 61126 -35220
rect 55020 -35528 55030 -35448
rect 55030 -35528 55110 -35448
rect 55110 -35528 55120 -35448
rect 55880 -35528 55970 -35438
rect 56480 -35528 56550 -35438
rect 57800 -35540 58240 -35420
rect 58556 -35480 58756 -35460
rect 58556 -35640 58576 -35480
rect 58576 -35640 58736 -35480
rect 58736 -35640 58756 -35480
rect 58556 -35660 58756 -35640
rect 59076 -35480 59166 -35410
rect 59316 -35490 59376 -35430
rect 59076 -35640 59166 -35570
rect 60096 -35640 60176 -35480
rect 61276 -35660 61356 -35450
rect 59266 -35810 59366 -35720
rect 56480 -35988 56550 -35928
rect 57098 -36014 57368 -35874
rect 59916 -35880 60006 -35690
rect 60476 -35770 60536 -35710
rect 59266 -36050 59366 -35960
rect 59516 -35920 59596 -35910
rect 59516 -35980 59596 -35920
rect 61336 -35960 61456 -35830
rect 55220 -36318 55310 -36148
rect 55410 -36328 55500 -36158
rect 59076 -36200 59166 -36140
rect 59316 -36180 59376 -36120
rect 59996 -36180 60106 -36120
rect 53510 -36648 53630 -36528
rect 55880 -36558 55970 -36478
rect 55620 -36678 55710 -36588
rect 55220 -36918 55320 -36818
rect 56020 -36808 56080 -36658
rect 59256 -36490 59366 -36430
rect 59546 -36400 59606 -36390
rect 59546 -36460 59606 -36400
rect 59016 -36560 59076 -36500
rect 59546 -36570 59606 -36510
rect 59806 -36520 59916 -36410
rect 60446 -36550 60526 -36430
rect 55320 -37268 55470 -37128
rect 56654 -36886 56998 -36668
rect 59016 -36910 59076 -36840
rect 59546 -36910 59606 -36840
rect 60266 -36930 60406 -36800
rect 58966 -37020 59146 -37000
rect 58966 -37160 58986 -37020
rect 58986 -37160 59126 -37020
rect 59126 -37160 59146 -37020
rect 58966 -37180 59146 -37160
rect 59996 -37100 60106 -36990
rect 59900 -37400 60200 -37200
rect 55400 -38100 56100 -37700
rect 62000 -37700 62500 -37100
rect 51500 -38900 52500 -38700
rect 55460 -38960 55720 -38680
rect 53480 -39540 53780 -39340
rect 53520 -39768 53640 -39658
rect 55960 -39688 56040 -39538
rect 55280 -39728 55400 -39718
rect 55280 -39798 55290 -39728
rect 55290 -39798 55390 -39728
rect 55390 -39798 55400 -39728
rect 55280 -39808 55400 -39798
rect 56506 -39630 57016 -39380
rect 58966 -39430 59126 -39270
rect 59336 -39450 59416 -39310
rect 60046 -39440 60126 -39320
rect 58996 -39640 59106 -39530
rect 59516 -39640 59616 -39540
rect 61056 -39650 61126 -39520
rect 53050 -41708 53250 -39958
rect 55880 -39898 55970 -39818
rect 55230 -40228 55320 -40058
rect 55600 -40198 55710 -40068
rect 58486 -40090 58816 -39730
rect 59286 -39990 59346 -39930
rect 59546 -39950 59606 -39890
rect 59006 -40060 59016 -40000
rect 59016 -40060 59066 -40000
rect 59546 -40070 59606 -40010
rect 59866 -40030 59966 -39940
rect 60446 -40020 60526 -39920
rect 60046 -40140 60126 -40120
rect 60046 -40200 60126 -40140
rect 59076 -40310 59166 -40240
rect 60556 -40290 60626 -40210
rect 59976 -40352 60316 -40300
rect 59976 -40360 60316 -40352
rect 56480 -40448 56550 -40388
rect 57098 -40504 57368 -40364
rect 59286 -40520 59366 -40430
rect 59576 -40530 59636 -40470
rect 61206 -40500 61346 -40320
rect 59286 -40730 59356 -40640
rect 59916 -40760 60006 -40580
rect 60306 -40690 60456 -40550
rect 61036 -40730 61126 -40620
rect 55020 -40928 55030 -40848
rect 55030 -40928 55110 -40848
rect 55110 -40928 55120 -40848
rect 55880 -40928 55970 -40838
rect 56480 -40928 56550 -40838
rect 57800 -40940 58240 -40820
rect 58556 -40880 58756 -40860
rect 58556 -41040 58576 -40880
rect 58576 -41040 58736 -40880
rect 58736 -41040 58756 -40880
rect 58556 -41060 58756 -41040
rect 59076 -40880 59166 -40810
rect 59316 -40890 59376 -40830
rect 59076 -41040 59166 -40970
rect 60096 -41040 60176 -40880
rect 61276 -41060 61356 -40850
rect 59266 -41210 59366 -41120
rect 56480 -41388 56550 -41328
rect 57098 -41414 57368 -41274
rect 59916 -41280 60006 -41090
rect 60476 -41170 60536 -41110
rect 59266 -41450 59366 -41360
rect 59516 -41320 59596 -41310
rect 59516 -41380 59596 -41320
rect 61336 -41360 61456 -41230
rect 72000 -35500 74000 -34100
rect 75390 -38270 75550 -38150
rect 78770 -38270 78890 -38150
rect 72820 -38920 73040 -38740
rect 68100 -39200 68600 -39000
rect 72820 -39250 73040 -39070
rect 66900 -39600 67400 -39400
rect 72820 -39740 73040 -39560
rect 65900 -40000 66400 -39800
rect 72820 -40020 73040 -39840
rect 64900 -40400 65400 -40200
rect 72820 -40480 73040 -40300
rect 63640 -40800 64160 -40660
rect 72820 -40840 73040 -40660
rect 62900 -41300 63300 -41000
rect 72820 -41240 73040 -41060
rect 55220 -41718 55310 -41548
rect 55410 -41728 55500 -41558
rect 59076 -41600 59166 -41540
rect 59316 -41580 59376 -41520
rect 59996 -41580 60106 -41520
rect 53510 -42048 53630 -41928
rect 55880 -41958 55970 -41878
rect 55620 -42078 55710 -41988
rect 55220 -42318 55320 -42218
rect 56020 -42208 56080 -42058
rect 59256 -41890 59366 -41830
rect 59546 -41800 59606 -41790
rect 59546 -41860 59606 -41800
rect 59016 -41960 59076 -41900
rect 59546 -41970 59606 -41910
rect 62000 -41700 62500 -41500
rect 72820 -41690 73040 -41510
rect 59806 -41920 59916 -41810
rect 60446 -41950 60526 -41830
rect 55320 -42668 55470 -42528
rect 56654 -42286 56998 -42068
rect 72820 -42060 73040 -41880
rect 73220 -42040 73340 -41900
rect 73470 -41670 73590 -41530
rect 59016 -42310 59076 -42240
rect 59546 -42310 59606 -42240
rect 60266 -42330 60406 -42200
rect 58966 -42420 59146 -42400
rect 58966 -42560 58986 -42420
rect 58986 -42560 59126 -42420
rect 59126 -42560 59146 -42420
rect 58966 -42580 59146 -42560
rect 59996 -42500 60106 -42390
rect 55500 -43500 56100 -43100
rect 59800 -43400 60400 -42800
rect 51500 -44300 52500 -44100
rect 55500 -44360 55720 -44080
rect 73720 -41220 73840 -41090
rect 73720 -43000 73840 -42930
rect 73970 -39490 74090 -39430
rect 74220 -40450 74340 -40390
rect 74477 -38674 74594 -38570
rect 74470 -40000 74590 -39860
rect 74470 -40180 74590 -40110
rect 73970 -40820 74090 -40680
rect 73470 -44440 73590 -44380
rect 73970 -43830 74090 -43760
rect 53480 -44940 53780 -44740
rect 53520 -45168 53640 -45058
rect 55960 -45088 56040 -44938
rect 55280 -45128 55400 -45118
rect 55280 -45198 55290 -45128
rect 55290 -45198 55390 -45128
rect 55390 -45198 55400 -45128
rect 55280 -45208 55400 -45198
rect 56506 -45030 57016 -44780
rect 58966 -44830 59126 -44670
rect 59336 -44850 59416 -44710
rect 60046 -44840 60126 -44720
rect 73970 -44800 74090 -44740
rect 74470 -41380 74590 -41320
rect 58996 -45040 59106 -44930
rect 59516 -45040 59616 -44940
rect 61056 -45050 61126 -44920
rect 53050 -47108 53250 -45358
rect 55880 -45298 55970 -45218
rect 55230 -45628 55320 -45458
rect 55600 -45598 55710 -45468
rect 58486 -45490 58816 -45130
rect 59286 -45390 59346 -45330
rect 59546 -45350 59606 -45290
rect 59006 -45460 59016 -45400
rect 59016 -45460 59066 -45400
rect 59546 -45470 59606 -45410
rect 59866 -45430 59966 -45340
rect 60446 -45420 60526 -45320
rect 74724 -38830 74841 -38752
rect 74720 -39720 74840 -39580
rect 74720 -41690 74840 -41630
rect 74970 -39220 75090 -39100
rect 74980 -39850 75080 -39780
rect 74970 -42330 75090 -42270
rect 75231 -38492 75322 -38427
rect 76648 -38505 76726 -38440
rect 75220 -39020 75340 -38920
rect 76102 -38661 76167 -38583
rect 76167 -38661 76180 -38583
rect 76375 -38804 76440 -38726
rect 75220 -40610 75340 -40540
rect 75220 -41240 75340 -41160
rect 75220 -41860 75340 -41770
rect 60046 -45540 60126 -45520
rect 60046 -45600 60126 -45540
rect 74470 -45560 74590 -45480
rect 75220 -42500 75340 -42410
rect 75220 -43250 75340 -43190
rect 75220 -43680 75340 -43620
rect 76920 -38530 77060 -38410
rect 76780 -38674 76791 -38630
rect 76791 -38674 76843 -38630
rect 76843 -38674 76860 -38630
rect 76780 -38700 76860 -38674
rect 78280 -38700 78350 -38630
rect 76210 -43130 76340 -43070
rect 77170 -39040 77430 -38790
rect 77230 -39500 77310 -39440
rect 76920 -39720 77060 -39570
rect 77170 -39850 77260 -39780
rect 84960 -38480 85400 -38050
rect 88150 -38820 88590 -38390
rect 82780 -39100 82890 -39010
rect 79080 -39510 79250 -39350
rect 80080 -39580 80430 -39270
rect 83370 -39080 83740 -39010
rect 84870 -39070 85240 -39000
rect 86330 -39070 86700 -39000
rect 78580 -39900 78640 -39840
rect 80080 -40060 80430 -39680
rect 84230 -39810 84310 -39700
rect 87460 -39070 87750 -39000
rect 85710 -39810 85790 -39700
rect 87180 -39810 87260 -39700
rect 88650 -39810 88730 -39700
rect 77410 -40180 77480 -40110
rect 77780 -40450 77840 -40390
rect 79410 -40390 79680 -40150
rect 83150 -40180 83510 -39830
rect 91780 -39960 92130 -39580
rect 77450 -40610 77520 -40540
rect 76920 -40960 77060 -40820
rect 77450 -41240 77530 -41160
rect 77780 -41380 77840 -41320
rect 77780 -41690 77840 -41630
rect 77490 -41860 77580 -41770
rect 76920 -42210 77060 -42060
rect 77780 -42330 77840 -42270
rect 77470 -42500 77560 -42410
rect 78670 -41180 78780 -41030
rect 79410 -41620 79680 -41380
rect 78160 -42470 78260 -42370
rect 79050 -42470 79150 -42360
rect 77470 -42990 77540 -42930
rect 77860 -43110 77920 -43050
rect 76920 -43450 77060 -43310
rect 77960 -43250 78020 -43190
rect 78860 -43210 78980 -42920
rect 77970 -43680 78030 -43620
rect 77430 -43830 77500 -43760
rect 76490 -44310 76610 -44250
rect 77760 -44480 77820 -44420
rect 77970 -44470 78030 -44350
rect 76920 -44610 77060 -44520
rect 77760 -44800 77820 -44740
rect 76490 -44950 76610 -44880
rect 77960 -44920 78020 -44850
rect 59076 -45710 59166 -45640
rect 60556 -45690 60626 -45610
rect 59976 -45752 60316 -45700
rect 59976 -45760 60316 -45752
rect 56480 -45848 56550 -45788
rect 57098 -45904 57368 -45764
rect 59286 -45920 59366 -45830
rect 59576 -45930 59636 -45870
rect 61206 -45900 61346 -45720
rect 76920 -45740 77060 -45640
rect 77600 -45680 77710 -45610
rect 59286 -46130 59356 -46040
rect 59916 -46160 60006 -45980
rect 60306 -46090 60456 -45950
rect 75220 -45950 75340 -45890
rect 78780 -44890 78920 -44770
rect 79410 -42880 79680 -42640
rect 79410 -44100 79680 -43860
rect 79070 -44870 79140 -44800
rect 79410 -45360 79680 -45120
rect 79080 -45680 79190 -45560
rect 78070 -45950 78140 -45890
rect 61036 -46130 61126 -46020
rect 55020 -46328 55030 -46248
rect 55030 -46328 55110 -46248
rect 55110 -46328 55120 -46248
rect 55880 -46328 55970 -46238
rect 56480 -46328 56550 -46238
rect 57800 -46340 58240 -46220
rect 58556 -46280 58756 -46260
rect 58556 -46440 58576 -46280
rect 58576 -46440 58736 -46280
rect 58736 -46440 58756 -46280
rect 58556 -46460 58756 -46440
rect 59076 -46280 59166 -46210
rect 59316 -46290 59376 -46230
rect 59076 -46440 59166 -46370
rect 60096 -46440 60176 -46280
rect 61276 -46460 61356 -46250
rect 75390 -46310 75550 -46190
rect 78770 -46310 78890 -46190
rect 81140 -40510 81570 -40250
rect 87830 -40590 88190 -40240
rect 80080 -41290 80430 -40910
rect 82460 -41290 82950 -40910
rect 80010 -43290 80360 -42910
rect 82120 -43290 82490 -42910
rect 80010 -45810 80360 -45430
rect 81510 -45810 81930 -45430
rect 79740 -46310 79910 -46190
rect 59266 -46610 59366 -46520
rect 56480 -46788 56550 -46728
rect 57098 -46814 57368 -46674
rect 59916 -46680 60006 -46490
rect 60476 -46570 60536 -46510
rect 59266 -46850 59366 -46760
rect 59516 -46720 59596 -46710
rect 59516 -46780 59596 -46720
rect 61336 -46760 61456 -46630
rect 55220 -47118 55310 -46948
rect 55410 -47128 55500 -46958
rect 59076 -47000 59166 -46940
rect 59316 -46980 59376 -46920
rect 59996 -46980 60106 -46920
rect 72820 -47080 73040 -46900
rect 53510 -47448 53630 -47328
rect 55880 -47358 55970 -47278
rect 55620 -47478 55710 -47388
rect 55220 -47718 55320 -47618
rect 56020 -47608 56080 -47458
rect 59256 -47290 59366 -47230
rect 59546 -47200 59606 -47190
rect 59546 -47260 59606 -47200
rect 59016 -47360 59076 -47300
rect 59546 -47370 59606 -47310
rect 59806 -47320 59916 -47210
rect 60446 -47350 60526 -47230
rect 55320 -48068 55470 -47928
rect 56654 -47686 56998 -47468
rect 62500 -47500 62900 -47200
rect 72820 -47410 73040 -47230
rect 59016 -47710 59076 -47640
rect 59546 -47710 59606 -47640
rect 60266 -47730 60406 -47600
rect 58966 -47820 59146 -47800
rect 58966 -47960 58986 -47820
rect 58986 -47960 59126 -47820
rect 59126 -47960 59146 -47820
rect 58966 -47980 59146 -47960
rect 59996 -47900 60106 -47790
rect 59700 -48400 60400 -48000
rect 62500 -48400 62900 -48000
rect 64200 -47900 64500 -47700
rect 55500 -48900 56100 -48500
rect 51500 -49700 52500 -49500
rect 55460 -49760 55720 -49480
rect 53460 -50340 53780 -50140
rect 53520 -50568 53640 -50458
rect 55960 -50488 56040 -50338
rect 55280 -50528 55400 -50518
rect 55280 -50598 55290 -50528
rect 55290 -50598 55390 -50528
rect 55390 -50598 55400 -50528
rect 55280 -50608 55400 -50598
rect 56506 -50430 57016 -50180
rect 58966 -50230 59126 -50070
rect 59336 -50250 59416 -50110
rect 60046 -50240 60126 -50120
rect 58996 -50440 59106 -50330
rect 59516 -50440 59616 -50340
rect 61056 -50450 61126 -50320
rect 53050 -52508 53250 -50758
rect 55880 -50698 55970 -50618
rect 55230 -51028 55320 -50858
rect 55600 -50998 55710 -50868
rect 58486 -50890 58816 -50530
rect 59286 -50790 59346 -50730
rect 59546 -50750 59606 -50690
rect 59006 -50860 59016 -50800
rect 59016 -50860 59066 -50800
rect 59546 -50870 59606 -50810
rect 59866 -50830 59966 -50740
rect 60446 -50820 60526 -50720
rect 60046 -50940 60126 -50920
rect 60046 -51000 60126 -50940
rect 59076 -51110 59166 -51040
rect 60556 -51090 60626 -51010
rect 59976 -51152 60316 -51100
rect 59976 -51160 60316 -51152
rect 56480 -51248 56550 -51188
rect 57098 -51304 57368 -51164
rect 59286 -51320 59366 -51230
rect 59576 -51330 59636 -51270
rect 61206 -51300 61346 -51120
rect 59286 -51530 59356 -51440
rect 59916 -51560 60006 -51380
rect 60306 -51490 60456 -51350
rect 61036 -51530 61126 -51420
rect 55020 -51728 55030 -51648
rect 55030 -51728 55110 -51648
rect 55110 -51728 55120 -51648
rect 55880 -51728 55970 -51638
rect 56480 -51728 56550 -51638
rect 57800 -51740 58240 -51620
rect 58556 -51680 58756 -51660
rect 58556 -51840 58576 -51680
rect 58576 -51840 58736 -51680
rect 58736 -51840 58756 -51680
rect 58556 -51860 58756 -51840
rect 59076 -51680 59166 -51610
rect 59316 -51690 59376 -51630
rect 59076 -51840 59166 -51770
rect 60096 -51840 60176 -51680
rect 61276 -51860 61356 -51650
rect 59266 -52010 59366 -51920
rect 56480 -52188 56550 -52128
rect 57098 -52214 57368 -52074
rect 59916 -52080 60006 -51890
rect 60476 -51970 60536 -51910
rect 59266 -52250 59366 -52160
rect 59516 -52120 59596 -52110
rect 59516 -52180 59596 -52120
rect 61336 -52160 61456 -52030
rect 55220 -52518 55310 -52348
rect 55410 -52528 55500 -52358
rect 59076 -52400 59166 -52340
rect 59316 -52380 59376 -52320
rect 59996 -52380 60106 -52320
rect 53510 -52848 53630 -52728
rect 55880 -52758 55970 -52678
rect 55620 -52878 55710 -52788
rect 55220 -53118 55320 -53018
rect 56020 -53008 56080 -52858
rect 59256 -52690 59366 -52630
rect 59546 -52600 59606 -52590
rect 59546 -52660 59606 -52600
rect 59016 -52760 59076 -52700
rect 59546 -52770 59606 -52710
rect 59806 -52720 59916 -52610
rect 60446 -52750 60526 -52630
rect 55320 -53468 55470 -53328
rect 56654 -53086 56998 -52868
rect 59016 -53110 59076 -53040
rect 59546 -53110 59606 -53040
rect 60266 -53130 60406 -53000
rect 58966 -53220 59146 -53200
rect 58966 -53360 58986 -53220
rect 58986 -53360 59126 -53220
rect 59126 -53360 59146 -53220
rect 58966 -53380 59146 -53360
rect 59996 -53300 60106 -53190
rect 59700 -53800 60400 -53400
rect 72820 -47900 73040 -47720
rect 64200 -53800 64500 -53400
rect 65100 -48300 65400 -48100
rect 72820 -48180 73040 -48000
rect 55400 -54300 56100 -53900
rect 51500 -55100 52500 -54900
rect 55460 -55160 55720 -54880
rect 53480 -55740 53780 -55540
rect 53520 -55968 53640 -55858
rect 55960 -55888 56040 -55738
rect 55280 -55928 55400 -55918
rect 55280 -55998 55290 -55928
rect 55290 -55998 55390 -55928
rect 55390 -55998 55400 -55928
rect 55280 -56008 55400 -55998
rect 56506 -55830 57016 -55580
rect 58966 -55630 59126 -55470
rect 59336 -55650 59416 -55510
rect 60046 -55640 60126 -55520
rect 58996 -55840 59106 -55730
rect 59516 -55840 59616 -55740
rect 61056 -55850 61126 -55720
rect 53050 -57908 53250 -56158
rect 55880 -56098 55970 -56018
rect 55230 -56428 55320 -56258
rect 55600 -56398 55710 -56268
rect 58486 -56290 58816 -55930
rect 59286 -56190 59346 -56130
rect 59546 -56150 59606 -56090
rect 59006 -56260 59016 -56200
rect 59016 -56260 59066 -56200
rect 59546 -56270 59606 -56210
rect 59866 -56230 59966 -56140
rect 60446 -56220 60526 -56120
rect 60046 -56340 60126 -56320
rect 60046 -56400 60126 -56340
rect 59076 -56510 59166 -56440
rect 60556 -56490 60626 -56410
rect 59976 -56552 60316 -56500
rect 59976 -56560 60316 -56552
rect 56480 -56648 56550 -56588
rect 57098 -56704 57368 -56564
rect 59286 -56720 59366 -56630
rect 59576 -56730 59636 -56670
rect 61206 -56700 61346 -56520
rect 59286 -56930 59356 -56840
rect 59916 -56960 60006 -56780
rect 60306 -56890 60456 -56750
rect 61036 -56930 61126 -56820
rect 55020 -57128 55030 -57048
rect 55030 -57128 55110 -57048
rect 55110 -57128 55120 -57048
rect 55880 -57128 55970 -57038
rect 56480 -57128 56550 -57038
rect 57800 -57140 58240 -57020
rect 58556 -57080 58756 -57060
rect 58556 -57240 58576 -57080
rect 58576 -57240 58736 -57080
rect 58736 -57240 58756 -57080
rect 58556 -57260 58756 -57240
rect 59076 -57080 59166 -57010
rect 59316 -57090 59376 -57030
rect 59076 -57240 59166 -57170
rect 60096 -57240 60176 -57080
rect 61276 -57260 61356 -57050
rect 59266 -57410 59366 -57320
rect 56480 -57588 56550 -57528
rect 57098 -57614 57368 -57474
rect 59916 -57480 60006 -57290
rect 60476 -57370 60536 -57310
rect 59266 -57650 59366 -57560
rect 59516 -57520 59596 -57510
rect 59516 -57580 59596 -57520
rect 61336 -57560 61456 -57430
rect 55220 -57918 55310 -57748
rect 55410 -57928 55500 -57758
rect 59076 -57800 59166 -57740
rect 59316 -57780 59376 -57720
rect 59996 -57780 60106 -57720
rect 53510 -58248 53630 -58128
rect 55880 -58158 55970 -58078
rect 55620 -58278 55710 -58188
rect 55220 -58518 55320 -58418
rect 56020 -58408 56080 -58258
rect 59256 -58090 59366 -58030
rect 59546 -58000 59606 -57990
rect 59546 -58060 59606 -58000
rect 59016 -58160 59076 -58100
rect 59546 -58170 59606 -58110
rect 59806 -58120 59916 -58010
rect 60446 -58150 60526 -58030
rect 55320 -58868 55470 -58728
rect 56654 -58486 56998 -58268
rect 59016 -58510 59076 -58440
rect 59546 -58510 59606 -58440
rect 60266 -58530 60406 -58400
rect 58966 -58620 59146 -58600
rect 58966 -58760 58986 -58620
rect 58986 -58760 59126 -58620
rect 59126 -58760 59146 -58620
rect 58966 -58780 59146 -58760
rect 59996 -58700 60106 -58590
rect 59700 -59200 60400 -58800
rect 65100 -59200 65400 -58800
rect 66100 -48700 66400 -48500
rect 72820 -48640 73040 -48460
rect 55500 -59700 56100 -59300
rect 51500 -60500 52500 -60300
rect 55460 -60560 55720 -60280
rect 53480 -61140 53780 -60940
rect 53520 -61368 53640 -61258
rect 55960 -61288 56040 -61138
rect 55280 -61328 55400 -61318
rect 55280 -61398 55290 -61328
rect 55290 -61398 55390 -61328
rect 55390 -61398 55400 -61328
rect 55280 -61408 55400 -61398
rect 56506 -61230 57016 -60980
rect 58966 -61030 59126 -60870
rect 59336 -61050 59416 -60910
rect 60046 -61040 60126 -60920
rect 58996 -61240 59106 -61130
rect 59516 -61240 59616 -61140
rect 61056 -61250 61126 -61120
rect 53050 -63308 53250 -61558
rect 55880 -61498 55970 -61418
rect 55230 -61828 55320 -61658
rect 55600 -61798 55710 -61668
rect 58486 -61690 58816 -61330
rect 59286 -61590 59346 -61530
rect 59546 -61550 59606 -61490
rect 59006 -61660 59016 -61600
rect 59016 -61660 59066 -61600
rect 59546 -61670 59606 -61610
rect 59866 -61630 59966 -61540
rect 60446 -61620 60526 -61520
rect 60046 -61740 60126 -61720
rect 60046 -61800 60126 -61740
rect 59076 -61910 59166 -61840
rect 60556 -61890 60626 -61810
rect 59976 -61952 60316 -61900
rect 59976 -61960 60316 -61952
rect 56480 -62048 56550 -61988
rect 57098 -62104 57368 -61964
rect 59286 -62120 59366 -62030
rect 59576 -62130 59636 -62070
rect 61206 -62100 61346 -61920
rect 59286 -62330 59356 -62240
rect 59916 -62360 60006 -62180
rect 60306 -62290 60456 -62150
rect 61036 -62330 61126 -62220
rect 55020 -62528 55030 -62448
rect 55030 -62528 55110 -62448
rect 55110 -62528 55120 -62448
rect 55880 -62528 55970 -62438
rect 56480 -62528 56550 -62438
rect 57800 -62540 58240 -62420
rect 58556 -62480 58756 -62460
rect 58556 -62640 58576 -62480
rect 58576 -62640 58736 -62480
rect 58736 -62640 58756 -62480
rect 58556 -62660 58756 -62640
rect 59076 -62480 59166 -62410
rect 59316 -62490 59376 -62430
rect 59076 -62640 59166 -62570
rect 60096 -62640 60176 -62480
rect 61276 -62660 61356 -62450
rect 59266 -62810 59366 -62720
rect 56480 -62988 56550 -62928
rect 57098 -63014 57368 -62874
rect 59916 -62880 60006 -62690
rect 60476 -62770 60536 -62710
rect 59266 -63050 59366 -62960
rect 59516 -62920 59596 -62910
rect 59516 -62980 59596 -62920
rect 61336 -62960 61456 -62830
rect 55220 -63318 55310 -63148
rect 55410 -63328 55500 -63158
rect 59076 -63200 59166 -63140
rect 59316 -63180 59376 -63120
rect 59996 -63180 60106 -63120
rect 53510 -63648 53630 -63528
rect 55880 -63558 55970 -63478
rect 55620 -63678 55710 -63588
rect 55220 -63918 55320 -63818
rect 56020 -63808 56080 -63658
rect 59256 -63490 59366 -63430
rect 59546 -63400 59606 -63390
rect 59546 -63460 59606 -63400
rect 59016 -63560 59076 -63500
rect 59546 -63570 59606 -63510
rect 59806 -63520 59916 -63410
rect 60446 -63550 60526 -63430
rect 55320 -64268 55470 -64128
rect 56654 -63886 56998 -63668
rect 59016 -63910 59076 -63840
rect 59546 -63910 59606 -63840
rect 60266 -63930 60406 -63800
rect 58966 -64020 59146 -64000
rect 58966 -64160 58986 -64020
rect 58986 -64160 59126 -64020
rect 59126 -64160 59146 -64020
rect 58966 -64180 59146 -64160
rect 59996 -64100 60106 -63990
rect 59700 -64600 60400 -64200
rect 66100 -64600 66400 -64200
rect 67100 -49100 67400 -48900
rect 72820 -49000 73040 -48820
rect 55500 -65100 56100 -64700
rect 51500 -65900 52500 -65700
rect 55440 -65960 55720 -65680
rect 53480 -66540 53780 -66340
rect 53520 -66768 53640 -66658
rect 55960 -66688 56040 -66538
rect 55280 -66728 55400 -66718
rect 55280 -66798 55290 -66728
rect 55290 -66798 55390 -66728
rect 55390 -66798 55400 -66728
rect 55280 -66808 55400 -66798
rect 56506 -66630 57016 -66380
rect 58966 -66430 59126 -66270
rect 59336 -66450 59416 -66310
rect 60046 -66440 60126 -66320
rect 58996 -66640 59106 -66530
rect 59516 -66640 59616 -66540
rect 61056 -66650 61126 -66520
rect 53050 -68708 53250 -66958
rect 55880 -66898 55970 -66818
rect 55230 -67228 55320 -67058
rect 55600 -67198 55710 -67068
rect 58486 -67090 58816 -66730
rect 59286 -66990 59346 -66930
rect 59546 -66950 59606 -66890
rect 59006 -67060 59016 -67000
rect 59016 -67060 59066 -67000
rect 59546 -67070 59606 -67010
rect 59866 -67030 59966 -66940
rect 60446 -67020 60526 -66920
rect 60046 -67140 60126 -67120
rect 60046 -67200 60126 -67140
rect 59076 -67310 59166 -67240
rect 60556 -67290 60626 -67210
rect 59976 -67352 60316 -67300
rect 59976 -67360 60316 -67352
rect 56480 -67448 56550 -67388
rect 57098 -67504 57368 -67364
rect 59286 -67520 59366 -67430
rect 59576 -67530 59636 -67470
rect 61206 -67500 61346 -67320
rect 59286 -67730 59356 -67640
rect 59916 -67760 60006 -67580
rect 60306 -67690 60456 -67550
rect 61036 -67730 61126 -67620
rect 55020 -67928 55030 -67848
rect 55030 -67928 55110 -67848
rect 55110 -67928 55120 -67848
rect 55880 -67928 55970 -67838
rect 56480 -67928 56550 -67838
rect 57800 -67940 58240 -67820
rect 58556 -67880 58756 -67860
rect 58556 -68040 58576 -67880
rect 58576 -68040 58736 -67880
rect 58736 -68040 58756 -67880
rect 58556 -68060 58756 -68040
rect 59076 -67880 59166 -67810
rect 59316 -67890 59376 -67830
rect 59076 -68040 59166 -67970
rect 60096 -68040 60176 -67880
rect 61276 -68060 61356 -67850
rect 59266 -68210 59366 -68120
rect 56480 -68388 56550 -68328
rect 57098 -68414 57368 -68274
rect 59916 -68280 60006 -68090
rect 60476 -68170 60536 -68110
rect 59266 -68450 59366 -68360
rect 59516 -68320 59596 -68310
rect 59516 -68380 59596 -68320
rect 61336 -68360 61456 -68230
rect 55220 -68718 55310 -68548
rect 55410 -68728 55500 -68558
rect 59076 -68600 59166 -68540
rect 59316 -68580 59376 -68520
rect 59996 -68580 60106 -68520
rect 53510 -69048 53630 -68928
rect 55880 -68958 55970 -68878
rect 55620 -69078 55710 -68988
rect 55220 -69318 55320 -69218
rect 56020 -69208 56080 -69058
rect 59256 -68890 59366 -68830
rect 59546 -68800 59606 -68790
rect 59546 -68860 59606 -68800
rect 59016 -68960 59076 -68900
rect 59546 -68970 59606 -68910
rect 59806 -68920 59916 -68810
rect 60446 -68950 60526 -68830
rect 55320 -69668 55470 -69528
rect 56654 -69286 56998 -69068
rect 59016 -69310 59076 -69240
rect 59546 -69310 59606 -69240
rect 60266 -69330 60406 -69200
rect 58966 -69420 59146 -69400
rect 58966 -69560 58986 -69420
rect 58986 -69560 59126 -69420
rect 59126 -69560 59146 -69420
rect 58966 -69580 59146 -69560
rect 59996 -69500 60106 -69390
rect 59700 -70000 60400 -69600
rect 67100 -70000 67400 -69600
rect 68000 -49500 68300 -49300
rect 72820 -49400 73040 -49220
rect 55500 -70500 56100 -70100
rect 51500 -71300 52500 -71100
rect 55460 -71360 55720 -71080
rect 53480 -71940 53780 -71740
rect 53520 -72168 53640 -72058
rect 55960 -72088 56040 -71938
rect 55280 -72128 55400 -72118
rect 55280 -72198 55290 -72128
rect 55290 -72198 55390 -72128
rect 55390 -72198 55400 -72128
rect 55280 -72208 55400 -72198
rect 56506 -72030 57016 -71780
rect 58966 -71830 59126 -71670
rect 59336 -71850 59416 -71710
rect 60046 -71840 60126 -71720
rect 58996 -72040 59106 -71930
rect 59516 -72040 59616 -71940
rect 61056 -72050 61126 -71920
rect 53050 -74108 53250 -72358
rect 55880 -72298 55970 -72218
rect 55230 -72628 55320 -72458
rect 55600 -72598 55710 -72468
rect 58486 -72490 58816 -72130
rect 59286 -72390 59346 -72330
rect 59546 -72350 59606 -72290
rect 59006 -72460 59016 -72400
rect 59016 -72460 59066 -72400
rect 59546 -72470 59606 -72410
rect 59866 -72430 59966 -72340
rect 60446 -72420 60526 -72320
rect 60046 -72540 60126 -72520
rect 60046 -72600 60126 -72540
rect 59076 -72710 59166 -72640
rect 60556 -72690 60626 -72610
rect 59976 -72752 60316 -72700
rect 59976 -72760 60316 -72752
rect 56480 -72848 56550 -72788
rect 57098 -72904 57368 -72764
rect 59286 -72920 59366 -72830
rect 59576 -72930 59636 -72870
rect 61206 -72900 61346 -72720
rect 59286 -73130 59356 -73040
rect 59916 -73160 60006 -72980
rect 60306 -73090 60456 -72950
rect 61036 -73130 61126 -73020
rect 55020 -73328 55030 -73248
rect 55030 -73328 55110 -73248
rect 55110 -73328 55120 -73248
rect 55880 -73328 55970 -73238
rect 56480 -73328 56550 -73238
rect 57800 -73340 58240 -73220
rect 58556 -73280 58756 -73260
rect 58556 -73440 58576 -73280
rect 58576 -73440 58736 -73280
rect 58736 -73440 58756 -73280
rect 58556 -73460 58756 -73440
rect 59076 -73280 59166 -73210
rect 59316 -73290 59376 -73230
rect 59076 -73440 59166 -73370
rect 60096 -73440 60176 -73280
rect 61276 -73460 61356 -73250
rect 59266 -73610 59366 -73520
rect 56480 -73788 56550 -73728
rect 57098 -73814 57368 -73674
rect 59916 -73680 60006 -73490
rect 60476 -73570 60536 -73510
rect 59266 -73850 59366 -73760
rect 59516 -73720 59596 -73710
rect 59516 -73780 59596 -73720
rect 61336 -73760 61456 -73630
rect 55220 -74118 55310 -73948
rect 55410 -74128 55500 -73958
rect 59076 -74000 59166 -73940
rect 59316 -73980 59376 -73920
rect 59996 -73980 60106 -73920
rect 53510 -74448 53630 -74328
rect 55880 -74358 55970 -74278
rect 55620 -74478 55710 -74388
rect 55220 -74718 55320 -74618
rect 56020 -74608 56080 -74458
rect 59256 -74290 59366 -74230
rect 59546 -74200 59606 -74190
rect 59546 -74260 59606 -74200
rect 59016 -74360 59076 -74300
rect 59546 -74370 59606 -74310
rect 59806 -74320 59916 -74210
rect 60446 -74350 60526 -74230
rect 55320 -75068 55470 -74928
rect 56654 -74686 56998 -74468
rect 59016 -74710 59076 -74640
rect 59546 -74710 59606 -74640
rect 60266 -74730 60406 -74600
rect 58966 -74820 59146 -74800
rect 58966 -74960 58986 -74820
rect 58986 -74960 59126 -74820
rect 59126 -74960 59146 -74820
rect 58966 -74980 59146 -74960
rect 59996 -74900 60106 -74790
rect 59700 -75400 60400 -75000
rect 68000 -75400 68300 -75000
rect 69000 -49900 69300 -49700
rect 72820 -49850 73040 -49670
rect 55500 -75900 56100 -75500
rect 51500 -76700 52500 -76500
rect 55400 -76760 55720 -76480
rect 53480 -77340 53780 -77140
rect 53520 -77568 53640 -77458
rect 55960 -77488 56040 -77338
rect 55280 -77528 55400 -77518
rect 55280 -77598 55290 -77528
rect 55290 -77598 55390 -77528
rect 55390 -77598 55400 -77528
rect 55280 -77608 55400 -77598
rect 56506 -77430 57016 -77180
rect 58966 -77230 59126 -77070
rect 59336 -77250 59416 -77110
rect 60046 -77240 60126 -77120
rect 58996 -77440 59106 -77330
rect 59516 -77440 59616 -77340
rect 61056 -77450 61126 -77320
rect 53050 -79508 53250 -77758
rect 55880 -77698 55970 -77618
rect 55230 -78028 55320 -77858
rect 55600 -77998 55710 -77868
rect 58486 -77890 58816 -77530
rect 59286 -77790 59346 -77730
rect 59546 -77750 59606 -77690
rect 59006 -77860 59016 -77800
rect 59016 -77860 59066 -77800
rect 59546 -77870 59606 -77810
rect 59866 -77830 59966 -77740
rect 60446 -77820 60526 -77720
rect 60046 -77940 60126 -77920
rect 60046 -78000 60126 -77940
rect 59076 -78110 59166 -78040
rect 60556 -78090 60626 -78010
rect 59976 -78152 60316 -78100
rect 59976 -78160 60316 -78152
rect 56480 -78248 56550 -78188
rect 57098 -78304 57368 -78164
rect 59286 -78320 59366 -78230
rect 59576 -78330 59636 -78270
rect 61206 -78300 61346 -78120
rect 59286 -78530 59356 -78440
rect 59916 -78560 60006 -78380
rect 60306 -78490 60456 -78350
rect 61036 -78530 61126 -78420
rect 55020 -78728 55030 -78648
rect 55030 -78728 55110 -78648
rect 55110 -78728 55120 -78648
rect 55880 -78728 55970 -78638
rect 56480 -78728 56550 -78638
rect 57800 -78740 58240 -78620
rect 58556 -78680 58756 -78660
rect 58556 -78840 58576 -78680
rect 58576 -78840 58736 -78680
rect 58736 -78840 58756 -78680
rect 58556 -78860 58756 -78840
rect 59076 -78680 59166 -78610
rect 59316 -78690 59376 -78630
rect 59076 -78840 59166 -78770
rect 60096 -78840 60176 -78680
rect 61276 -78860 61356 -78650
rect 59266 -79010 59366 -78920
rect 56480 -79188 56550 -79128
rect 57098 -79214 57368 -79074
rect 59916 -79080 60006 -78890
rect 60476 -78970 60536 -78910
rect 59266 -79250 59366 -79160
rect 59516 -79120 59596 -79110
rect 59516 -79180 59596 -79120
rect 61336 -79160 61456 -79030
rect 55220 -79518 55310 -79348
rect 55410 -79528 55500 -79358
rect 59076 -79400 59166 -79340
rect 59316 -79380 59376 -79320
rect 59996 -79380 60106 -79320
rect 53510 -79848 53630 -79728
rect 55880 -79758 55970 -79678
rect 55620 -79878 55710 -79788
rect 55220 -80118 55320 -80018
rect 56020 -80008 56080 -79858
rect 59256 -79690 59366 -79630
rect 59546 -79600 59606 -79590
rect 59546 -79660 59606 -79600
rect 59016 -79760 59076 -79700
rect 59546 -79770 59606 -79710
rect 59806 -79720 59916 -79610
rect 60446 -79750 60526 -79630
rect 55320 -80468 55470 -80328
rect 56654 -80086 56998 -79868
rect 59016 -80110 59076 -80040
rect 59546 -80110 59606 -80040
rect 60266 -80130 60406 -80000
rect 58966 -80220 59146 -80200
rect 58966 -80360 58986 -80220
rect 58986 -80360 59126 -80220
rect 59126 -80360 59146 -80220
rect 58966 -80380 59146 -80360
rect 59996 -80300 60106 -80190
rect 59700 -80800 60400 -80400
rect 69000 -80800 69300 -80400
rect 70000 -50300 70300 -50100
rect 72820 -50220 73040 -50040
rect 73220 -50200 73340 -50060
rect 73470 -49830 73590 -49690
rect 55500 -81300 56200 -80900
rect 51500 -82100 52500 -81900
rect 37200 -86700 37700 -86200
rect 55440 -82160 55720 -81880
rect 53480 -82740 53780 -82540
rect 53520 -82968 53640 -82858
rect 55960 -82888 56040 -82738
rect 55280 -82928 55400 -82918
rect 55280 -82998 55290 -82928
rect 55290 -82998 55390 -82928
rect 55390 -82998 55400 -82928
rect 55280 -83008 55400 -82998
rect 56506 -82830 57016 -82580
rect 58966 -82630 59126 -82470
rect 59336 -82650 59416 -82510
rect 60046 -82640 60126 -82520
rect 58996 -82840 59106 -82730
rect 59516 -82840 59616 -82740
rect 61056 -82850 61126 -82720
rect 53050 -84908 53250 -83158
rect 55880 -83098 55970 -83018
rect 55230 -83428 55320 -83258
rect 55600 -83398 55710 -83268
rect 58486 -83290 58816 -82930
rect 59286 -83190 59346 -83130
rect 59546 -83150 59606 -83090
rect 59006 -83260 59016 -83200
rect 59016 -83260 59066 -83200
rect 59546 -83270 59606 -83210
rect 59866 -83230 59966 -83140
rect 60446 -83220 60526 -83120
rect 60046 -83340 60126 -83320
rect 60046 -83400 60126 -83340
rect 59076 -83510 59166 -83440
rect 60556 -83490 60626 -83410
rect 59976 -83552 60316 -83500
rect 59976 -83560 60316 -83552
rect 56480 -83648 56550 -83588
rect 57098 -83704 57368 -83564
rect 59286 -83720 59366 -83630
rect 59576 -83730 59636 -83670
rect 61206 -83700 61346 -83520
rect 59286 -83930 59356 -83840
rect 59916 -83960 60006 -83780
rect 60306 -83890 60456 -83750
rect 61036 -83930 61126 -83820
rect 55020 -84128 55030 -84048
rect 55030 -84128 55110 -84048
rect 55110 -84128 55120 -84048
rect 55880 -84128 55970 -84038
rect 56480 -84128 56550 -84038
rect 57800 -84140 58240 -84020
rect 58556 -84080 58756 -84060
rect 58556 -84240 58576 -84080
rect 58576 -84240 58736 -84080
rect 58736 -84240 58756 -84080
rect 58556 -84260 58756 -84240
rect 59076 -84080 59166 -84010
rect 59316 -84090 59376 -84030
rect 59076 -84240 59166 -84170
rect 60096 -84240 60176 -84080
rect 61276 -84260 61356 -84050
rect 59266 -84410 59366 -84320
rect 56480 -84588 56550 -84528
rect 57098 -84614 57368 -84474
rect 59916 -84480 60006 -84290
rect 60476 -84370 60536 -84310
rect 59266 -84650 59366 -84560
rect 59516 -84520 59596 -84510
rect 59516 -84580 59596 -84520
rect 61336 -84560 61456 -84430
rect 55220 -84918 55310 -84748
rect 55410 -84928 55500 -84758
rect 59076 -84800 59166 -84740
rect 59316 -84780 59376 -84720
rect 59996 -84780 60106 -84720
rect 53510 -85248 53630 -85128
rect 55880 -85158 55970 -85078
rect 55620 -85278 55710 -85188
rect 55220 -85518 55320 -85418
rect 56020 -85408 56080 -85258
rect 59256 -85090 59366 -85030
rect 59546 -85000 59606 -84990
rect 59546 -85060 59606 -85000
rect 59016 -85160 59076 -85100
rect 59546 -85170 59606 -85110
rect 59806 -85120 59916 -85010
rect 60446 -85150 60526 -85030
rect 55320 -85868 55470 -85728
rect 56654 -85486 56998 -85268
rect 59016 -85510 59076 -85440
rect 59546 -85510 59606 -85440
rect 60266 -85530 60406 -85400
rect 58966 -85620 59146 -85600
rect 58966 -85760 58986 -85620
rect 58986 -85760 59126 -85620
rect 59126 -85760 59146 -85620
rect 58966 -85780 59146 -85760
rect 59996 -85700 60106 -85590
rect 59700 -86200 60400 -85800
rect 73720 -49380 73840 -49240
rect 73720 -51040 73840 -50970
rect 73970 -47530 74090 -47470
rect 74220 -48490 74340 -48430
rect 74477 -46714 74594 -46610
rect 74470 -48220 74590 -48150
rect 73970 -48980 74090 -48840
rect 73470 -52480 73590 -52420
rect 73970 -51870 74090 -51800
rect 73970 -52840 74090 -52780
rect 74470 -49420 74590 -49360
rect 74724 -46870 74841 -46792
rect 74720 -47880 74840 -47740
rect 74720 -49730 74840 -49670
rect 74970 -47380 75090 -47260
rect 74980 -47890 75080 -47820
rect 74970 -50370 75090 -50310
rect 75231 -46532 75322 -46467
rect 76648 -46545 76726 -46480
rect 75220 -47180 75340 -47080
rect 76102 -46701 76167 -46623
rect 76167 -46701 76180 -46623
rect 76375 -46844 76440 -46766
rect 75220 -48650 75340 -48580
rect 75220 -49280 75340 -49200
rect 75220 -49900 75340 -49810
rect 74470 -53600 74590 -53520
rect 75220 -50540 75340 -50450
rect 75220 -51290 75340 -51230
rect 75220 -51720 75340 -51660
rect 76920 -46570 77060 -46450
rect 76780 -46714 76791 -46670
rect 76791 -46714 76843 -46670
rect 76843 -46714 76860 -46670
rect 76780 -46740 76860 -46714
rect 78280 -46740 78350 -46670
rect 76210 -51170 76340 -51110
rect 77170 -47080 77430 -46830
rect 77230 -47540 77310 -47480
rect 76920 -47760 77060 -47610
rect 77170 -47890 77260 -47820
rect 79080 -47550 79250 -47390
rect 80080 -47620 80430 -47310
rect 78580 -47940 78640 -47880
rect 80080 -48100 80430 -47720
rect 77410 -48220 77480 -48150
rect 77780 -48490 77840 -48430
rect 79410 -48430 79680 -48190
rect 77450 -48650 77520 -48580
rect 76920 -49000 77060 -48860
rect 77450 -49280 77530 -49200
rect 77780 -49420 77840 -49360
rect 77780 -49730 77840 -49670
rect 77490 -49900 77580 -49810
rect 76920 -50250 77060 -50100
rect 77780 -50370 77840 -50310
rect 77470 -50540 77560 -50450
rect 78670 -49220 78780 -49070
rect 80080 -49330 80430 -48950
rect 79410 -49660 79680 -49420
rect 78160 -50510 78260 -50410
rect 79050 -50510 79150 -50400
rect 77470 -51030 77540 -50970
rect 77860 -51150 77920 -51090
rect 76920 -51490 77060 -51350
rect 77960 -51290 78020 -51230
rect 78860 -51250 78980 -50960
rect 77970 -51720 78030 -51660
rect 77430 -51870 77500 -51800
rect 76490 -52350 76610 -52290
rect 77760 -52520 77820 -52460
rect 77970 -52510 78030 -52390
rect 76920 -52650 77060 -52560
rect 77760 -52840 77820 -52780
rect 76490 -52990 76610 -52920
rect 77960 -52960 78020 -52890
rect 76920 -53780 77060 -53680
rect 77600 -53720 77710 -53650
rect 75220 -53990 75340 -53930
rect 78780 -52930 78920 -52810
rect 79410 -50920 79680 -50680
rect 80010 -51330 80360 -50950
rect 82220 -48140 82340 -48020
rect 82820 -43310 91410 -42740
rect 85320 -43540 85390 -43450
rect 82640 -44000 82720 -43890
rect 83040 -44000 83100 -43890
rect 85590 -43540 86480 -43450
rect 87040 -43540 87920 -43450
rect 88510 -43540 89390 -43450
rect 86800 -44310 86870 -44230
rect 89980 -43540 90760 -43450
rect 88270 -44310 88340 -44230
rect 89750 -44310 89810 -44230
rect 91210 -44310 91280 -44230
rect 82820 -45010 91410 -44440
rect 91780 -44460 92130 -44080
rect 82824 -47448 91414 -46878
rect 85324 -47678 85394 -47588
rect 83040 -48140 83100 -48020
rect 85594 -47678 86484 -47588
rect 87044 -47678 87924 -47588
rect 88514 -47678 89394 -47588
rect 86804 -48448 86874 -48368
rect 89984 -47678 90764 -47588
rect 88274 -48448 88344 -48368
rect 89754 -48448 89814 -48368
rect 91214 -48448 91284 -48368
rect 82450 -49330 82610 -48950
rect 82824 -49148 91414 -48578
rect 91780 -48620 92130 -48240
rect 82820 -51100 91410 -50530
rect 81950 -51350 82070 -51140
rect 85320 -51330 85390 -51240
rect 81640 -51790 81760 -51680
rect 79410 -52140 79680 -51900
rect 79070 -52910 79140 -52840
rect 79410 -53400 79680 -53160
rect 79080 -53720 79190 -53600
rect 83030 -51790 83100 -51680
rect 85590 -51330 86480 -51240
rect 87040 -51330 87920 -51240
rect 88510 -51330 89390 -51240
rect 86800 -52100 86870 -52020
rect 89980 -51330 90760 -51240
rect 88270 -52100 88340 -52020
rect 89750 -52100 89810 -52020
rect 91210 -52100 91280 -52020
rect 82820 -52800 91410 -52230
rect 91780 -52250 92130 -51870
rect 80010 -53850 80360 -53470
rect 82140 -53850 82750 -53470
rect 78070 -53990 78140 -53930
rect 70000 -86200 70300 -85800
rect 55500 -86600 56100 -86300
<< metal3 >>
rect 37800 2800 41600 3000
rect 37800 1400 38000 2800
rect 41400 1400 41600 2800
rect 37800 1200 41600 1400
rect 42800 2400 46600 2600
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 800 46600 1000
rect 56870 1020 59090 1025
rect 42800 0 46600 200
rect 37800 -400 41600 -300
rect 37800 -3600 37900 -400
rect 41500 -3600 41600 -400
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 56870 -40 56880 1020
rect 59080 -40 59090 1020
rect 56870 -45 59090 -40
rect 55300 -600 55800 -500
rect 55300 -700 55400 -600
rect 51400 -800 55400 -700
rect 51400 -1000 51500 -800
rect 52500 -1000 55400 -800
rect 55700 -1000 55800 -600
rect 51400 -1100 55800 -1000
rect 42800 -1600 46600 -1400
rect 47600 -1300 48100 -1200
rect 47600 -1700 47700 -1300
rect 48000 -1400 53800 -1300
rect 48000 -1600 53400 -1400
rect 53700 -1600 53800 -1400
rect 48000 -1700 53800 -1600
rect 56496 -1580 57026 -1575
rect 47600 -1800 48100 -1700
rect 55955 -1738 56045 -1728
rect 53515 -1858 53645 -1848
rect 53510 -1968 53520 -1858
rect 53640 -1968 53645 -1858
rect 55955 -1888 55960 -1738
rect 56040 -1888 56200 -1738
rect 56496 -1830 56506 -1580
rect 57016 -1830 57026 -1580
rect 56496 -1835 57026 -1830
rect 55955 -1898 56200 -1888
rect 53510 -1978 53645 -1968
rect 55275 -1918 55490 -1908
rect 37800 -3700 41600 -3600
rect 53045 -2158 53255 -2148
rect 53045 -3908 53050 -2158
rect 53250 -3908 53255 -2158
rect 53045 -3918 53255 -3908
rect 53510 -4118 53630 -1978
rect 55275 -2008 55280 -1918
rect 55400 -2008 55490 -1918
rect 56060 -1938 56200 -1898
rect 56060 -1948 56220 -1938
rect 55275 -2018 55490 -2008
rect 55220 -2258 55325 -2248
rect 55220 -2428 55230 -2258
rect 55320 -2428 55325 -2258
rect 55220 -2438 55325 -2428
rect 55015 -3048 55125 -3038
rect 55015 -3128 55020 -3048
rect 55120 -3128 55125 -3048
rect 55015 -3138 55125 -3128
rect 55220 -3738 55310 -2438
rect 55215 -3748 55315 -3738
rect 55215 -3918 55220 -3748
rect 55310 -3838 55315 -3748
rect 55400 -3748 55490 -2018
rect 55875 -2018 55990 -2008
rect 55875 -2058 55880 -2018
rect 55870 -2098 55880 -2058
rect 55970 -2098 55990 -2018
rect 55870 -2178 55990 -2098
rect 56060 -2118 56220 -2108
rect 55590 -2268 55720 -2258
rect 55590 -2398 55600 -2268
rect 55710 -2398 55720 -2268
rect 55400 -3758 55510 -3748
rect 55310 -3918 55320 -3838
rect 55400 -3918 55410 -3758
rect 55215 -3928 55320 -3918
rect 53505 -4128 53635 -4118
rect 53505 -4248 53510 -4128
rect 53630 -4248 53635 -4128
rect 53505 -4258 53635 -4248
rect 55220 -4408 55320 -3928
rect 55405 -3928 55410 -3918
rect 55500 -3928 55510 -3758
rect 55405 -3938 55510 -3928
rect 55590 -4188 55720 -2398
rect 55870 -2558 55980 -2178
rect 57093 -2564 57373 -2554
rect 56475 -2588 56555 -2578
rect 56470 -2648 56480 -2588
rect 56550 -2648 56555 -2588
rect 56470 -2658 56555 -2648
rect 55870 -3038 55980 -2668
rect 55870 -3128 55880 -3038
rect 55970 -3128 55980 -3038
rect 55870 -3528 55980 -3128
rect 56470 -3028 56550 -2658
rect 57093 -2704 57098 -2564
rect 57368 -2704 57373 -2564
rect 57093 -2714 57373 -2704
rect 57760 -3020 58280 -45
rect 58946 -1470 59146 -1450
rect 58946 -1630 58966 -1470
rect 59126 -1630 59146 -1470
rect 58946 -1650 59146 -1630
rect 59316 -1510 59426 -1450
rect 59316 -1650 59336 -1510
rect 59416 -1650 59426 -1510
rect 58956 -1730 59136 -1650
rect 58956 -1840 58996 -1730
rect 59106 -1840 59136 -1730
rect 58396 -1930 58896 -1840
rect 58956 -1900 59136 -1840
rect 59316 -1880 59426 -1650
rect 59946 -1520 60386 -1400
rect 59946 -1640 60046 -1520
rect 60126 -1640 60386 -1520
rect 59946 -1690 60386 -1640
rect 58396 -2290 58486 -1930
rect 58816 -2290 58896 -1930
rect 58996 -2200 59086 -1900
rect 58996 -2260 59006 -2200
rect 59066 -2260 59086 -2200
rect 58996 -2270 59086 -2260
rect 59266 -1930 59426 -1880
rect 59506 -1740 59796 -1700
rect 59506 -1840 59516 -1740
rect 59616 -1840 59796 -1740
rect 59506 -1900 59796 -1840
rect 59266 -2130 59366 -1930
rect 59266 -2190 59286 -2130
rect 59346 -2190 59366 -2130
rect 58396 -2400 58896 -2290
rect 59066 -2440 59176 -2430
rect 59066 -2510 59076 -2440
rect 59166 -2510 59176 -2440
rect 56470 -3038 56555 -3028
rect 56470 -3128 56480 -3038
rect 56550 -3128 56555 -3038
rect 56470 -3138 56555 -3128
rect 56470 -3518 56550 -3138
rect 57760 -3140 57800 -3020
rect 58240 -3140 58280 -3020
rect 57093 -3474 57373 -3464
rect 56470 -3528 56555 -3518
rect 56470 -3578 56480 -3528
rect 56475 -3588 56480 -3578
rect 56550 -3588 56555 -3528
rect 56475 -3598 56555 -3588
rect 57093 -3614 57098 -3474
rect 57368 -3614 57373 -3474
rect 57093 -3624 57373 -3614
rect 55870 -4078 55980 -3638
rect 55870 -4118 55880 -4078
rect 55875 -4158 55880 -4118
rect 55970 -4118 55980 -4078
rect 56060 -4068 56220 -4058
rect 55970 -4158 55975 -4118
rect 55875 -4168 55975 -4158
rect 55590 -4278 55620 -4188
rect 55710 -4278 55720 -4188
rect 56060 -4238 56220 -4228
rect 56060 -4248 56200 -4238
rect 55590 -4288 55720 -4278
rect 56015 -4258 56200 -4248
rect 56015 -4408 56020 -4258
rect 56080 -4408 56200 -4258
rect 56644 -4268 57008 -4263
rect 55215 -4418 55325 -4408
rect 56015 -4418 56085 -4408
rect 55215 -4518 55220 -4418
rect 55320 -4518 55325 -4418
rect 56644 -4486 56654 -4268
rect 56998 -4486 57008 -4268
rect 56644 -4491 57008 -4486
rect 55215 -4528 55325 -4518
rect 55315 -4728 55475 -4718
rect 36200 -5000 37200 -4800
rect 55315 -4868 55320 -4728
rect 55470 -4868 55475 -4728
rect 55315 -4878 55475 -4868
rect 36200 -5800 36400 -5000
rect 37000 -5200 37200 -5000
rect 37000 -5300 56000 -5200
rect 37000 -5600 55600 -5300
rect 55900 -5600 56000 -5300
rect 37000 -5700 56000 -5600
rect 37000 -5800 37200 -5700
rect 36200 -6000 37200 -5800
rect 55300 -6200 55800 -6100
rect 51400 -6300 55400 -6200
rect 20800 -6600 22200 -6400
rect 51400 -6500 51500 -6300
rect 52500 -6500 55400 -6300
rect 55700 -6500 55800 -6200
rect 51400 -6600 55800 -6500
rect 20800 -7400 21000 -6600
rect 22000 -7400 22200 -6600
rect 47620 -6780 48100 -6760
rect 47620 -7200 47640 -6780
rect 48080 -6840 48100 -6780
rect 48080 -6860 53800 -6840
rect 48080 -7120 53520 -6860
rect 53780 -7120 53800 -6860
rect 48080 -7140 53800 -7120
rect 56496 -6980 57026 -6975
rect 55955 -7138 56045 -7128
rect 48080 -7200 48100 -7140
rect 47620 -7220 48100 -7200
rect 53515 -7258 53645 -7248
rect 20800 -7600 22200 -7400
rect 53510 -7368 53520 -7258
rect 53640 -7368 53645 -7258
rect 55955 -7288 55960 -7138
rect 56040 -7288 56200 -7138
rect 56496 -7230 56506 -6980
rect 57016 -7230 57026 -6980
rect 56496 -7235 57026 -7230
rect 55955 -7298 56200 -7288
rect 53510 -7378 53645 -7368
rect 55275 -7318 55490 -7308
rect 53045 -7558 53255 -7548
rect 20794 -7875 20888 -7870
rect 20794 -11629 20804 -7875
rect 20878 -11629 20888 -7875
rect 24600 -8700 47900 -8600
rect 24600 -9400 24700 -8700
rect 25700 -9400 46700 -8700
rect 47800 -9400 47900 -8700
rect 53045 -9308 53050 -7558
rect 53250 -9308 53255 -7558
rect 53045 -9318 53255 -9308
rect 24600 -9500 47900 -9400
rect 53510 -9518 53630 -7378
rect 55275 -7408 55280 -7318
rect 55400 -7408 55490 -7318
rect 56060 -7338 56200 -7298
rect 56060 -7348 56220 -7338
rect 55275 -7418 55490 -7408
rect 55220 -7658 55325 -7648
rect 55220 -7828 55230 -7658
rect 55320 -7828 55325 -7658
rect 55220 -7838 55325 -7828
rect 55015 -8448 55125 -8438
rect 55015 -8528 55020 -8448
rect 55120 -8528 55125 -8448
rect 55015 -8538 55125 -8528
rect 55220 -9138 55310 -7838
rect 55215 -9148 55315 -9138
rect 55215 -9318 55220 -9148
rect 55310 -9238 55315 -9148
rect 55400 -9148 55490 -7418
rect 55875 -7418 55990 -7408
rect 55875 -7458 55880 -7418
rect 55870 -7498 55880 -7458
rect 55970 -7498 55990 -7418
rect 55870 -7578 55990 -7498
rect 56060 -7518 56220 -7508
rect 55590 -7668 55720 -7658
rect 55590 -7798 55600 -7668
rect 55710 -7798 55720 -7668
rect 55400 -9158 55510 -9148
rect 55310 -9318 55320 -9238
rect 55400 -9318 55410 -9158
rect 55215 -9328 55320 -9318
rect 53505 -9528 53635 -9518
rect 53505 -9648 53510 -9528
rect 53630 -9648 53635 -9528
rect 53505 -9658 53635 -9648
rect 55220 -9808 55320 -9328
rect 55405 -9328 55410 -9318
rect 55500 -9328 55510 -9158
rect 55405 -9338 55510 -9328
rect 55590 -9588 55720 -7798
rect 55870 -7958 55980 -7578
rect 57093 -7964 57373 -7954
rect 56475 -7988 56555 -7978
rect 56470 -8048 56480 -7988
rect 56550 -8048 56555 -7988
rect 56470 -8058 56555 -8048
rect 55870 -8438 55980 -8068
rect 55870 -8528 55880 -8438
rect 55970 -8528 55980 -8438
rect 55870 -8928 55980 -8528
rect 56470 -8428 56550 -8058
rect 57093 -8104 57098 -7964
rect 57368 -8104 57373 -7964
rect 57093 -8114 57373 -8104
rect 57760 -8420 58280 -3140
rect 58516 -3060 58796 -2990
rect 58516 -3260 58556 -3060
rect 58756 -3260 58796 -3060
rect 59066 -3010 59176 -2510
rect 59266 -2620 59366 -2190
rect 59536 -2090 59616 -1900
rect 59536 -2150 59546 -2090
rect 59606 -2150 59616 -2090
rect 59536 -2210 59616 -2150
rect 59536 -2270 59546 -2210
rect 59606 -2270 59616 -2210
rect 59536 -2280 59616 -2270
rect 59266 -2630 59376 -2620
rect 59266 -2720 59286 -2630
rect 59366 -2720 59376 -2630
rect 59736 -2650 59796 -1900
rect 59856 -2140 59976 -2130
rect 59856 -2230 59866 -2140
rect 59966 -2230 59976 -2140
rect 59856 -2240 59976 -2230
rect 60036 -2320 60136 -1690
rect 61026 -1720 61136 -1710
rect 61026 -1850 61056 -1720
rect 61126 -1850 61136 -1720
rect 60436 -2120 60536 -2110
rect 60436 -2220 60446 -2120
rect 60526 -2220 60536 -2120
rect 60436 -2230 60536 -2220
rect 60036 -2400 60046 -2320
rect 60126 -2400 60136 -2320
rect 60036 -2410 60136 -2400
rect 60546 -2410 60636 -2400
rect 60386 -2490 60556 -2410
rect 60626 -2490 60636 -2410
rect 59966 -2500 60326 -2490
rect 59966 -2570 59976 -2500
rect 60316 -2570 60326 -2500
rect 60546 -2510 60636 -2490
rect 59966 -2580 60326 -2570
rect 59566 -2670 59796 -2650
rect 59566 -2680 59576 -2670
rect 59266 -2730 59376 -2720
rect 59516 -2730 59576 -2680
rect 59636 -2730 59796 -2670
rect 59266 -2840 59366 -2730
rect 59266 -2930 59286 -2840
rect 59356 -2930 59366 -2840
rect 59266 -2960 59366 -2930
rect 59516 -2740 59796 -2730
rect 59066 -3080 59076 -3010
rect 59166 -3080 59176 -3010
rect 59066 -3090 59176 -3080
rect 59306 -3030 59386 -3020
rect 59306 -3090 59316 -3030
rect 59376 -3090 59386 -3030
rect 59516 -3070 59596 -2740
rect 60286 -2750 60476 -2740
rect 59906 -2780 60016 -2770
rect 59906 -2960 59916 -2780
rect 60006 -2960 60016 -2780
rect 59906 -2970 60016 -2960
rect 60286 -2890 60306 -2750
rect 60456 -2890 60476 -2750
rect 60286 -2900 60476 -2890
rect 58516 -3340 58796 -3260
rect 59066 -3170 59176 -3160
rect 59066 -3240 59076 -3170
rect 59166 -3240 59176 -3170
rect 59066 -3740 59176 -3240
rect 59306 -3290 59386 -3090
rect 60076 -3080 60196 -3040
rect 60076 -3240 60096 -3080
rect 60176 -3240 60196 -3080
rect 60076 -3280 60196 -3240
rect 59066 -3800 59076 -3740
rect 59166 -3800 59176 -3740
rect 59066 -3810 59176 -3800
rect 59236 -3320 59386 -3290
rect 59236 -3410 59266 -3320
rect 59366 -3410 59386 -3320
rect 59236 -3430 59386 -3410
rect 59906 -3290 60016 -3280
rect 59236 -3560 59376 -3430
rect 59906 -3480 59916 -3290
rect 60006 -3480 60016 -3290
rect 59906 -3490 60016 -3480
rect 60286 -3310 60376 -2900
rect 60556 -3300 60626 -2510
rect 61026 -2820 61136 -1850
rect 61196 -2520 61356 -2510
rect 61196 -2700 61206 -2520
rect 61346 -2700 61356 -2520
rect 61196 -2710 61356 -2700
rect 61026 -2930 61036 -2820
rect 61126 -2930 61136 -2820
rect 61026 -2940 61136 -2930
rect 61246 -3050 61366 -3040
rect 61246 -3060 61276 -3050
rect 61246 -3260 61256 -3060
rect 61356 -3260 61366 -3050
rect 61246 -3270 61366 -3260
rect 60466 -3310 60626 -3300
rect 60286 -3370 60406 -3310
rect 60466 -3370 60476 -3310
rect 60536 -3370 60626 -3310
rect 59236 -3650 59266 -3560
rect 59366 -3650 59376 -3560
rect 59236 -3700 59376 -3650
rect 59506 -3510 59606 -3500
rect 59506 -3580 59516 -3510
rect 59596 -3580 59606 -3510
rect 59506 -3590 59606 -3580
rect 59236 -3720 59386 -3700
rect 59236 -3780 59316 -3720
rect 59376 -3780 59386 -3720
rect 58396 -4350 58896 -3850
rect 59236 -4030 59386 -3780
rect 59006 -4100 59086 -4080
rect 59236 -4090 59256 -4030
rect 59366 -4090 59386 -4030
rect 59236 -4100 59386 -4090
rect 59506 -3980 59596 -3590
rect 59986 -3720 60116 -3710
rect 59986 -3780 59996 -3720
rect 60106 -3780 60116 -3720
rect 59506 -3990 59616 -3980
rect 59506 -4060 59546 -3990
rect 59606 -4060 59616 -3990
rect 59006 -4160 59016 -4100
rect 59076 -4160 59086 -4100
rect 59006 -4350 59086 -4160
rect 59506 -4110 59616 -4060
rect 59506 -4170 59546 -4110
rect 59606 -4170 59616 -4110
rect 59796 -4010 59926 -4000
rect 59796 -4120 59806 -4010
rect 59916 -4120 59926 -4010
rect 59796 -4130 59926 -4120
rect 59006 -4440 59126 -4350
rect 59006 -4510 59016 -4440
rect 59076 -4510 59126 -4440
rect 59006 -4590 59126 -4510
rect 59506 -4440 59616 -4170
rect 59506 -4510 59546 -4440
rect 59606 -4510 59616 -4440
rect 59506 -4520 59616 -4510
rect 59986 -4590 60116 -3780
rect 60286 -4270 60376 -3370
rect 60466 -3380 60626 -3370
rect 61486 -3370 61726 -3340
rect 61486 -3420 61496 -3370
rect 61326 -3430 61496 -3420
rect 61326 -3550 61336 -3430
rect 61196 -3560 61336 -3550
rect 61456 -3540 61496 -3430
rect 61696 -3540 61726 -3370
rect 61456 -3560 61726 -3540
rect 61196 -3570 61726 -3560
rect 61196 -3740 61426 -3570
rect 60436 -4030 60536 -4010
rect 60436 -4150 60446 -4030
rect 60526 -4150 60536 -4030
rect 60436 -4160 60536 -4150
rect 60256 -4400 60416 -4270
rect 60256 -4530 60266 -4400
rect 60406 -4530 60416 -4400
rect 60256 -4550 60416 -4530
rect 58956 -4600 59156 -4590
rect 58956 -4780 58966 -4600
rect 59146 -4780 59156 -4600
rect 59986 -4700 59996 -4590
rect 60106 -4700 60116 -4590
rect 59986 -4710 60116 -4700
rect 58956 -4790 59156 -4780
rect 59600 -4900 68700 -4800
rect 59600 -5200 59700 -4900
rect 60400 -5200 68100 -4900
rect 68600 -5200 68700 -4900
rect 59600 -5300 68700 -5200
rect 58946 -6870 59146 -6850
rect 58946 -7030 58966 -6870
rect 59126 -7030 59146 -6870
rect 58946 -7050 59146 -7030
rect 59316 -6910 59426 -6850
rect 59316 -7050 59336 -6910
rect 59416 -7050 59426 -6910
rect 58956 -7130 59136 -7050
rect 58956 -7240 58996 -7130
rect 59106 -7240 59136 -7130
rect 58396 -7330 58896 -7240
rect 58956 -7300 59136 -7240
rect 59316 -7280 59426 -7050
rect 59946 -6920 60386 -6800
rect 59946 -7040 60046 -6920
rect 60126 -7040 60386 -6920
rect 59946 -7090 60386 -7040
rect 58396 -7690 58486 -7330
rect 58816 -7690 58896 -7330
rect 58996 -7600 59086 -7300
rect 58996 -7660 59006 -7600
rect 59066 -7660 59086 -7600
rect 58996 -7670 59086 -7660
rect 59266 -7330 59426 -7280
rect 59506 -7140 59796 -7100
rect 59506 -7240 59516 -7140
rect 59616 -7240 59796 -7140
rect 59506 -7300 59796 -7240
rect 59266 -7530 59366 -7330
rect 59266 -7590 59286 -7530
rect 59346 -7590 59366 -7530
rect 58396 -7800 58896 -7690
rect 59066 -7840 59176 -7830
rect 59066 -7910 59076 -7840
rect 59166 -7910 59176 -7840
rect 56470 -8438 56555 -8428
rect 56470 -8528 56480 -8438
rect 56550 -8528 56555 -8438
rect 56470 -8538 56555 -8528
rect 56470 -8918 56550 -8538
rect 57760 -8540 57800 -8420
rect 58240 -8540 58280 -8420
rect 57093 -8874 57373 -8864
rect 56470 -8928 56555 -8918
rect 56470 -8978 56480 -8928
rect 56475 -8988 56480 -8978
rect 56550 -8988 56555 -8928
rect 56475 -8998 56555 -8988
rect 57093 -9014 57098 -8874
rect 57368 -9014 57373 -8874
rect 57093 -9024 57373 -9014
rect 55870 -9478 55980 -9038
rect 55870 -9518 55880 -9478
rect 55875 -9558 55880 -9518
rect 55970 -9518 55980 -9478
rect 56060 -9468 56220 -9458
rect 55970 -9558 55975 -9518
rect 55875 -9568 55975 -9558
rect 55590 -9678 55620 -9588
rect 55710 -9678 55720 -9588
rect 56060 -9638 56220 -9628
rect 56060 -9648 56200 -9638
rect 55590 -9688 55720 -9678
rect 56015 -9658 56200 -9648
rect 56015 -9808 56020 -9658
rect 56080 -9808 56200 -9658
rect 56644 -9668 57008 -9663
rect 55215 -9818 55325 -9808
rect 56015 -9818 56085 -9808
rect 55215 -9918 55220 -9818
rect 55320 -9918 55325 -9818
rect 56644 -9886 56654 -9668
rect 56998 -9886 57008 -9668
rect 56644 -9891 57008 -9886
rect 55215 -9928 55325 -9918
rect 55315 -10128 55475 -10118
rect 55315 -10268 55320 -10128
rect 55470 -10268 55475 -10128
rect 55315 -10278 55475 -10268
rect 20794 -11634 20888 -11629
rect 27000 -10600 34600 -10400
rect 20801 -11997 20877 -11634
rect 20790 -12002 20890 -11997
rect 20790 -12092 20800 -12002
rect 20880 -12092 20890 -12002
rect 20790 -12097 20890 -12092
rect 20801 -12232 20877 -12097
rect 20800 -12346 20880 -12232
rect 20570 -12352 20650 -12347
rect 20570 -13042 20580 -12352
rect 20640 -13042 20650 -12352
rect 20570 -13047 20650 -13042
rect 20791 -12351 20880 -12346
rect 20791 -13041 20801 -12351
rect 20861 -12402 20880 -12351
rect 20861 -13041 20877 -12402
rect 27000 -13000 27200 -10600
rect 34400 -13000 34600 -10600
rect 37500 -10700 56100 -10600
rect 37500 -11100 37600 -10700
rect 38100 -11100 55500 -10700
rect 56000 -11100 56100 -10700
rect 37500 -11200 56100 -11100
rect 51400 -11660 55800 -11600
rect 51400 -11700 55380 -11660
rect 51400 -11900 51500 -11700
rect 52500 -11900 55380 -11700
rect 51400 -11980 55380 -11900
rect 55740 -11980 55800 -11660
rect 51400 -12000 55800 -11980
rect 55320 -12040 55800 -12000
rect 47680 -12220 48100 -12200
rect 47680 -12640 47700 -12220
rect 48080 -12320 48100 -12220
rect 48080 -12340 53800 -12320
rect 48080 -12540 53480 -12340
rect 53780 -12540 53800 -12340
rect 56496 -12380 57026 -12375
rect 48080 -12560 53800 -12540
rect 55955 -12538 56045 -12528
rect 48080 -12640 48100 -12560
rect 47680 -12660 48100 -12640
rect 53515 -12658 53645 -12648
rect 53510 -12768 53520 -12658
rect 53640 -12768 53645 -12658
rect 55955 -12688 55960 -12538
rect 56040 -12688 56200 -12538
rect 56496 -12630 56506 -12380
rect 57016 -12630 57026 -12380
rect 56496 -12635 57026 -12630
rect 55955 -12698 56200 -12688
rect 53510 -12778 53645 -12768
rect 55275 -12718 55490 -12708
rect 20791 -13046 20871 -13041
rect 20570 -13307 20640 -13047
rect 27000 -13200 34600 -13000
rect 53045 -12958 53255 -12948
rect 20560 -13312 20680 -13307
rect 20560 -13392 20570 -13312
rect 20670 -13392 20680 -13312
rect 20560 -13397 20680 -13392
rect 53045 -14708 53050 -12958
rect 53250 -14708 53255 -12958
rect 53045 -14718 53255 -14708
rect 53510 -14918 53630 -12778
rect 55275 -12808 55280 -12718
rect 55400 -12808 55490 -12718
rect 56060 -12738 56200 -12698
rect 56060 -12748 56220 -12738
rect 55275 -12818 55490 -12808
rect 55220 -13058 55325 -13048
rect 55220 -13228 55230 -13058
rect 55320 -13228 55325 -13058
rect 55220 -13238 55325 -13228
rect 55015 -13848 55125 -13838
rect 55015 -13928 55020 -13848
rect 55120 -13928 55125 -13848
rect 55015 -13938 55125 -13928
rect 55220 -14538 55310 -13238
rect 55215 -14548 55315 -14538
rect 55215 -14718 55220 -14548
rect 55310 -14638 55315 -14548
rect 55400 -14548 55490 -12818
rect 55875 -12818 55990 -12808
rect 55875 -12858 55880 -12818
rect 55870 -12898 55880 -12858
rect 55970 -12898 55990 -12818
rect 55870 -12978 55990 -12898
rect 56060 -12918 56220 -12908
rect 55590 -13068 55720 -13058
rect 55590 -13198 55600 -13068
rect 55710 -13198 55720 -13068
rect 55400 -14558 55510 -14548
rect 55310 -14718 55320 -14638
rect 55400 -14718 55410 -14558
rect 55215 -14728 55320 -14718
rect 53505 -14928 53635 -14918
rect 53505 -15048 53510 -14928
rect 53630 -15048 53635 -14928
rect 53505 -15058 53635 -15048
rect 55220 -15208 55320 -14728
rect 55405 -14728 55410 -14718
rect 55500 -14728 55510 -14558
rect 55405 -14738 55510 -14728
rect 55590 -14988 55720 -13198
rect 55870 -13358 55980 -12978
rect 57093 -13364 57373 -13354
rect 56475 -13388 56555 -13378
rect 56470 -13448 56480 -13388
rect 56550 -13448 56555 -13388
rect 56470 -13458 56555 -13448
rect 55870 -13838 55980 -13468
rect 55870 -13928 55880 -13838
rect 55970 -13928 55980 -13838
rect 55870 -14328 55980 -13928
rect 56470 -13828 56550 -13458
rect 57093 -13504 57098 -13364
rect 57368 -13504 57373 -13364
rect 57093 -13514 57373 -13504
rect 57760 -13820 58280 -8540
rect 58516 -8460 58796 -8390
rect 58516 -8660 58556 -8460
rect 58756 -8660 58796 -8460
rect 59066 -8410 59176 -7910
rect 59266 -8020 59366 -7590
rect 59536 -7490 59616 -7300
rect 59536 -7550 59546 -7490
rect 59606 -7550 59616 -7490
rect 59536 -7610 59616 -7550
rect 59536 -7670 59546 -7610
rect 59606 -7670 59616 -7610
rect 59536 -7680 59616 -7670
rect 59266 -8030 59376 -8020
rect 59266 -8120 59286 -8030
rect 59366 -8120 59376 -8030
rect 59736 -8050 59796 -7300
rect 59856 -7540 59976 -7530
rect 59856 -7630 59866 -7540
rect 59966 -7630 59976 -7540
rect 59856 -7640 59976 -7630
rect 60036 -7720 60136 -7090
rect 61026 -7120 61136 -7110
rect 61026 -7250 61056 -7120
rect 61126 -7250 61136 -7120
rect 60436 -7520 60536 -7510
rect 60436 -7620 60446 -7520
rect 60526 -7620 60536 -7520
rect 60436 -7630 60536 -7620
rect 60036 -7800 60046 -7720
rect 60126 -7800 60136 -7720
rect 60036 -7810 60136 -7800
rect 60546 -7810 60636 -7800
rect 60386 -7890 60556 -7810
rect 60626 -7890 60636 -7810
rect 59966 -7900 60326 -7890
rect 59966 -7970 59976 -7900
rect 60316 -7970 60326 -7900
rect 60546 -7910 60636 -7890
rect 59966 -7980 60326 -7970
rect 59566 -8070 59796 -8050
rect 59566 -8080 59576 -8070
rect 59266 -8130 59376 -8120
rect 59516 -8130 59576 -8080
rect 59636 -8130 59796 -8070
rect 59266 -8240 59366 -8130
rect 59266 -8330 59286 -8240
rect 59356 -8330 59366 -8240
rect 59266 -8360 59366 -8330
rect 59516 -8140 59796 -8130
rect 59066 -8480 59076 -8410
rect 59166 -8480 59176 -8410
rect 59066 -8490 59176 -8480
rect 59306 -8430 59386 -8420
rect 59306 -8490 59316 -8430
rect 59376 -8490 59386 -8430
rect 59516 -8470 59596 -8140
rect 60286 -8150 60476 -8140
rect 59906 -8180 60016 -8170
rect 59906 -8360 59916 -8180
rect 60006 -8360 60016 -8180
rect 59906 -8370 60016 -8360
rect 60286 -8290 60306 -8150
rect 60456 -8290 60476 -8150
rect 60286 -8300 60476 -8290
rect 58516 -8740 58796 -8660
rect 59066 -8570 59176 -8560
rect 59066 -8640 59076 -8570
rect 59166 -8640 59176 -8570
rect 59066 -9140 59176 -8640
rect 59306 -8690 59386 -8490
rect 60076 -8480 60196 -8440
rect 60076 -8640 60096 -8480
rect 60176 -8640 60196 -8480
rect 60076 -8680 60196 -8640
rect 59066 -9200 59076 -9140
rect 59166 -9200 59176 -9140
rect 59066 -9210 59176 -9200
rect 59236 -8720 59386 -8690
rect 59236 -8810 59266 -8720
rect 59366 -8810 59386 -8720
rect 59236 -8830 59386 -8810
rect 59906 -8690 60016 -8680
rect 59236 -8960 59376 -8830
rect 59906 -8880 59916 -8690
rect 60006 -8880 60016 -8690
rect 59906 -8890 60016 -8880
rect 60286 -8710 60376 -8300
rect 60556 -8700 60626 -7910
rect 61026 -8220 61136 -7250
rect 61196 -7920 61356 -7910
rect 61196 -8100 61206 -7920
rect 61346 -8100 61356 -7920
rect 61196 -8110 61356 -8100
rect 61026 -8330 61036 -8220
rect 61126 -8330 61136 -8220
rect 61026 -8340 61136 -8330
rect 61246 -8450 61366 -8440
rect 61246 -8460 61276 -8450
rect 61246 -8660 61256 -8460
rect 61356 -8660 61366 -8450
rect 61246 -8670 61366 -8660
rect 60466 -8710 60626 -8700
rect 60286 -8770 60406 -8710
rect 60466 -8770 60476 -8710
rect 60536 -8770 60626 -8710
rect 59236 -9050 59266 -8960
rect 59366 -9050 59376 -8960
rect 59236 -9100 59376 -9050
rect 59506 -8910 59606 -8900
rect 59506 -8980 59516 -8910
rect 59596 -8980 59606 -8910
rect 59506 -8990 59606 -8980
rect 59236 -9120 59386 -9100
rect 59236 -9180 59316 -9120
rect 59376 -9180 59386 -9120
rect 58396 -9750 58896 -9250
rect 59236 -9430 59386 -9180
rect 59006 -9500 59086 -9480
rect 59236 -9490 59256 -9430
rect 59366 -9490 59386 -9430
rect 59236 -9500 59386 -9490
rect 59506 -9380 59596 -8990
rect 59986 -9120 60116 -9110
rect 59986 -9180 59996 -9120
rect 60106 -9180 60116 -9120
rect 59506 -9390 59616 -9380
rect 59506 -9460 59546 -9390
rect 59606 -9460 59616 -9390
rect 59006 -9560 59016 -9500
rect 59076 -9560 59086 -9500
rect 59006 -9750 59086 -9560
rect 59506 -9510 59616 -9460
rect 59506 -9570 59546 -9510
rect 59606 -9570 59616 -9510
rect 59796 -9410 59926 -9400
rect 59796 -9520 59806 -9410
rect 59916 -9520 59926 -9410
rect 59796 -9530 59926 -9520
rect 59006 -9840 59126 -9750
rect 59006 -9910 59016 -9840
rect 59076 -9910 59126 -9840
rect 59006 -9990 59126 -9910
rect 59506 -9840 59616 -9570
rect 59506 -9910 59546 -9840
rect 59606 -9910 59616 -9840
rect 59506 -9920 59616 -9910
rect 59986 -9990 60116 -9180
rect 60286 -9670 60376 -8770
rect 60466 -8780 60626 -8770
rect 61486 -8770 61726 -8740
rect 61486 -8820 61496 -8770
rect 61326 -8830 61496 -8820
rect 61326 -8950 61336 -8830
rect 61196 -8960 61336 -8950
rect 61456 -8940 61496 -8830
rect 61696 -8940 61726 -8770
rect 61456 -8960 61726 -8940
rect 61196 -8970 61726 -8960
rect 61196 -9140 61426 -8970
rect 60436 -9430 60536 -9410
rect 60436 -9550 60446 -9430
rect 60526 -9550 60536 -9430
rect 60436 -9560 60536 -9550
rect 60256 -9800 60416 -9670
rect 60256 -9930 60266 -9800
rect 60406 -9930 60416 -9800
rect 60256 -9950 60416 -9930
rect 58956 -10000 59156 -9990
rect 58956 -10180 58966 -10000
rect 59146 -10180 59156 -10000
rect 59986 -10100 59996 -9990
rect 60106 -10100 60116 -9990
rect 59986 -10110 60116 -10100
rect 58956 -10190 59156 -10180
rect 59600 -10300 67500 -10200
rect 59600 -10700 59700 -10300
rect 60400 -10700 66900 -10300
rect 67400 -10700 67500 -10300
rect 59600 -10800 67500 -10700
rect 58946 -12270 59146 -12250
rect 58946 -12430 58966 -12270
rect 59126 -12430 59146 -12270
rect 58946 -12450 59146 -12430
rect 59316 -12310 59426 -12250
rect 59316 -12450 59336 -12310
rect 59416 -12450 59426 -12310
rect 58956 -12530 59136 -12450
rect 58956 -12640 58996 -12530
rect 59106 -12640 59136 -12530
rect 58396 -12730 58896 -12640
rect 58956 -12700 59136 -12640
rect 59316 -12680 59426 -12450
rect 59946 -12320 60386 -12200
rect 59946 -12440 60046 -12320
rect 60126 -12440 60386 -12320
rect 59946 -12490 60386 -12440
rect 58396 -13090 58486 -12730
rect 58816 -13090 58896 -12730
rect 58996 -13000 59086 -12700
rect 58996 -13060 59006 -13000
rect 59066 -13060 59086 -13000
rect 58996 -13070 59086 -13060
rect 59266 -12730 59426 -12680
rect 59506 -12540 59796 -12500
rect 59506 -12640 59516 -12540
rect 59616 -12640 59796 -12540
rect 59506 -12700 59796 -12640
rect 59266 -12930 59366 -12730
rect 59266 -12990 59286 -12930
rect 59346 -12990 59366 -12930
rect 58396 -13200 58896 -13090
rect 59066 -13240 59176 -13230
rect 59066 -13310 59076 -13240
rect 59166 -13310 59176 -13240
rect 56470 -13838 56555 -13828
rect 56470 -13928 56480 -13838
rect 56550 -13928 56555 -13838
rect 56470 -13938 56555 -13928
rect 56470 -14318 56550 -13938
rect 57760 -13940 57800 -13820
rect 58240 -13940 58280 -13820
rect 57093 -14274 57373 -14264
rect 56470 -14328 56555 -14318
rect 56470 -14378 56480 -14328
rect 56475 -14388 56480 -14378
rect 56550 -14388 56555 -14328
rect 56475 -14398 56555 -14388
rect 57093 -14414 57098 -14274
rect 57368 -14414 57373 -14274
rect 57093 -14424 57373 -14414
rect 55870 -14878 55980 -14438
rect 55870 -14918 55880 -14878
rect 55875 -14958 55880 -14918
rect 55970 -14918 55980 -14878
rect 56060 -14868 56220 -14858
rect 55970 -14958 55975 -14918
rect 55875 -14968 55975 -14958
rect 55590 -15078 55620 -14988
rect 55710 -15078 55720 -14988
rect 56060 -15038 56220 -15028
rect 56060 -15048 56200 -15038
rect 55590 -15088 55720 -15078
rect 56015 -15058 56200 -15048
rect 56015 -15208 56020 -15058
rect 56080 -15208 56200 -15058
rect 56644 -15068 57008 -15063
rect 55215 -15218 55325 -15208
rect 56015 -15218 56085 -15208
rect 55215 -15318 55220 -15218
rect 55320 -15318 55325 -15218
rect 56644 -15286 56654 -15068
rect 56998 -15286 57008 -15068
rect 56644 -15291 57008 -15286
rect 55215 -15328 55325 -15318
rect 55315 -15528 55475 -15518
rect 55315 -15668 55320 -15528
rect 55470 -15668 55475 -15528
rect 55315 -15678 55475 -15668
rect 38400 -16000 39100 -15900
rect 38400 -16600 38500 -16000
rect 39000 -16100 56100 -16000
rect 39000 -16500 55500 -16100
rect 56000 -16500 56100 -16100
rect 39000 -16600 56100 -16500
rect 38400 -16700 39100 -16600
rect 51400 -17100 55800 -17000
rect 51400 -17300 51500 -17100
rect 52500 -17300 55400 -17100
rect 51400 -17400 55400 -17300
rect 55700 -17400 55800 -17100
rect 55300 -17500 55800 -17400
rect 47620 -17620 48100 -17600
rect 47620 -18100 47640 -17620
rect 48080 -17720 48100 -17620
rect 48080 -17740 53800 -17720
rect 48080 -17940 53500 -17740
rect 53780 -17940 53800 -17740
rect 56496 -17780 57026 -17775
rect 48080 -17960 53800 -17940
rect 55955 -17938 56045 -17928
rect 48080 -18100 48100 -17960
rect 53515 -18058 53645 -18048
rect 47620 -18120 48100 -18100
rect 53510 -18168 53520 -18058
rect 53640 -18168 53645 -18058
rect 55955 -18088 55960 -17938
rect 56040 -18088 56200 -17938
rect 56496 -18030 56506 -17780
rect 57016 -18030 57026 -17780
rect 56496 -18035 57026 -18030
rect 55955 -18098 56200 -18088
rect 53510 -18178 53645 -18168
rect 55275 -18118 55490 -18108
rect 53045 -18358 53255 -18348
rect 53045 -20108 53050 -18358
rect 53250 -20108 53255 -18358
rect 53045 -20118 53255 -20108
rect 53510 -20318 53630 -18178
rect 55275 -18208 55280 -18118
rect 55400 -18208 55490 -18118
rect 56060 -18138 56200 -18098
rect 56060 -18148 56220 -18138
rect 55275 -18218 55490 -18208
rect 55220 -18458 55325 -18448
rect 55220 -18628 55230 -18458
rect 55320 -18628 55325 -18458
rect 55220 -18638 55325 -18628
rect 55015 -19248 55125 -19238
rect 55015 -19328 55020 -19248
rect 55120 -19328 55125 -19248
rect 55015 -19338 55125 -19328
rect 55220 -19938 55310 -18638
rect 55215 -19948 55315 -19938
rect 55215 -20118 55220 -19948
rect 55310 -20038 55315 -19948
rect 55400 -19948 55490 -18218
rect 55875 -18218 55990 -18208
rect 55875 -18258 55880 -18218
rect 55870 -18298 55880 -18258
rect 55970 -18298 55990 -18218
rect 55870 -18378 55990 -18298
rect 56060 -18318 56220 -18308
rect 55590 -18468 55720 -18458
rect 55590 -18598 55600 -18468
rect 55710 -18598 55720 -18468
rect 55400 -19958 55510 -19948
rect 55310 -20118 55320 -20038
rect 55400 -20118 55410 -19958
rect 55215 -20128 55320 -20118
rect 53505 -20328 53635 -20318
rect 53505 -20448 53510 -20328
rect 53630 -20448 53635 -20328
rect 53505 -20458 53635 -20448
rect 55220 -20608 55320 -20128
rect 55405 -20128 55410 -20118
rect 55500 -20128 55510 -19958
rect 55405 -20138 55510 -20128
rect 55590 -20388 55720 -18598
rect 55870 -18758 55980 -18378
rect 57093 -18764 57373 -18754
rect 56475 -18788 56555 -18778
rect 56470 -18848 56480 -18788
rect 56550 -18848 56555 -18788
rect 56470 -18858 56555 -18848
rect 55870 -19238 55980 -18868
rect 55870 -19328 55880 -19238
rect 55970 -19328 55980 -19238
rect 55870 -19728 55980 -19328
rect 56470 -19228 56550 -18858
rect 57093 -18904 57098 -18764
rect 57368 -18904 57373 -18764
rect 57093 -18914 57373 -18904
rect 57760 -19220 58280 -13940
rect 58516 -13860 58796 -13790
rect 58516 -14060 58556 -13860
rect 58756 -14060 58796 -13860
rect 59066 -13810 59176 -13310
rect 59266 -13420 59366 -12990
rect 59536 -12890 59616 -12700
rect 59536 -12950 59546 -12890
rect 59606 -12950 59616 -12890
rect 59536 -13010 59616 -12950
rect 59536 -13070 59546 -13010
rect 59606 -13070 59616 -13010
rect 59536 -13080 59616 -13070
rect 59266 -13430 59376 -13420
rect 59266 -13520 59286 -13430
rect 59366 -13520 59376 -13430
rect 59736 -13450 59796 -12700
rect 59856 -12940 59976 -12930
rect 59856 -13030 59866 -12940
rect 59966 -13030 59976 -12940
rect 59856 -13040 59976 -13030
rect 60036 -13120 60136 -12490
rect 61026 -12520 61136 -12510
rect 61026 -12650 61056 -12520
rect 61126 -12650 61136 -12520
rect 60436 -12920 60536 -12910
rect 60436 -13020 60446 -12920
rect 60526 -13020 60536 -12920
rect 60436 -13030 60536 -13020
rect 60036 -13200 60046 -13120
rect 60126 -13200 60136 -13120
rect 60036 -13210 60136 -13200
rect 60546 -13210 60636 -13200
rect 60386 -13290 60556 -13210
rect 60626 -13290 60636 -13210
rect 59966 -13300 60326 -13290
rect 59966 -13370 59976 -13300
rect 60316 -13370 60326 -13300
rect 60546 -13310 60636 -13290
rect 59966 -13380 60326 -13370
rect 59566 -13470 59796 -13450
rect 59566 -13480 59576 -13470
rect 59266 -13530 59376 -13520
rect 59516 -13530 59576 -13480
rect 59636 -13530 59796 -13470
rect 59266 -13640 59366 -13530
rect 59266 -13730 59286 -13640
rect 59356 -13730 59366 -13640
rect 59266 -13760 59366 -13730
rect 59516 -13540 59796 -13530
rect 59066 -13880 59076 -13810
rect 59166 -13880 59176 -13810
rect 59066 -13890 59176 -13880
rect 59306 -13830 59386 -13820
rect 59306 -13890 59316 -13830
rect 59376 -13890 59386 -13830
rect 59516 -13870 59596 -13540
rect 60286 -13550 60476 -13540
rect 59906 -13580 60016 -13570
rect 59906 -13760 59916 -13580
rect 60006 -13760 60016 -13580
rect 59906 -13770 60016 -13760
rect 60286 -13690 60306 -13550
rect 60456 -13690 60476 -13550
rect 60286 -13700 60476 -13690
rect 58516 -14140 58796 -14060
rect 59066 -13970 59176 -13960
rect 59066 -14040 59076 -13970
rect 59166 -14040 59176 -13970
rect 59066 -14540 59176 -14040
rect 59306 -14090 59386 -13890
rect 60076 -13880 60196 -13840
rect 60076 -14040 60096 -13880
rect 60176 -14040 60196 -13880
rect 60076 -14080 60196 -14040
rect 59066 -14600 59076 -14540
rect 59166 -14600 59176 -14540
rect 59066 -14610 59176 -14600
rect 59236 -14120 59386 -14090
rect 59236 -14210 59266 -14120
rect 59366 -14210 59386 -14120
rect 59236 -14230 59386 -14210
rect 59906 -14090 60016 -14080
rect 59236 -14360 59376 -14230
rect 59906 -14280 59916 -14090
rect 60006 -14280 60016 -14090
rect 59906 -14290 60016 -14280
rect 60286 -14110 60376 -13700
rect 60556 -14100 60626 -13310
rect 61026 -13620 61136 -12650
rect 61196 -13320 61356 -13310
rect 61196 -13500 61206 -13320
rect 61346 -13500 61356 -13320
rect 61196 -13510 61356 -13500
rect 61026 -13730 61036 -13620
rect 61126 -13730 61136 -13620
rect 61026 -13740 61136 -13730
rect 61246 -13850 61366 -13840
rect 61246 -13860 61276 -13850
rect 61246 -14060 61256 -13860
rect 61356 -14060 61366 -13850
rect 61246 -14070 61366 -14060
rect 60466 -14110 60626 -14100
rect 60286 -14170 60406 -14110
rect 60466 -14170 60476 -14110
rect 60536 -14170 60626 -14110
rect 59236 -14450 59266 -14360
rect 59366 -14450 59376 -14360
rect 59236 -14500 59376 -14450
rect 59506 -14310 59606 -14300
rect 59506 -14380 59516 -14310
rect 59596 -14380 59606 -14310
rect 59506 -14390 59606 -14380
rect 59236 -14520 59386 -14500
rect 59236 -14580 59316 -14520
rect 59376 -14580 59386 -14520
rect 58396 -15150 58896 -14650
rect 59236 -14830 59386 -14580
rect 59006 -14900 59086 -14880
rect 59236 -14890 59256 -14830
rect 59366 -14890 59386 -14830
rect 59236 -14900 59386 -14890
rect 59506 -14780 59596 -14390
rect 59986 -14520 60116 -14510
rect 59986 -14580 59996 -14520
rect 60106 -14580 60116 -14520
rect 59506 -14790 59616 -14780
rect 59506 -14860 59546 -14790
rect 59606 -14860 59616 -14790
rect 59006 -14960 59016 -14900
rect 59076 -14960 59086 -14900
rect 59006 -15150 59086 -14960
rect 59506 -14910 59616 -14860
rect 59506 -14970 59546 -14910
rect 59606 -14970 59616 -14910
rect 59796 -14810 59926 -14800
rect 59796 -14920 59806 -14810
rect 59916 -14920 59926 -14810
rect 59796 -14930 59926 -14920
rect 59006 -15240 59126 -15150
rect 59006 -15310 59016 -15240
rect 59076 -15310 59126 -15240
rect 59006 -15390 59126 -15310
rect 59506 -15240 59616 -14970
rect 59506 -15310 59546 -15240
rect 59606 -15310 59616 -15240
rect 59506 -15320 59616 -15310
rect 59986 -15390 60116 -14580
rect 60286 -15070 60376 -14170
rect 60466 -14180 60626 -14170
rect 61486 -14170 61726 -14140
rect 61486 -14220 61496 -14170
rect 61326 -14230 61496 -14220
rect 61326 -14350 61336 -14230
rect 61196 -14360 61336 -14350
rect 61456 -14340 61496 -14230
rect 61696 -14340 61726 -14170
rect 61456 -14360 61726 -14340
rect 61196 -14370 61726 -14360
rect 61196 -14540 61426 -14370
rect 60436 -14830 60536 -14810
rect 60436 -14950 60446 -14830
rect 60526 -14950 60536 -14830
rect 60436 -14960 60536 -14950
rect 60256 -15200 60416 -15070
rect 60256 -15330 60266 -15200
rect 60406 -15330 60416 -15200
rect 60256 -15350 60416 -15330
rect 58956 -15400 59156 -15390
rect 58956 -15580 58966 -15400
rect 59146 -15580 59156 -15400
rect 59986 -15500 59996 -15390
rect 60106 -15500 60116 -15390
rect 58956 -15590 59156 -15580
rect 59700 -15600 66500 -15500
rect 59700 -15900 59800 -15600
rect 60300 -15900 65900 -15600
rect 66400 -15900 66500 -15600
rect 59700 -16000 66500 -15900
rect 58946 -17670 59146 -17650
rect 58946 -17830 58966 -17670
rect 59126 -17830 59146 -17670
rect 58946 -17850 59146 -17830
rect 59316 -17710 59426 -17650
rect 59316 -17850 59336 -17710
rect 59416 -17850 59426 -17710
rect 58956 -17930 59136 -17850
rect 58956 -18040 58996 -17930
rect 59106 -18040 59136 -17930
rect 58396 -18130 58896 -18040
rect 58956 -18100 59136 -18040
rect 59316 -18080 59426 -17850
rect 59946 -17720 60386 -17600
rect 59946 -17840 60046 -17720
rect 60126 -17840 60386 -17720
rect 59946 -17890 60386 -17840
rect 58396 -18490 58486 -18130
rect 58816 -18490 58896 -18130
rect 58996 -18400 59086 -18100
rect 58996 -18460 59006 -18400
rect 59066 -18460 59086 -18400
rect 58996 -18470 59086 -18460
rect 59266 -18130 59426 -18080
rect 59506 -17940 59796 -17900
rect 59506 -18040 59516 -17940
rect 59616 -18040 59796 -17940
rect 59506 -18100 59796 -18040
rect 59266 -18330 59366 -18130
rect 59266 -18390 59286 -18330
rect 59346 -18390 59366 -18330
rect 58396 -18600 58896 -18490
rect 59066 -18640 59176 -18630
rect 59066 -18710 59076 -18640
rect 59166 -18710 59176 -18640
rect 56470 -19238 56555 -19228
rect 56470 -19328 56480 -19238
rect 56550 -19328 56555 -19238
rect 56470 -19338 56555 -19328
rect 56470 -19718 56550 -19338
rect 57760 -19340 57800 -19220
rect 58240 -19340 58280 -19220
rect 57093 -19674 57373 -19664
rect 56470 -19728 56555 -19718
rect 56470 -19778 56480 -19728
rect 56475 -19788 56480 -19778
rect 56550 -19788 56555 -19728
rect 56475 -19798 56555 -19788
rect 57093 -19814 57098 -19674
rect 57368 -19814 57373 -19674
rect 57093 -19824 57373 -19814
rect 55870 -20278 55980 -19838
rect 55870 -20318 55880 -20278
rect 55875 -20358 55880 -20318
rect 55970 -20318 55980 -20278
rect 56060 -20268 56220 -20258
rect 55970 -20358 55975 -20318
rect 55875 -20368 55975 -20358
rect 55590 -20478 55620 -20388
rect 55710 -20478 55720 -20388
rect 56060 -20438 56220 -20428
rect 56060 -20448 56200 -20438
rect 55590 -20488 55720 -20478
rect 56015 -20458 56200 -20448
rect 56015 -20608 56020 -20458
rect 56080 -20608 56200 -20458
rect 56644 -20468 57008 -20463
rect 55215 -20618 55325 -20608
rect 56015 -20618 56085 -20608
rect 55215 -20718 55220 -20618
rect 55320 -20718 55325 -20618
rect 56644 -20686 56654 -20468
rect 56998 -20686 57008 -20468
rect 56644 -20691 57008 -20686
rect 55215 -20728 55325 -20718
rect 55315 -20928 55475 -20918
rect 55315 -21068 55320 -20928
rect 55470 -21068 55475 -20928
rect 55315 -21078 55475 -21068
rect 39400 -21400 40100 -21300
rect 39400 -22000 39500 -21400
rect 40000 -21500 56200 -21400
rect 40000 -21900 55500 -21500
rect 56100 -21900 56200 -21500
rect 40000 -22000 56200 -21900
rect 39400 -22100 40100 -22000
rect 51400 -22480 55800 -22400
rect 51400 -22500 55440 -22480
rect 51400 -22700 51500 -22500
rect 52500 -22700 55440 -22500
rect 51400 -22760 55440 -22700
rect 55720 -22760 55800 -22480
rect 51400 -22800 55800 -22760
rect 55360 -22840 55800 -22800
rect 47660 -23020 48100 -23000
rect 47660 -23440 47680 -23020
rect 48080 -23120 48100 -23020
rect 48080 -23140 53800 -23120
rect 48080 -23340 53480 -23140
rect 53780 -23340 53800 -23140
rect 56496 -23180 57026 -23175
rect 48080 -23360 53800 -23340
rect 55955 -23338 56045 -23328
rect 48080 -23440 48100 -23360
rect 47660 -23460 48100 -23440
rect 53515 -23458 53645 -23448
rect 53510 -23568 53520 -23458
rect 53640 -23568 53645 -23458
rect 55955 -23488 55960 -23338
rect 56040 -23488 56200 -23338
rect 56496 -23430 56506 -23180
rect 57016 -23430 57026 -23180
rect 56496 -23435 57026 -23430
rect 55955 -23498 56200 -23488
rect 53510 -23578 53645 -23568
rect 55275 -23518 55490 -23508
rect 53045 -23758 53255 -23748
rect 53045 -25508 53050 -23758
rect 53250 -25508 53255 -23758
rect 53045 -25518 53255 -25508
rect 53510 -25718 53630 -23578
rect 55275 -23608 55280 -23518
rect 55400 -23608 55490 -23518
rect 56060 -23538 56200 -23498
rect 56060 -23548 56220 -23538
rect 55275 -23618 55490 -23608
rect 55220 -23858 55325 -23848
rect 55220 -24028 55230 -23858
rect 55320 -24028 55325 -23858
rect 55220 -24038 55325 -24028
rect 55015 -24648 55125 -24638
rect 55015 -24728 55020 -24648
rect 55120 -24728 55125 -24648
rect 55015 -24738 55125 -24728
rect 55220 -25338 55310 -24038
rect 55215 -25348 55315 -25338
rect 55215 -25518 55220 -25348
rect 55310 -25438 55315 -25348
rect 55400 -25348 55490 -23618
rect 55875 -23618 55990 -23608
rect 55875 -23658 55880 -23618
rect 55870 -23698 55880 -23658
rect 55970 -23698 55990 -23618
rect 55870 -23778 55990 -23698
rect 56060 -23718 56220 -23708
rect 55590 -23868 55720 -23858
rect 55590 -23998 55600 -23868
rect 55710 -23998 55720 -23868
rect 55400 -25358 55510 -25348
rect 55310 -25518 55320 -25438
rect 55400 -25518 55410 -25358
rect 55215 -25528 55320 -25518
rect 53505 -25728 53635 -25718
rect 14400 -26400 36000 -25800
rect 53505 -25848 53510 -25728
rect 53630 -25848 53635 -25728
rect 53505 -25858 53635 -25848
rect 55220 -26008 55320 -25528
rect 55405 -25528 55410 -25518
rect 55500 -25528 55510 -25358
rect 55405 -25538 55510 -25528
rect 55590 -25788 55720 -23998
rect 55870 -24158 55980 -23778
rect 57093 -24164 57373 -24154
rect 56475 -24188 56555 -24178
rect 56470 -24248 56480 -24188
rect 56550 -24248 56555 -24188
rect 56470 -24258 56555 -24248
rect 55870 -24638 55980 -24268
rect 55870 -24728 55880 -24638
rect 55970 -24728 55980 -24638
rect 55870 -25128 55980 -24728
rect 56470 -24628 56550 -24258
rect 57093 -24304 57098 -24164
rect 57368 -24304 57373 -24164
rect 57093 -24314 57373 -24304
rect 57760 -24620 58280 -19340
rect 58516 -19260 58796 -19190
rect 58516 -19460 58556 -19260
rect 58756 -19460 58796 -19260
rect 59066 -19210 59176 -18710
rect 59266 -18820 59366 -18390
rect 59536 -18290 59616 -18100
rect 59536 -18350 59546 -18290
rect 59606 -18350 59616 -18290
rect 59536 -18410 59616 -18350
rect 59536 -18470 59546 -18410
rect 59606 -18470 59616 -18410
rect 59536 -18480 59616 -18470
rect 59266 -18830 59376 -18820
rect 59266 -18920 59286 -18830
rect 59366 -18920 59376 -18830
rect 59736 -18850 59796 -18100
rect 59856 -18340 59976 -18330
rect 59856 -18430 59866 -18340
rect 59966 -18430 59976 -18340
rect 59856 -18440 59976 -18430
rect 60036 -18520 60136 -17890
rect 61026 -17920 61136 -17910
rect 61026 -18050 61056 -17920
rect 61126 -18050 61136 -17920
rect 60436 -18320 60536 -18310
rect 60436 -18420 60446 -18320
rect 60526 -18420 60536 -18320
rect 60436 -18430 60536 -18420
rect 60036 -18600 60046 -18520
rect 60126 -18600 60136 -18520
rect 60036 -18610 60136 -18600
rect 60546 -18610 60636 -18600
rect 60386 -18690 60556 -18610
rect 60626 -18690 60636 -18610
rect 59966 -18700 60326 -18690
rect 59966 -18770 59976 -18700
rect 60316 -18770 60326 -18700
rect 60546 -18710 60636 -18690
rect 59966 -18780 60326 -18770
rect 59566 -18870 59796 -18850
rect 59566 -18880 59576 -18870
rect 59266 -18930 59376 -18920
rect 59516 -18930 59576 -18880
rect 59636 -18930 59796 -18870
rect 59266 -19040 59366 -18930
rect 59266 -19130 59286 -19040
rect 59356 -19130 59366 -19040
rect 59266 -19160 59366 -19130
rect 59516 -18940 59796 -18930
rect 59066 -19280 59076 -19210
rect 59166 -19280 59176 -19210
rect 59066 -19290 59176 -19280
rect 59306 -19230 59386 -19220
rect 59306 -19290 59316 -19230
rect 59376 -19290 59386 -19230
rect 59516 -19270 59596 -18940
rect 60286 -18950 60476 -18940
rect 59906 -18980 60016 -18970
rect 59906 -19160 59916 -18980
rect 60006 -19160 60016 -18980
rect 59906 -19170 60016 -19160
rect 60286 -19090 60306 -18950
rect 60456 -19090 60476 -18950
rect 60286 -19100 60476 -19090
rect 58516 -19540 58796 -19460
rect 59066 -19370 59176 -19360
rect 59066 -19440 59076 -19370
rect 59166 -19440 59176 -19370
rect 59066 -19940 59176 -19440
rect 59306 -19490 59386 -19290
rect 60076 -19280 60196 -19240
rect 60076 -19440 60096 -19280
rect 60176 -19440 60196 -19280
rect 60076 -19480 60196 -19440
rect 59066 -20000 59076 -19940
rect 59166 -20000 59176 -19940
rect 59066 -20010 59176 -20000
rect 59236 -19520 59386 -19490
rect 59236 -19610 59266 -19520
rect 59366 -19610 59386 -19520
rect 59236 -19630 59386 -19610
rect 59906 -19490 60016 -19480
rect 59236 -19760 59376 -19630
rect 59906 -19680 59916 -19490
rect 60006 -19680 60016 -19490
rect 59906 -19690 60016 -19680
rect 60286 -19510 60376 -19100
rect 60556 -19500 60626 -18710
rect 61026 -19020 61136 -18050
rect 61196 -18720 61356 -18710
rect 61196 -18900 61206 -18720
rect 61346 -18900 61356 -18720
rect 61196 -18910 61356 -18900
rect 61026 -19130 61036 -19020
rect 61126 -19130 61136 -19020
rect 61026 -19140 61136 -19130
rect 61246 -19250 61366 -19240
rect 61246 -19260 61276 -19250
rect 61246 -19460 61256 -19260
rect 61356 -19460 61366 -19250
rect 61246 -19470 61366 -19460
rect 60466 -19510 60626 -19500
rect 60286 -19570 60406 -19510
rect 60466 -19570 60476 -19510
rect 60536 -19570 60626 -19510
rect 59236 -19850 59266 -19760
rect 59366 -19850 59376 -19760
rect 59236 -19900 59376 -19850
rect 59506 -19710 59606 -19700
rect 59506 -19780 59516 -19710
rect 59596 -19780 59606 -19710
rect 59506 -19790 59606 -19780
rect 59236 -19920 59386 -19900
rect 59236 -19980 59316 -19920
rect 59376 -19980 59386 -19920
rect 58396 -20550 58896 -20050
rect 59236 -20230 59386 -19980
rect 59006 -20300 59086 -20280
rect 59236 -20290 59256 -20230
rect 59366 -20290 59386 -20230
rect 59236 -20300 59386 -20290
rect 59506 -20180 59596 -19790
rect 59986 -19920 60116 -19910
rect 59986 -19980 59996 -19920
rect 60106 -19980 60116 -19920
rect 59506 -20190 59616 -20180
rect 59506 -20260 59546 -20190
rect 59606 -20260 59616 -20190
rect 59006 -20360 59016 -20300
rect 59076 -20360 59086 -20300
rect 59006 -20550 59086 -20360
rect 59506 -20310 59616 -20260
rect 59506 -20370 59546 -20310
rect 59606 -20370 59616 -20310
rect 59796 -20210 59926 -20200
rect 59796 -20320 59806 -20210
rect 59916 -20320 59926 -20210
rect 59796 -20330 59926 -20320
rect 59006 -20640 59126 -20550
rect 59006 -20710 59016 -20640
rect 59076 -20710 59126 -20640
rect 59006 -20790 59126 -20710
rect 59506 -20640 59616 -20370
rect 59506 -20710 59546 -20640
rect 59606 -20710 59616 -20640
rect 59506 -20720 59616 -20710
rect 59986 -20790 60116 -19980
rect 60286 -20470 60376 -19570
rect 60466 -19580 60626 -19570
rect 61486 -19570 61726 -19540
rect 61486 -19620 61496 -19570
rect 61326 -19630 61496 -19620
rect 61326 -19750 61336 -19630
rect 61196 -19760 61336 -19750
rect 61456 -19740 61496 -19630
rect 61696 -19740 61726 -19570
rect 61456 -19760 61726 -19740
rect 61196 -19770 61726 -19760
rect 61196 -19940 61426 -19770
rect 60436 -20230 60536 -20210
rect 60436 -20350 60446 -20230
rect 60526 -20350 60536 -20230
rect 60436 -20360 60536 -20350
rect 60256 -20600 60416 -20470
rect 60256 -20730 60266 -20600
rect 60406 -20730 60416 -20600
rect 60256 -20750 60416 -20730
rect 58956 -20800 59156 -20790
rect 58956 -20980 58966 -20800
rect 59146 -20980 59156 -20800
rect 59986 -20900 59996 -20790
rect 60106 -20900 60116 -20790
rect 58956 -20990 59156 -20980
rect 59700 -21000 65500 -20900
rect 59700 -21300 59800 -21000
rect 60300 -21300 64900 -21000
rect 65400 -21300 65500 -21000
rect 59700 -21400 65500 -21300
rect 58946 -23070 59146 -23050
rect 58946 -23230 58966 -23070
rect 59126 -23230 59146 -23070
rect 58946 -23250 59146 -23230
rect 59316 -23110 59426 -23050
rect 59316 -23250 59336 -23110
rect 59416 -23250 59426 -23110
rect 58956 -23330 59136 -23250
rect 58956 -23440 58996 -23330
rect 59106 -23440 59136 -23330
rect 58396 -23530 58896 -23440
rect 58956 -23500 59136 -23440
rect 59316 -23480 59426 -23250
rect 59946 -23120 60386 -23000
rect 59946 -23240 60046 -23120
rect 60126 -23240 60386 -23120
rect 59946 -23290 60386 -23240
rect 58396 -23890 58486 -23530
rect 58816 -23890 58896 -23530
rect 58996 -23800 59086 -23500
rect 58996 -23860 59006 -23800
rect 59066 -23860 59086 -23800
rect 58996 -23870 59086 -23860
rect 59266 -23530 59426 -23480
rect 59506 -23340 59796 -23300
rect 59506 -23440 59516 -23340
rect 59616 -23440 59796 -23340
rect 59506 -23500 59796 -23440
rect 59266 -23730 59366 -23530
rect 59266 -23790 59286 -23730
rect 59346 -23790 59366 -23730
rect 58396 -24000 58896 -23890
rect 59066 -24040 59176 -24030
rect 59066 -24110 59076 -24040
rect 59166 -24110 59176 -24040
rect 56470 -24638 56555 -24628
rect 56470 -24728 56480 -24638
rect 56550 -24728 56555 -24638
rect 56470 -24738 56555 -24728
rect 56470 -25118 56550 -24738
rect 57760 -24740 57800 -24620
rect 58240 -24740 58280 -24620
rect 57093 -25074 57373 -25064
rect 56470 -25128 56555 -25118
rect 56470 -25178 56480 -25128
rect 56475 -25188 56480 -25178
rect 56550 -25188 56555 -25128
rect 56475 -25198 56555 -25188
rect 57093 -25214 57098 -25074
rect 57368 -25214 57373 -25074
rect 57093 -25224 57373 -25214
rect 55870 -25678 55980 -25238
rect 55870 -25718 55880 -25678
rect 55875 -25758 55880 -25718
rect 55970 -25718 55980 -25678
rect 56060 -25668 56220 -25658
rect 55970 -25758 55975 -25718
rect 55875 -25768 55975 -25758
rect 55590 -25878 55620 -25788
rect 55710 -25878 55720 -25788
rect 56060 -25838 56220 -25828
rect 56060 -25848 56200 -25838
rect 55590 -25888 55720 -25878
rect 56015 -25858 56200 -25848
rect 56015 -26008 56020 -25858
rect 56080 -26008 56200 -25858
rect 56644 -25868 57008 -25863
rect 55215 -26018 55325 -26008
rect 56015 -26018 56085 -26008
rect 55215 -26118 55220 -26018
rect 55320 -26118 55325 -26018
rect 56644 -26086 56654 -25868
rect 56998 -26086 57008 -25868
rect 56644 -26091 57008 -26086
rect 55215 -26128 55325 -26118
rect 14400 -31200 15000 -26400
rect 19400 -30400 26600 -26400
rect 35200 -30400 36000 -26400
rect 55315 -26328 55475 -26318
rect 55315 -26468 55320 -26328
rect 55470 -26468 55475 -26328
rect 55315 -26478 55475 -26468
rect 40300 -26800 41100 -26700
rect 40300 -27400 40400 -26800
rect 41000 -26900 56200 -26800
rect 41000 -27300 55500 -26900
rect 56100 -27300 56200 -26900
rect 41000 -27400 56200 -27300
rect 40300 -27500 41100 -27400
rect 51400 -27880 55800 -27800
rect 51400 -27900 55460 -27880
rect 51400 -28100 51500 -27900
rect 52500 -28100 55460 -27900
rect 51400 -28160 55460 -28100
rect 55720 -28160 55800 -27880
rect 51400 -28200 55800 -28160
rect 55380 -28240 55800 -28200
rect 47780 -28460 48100 -28440
rect 47780 -28840 47800 -28460
rect 48080 -28520 48100 -28460
rect 48080 -28540 53800 -28520
rect 48080 -28740 53480 -28540
rect 53780 -28740 53800 -28540
rect 56496 -28580 57026 -28575
rect 48080 -28760 53800 -28740
rect 55955 -28738 56045 -28728
rect 48080 -28840 48100 -28760
rect 47780 -28860 48100 -28840
rect 53515 -28858 53645 -28848
rect 53510 -28968 53520 -28858
rect 53640 -28968 53645 -28858
rect 55955 -28888 55960 -28738
rect 56040 -28888 56200 -28738
rect 56496 -28830 56506 -28580
rect 57016 -28830 57026 -28580
rect 56496 -28835 57026 -28830
rect 55955 -28898 56200 -28888
rect 53510 -28978 53645 -28968
rect 55275 -28918 55490 -28908
rect 19400 -31200 36000 -30400
rect 53045 -29158 53255 -29148
rect 53045 -30908 53050 -29158
rect 53250 -30908 53255 -29158
rect 53045 -30918 53255 -30908
rect 53510 -31118 53630 -28978
rect 55275 -29008 55280 -28918
rect 55400 -29008 55490 -28918
rect 56060 -28938 56200 -28898
rect 56060 -28948 56220 -28938
rect 55275 -29018 55490 -29008
rect 55220 -29258 55325 -29248
rect 55220 -29428 55230 -29258
rect 55320 -29428 55325 -29258
rect 55220 -29438 55325 -29428
rect 55015 -30048 55125 -30038
rect 55015 -30128 55020 -30048
rect 55120 -30128 55125 -30048
rect 55015 -30138 55125 -30128
rect 55220 -30738 55310 -29438
rect 55215 -30748 55315 -30738
rect 55215 -30918 55220 -30748
rect 55310 -30838 55315 -30748
rect 55400 -30748 55490 -29018
rect 55875 -29018 55990 -29008
rect 55875 -29058 55880 -29018
rect 55870 -29098 55880 -29058
rect 55970 -29098 55990 -29018
rect 55870 -29178 55990 -29098
rect 56060 -29118 56220 -29108
rect 55590 -29268 55720 -29258
rect 55590 -29398 55600 -29268
rect 55710 -29398 55720 -29268
rect 55400 -30758 55510 -30748
rect 55310 -30918 55320 -30838
rect 55400 -30918 55410 -30758
rect 55215 -30928 55320 -30918
rect 14400 -31800 36000 -31200
rect 53505 -31128 53635 -31118
rect 53505 -31248 53510 -31128
rect 53630 -31248 53635 -31128
rect 53505 -31258 53635 -31248
rect 55220 -31408 55320 -30928
rect 55405 -30928 55410 -30918
rect 55500 -30928 55510 -30758
rect 55405 -30938 55510 -30928
rect 55590 -31188 55720 -29398
rect 55870 -29558 55980 -29178
rect 57093 -29564 57373 -29554
rect 56475 -29588 56555 -29578
rect 56470 -29648 56480 -29588
rect 56550 -29648 56555 -29588
rect 56470 -29658 56555 -29648
rect 55870 -30038 55980 -29668
rect 55870 -30128 55880 -30038
rect 55970 -30128 55980 -30038
rect 55870 -30528 55980 -30128
rect 56470 -30028 56550 -29658
rect 57093 -29704 57098 -29564
rect 57368 -29704 57373 -29564
rect 57093 -29714 57373 -29704
rect 57760 -30020 58280 -24740
rect 58516 -24660 58796 -24590
rect 58516 -24860 58556 -24660
rect 58756 -24860 58796 -24660
rect 59066 -24610 59176 -24110
rect 59266 -24220 59366 -23790
rect 59536 -23690 59616 -23500
rect 59536 -23750 59546 -23690
rect 59606 -23750 59616 -23690
rect 59536 -23810 59616 -23750
rect 59536 -23870 59546 -23810
rect 59606 -23870 59616 -23810
rect 59536 -23880 59616 -23870
rect 59266 -24230 59376 -24220
rect 59266 -24320 59286 -24230
rect 59366 -24320 59376 -24230
rect 59736 -24250 59796 -23500
rect 59856 -23740 59976 -23730
rect 59856 -23830 59866 -23740
rect 59966 -23830 59976 -23740
rect 59856 -23840 59976 -23830
rect 60036 -23920 60136 -23290
rect 61026 -23320 61136 -23310
rect 61026 -23450 61056 -23320
rect 61126 -23450 61136 -23320
rect 60436 -23720 60536 -23710
rect 60436 -23820 60446 -23720
rect 60526 -23820 60536 -23720
rect 60436 -23830 60536 -23820
rect 60036 -24000 60046 -23920
rect 60126 -24000 60136 -23920
rect 60036 -24010 60136 -24000
rect 60546 -24010 60636 -24000
rect 60386 -24090 60556 -24010
rect 60626 -24090 60636 -24010
rect 59966 -24100 60326 -24090
rect 59966 -24170 59976 -24100
rect 60316 -24170 60326 -24100
rect 60546 -24110 60636 -24090
rect 59966 -24180 60326 -24170
rect 59566 -24270 59796 -24250
rect 59566 -24280 59576 -24270
rect 59266 -24330 59376 -24320
rect 59516 -24330 59576 -24280
rect 59636 -24330 59796 -24270
rect 59266 -24440 59366 -24330
rect 59266 -24530 59286 -24440
rect 59356 -24530 59366 -24440
rect 59266 -24560 59366 -24530
rect 59516 -24340 59796 -24330
rect 59066 -24680 59076 -24610
rect 59166 -24680 59176 -24610
rect 59066 -24690 59176 -24680
rect 59306 -24630 59386 -24620
rect 59306 -24690 59316 -24630
rect 59376 -24690 59386 -24630
rect 59516 -24670 59596 -24340
rect 60286 -24350 60476 -24340
rect 59906 -24380 60016 -24370
rect 59906 -24560 59916 -24380
rect 60006 -24560 60016 -24380
rect 59906 -24570 60016 -24560
rect 60286 -24490 60306 -24350
rect 60456 -24490 60476 -24350
rect 60286 -24500 60476 -24490
rect 58516 -24940 58796 -24860
rect 59066 -24770 59176 -24760
rect 59066 -24840 59076 -24770
rect 59166 -24840 59176 -24770
rect 59066 -25340 59176 -24840
rect 59306 -24890 59386 -24690
rect 60076 -24680 60196 -24640
rect 60076 -24840 60096 -24680
rect 60176 -24840 60196 -24680
rect 60076 -24880 60196 -24840
rect 59066 -25400 59076 -25340
rect 59166 -25400 59176 -25340
rect 59066 -25410 59176 -25400
rect 59236 -24920 59386 -24890
rect 59236 -25010 59266 -24920
rect 59366 -25010 59386 -24920
rect 59236 -25030 59386 -25010
rect 59906 -24890 60016 -24880
rect 59236 -25160 59376 -25030
rect 59906 -25080 59916 -24890
rect 60006 -25080 60016 -24890
rect 59906 -25090 60016 -25080
rect 60286 -24910 60376 -24500
rect 60556 -24900 60626 -24110
rect 61026 -24420 61136 -23450
rect 61196 -24120 61356 -24110
rect 61196 -24300 61206 -24120
rect 61346 -24300 61356 -24120
rect 61196 -24310 61356 -24300
rect 61026 -24530 61036 -24420
rect 61126 -24530 61136 -24420
rect 61026 -24540 61136 -24530
rect 61246 -24650 61366 -24640
rect 61246 -24660 61276 -24650
rect 61246 -24860 61256 -24660
rect 61356 -24860 61366 -24650
rect 61246 -24870 61366 -24860
rect 60466 -24910 60626 -24900
rect 60286 -24970 60406 -24910
rect 60466 -24970 60476 -24910
rect 60536 -24970 60626 -24910
rect 59236 -25250 59266 -25160
rect 59366 -25250 59376 -25160
rect 59236 -25300 59376 -25250
rect 59506 -25110 59606 -25100
rect 59506 -25180 59516 -25110
rect 59596 -25180 59606 -25110
rect 59506 -25190 59606 -25180
rect 59236 -25320 59386 -25300
rect 59236 -25380 59316 -25320
rect 59376 -25380 59386 -25320
rect 58396 -25950 58896 -25450
rect 59236 -25630 59386 -25380
rect 59006 -25700 59086 -25680
rect 59236 -25690 59256 -25630
rect 59366 -25690 59386 -25630
rect 59236 -25700 59386 -25690
rect 59506 -25580 59596 -25190
rect 59986 -25320 60116 -25310
rect 59986 -25380 59996 -25320
rect 60106 -25380 60116 -25320
rect 59506 -25590 59616 -25580
rect 59506 -25660 59546 -25590
rect 59606 -25660 59616 -25590
rect 59006 -25760 59016 -25700
rect 59076 -25760 59086 -25700
rect 59006 -25950 59086 -25760
rect 59506 -25710 59616 -25660
rect 59506 -25770 59546 -25710
rect 59606 -25770 59616 -25710
rect 59796 -25610 59926 -25600
rect 59796 -25720 59806 -25610
rect 59916 -25720 59926 -25610
rect 59796 -25730 59926 -25720
rect 59006 -26040 59126 -25950
rect 59006 -26110 59016 -26040
rect 59076 -26110 59126 -26040
rect 59006 -26190 59126 -26110
rect 59506 -26040 59616 -25770
rect 59506 -26110 59546 -26040
rect 59606 -26110 59616 -26040
rect 59506 -26120 59616 -26110
rect 59986 -26190 60116 -25380
rect 60286 -25870 60376 -24970
rect 60466 -24980 60626 -24970
rect 61486 -24970 61726 -24940
rect 61486 -25020 61496 -24970
rect 61326 -25030 61496 -25020
rect 61326 -25150 61336 -25030
rect 61196 -25160 61336 -25150
rect 61456 -25140 61496 -25030
rect 61696 -25140 61726 -24970
rect 61456 -25160 61726 -25140
rect 61196 -25170 61726 -25160
rect 61196 -25340 61426 -25170
rect 60436 -25630 60536 -25610
rect 60436 -25750 60446 -25630
rect 60526 -25750 60536 -25630
rect 60436 -25760 60536 -25750
rect 60256 -26000 60416 -25870
rect 60256 -26130 60266 -26000
rect 60406 -26130 60416 -26000
rect 60256 -26150 60416 -26130
rect 58956 -26200 59156 -26190
rect 58956 -26380 58966 -26200
rect 59146 -26380 59156 -26200
rect 59986 -26300 59996 -26190
rect 60106 -26300 60116 -26190
rect 58956 -26390 59156 -26380
rect 59600 -26400 64200 -26300
rect 59600 -26800 59700 -26400
rect 60400 -26800 63700 -26400
rect 64100 -26800 64200 -26400
rect 59600 -26900 64200 -26800
rect 58946 -28470 59146 -28450
rect 58946 -28630 58966 -28470
rect 59126 -28630 59146 -28470
rect 58946 -28650 59146 -28630
rect 59316 -28510 59426 -28450
rect 59316 -28650 59336 -28510
rect 59416 -28650 59426 -28510
rect 58956 -28730 59136 -28650
rect 58956 -28840 58996 -28730
rect 59106 -28840 59136 -28730
rect 58396 -28930 58896 -28840
rect 58956 -28900 59136 -28840
rect 59316 -28880 59426 -28650
rect 59946 -28520 60386 -28400
rect 59946 -28640 60046 -28520
rect 60126 -28640 60386 -28520
rect 59946 -28690 60386 -28640
rect 58396 -29290 58486 -28930
rect 58816 -29290 58896 -28930
rect 58996 -29200 59086 -28900
rect 58996 -29260 59006 -29200
rect 59066 -29260 59086 -29200
rect 58996 -29270 59086 -29260
rect 59266 -28930 59426 -28880
rect 59506 -28740 59796 -28700
rect 59506 -28840 59516 -28740
rect 59616 -28840 59796 -28740
rect 59506 -28900 59796 -28840
rect 59266 -29130 59366 -28930
rect 59266 -29190 59286 -29130
rect 59346 -29190 59366 -29130
rect 58396 -29400 58896 -29290
rect 59066 -29440 59176 -29430
rect 59066 -29510 59076 -29440
rect 59166 -29510 59176 -29440
rect 56470 -30038 56555 -30028
rect 56470 -30128 56480 -30038
rect 56550 -30128 56555 -30038
rect 56470 -30138 56555 -30128
rect 56470 -30518 56550 -30138
rect 57760 -30140 57800 -30020
rect 58240 -30140 58280 -30020
rect 57093 -30474 57373 -30464
rect 56470 -30528 56555 -30518
rect 56470 -30578 56480 -30528
rect 56475 -30588 56480 -30578
rect 56550 -30588 56555 -30528
rect 56475 -30598 56555 -30588
rect 57093 -30614 57098 -30474
rect 57368 -30614 57373 -30474
rect 57093 -30624 57373 -30614
rect 55870 -31078 55980 -30638
rect 55870 -31118 55880 -31078
rect 55875 -31158 55880 -31118
rect 55970 -31118 55980 -31078
rect 56060 -31068 56220 -31058
rect 55970 -31158 55975 -31118
rect 55875 -31168 55975 -31158
rect 55590 -31278 55620 -31188
rect 55710 -31278 55720 -31188
rect 56060 -31238 56220 -31228
rect 56060 -31248 56200 -31238
rect 55590 -31288 55720 -31278
rect 56015 -31258 56200 -31248
rect 56015 -31408 56020 -31258
rect 56080 -31408 56200 -31258
rect 56644 -31268 57008 -31263
rect 55215 -31418 55325 -31408
rect 56015 -31418 56085 -31408
rect 55215 -31518 55220 -31418
rect 55320 -31518 55325 -31418
rect 56644 -31486 56654 -31268
rect 56998 -31486 57008 -31268
rect 56644 -31491 57008 -31486
rect 55215 -31528 55325 -31518
rect 55315 -31728 55475 -31718
rect 55315 -31868 55320 -31728
rect 55470 -31868 55475 -31728
rect 55315 -31878 55475 -31868
rect 41400 -32200 42200 -32100
rect 41400 -32800 41500 -32200
rect 42100 -32300 56200 -32200
rect 42100 -32700 55500 -32300
rect 56100 -32700 56200 -32300
rect 42100 -32800 56200 -32700
rect 41400 -32900 42200 -32800
rect 51400 -33280 55800 -33200
rect 51400 -33300 55460 -33280
rect 51400 -33500 51500 -33300
rect 52500 -33500 55460 -33300
rect 51400 -33560 55460 -33500
rect 55720 -33560 55800 -33280
rect 51400 -33600 55800 -33560
rect 55380 -33640 55800 -33600
rect 47740 -33860 48100 -33840
rect 47740 -34200 47760 -33860
rect 48080 -33920 48100 -33860
rect 48080 -33940 53800 -33920
rect 48080 -34140 53480 -33940
rect 53780 -34140 53800 -33940
rect 56496 -33980 57026 -33975
rect 48080 -34160 53800 -34140
rect 55955 -34138 56045 -34128
rect 48080 -34200 48100 -34160
rect 47740 -34220 48100 -34200
rect 53515 -34258 53645 -34248
rect 53510 -34368 53520 -34258
rect 53640 -34368 53645 -34258
rect 55955 -34288 55960 -34138
rect 56040 -34288 56200 -34138
rect 56496 -34230 56506 -33980
rect 57016 -34230 57026 -33980
rect 56496 -34235 57026 -34230
rect 55955 -34298 56200 -34288
rect 53510 -34378 53645 -34368
rect 55275 -34318 55490 -34308
rect 53045 -34558 53255 -34548
rect 53045 -36308 53050 -34558
rect 53250 -36308 53255 -34558
rect 53045 -36318 53255 -36308
rect 53510 -36518 53630 -34378
rect 55275 -34408 55280 -34318
rect 55400 -34408 55490 -34318
rect 56060 -34338 56200 -34298
rect 56060 -34348 56220 -34338
rect 55275 -34418 55490 -34408
rect 55220 -34658 55325 -34648
rect 55220 -34828 55230 -34658
rect 55320 -34828 55325 -34658
rect 55220 -34838 55325 -34828
rect 55015 -35448 55125 -35438
rect 55015 -35528 55020 -35448
rect 55120 -35528 55125 -35448
rect 55015 -35538 55125 -35528
rect 55220 -36138 55310 -34838
rect 55215 -36148 55315 -36138
rect 55215 -36318 55220 -36148
rect 55310 -36238 55315 -36148
rect 55400 -36148 55490 -34418
rect 55875 -34418 55990 -34408
rect 55875 -34458 55880 -34418
rect 55870 -34498 55880 -34458
rect 55970 -34498 55990 -34418
rect 55870 -34578 55990 -34498
rect 56060 -34518 56220 -34508
rect 55590 -34668 55720 -34658
rect 55590 -34798 55600 -34668
rect 55710 -34798 55720 -34668
rect 55400 -36158 55510 -36148
rect 55310 -36318 55320 -36238
rect 55400 -36318 55410 -36158
rect 55215 -36328 55320 -36318
rect 53505 -36528 53635 -36518
rect 53505 -36648 53510 -36528
rect 53630 -36648 53635 -36528
rect 53505 -36658 53635 -36648
rect 55220 -36808 55320 -36328
rect 55405 -36328 55410 -36318
rect 55500 -36328 55510 -36158
rect 55405 -36338 55510 -36328
rect 55590 -36588 55720 -34798
rect 55870 -34958 55980 -34578
rect 57093 -34964 57373 -34954
rect 56475 -34988 56555 -34978
rect 56470 -35048 56480 -34988
rect 56550 -35048 56555 -34988
rect 56470 -35058 56555 -35048
rect 55870 -35438 55980 -35068
rect 55870 -35528 55880 -35438
rect 55970 -35528 55980 -35438
rect 55870 -35928 55980 -35528
rect 56470 -35428 56550 -35058
rect 57093 -35104 57098 -34964
rect 57368 -35104 57373 -34964
rect 57093 -35114 57373 -35104
rect 57760 -35420 58280 -30140
rect 58516 -30060 58796 -29990
rect 58516 -30260 58556 -30060
rect 58756 -30260 58796 -30060
rect 59066 -30010 59176 -29510
rect 59266 -29620 59366 -29190
rect 59536 -29090 59616 -28900
rect 59536 -29150 59546 -29090
rect 59606 -29150 59616 -29090
rect 59536 -29210 59616 -29150
rect 59536 -29270 59546 -29210
rect 59606 -29270 59616 -29210
rect 59536 -29280 59616 -29270
rect 59266 -29630 59376 -29620
rect 59266 -29720 59286 -29630
rect 59366 -29720 59376 -29630
rect 59736 -29650 59796 -28900
rect 59856 -29140 59976 -29130
rect 59856 -29230 59866 -29140
rect 59966 -29230 59976 -29140
rect 59856 -29240 59976 -29230
rect 60036 -29320 60136 -28690
rect 61026 -28720 61136 -28710
rect 61026 -28850 61056 -28720
rect 61126 -28850 61136 -28720
rect 60436 -29120 60536 -29110
rect 60436 -29220 60446 -29120
rect 60526 -29220 60536 -29120
rect 60436 -29230 60536 -29220
rect 60036 -29400 60046 -29320
rect 60126 -29400 60136 -29320
rect 60036 -29410 60136 -29400
rect 60546 -29410 60636 -29400
rect 60386 -29490 60556 -29410
rect 60626 -29490 60636 -29410
rect 59966 -29500 60326 -29490
rect 59966 -29570 59976 -29500
rect 60316 -29570 60326 -29500
rect 60546 -29510 60636 -29490
rect 59966 -29580 60326 -29570
rect 59566 -29670 59796 -29650
rect 59566 -29680 59576 -29670
rect 59266 -29730 59376 -29720
rect 59516 -29730 59576 -29680
rect 59636 -29730 59796 -29670
rect 59266 -29840 59366 -29730
rect 59266 -29930 59286 -29840
rect 59356 -29930 59366 -29840
rect 59266 -29960 59366 -29930
rect 59516 -29740 59796 -29730
rect 59066 -30080 59076 -30010
rect 59166 -30080 59176 -30010
rect 59066 -30090 59176 -30080
rect 59306 -30030 59386 -30020
rect 59306 -30090 59316 -30030
rect 59376 -30090 59386 -30030
rect 59516 -30070 59596 -29740
rect 60286 -29750 60476 -29740
rect 59906 -29780 60016 -29770
rect 59906 -29960 59916 -29780
rect 60006 -29960 60016 -29780
rect 59906 -29970 60016 -29960
rect 60286 -29890 60306 -29750
rect 60456 -29890 60476 -29750
rect 60286 -29900 60476 -29890
rect 58516 -30340 58796 -30260
rect 59066 -30170 59176 -30160
rect 59066 -30240 59076 -30170
rect 59166 -30240 59176 -30170
rect 59066 -30740 59176 -30240
rect 59306 -30290 59386 -30090
rect 60076 -30080 60196 -30040
rect 60076 -30240 60096 -30080
rect 60176 -30240 60196 -30080
rect 60076 -30280 60196 -30240
rect 59066 -30800 59076 -30740
rect 59166 -30800 59176 -30740
rect 59066 -30810 59176 -30800
rect 59236 -30320 59386 -30290
rect 59236 -30410 59266 -30320
rect 59366 -30410 59386 -30320
rect 59236 -30430 59386 -30410
rect 59906 -30290 60016 -30280
rect 59236 -30560 59376 -30430
rect 59906 -30480 59916 -30290
rect 60006 -30480 60016 -30290
rect 59906 -30490 60016 -30480
rect 60286 -30310 60376 -29900
rect 60556 -30300 60626 -29510
rect 61026 -29820 61136 -28850
rect 61196 -29520 61356 -29510
rect 61196 -29700 61206 -29520
rect 61346 -29700 61356 -29520
rect 61196 -29710 61356 -29700
rect 61026 -29930 61036 -29820
rect 61126 -29930 61136 -29820
rect 61026 -29940 61136 -29930
rect 61246 -30050 61366 -30040
rect 61246 -30060 61276 -30050
rect 61246 -30260 61256 -30060
rect 61356 -30260 61366 -30050
rect 61246 -30270 61366 -30260
rect 60466 -30310 60626 -30300
rect 60286 -30370 60406 -30310
rect 60466 -30370 60476 -30310
rect 60536 -30370 60626 -30310
rect 59236 -30650 59266 -30560
rect 59366 -30650 59376 -30560
rect 59236 -30700 59376 -30650
rect 59506 -30510 59606 -30500
rect 59506 -30580 59516 -30510
rect 59596 -30580 59606 -30510
rect 59506 -30590 59606 -30580
rect 59236 -30720 59386 -30700
rect 59236 -30780 59316 -30720
rect 59376 -30780 59386 -30720
rect 58396 -31350 58896 -30850
rect 59236 -31030 59386 -30780
rect 59006 -31100 59086 -31080
rect 59236 -31090 59256 -31030
rect 59366 -31090 59386 -31030
rect 59236 -31100 59386 -31090
rect 59506 -30980 59596 -30590
rect 59986 -30720 60116 -30710
rect 59986 -30780 59996 -30720
rect 60106 -30780 60116 -30720
rect 59506 -30990 59616 -30980
rect 59506 -31060 59546 -30990
rect 59606 -31060 59616 -30990
rect 59006 -31160 59016 -31100
rect 59076 -31160 59086 -31100
rect 59006 -31350 59086 -31160
rect 59506 -31110 59616 -31060
rect 59506 -31170 59546 -31110
rect 59606 -31170 59616 -31110
rect 59796 -31010 59926 -31000
rect 59796 -31120 59806 -31010
rect 59916 -31120 59926 -31010
rect 59796 -31130 59926 -31120
rect 59006 -31440 59126 -31350
rect 59006 -31510 59016 -31440
rect 59076 -31510 59126 -31440
rect 59006 -31590 59126 -31510
rect 59506 -31440 59616 -31170
rect 59506 -31510 59546 -31440
rect 59606 -31510 59616 -31440
rect 59506 -31520 59616 -31510
rect 59986 -31590 60116 -30780
rect 60286 -31270 60376 -30370
rect 60466 -30380 60626 -30370
rect 61486 -30370 61726 -30340
rect 61486 -30420 61496 -30370
rect 61326 -30430 61496 -30420
rect 61326 -30550 61336 -30430
rect 61196 -30560 61336 -30550
rect 61456 -30540 61496 -30430
rect 61696 -30540 61726 -30370
rect 61456 -30560 61726 -30540
rect 61196 -30570 61726 -30560
rect 61196 -30740 61426 -30570
rect 60436 -31030 60536 -31010
rect 60436 -31150 60446 -31030
rect 60526 -31150 60536 -31030
rect 60436 -31160 60536 -31150
rect 60256 -31400 60416 -31270
rect 60256 -31530 60266 -31400
rect 60406 -31530 60416 -31400
rect 60256 -31550 60416 -31530
rect 58956 -31600 59156 -31590
rect 58956 -31780 58966 -31600
rect 59146 -31780 59156 -31600
rect 59986 -31700 59996 -31590
rect 60106 -31700 60116 -31590
rect 58956 -31790 59156 -31780
rect 59700 -31800 63400 -31700
rect 59700 -32100 59800 -31800
rect 60300 -32100 62900 -31800
rect 63300 -32100 63400 -31800
rect 59700 -32200 63400 -32100
rect 58946 -33870 59146 -33850
rect 58946 -34030 58966 -33870
rect 59126 -34030 59146 -33870
rect 58946 -34050 59146 -34030
rect 59316 -33910 59426 -33850
rect 59316 -34050 59336 -33910
rect 59416 -34050 59426 -33910
rect 58956 -34130 59136 -34050
rect 58956 -34240 58996 -34130
rect 59106 -34240 59136 -34130
rect 58396 -34330 58896 -34240
rect 58956 -34300 59136 -34240
rect 59316 -34280 59426 -34050
rect 59946 -33920 60386 -33800
rect 59946 -34040 60046 -33920
rect 60126 -34040 60386 -33920
rect 59946 -34090 60386 -34040
rect 58396 -34690 58486 -34330
rect 58816 -34690 58896 -34330
rect 58996 -34600 59086 -34300
rect 58996 -34660 59006 -34600
rect 59066 -34660 59086 -34600
rect 58996 -34670 59086 -34660
rect 59266 -34330 59426 -34280
rect 59506 -34140 59796 -34100
rect 59506 -34240 59516 -34140
rect 59616 -34240 59796 -34140
rect 59506 -34300 59796 -34240
rect 59266 -34530 59366 -34330
rect 59266 -34590 59286 -34530
rect 59346 -34590 59366 -34530
rect 58396 -34800 58896 -34690
rect 59066 -34840 59176 -34830
rect 59066 -34910 59076 -34840
rect 59166 -34910 59176 -34840
rect 56470 -35438 56555 -35428
rect 56470 -35528 56480 -35438
rect 56550 -35528 56555 -35438
rect 56470 -35538 56555 -35528
rect 56470 -35918 56550 -35538
rect 57760 -35540 57800 -35420
rect 58240 -35540 58280 -35420
rect 57093 -35874 57373 -35864
rect 56470 -35928 56555 -35918
rect 56470 -35978 56480 -35928
rect 56475 -35988 56480 -35978
rect 56550 -35988 56555 -35928
rect 56475 -35998 56555 -35988
rect 57093 -36014 57098 -35874
rect 57368 -36014 57373 -35874
rect 57093 -36024 57373 -36014
rect 55870 -36478 55980 -36038
rect 55870 -36518 55880 -36478
rect 55875 -36558 55880 -36518
rect 55970 -36518 55980 -36478
rect 56060 -36468 56220 -36458
rect 55970 -36558 55975 -36518
rect 55875 -36568 55975 -36558
rect 55590 -36678 55620 -36588
rect 55710 -36678 55720 -36588
rect 56060 -36638 56220 -36628
rect 56060 -36648 56200 -36638
rect 55590 -36688 55720 -36678
rect 56015 -36658 56200 -36648
rect 56015 -36808 56020 -36658
rect 56080 -36808 56200 -36658
rect 56644 -36668 57008 -36663
rect 55215 -36818 55325 -36808
rect 56015 -36818 56085 -36808
rect 55215 -36918 55220 -36818
rect 55320 -36918 55325 -36818
rect 56644 -36886 56654 -36668
rect 56998 -36886 57008 -36668
rect 56644 -36891 57008 -36886
rect 55215 -36928 55325 -36918
rect 14000 -38000 25000 -37000
rect 55315 -37128 55475 -37118
rect 55315 -37268 55320 -37128
rect 55470 -37268 55475 -37128
rect 55315 -37278 55475 -37268
rect 14000 -49000 15000 -38000
rect 24000 -49000 25000 -38000
rect 42400 -37600 43200 -37500
rect 42400 -38200 42500 -37600
rect 43100 -37700 56200 -37600
rect 43100 -38100 55400 -37700
rect 56100 -38100 56200 -37700
rect 43100 -38200 56200 -38100
rect 42400 -38300 43200 -38200
rect 51400 -38680 55800 -38600
rect 51400 -38700 55460 -38680
rect 51400 -38900 51500 -38700
rect 52500 -38900 55460 -38700
rect 51400 -38960 55460 -38900
rect 55720 -38960 55800 -38680
rect 51400 -39000 55800 -38960
rect 55380 -39040 55800 -39000
rect 47740 -39220 48100 -39200
rect 47740 -39640 47760 -39220
rect 48080 -39320 48100 -39220
rect 48080 -39340 53800 -39320
rect 48080 -39540 53480 -39340
rect 53780 -39540 53800 -39340
rect 56496 -39380 57026 -39375
rect 48080 -39560 53800 -39540
rect 55955 -39538 56045 -39528
rect 48080 -39640 48100 -39560
rect 47740 -39660 48100 -39640
rect 53515 -39658 53645 -39648
rect 53510 -39768 53520 -39658
rect 53640 -39768 53645 -39658
rect 55955 -39688 55960 -39538
rect 56040 -39688 56200 -39538
rect 56496 -39630 56506 -39380
rect 57016 -39630 57026 -39380
rect 56496 -39635 57026 -39630
rect 55955 -39698 56200 -39688
rect 53510 -39778 53645 -39768
rect 55275 -39718 55490 -39708
rect 53045 -39958 53255 -39948
rect 53045 -41708 53050 -39958
rect 53250 -41708 53255 -39958
rect 53045 -41718 53255 -41708
rect 53510 -41918 53630 -39778
rect 55275 -39808 55280 -39718
rect 55400 -39808 55490 -39718
rect 56060 -39738 56200 -39698
rect 56060 -39748 56220 -39738
rect 55275 -39818 55490 -39808
rect 55220 -40058 55325 -40048
rect 55220 -40228 55230 -40058
rect 55320 -40228 55325 -40058
rect 55220 -40238 55325 -40228
rect 55015 -40848 55125 -40838
rect 55015 -40928 55020 -40848
rect 55120 -40928 55125 -40848
rect 55015 -40938 55125 -40928
rect 55220 -41538 55310 -40238
rect 55215 -41548 55315 -41538
rect 55215 -41718 55220 -41548
rect 55310 -41638 55315 -41548
rect 55400 -41548 55490 -39818
rect 55875 -39818 55990 -39808
rect 55875 -39858 55880 -39818
rect 55870 -39898 55880 -39858
rect 55970 -39898 55990 -39818
rect 55870 -39978 55990 -39898
rect 56060 -39918 56220 -39908
rect 55590 -40068 55720 -40058
rect 55590 -40198 55600 -40068
rect 55710 -40198 55720 -40068
rect 55400 -41558 55510 -41548
rect 55310 -41718 55320 -41638
rect 55400 -41718 55410 -41558
rect 55215 -41728 55320 -41718
rect 53505 -41928 53635 -41918
rect 53505 -42048 53510 -41928
rect 53630 -42048 53635 -41928
rect 53505 -42058 53635 -42048
rect 55220 -42208 55320 -41728
rect 55405 -41728 55410 -41718
rect 55500 -41728 55510 -41558
rect 55405 -41738 55510 -41728
rect 55590 -41988 55720 -40198
rect 55870 -40358 55980 -39978
rect 57093 -40364 57373 -40354
rect 56475 -40388 56555 -40378
rect 56470 -40448 56480 -40388
rect 56550 -40448 56555 -40388
rect 56470 -40458 56555 -40448
rect 55870 -40838 55980 -40468
rect 55870 -40928 55880 -40838
rect 55970 -40928 55980 -40838
rect 55870 -41328 55980 -40928
rect 56470 -40828 56550 -40458
rect 57093 -40504 57098 -40364
rect 57368 -40504 57373 -40364
rect 57093 -40514 57373 -40504
rect 57760 -40820 58280 -35540
rect 58516 -35460 58796 -35390
rect 58516 -35660 58556 -35460
rect 58756 -35660 58796 -35460
rect 59066 -35410 59176 -34910
rect 59266 -35020 59366 -34590
rect 59536 -34490 59616 -34300
rect 59536 -34550 59546 -34490
rect 59606 -34550 59616 -34490
rect 59536 -34610 59616 -34550
rect 59536 -34670 59546 -34610
rect 59606 -34670 59616 -34610
rect 59536 -34680 59616 -34670
rect 59266 -35030 59376 -35020
rect 59266 -35120 59286 -35030
rect 59366 -35120 59376 -35030
rect 59736 -35050 59796 -34300
rect 59856 -34540 59976 -34530
rect 59856 -34630 59866 -34540
rect 59966 -34630 59976 -34540
rect 59856 -34640 59976 -34630
rect 60036 -34720 60136 -34090
rect 71900 -34100 74100 -34000
rect 61026 -34120 61136 -34110
rect 61026 -34250 61056 -34120
rect 61126 -34250 61136 -34120
rect 60436 -34520 60536 -34510
rect 60436 -34620 60446 -34520
rect 60526 -34620 60536 -34520
rect 60436 -34630 60536 -34620
rect 60036 -34800 60046 -34720
rect 60126 -34800 60136 -34720
rect 60036 -34810 60136 -34800
rect 60546 -34810 60636 -34800
rect 60386 -34890 60556 -34810
rect 60626 -34890 60636 -34810
rect 59966 -34900 60326 -34890
rect 59966 -34970 59976 -34900
rect 60316 -34970 60326 -34900
rect 60546 -34910 60636 -34890
rect 59966 -34980 60326 -34970
rect 59566 -35070 59796 -35050
rect 59566 -35080 59576 -35070
rect 59266 -35130 59376 -35120
rect 59516 -35130 59576 -35080
rect 59636 -35130 59796 -35070
rect 59266 -35240 59366 -35130
rect 59266 -35330 59286 -35240
rect 59356 -35330 59366 -35240
rect 59266 -35360 59366 -35330
rect 59516 -35140 59796 -35130
rect 59066 -35480 59076 -35410
rect 59166 -35480 59176 -35410
rect 59066 -35490 59176 -35480
rect 59306 -35430 59386 -35420
rect 59306 -35490 59316 -35430
rect 59376 -35490 59386 -35430
rect 59516 -35470 59596 -35140
rect 60286 -35150 60476 -35140
rect 59906 -35180 60016 -35170
rect 59906 -35360 59916 -35180
rect 60006 -35360 60016 -35180
rect 59906 -35370 60016 -35360
rect 60286 -35290 60306 -35150
rect 60456 -35290 60476 -35150
rect 60286 -35300 60476 -35290
rect 58516 -35740 58796 -35660
rect 59066 -35570 59176 -35560
rect 59066 -35640 59076 -35570
rect 59166 -35640 59176 -35570
rect 59066 -36140 59176 -35640
rect 59306 -35690 59386 -35490
rect 60076 -35480 60196 -35440
rect 60076 -35640 60096 -35480
rect 60176 -35640 60196 -35480
rect 60076 -35680 60196 -35640
rect 59066 -36200 59076 -36140
rect 59166 -36200 59176 -36140
rect 59066 -36210 59176 -36200
rect 59236 -35720 59386 -35690
rect 59236 -35810 59266 -35720
rect 59366 -35810 59386 -35720
rect 59236 -35830 59386 -35810
rect 59906 -35690 60016 -35680
rect 59236 -35960 59376 -35830
rect 59906 -35880 59916 -35690
rect 60006 -35880 60016 -35690
rect 59906 -35890 60016 -35880
rect 60286 -35710 60376 -35300
rect 60556 -35700 60626 -34910
rect 61026 -35220 61136 -34250
rect 61196 -34920 61356 -34910
rect 61196 -35100 61206 -34920
rect 61346 -35100 61356 -34920
rect 61196 -35110 61356 -35100
rect 61026 -35330 61036 -35220
rect 61126 -35330 61136 -35220
rect 61026 -35340 61136 -35330
rect 61246 -35450 61366 -35440
rect 61246 -35460 61276 -35450
rect 61246 -35660 61256 -35460
rect 61356 -35660 61366 -35450
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 61246 -35670 61366 -35660
rect 60466 -35710 60626 -35700
rect 60286 -35770 60406 -35710
rect 60466 -35770 60476 -35710
rect 60536 -35770 60626 -35710
rect 59236 -36050 59266 -35960
rect 59366 -36050 59376 -35960
rect 59236 -36100 59376 -36050
rect 59506 -35910 59606 -35900
rect 59506 -35980 59516 -35910
rect 59596 -35980 59606 -35910
rect 59506 -35990 59606 -35980
rect 59236 -36120 59386 -36100
rect 59236 -36180 59316 -36120
rect 59376 -36180 59386 -36120
rect 58396 -36750 58896 -36250
rect 59236 -36430 59386 -36180
rect 59006 -36500 59086 -36480
rect 59236 -36490 59256 -36430
rect 59366 -36490 59386 -36430
rect 59236 -36500 59386 -36490
rect 59506 -36380 59596 -35990
rect 59986 -36120 60116 -36110
rect 59986 -36180 59996 -36120
rect 60106 -36180 60116 -36120
rect 59506 -36390 59616 -36380
rect 59506 -36460 59546 -36390
rect 59606 -36460 59616 -36390
rect 59006 -36560 59016 -36500
rect 59076 -36560 59086 -36500
rect 59006 -36750 59086 -36560
rect 59506 -36510 59616 -36460
rect 59506 -36570 59546 -36510
rect 59606 -36570 59616 -36510
rect 59796 -36410 59926 -36400
rect 59796 -36520 59806 -36410
rect 59916 -36520 59926 -36410
rect 59796 -36530 59926 -36520
rect 59006 -36840 59126 -36750
rect 59006 -36910 59016 -36840
rect 59076 -36910 59126 -36840
rect 59006 -36990 59126 -36910
rect 59506 -36840 59616 -36570
rect 59506 -36910 59546 -36840
rect 59606 -36910 59616 -36840
rect 59506 -36920 59616 -36910
rect 59986 -36990 60116 -36180
rect 60286 -36670 60376 -35770
rect 60466 -35780 60626 -35770
rect 61486 -35770 61726 -35740
rect 61486 -35820 61496 -35770
rect 61326 -35830 61496 -35820
rect 61326 -35950 61336 -35830
rect 61196 -35960 61336 -35950
rect 61456 -35940 61496 -35830
rect 61696 -35940 61726 -35770
rect 61456 -35960 61726 -35940
rect 61196 -35970 61726 -35960
rect 61196 -36140 61426 -35970
rect 60436 -36430 60536 -36410
rect 60436 -36550 60446 -36430
rect 60526 -36550 60536 -36430
rect 60436 -36560 60536 -36550
rect 60256 -36800 60416 -36670
rect 60256 -36930 60266 -36800
rect 60406 -36930 60416 -36800
rect 60256 -36950 60416 -36930
rect 58956 -37000 59156 -36990
rect 58956 -37180 58966 -37000
rect 59146 -37180 59156 -37000
rect 59986 -37100 59996 -36990
rect 60106 -37100 60116 -36990
rect 61900 -37100 62600 -37000
rect 58956 -37190 59156 -37180
rect 59800 -37200 60300 -37100
rect 61900 -37200 62000 -37100
rect 59800 -37400 59900 -37200
rect 60200 -37400 62000 -37200
rect 59800 -37500 62000 -37400
rect 61900 -37700 62000 -37500
rect 62500 -37700 62600 -37100
rect 61900 -37800 62600 -37700
rect 84700 -38050 85660 -37780
rect 75380 -38150 78900 -38140
rect 75380 -38270 75390 -38150
rect 75550 -38270 78770 -38150
rect 78890 -38270 78900 -38150
rect 75380 -38280 78900 -38270
rect 76900 -38400 77080 -38390
rect 75200 -38427 75380 -38410
rect 75200 -38492 75231 -38427
rect 75322 -38440 75380 -38427
rect 76635 -38440 76739 -38427
rect 75322 -38492 76648 -38440
rect 75200 -38505 76648 -38492
rect 76726 -38505 76739 -38440
rect 75200 -38510 76739 -38505
rect 76635 -38518 76739 -38510
rect 76900 -38540 76910 -38400
rect 77070 -38540 77080 -38400
rect 76900 -38550 77080 -38540
rect 84700 -38480 84960 -38050
rect 85400 -38480 85660 -38050
rect 74451 -38570 74620 -38557
rect 74451 -38674 74477 -38570
rect 74594 -38583 76193 -38570
rect 74594 -38661 76102 -38583
rect 76180 -38661 76193 -38583
rect 74594 -38674 76193 -38661
rect 76770 -38630 78360 -38620
rect 74451 -38687 74620 -38674
rect 76770 -38700 76780 -38630
rect 76860 -38700 78280 -38630
rect 78350 -38700 78360 -38630
rect 84700 -38690 85660 -38480
rect 87880 -38390 88840 -38140
rect 76770 -38710 78360 -38700
rect 76362 -38726 76453 -38713
rect 72810 -38740 73050 -38730
rect 76362 -38739 76375 -38726
rect 68000 -39000 68700 -38900
rect 72600 -38920 72820 -38740
rect 73040 -38750 73080 -38740
rect 73040 -38910 73370 -38750
rect 74711 -38752 76375 -38739
rect 74711 -38830 74724 -38752
rect 74841 -38804 76375 -38752
rect 76440 -38804 76453 -38726
rect 74841 -38817 76453 -38804
rect 77160 -38790 77440 -38780
rect 74841 -38830 74854 -38817
rect 74711 -38843 74854 -38830
rect 73040 -38920 73080 -38910
rect 73210 -38920 75350 -38910
rect 72810 -38930 73050 -38920
rect 68000 -39200 68100 -39000
rect 68600 -39060 68700 -39000
rect 73210 -39020 75220 -38920
rect 75340 -39020 75350 -38920
rect 73210 -39030 75350 -39020
rect 77160 -39040 77170 -38790
rect 77430 -39040 77440 -38790
rect 87880 -38820 88150 -38390
rect 88590 -38820 88840 -38390
rect 77160 -39050 77440 -39040
rect 82760 -39000 87770 -38990
rect 82760 -39010 84870 -39000
rect 68600 -39070 73080 -39060
rect 68600 -39200 72820 -39070
rect 58946 -39270 59146 -39250
rect 58946 -39430 58966 -39270
rect 59126 -39430 59146 -39270
rect 58946 -39450 59146 -39430
rect 59316 -39310 59426 -39250
rect 59316 -39450 59336 -39310
rect 59416 -39450 59426 -39310
rect 58956 -39530 59136 -39450
rect 58956 -39640 58996 -39530
rect 59106 -39640 59136 -39530
rect 58396 -39730 58896 -39640
rect 58956 -39700 59136 -39640
rect 59316 -39680 59426 -39450
rect 59946 -39320 60386 -39200
rect 68000 -39240 72820 -39200
rect 68000 -39300 68700 -39240
rect 72810 -39250 72820 -39240
rect 73040 -39090 73080 -39070
rect 73040 -39100 75100 -39090
rect 73040 -39220 74970 -39100
rect 75090 -39220 75100 -39100
rect 82760 -39100 82780 -39010
rect 82890 -39080 83370 -39010
rect 83740 -39070 84870 -39010
rect 85240 -39070 86330 -39000
rect 86700 -39070 87460 -39000
rect 87750 -39070 87770 -39000
rect 87880 -39050 88840 -38820
rect 83740 -39080 87770 -39070
rect 82890 -39090 87770 -39080
rect 82890 -39100 82910 -39090
rect 82760 -39120 82910 -39100
rect 73040 -39230 75100 -39220
rect 73040 -39240 73080 -39230
rect 73040 -39250 73050 -39240
rect 72810 -39260 73050 -39250
rect 80050 -39270 80460 -39240
rect 59946 -39440 60046 -39320
rect 60126 -39440 60386 -39320
rect 59946 -39490 60386 -39440
rect 66800 -39400 67500 -39300
rect 80050 -39330 80080 -39270
rect 58396 -40090 58486 -39730
rect 58816 -40090 58896 -39730
rect 58996 -40000 59086 -39700
rect 58996 -40060 59006 -40000
rect 59066 -40060 59086 -40000
rect 58996 -40070 59086 -40060
rect 59266 -39730 59426 -39680
rect 59506 -39540 59796 -39500
rect 59506 -39640 59516 -39540
rect 59616 -39640 59796 -39540
rect 59506 -39700 59796 -39640
rect 59266 -39930 59366 -39730
rect 59266 -39990 59286 -39930
rect 59346 -39990 59366 -39930
rect 58396 -40200 58896 -40090
rect 59066 -40240 59176 -40230
rect 59066 -40310 59076 -40240
rect 59166 -40310 59176 -40240
rect 56470 -40838 56555 -40828
rect 56470 -40928 56480 -40838
rect 56550 -40928 56555 -40838
rect 56470 -40938 56555 -40928
rect 56470 -41318 56550 -40938
rect 57760 -40940 57800 -40820
rect 58240 -40940 58280 -40820
rect 57093 -41274 57373 -41264
rect 56470 -41328 56555 -41318
rect 56470 -41378 56480 -41328
rect 56475 -41388 56480 -41378
rect 56550 -41388 56555 -41328
rect 56475 -41398 56555 -41388
rect 57093 -41414 57098 -41274
rect 57368 -41414 57373 -41274
rect 57093 -41424 57373 -41414
rect 55870 -41878 55980 -41438
rect 55870 -41918 55880 -41878
rect 55875 -41958 55880 -41918
rect 55970 -41918 55980 -41878
rect 56060 -41868 56220 -41858
rect 55970 -41958 55975 -41918
rect 55875 -41968 55975 -41958
rect 55590 -42078 55620 -41988
rect 55710 -42078 55720 -41988
rect 56060 -42038 56220 -42028
rect 56060 -42048 56200 -42038
rect 55590 -42088 55720 -42078
rect 56015 -42058 56200 -42048
rect 56015 -42208 56020 -42058
rect 56080 -42208 56200 -42058
rect 56644 -42068 57008 -42063
rect 55215 -42218 55325 -42208
rect 56015 -42218 56085 -42208
rect 55215 -42318 55220 -42218
rect 55320 -42318 55325 -42218
rect 56644 -42286 56654 -42068
rect 56998 -42286 57008 -42068
rect 56644 -42291 57008 -42286
rect 55215 -42328 55325 -42318
rect 55315 -42528 55475 -42518
rect 55315 -42668 55320 -42528
rect 55470 -42668 55475 -42528
rect 55315 -42678 55475 -42668
rect 43100 -43100 56200 -43000
rect 43100 -43800 43200 -43100
rect 44300 -43500 55500 -43100
rect 56100 -43500 56200 -43100
rect 44300 -43600 56200 -43500
rect 44300 -43800 44400 -43600
rect 43100 -43900 44400 -43800
rect 51400 -44080 55800 -44000
rect 51400 -44100 55500 -44080
rect 51400 -44300 51500 -44100
rect 52500 -44300 55500 -44100
rect 51400 -44360 55500 -44300
rect 55720 -44360 55800 -44080
rect 51400 -44400 55800 -44360
rect 55420 -44440 55800 -44400
rect 47800 -44640 48100 -44620
rect 47800 -45060 47820 -44640
rect 48080 -44720 48100 -44640
rect 48080 -44740 53800 -44720
rect 48080 -44940 53480 -44740
rect 53780 -44940 53800 -44740
rect 56496 -44780 57026 -44775
rect 48080 -44960 53800 -44940
rect 55955 -44938 56045 -44928
rect 48080 -45060 48100 -44960
rect 53515 -45058 53645 -45048
rect 47800 -45080 48100 -45060
rect 53510 -45168 53520 -45058
rect 53640 -45168 53645 -45058
rect 55955 -45088 55960 -44938
rect 56040 -45088 56200 -44938
rect 56496 -45030 56506 -44780
rect 57016 -45030 57026 -44780
rect 56496 -45035 57026 -45030
rect 55955 -45098 56200 -45088
rect 53510 -45178 53645 -45168
rect 55275 -45118 55490 -45108
rect 53045 -45358 53255 -45348
rect 53045 -47108 53050 -45358
rect 53250 -47108 53255 -45358
rect 53045 -47118 53255 -47108
rect 53510 -47318 53630 -45178
rect 55275 -45208 55280 -45118
rect 55400 -45208 55490 -45118
rect 56060 -45138 56200 -45098
rect 56060 -45148 56220 -45138
rect 55275 -45218 55490 -45208
rect 55220 -45458 55325 -45448
rect 55220 -45628 55230 -45458
rect 55320 -45628 55325 -45458
rect 55220 -45638 55325 -45628
rect 55015 -46248 55125 -46238
rect 55015 -46328 55020 -46248
rect 55120 -46328 55125 -46248
rect 55015 -46338 55125 -46328
rect 55220 -46938 55310 -45638
rect 55215 -46948 55315 -46938
rect 55215 -47118 55220 -46948
rect 55310 -47038 55315 -46948
rect 55400 -46948 55490 -45218
rect 55875 -45218 55990 -45208
rect 55875 -45258 55880 -45218
rect 55870 -45298 55880 -45258
rect 55970 -45298 55990 -45218
rect 55870 -45378 55990 -45298
rect 56060 -45318 56220 -45308
rect 55590 -45468 55720 -45458
rect 55590 -45598 55600 -45468
rect 55710 -45598 55720 -45468
rect 55400 -46958 55510 -46948
rect 55310 -47118 55320 -47038
rect 55400 -47118 55410 -46958
rect 55215 -47128 55320 -47118
rect 53505 -47328 53635 -47318
rect 53505 -47448 53510 -47328
rect 53630 -47448 53635 -47328
rect 53505 -47458 53635 -47448
rect 55220 -47608 55320 -47128
rect 55405 -47128 55410 -47118
rect 55500 -47128 55510 -46958
rect 55405 -47138 55510 -47128
rect 55590 -47388 55720 -45598
rect 55870 -45758 55980 -45378
rect 57093 -45764 57373 -45754
rect 56475 -45788 56555 -45778
rect 56470 -45848 56480 -45788
rect 56550 -45848 56555 -45788
rect 56470 -45858 56555 -45848
rect 55870 -46238 55980 -45868
rect 55870 -46328 55880 -46238
rect 55970 -46328 55980 -46238
rect 55870 -46728 55980 -46328
rect 56470 -46228 56550 -45858
rect 57093 -45904 57098 -45764
rect 57368 -45904 57373 -45764
rect 57093 -45914 57373 -45904
rect 57760 -46220 58280 -40940
rect 58516 -40860 58796 -40790
rect 58516 -41060 58556 -40860
rect 58756 -41060 58796 -40860
rect 59066 -40810 59176 -40310
rect 59266 -40420 59366 -39990
rect 59536 -39890 59616 -39700
rect 59536 -39950 59546 -39890
rect 59606 -39950 59616 -39890
rect 59536 -40010 59616 -39950
rect 59536 -40070 59546 -40010
rect 59606 -40070 59616 -40010
rect 59536 -40080 59616 -40070
rect 59266 -40430 59376 -40420
rect 59266 -40520 59286 -40430
rect 59366 -40520 59376 -40430
rect 59736 -40450 59796 -39700
rect 59856 -39940 59976 -39930
rect 59856 -40030 59866 -39940
rect 59966 -40030 59976 -39940
rect 59856 -40040 59976 -40030
rect 60036 -40120 60136 -39490
rect 61026 -39520 61136 -39510
rect 61026 -39650 61056 -39520
rect 61126 -39650 61136 -39520
rect 60436 -39920 60536 -39910
rect 60436 -40020 60446 -39920
rect 60526 -40020 60536 -39920
rect 60436 -40030 60536 -40020
rect 60036 -40200 60046 -40120
rect 60126 -40200 60136 -40120
rect 60036 -40210 60136 -40200
rect 60546 -40210 60636 -40200
rect 60386 -40290 60556 -40210
rect 60626 -40290 60636 -40210
rect 59966 -40300 60326 -40290
rect 59966 -40370 59976 -40300
rect 60316 -40370 60326 -40300
rect 60546 -40310 60636 -40290
rect 59966 -40380 60326 -40370
rect 59566 -40470 59796 -40450
rect 59566 -40480 59576 -40470
rect 59266 -40530 59376 -40520
rect 59516 -40530 59576 -40480
rect 59636 -40530 59796 -40470
rect 59266 -40640 59366 -40530
rect 59266 -40730 59286 -40640
rect 59356 -40730 59366 -40640
rect 59266 -40760 59366 -40730
rect 59516 -40540 59796 -40530
rect 59066 -40880 59076 -40810
rect 59166 -40880 59176 -40810
rect 59066 -40890 59176 -40880
rect 59306 -40830 59386 -40820
rect 59306 -40890 59316 -40830
rect 59376 -40890 59386 -40830
rect 59516 -40870 59596 -40540
rect 60286 -40550 60476 -40540
rect 59906 -40580 60016 -40570
rect 59906 -40760 59916 -40580
rect 60006 -40760 60016 -40580
rect 59906 -40770 60016 -40760
rect 60286 -40690 60306 -40550
rect 60456 -40690 60476 -40550
rect 60286 -40700 60476 -40690
rect 58516 -41140 58796 -41060
rect 59066 -40970 59176 -40960
rect 59066 -41040 59076 -40970
rect 59166 -41040 59176 -40970
rect 59066 -41540 59176 -41040
rect 59306 -41090 59386 -40890
rect 60076 -40880 60196 -40840
rect 60076 -41040 60096 -40880
rect 60176 -41040 60196 -40880
rect 60076 -41080 60196 -41040
rect 59066 -41600 59076 -41540
rect 59166 -41600 59176 -41540
rect 59066 -41610 59176 -41600
rect 59236 -41120 59386 -41090
rect 59236 -41210 59266 -41120
rect 59366 -41210 59386 -41120
rect 59236 -41230 59386 -41210
rect 59906 -41090 60016 -41080
rect 59236 -41360 59376 -41230
rect 59906 -41280 59916 -41090
rect 60006 -41280 60016 -41090
rect 59906 -41290 60016 -41280
rect 60286 -41110 60376 -40700
rect 60556 -41100 60626 -40310
rect 61026 -40620 61136 -39650
rect 66800 -39600 66900 -39400
rect 67400 -39560 67500 -39400
rect 79060 -39350 80080 -39330
rect 73960 -39430 77330 -39420
rect 73960 -39490 73970 -39430
rect 74090 -39440 77330 -39430
rect 74090 -39490 77230 -39440
rect 73960 -39500 77230 -39490
rect 77310 -39500 77330 -39440
rect 77200 -39520 77330 -39500
rect 79060 -39510 79080 -39350
rect 79250 -39510 80080 -39350
rect 79060 -39520 80080 -39510
rect 72810 -39560 73050 -39550
rect 67400 -39600 72820 -39560
rect 65800 -39800 66500 -39700
rect 66800 -39740 72820 -39600
rect 73040 -39570 73200 -39560
rect 76910 -39570 77070 -39560
rect 73040 -39580 74850 -39570
rect 73040 -39720 74720 -39580
rect 74840 -39720 74850 -39580
rect 73040 -39730 74850 -39720
rect 76910 -39720 76920 -39570
rect 77060 -39720 77070 -39570
rect 80050 -39580 80080 -39520
rect 80430 -39580 80460 -39270
rect 80050 -39590 80460 -39580
rect 89580 -39580 92160 -39550
rect 76910 -39730 77070 -39720
rect 80050 -39680 80460 -39650
rect 73040 -39740 73200 -39730
rect 72810 -39750 73050 -39740
rect 65800 -39839 65900 -39800
rect 65799 -40000 65900 -39839
rect 66400 -39839 66500 -39800
rect 74960 -39780 76620 -39770
rect 66400 -39840 72399 -39839
rect 72810 -39840 73050 -39830
rect 66400 -40000 72820 -39840
rect 65799 -40019 72820 -40000
rect 65800 -40100 66500 -40019
rect 66600 -40020 72820 -40019
rect 73040 -39850 73200 -39840
rect 74960 -39850 74980 -39780
rect 75080 -39790 76620 -39780
rect 77130 -39780 77270 -39770
rect 77130 -39790 77170 -39780
rect 75080 -39850 77170 -39790
rect 77260 -39850 77270 -39780
rect 80050 -39820 80080 -39680
rect 73040 -39860 74600 -39850
rect 74960 -39860 77270 -39850
rect 78570 -39840 80080 -39820
rect 73040 -40000 74470 -39860
rect 74590 -40000 74600 -39860
rect 78570 -39900 78580 -39840
rect 78640 -39900 80080 -39840
rect 78570 -39920 80080 -39900
rect 73040 -40010 74600 -40000
rect 73040 -40020 73200 -40010
rect 72810 -40030 73050 -40020
rect 80050 -40060 80080 -39920
rect 80430 -40060 80460 -39680
rect 89580 -39690 91780 -39580
rect 84220 -39700 91780 -39690
rect 80050 -40090 80460 -40060
rect 83000 -39830 83640 -39700
rect 84220 -39810 84230 -39700
rect 84310 -39810 85710 -39700
rect 85790 -39810 87180 -39700
rect 87260 -39810 88650 -39700
rect 88730 -39810 91780 -39700
rect 84220 -39820 91780 -39810
rect 64800 -40200 65500 -40100
rect 74460 -40110 77490 -40100
rect 74460 -40180 74470 -40110
rect 74590 -40180 77410 -40110
rect 77480 -40180 77490 -40110
rect 74460 -40190 77490 -40180
rect 79400 -40150 79690 -40140
rect 61196 -40320 61356 -40310
rect 61196 -40500 61206 -40320
rect 61346 -40500 61356 -40320
rect 64800 -40400 64900 -40200
rect 65400 -40300 65500 -40200
rect 72810 -40300 73050 -40290
rect 65400 -40400 72820 -40300
rect 64800 -40480 72820 -40400
rect 73040 -40310 73200 -40300
rect 73040 -40380 74350 -40310
rect 73040 -40390 77850 -40380
rect 73040 -40450 74220 -40390
rect 74340 -40450 77780 -40390
rect 77840 -40450 77850 -40390
rect 79400 -40390 79410 -40150
rect 79680 -40390 79690 -40150
rect 83000 -40180 83150 -39830
rect 83510 -40180 83640 -39830
rect 89580 -39960 91780 -39820
rect 92130 -39960 92160 -39580
rect 79400 -40400 79690 -40390
rect 81110 -40250 81600 -40220
rect 73040 -40460 77850 -40450
rect 73040 -40470 74350 -40460
rect 73040 -40480 73200 -40470
rect 64800 -40500 65500 -40480
rect 72810 -40490 73050 -40480
rect 61196 -40510 61356 -40500
rect 81110 -40510 81140 -40250
rect 81570 -40510 81600 -40250
rect 83000 -40290 83640 -40180
rect 87520 -40240 88480 -39980
rect 89580 -39990 92160 -39960
rect 75210 -40540 77530 -40530
rect 81110 -40540 81600 -40510
rect 75210 -40610 75220 -40540
rect 75340 -40610 77450 -40540
rect 77520 -40610 77530 -40540
rect 75210 -40620 77530 -40610
rect 87520 -40590 87830 -40240
rect 88190 -40590 88480 -40240
rect 61026 -40730 61036 -40620
rect 61126 -40730 61136 -40620
rect 61026 -40740 61136 -40730
rect 63600 -40660 64200 -40620
rect 72810 -40660 73050 -40650
rect 63600 -40800 63640 -40660
rect 64160 -40800 72820 -40660
rect 63600 -40840 72820 -40800
rect 73040 -40670 73200 -40660
rect 73040 -40680 74100 -40670
rect 73040 -40820 73970 -40680
rect 74090 -40820 74100 -40680
rect 73040 -40830 74100 -40820
rect 76910 -40820 77070 -40810
rect 73040 -40840 73200 -40830
rect 61246 -40850 61366 -40840
rect 72810 -40850 73050 -40840
rect 61246 -40860 61276 -40850
rect 61246 -41060 61256 -40860
rect 61356 -41060 61366 -40850
rect 61246 -41070 61366 -41060
rect 62800 -41000 63400 -40900
rect 76910 -40960 76920 -40820
rect 77060 -40960 77070 -40820
rect 76910 -40970 77070 -40960
rect 80050 -40910 82980 -40880
rect 87520 -40890 88480 -40590
rect 60466 -41110 60626 -41100
rect 60286 -41170 60406 -41110
rect 60466 -41170 60476 -41110
rect 60536 -41170 60626 -41110
rect 59236 -41450 59266 -41360
rect 59366 -41450 59376 -41360
rect 59236 -41500 59376 -41450
rect 59506 -41310 59606 -41300
rect 59506 -41380 59516 -41310
rect 59596 -41380 59606 -41310
rect 59506 -41390 59606 -41380
rect 59236 -41520 59386 -41500
rect 59236 -41580 59316 -41520
rect 59376 -41580 59386 -41520
rect 58396 -42150 58896 -41650
rect 59236 -41830 59386 -41580
rect 59006 -41900 59086 -41880
rect 59236 -41890 59256 -41830
rect 59366 -41890 59386 -41830
rect 59236 -41900 59386 -41890
rect 59506 -41780 59596 -41390
rect 59986 -41520 60116 -41510
rect 59986 -41580 59996 -41520
rect 60106 -41580 60116 -41520
rect 59506 -41790 59616 -41780
rect 59506 -41860 59546 -41790
rect 59606 -41860 59616 -41790
rect 59006 -41960 59016 -41900
rect 59076 -41960 59086 -41900
rect 59006 -42150 59086 -41960
rect 59506 -41910 59616 -41860
rect 59506 -41970 59546 -41910
rect 59606 -41970 59616 -41910
rect 59796 -41810 59926 -41800
rect 59796 -41920 59806 -41810
rect 59916 -41920 59926 -41810
rect 59796 -41930 59926 -41920
rect 59006 -42240 59126 -42150
rect 59006 -42310 59016 -42240
rect 59076 -42310 59126 -42240
rect 59006 -42390 59126 -42310
rect 59506 -42240 59616 -41970
rect 59506 -42310 59546 -42240
rect 59606 -42310 59616 -42240
rect 59506 -42320 59616 -42310
rect 59986 -42390 60116 -41580
rect 60286 -42070 60376 -41170
rect 60466 -41180 60626 -41170
rect 61486 -41170 61726 -41140
rect 61486 -41220 61496 -41170
rect 61326 -41230 61496 -41220
rect 61326 -41350 61336 -41230
rect 61196 -41360 61336 -41350
rect 61456 -41340 61496 -41230
rect 61696 -41340 61726 -41170
rect 61456 -41360 61726 -41340
rect 61196 -41370 61726 -41360
rect 62800 -41300 62900 -41000
rect 63300 -41060 73200 -41000
rect 80050 -41020 80080 -40910
rect 63300 -41240 72820 -41060
rect 73040 -41080 73200 -41060
rect 78660 -41030 80080 -41020
rect 73040 -41090 73850 -41080
rect 73040 -41220 73720 -41090
rect 73840 -41220 73850 -41090
rect 73040 -41230 73850 -41220
rect 75210 -41160 77540 -41150
rect 73040 -41240 73200 -41230
rect 63300 -41300 73200 -41240
rect 75210 -41240 75220 -41160
rect 75340 -41240 77450 -41160
rect 77530 -41240 77540 -41160
rect 78660 -41180 78670 -41030
rect 78780 -41180 80080 -41030
rect 78660 -41190 80080 -41180
rect 75210 -41250 77540 -41240
rect 80050 -41290 80080 -41190
rect 80430 -41290 82460 -40910
rect 82950 -41290 82980 -40910
rect 61196 -41540 61426 -41370
rect 62800 -41400 63400 -41300
rect 74460 -41320 77850 -41310
rect 80050 -41320 82980 -41290
rect 74460 -41380 74470 -41320
rect 74590 -41380 77780 -41320
rect 77840 -41380 77850 -41320
rect 74460 -41390 77850 -41380
rect 79400 -41380 79690 -41370
rect 61900 -41500 62600 -41400
rect 61900 -41700 62000 -41500
rect 62500 -41510 73100 -41500
rect 62500 -41690 72820 -41510
rect 73040 -41520 73100 -41510
rect 73040 -41530 73600 -41520
rect 73040 -41670 73470 -41530
rect 73590 -41670 73600 -41530
rect 79400 -41620 79410 -41380
rect 79680 -41620 79690 -41380
rect 73040 -41680 73600 -41670
rect 74710 -41630 77850 -41620
rect 79400 -41630 79690 -41620
rect 73040 -41690 73100 -41680
rect 62500 -41700 73100 -41690
rect 74710 -41690 74720 -41630
rect 74840 -41690 77780 -41630
rect 77840 -41690 77850 -41630
rect 74710 -41700 77850 -41690
rect 61900 -41800 62600 -41700
rect 75210 -41770 77590 -41760
rect 60436 -41830 60536 -41810
rect 60436 -41950 60446 -41830
rect 60526 -41950 60536 -41830
rect 75210 -41860 75220 -41770
rect 75340 -41860 77490 -41770
rect 77580 -41860 77590 -41770
rect 75210 -41870 77590 -41860
rect 72810 -41880 73050 -41870
rect 72810 -41900 72820 -41880
rect 60436 -41960 60536 -41950
rect 72600 -42060 72820 -41900
rect 73040 -41890 73050 -41880
rect 73040 -41900 73350 -41890
rect 73040 -42040 73220 -41900
rect 73340 -42040 73350 -41900
rect 73040 -42050 73350 -42040
rect 73040 -42060 73200 -42050
rect 60256 -42200 60416 -42070
rect 60256 -42330 60266 -42200
rect 60406 -42330 60416 -42200
rect 60256 -42350 60416 -42330
rect 58956 -42400 59156 -42390
rect 58956 -42580 58966 -42400
rect 59146 -42580 59156 -42400
rect 59986 -42500 59996 -42390
rect 60106 -42500 60116 -42390
rect 59986 -42510 60116 -42500
rect 58956 -42590 59156 -42580
rect 72600 -42600 73200 -42060
rect 76910 -42060 77070 -42050
rect 76910 -42220 76920 -42060
rect 77060 -42220 77070 -42060
rect 74960 -42270 76850 -42260
rect 74960 -42330 74970 -42270
rect 75090 -42280 76850 -42270
rect 77130 -42270 77850 -42260
rect 77130 -42280 77780 -42270
rect 75090 -42330 77780 -42280
rect 77840 -42330 77850 -42270
rect 74960 -42340 77850 -42330
rect 76850 -42350 77130 -42340
rect 78130 -42360 79170 -42340
rect 78130 -42370 79050 -42360
rect 75210 -42410 76790 -42400
rect 77190 -42410 77570 -42400
rect 75210 -42500 75220 -42410
rect 75340 -42500 77470 -42410
rect 77560 -42500 77570 -42410
rect 78130 -42470 78160 -42370
rect 78260 -42470 79050 -42370
rect 79150 -42470 79170 -42360
rect 78130 -42490 79170 -42470
rect 75210 -42510 77570 -42500
rect 59600 -42800 73200 -42600
rect 59600 -43400 59800 -42800
rect 60400 -43400 73200 -42800
rect 79400 -42640 79690 -42630
rect 79400 -42880 79410 -42640
rect 79680 -42880 79690 -42640
rect 82790 -42740 91440 -42710
rect 79400 -42890 79690 -42880
rect 78850 -42920 79000 -42900
rect 73710 -42930 77550 -42920
rect 73710 -43000 73720 -42930
rect 73840 -42990 77470 -42930
rect 77540 -42990 77550 -42930
rect 73840 -43000 77550 -42990
rect 73710 -43010 73850 -43000
rect 77740 -43050 77930 -43040
rect 77740 -43060 77860 -43050
rect 76200 -43070 77860 -43060
rect 76200 -43130 76210 -43070
rect 76340 -43110 77860 -43070
rect 77920 -43110 77930 -43050
rect 76340 -43120 77930 -43110
rect 76340 -43130 76350 -43120
rect 76200 -43140 76350 -43130
rect 75210 -43190 76140 -43180
rect 75210 -43250 75220 -43190
rect 75340 -43200 76140 -43190
rect 76410 -43190 78030 -43180
rect 76410 -43200 77960 -43190
rect 75340 -43240 77960 -43200
rect 75340 -43250 76840 -43240
rect 75210 -43260 76840 -43250
rect 77120 -43250 77960 -43240
rect 78020 -43250 78030 -43190
rect 78850 -43210 78860 -42920
rect 78980 -43000 79000 -42920
rect 79980 -42910 82520 -42880
rect 79980 -43000 80010 -42910
rect 78980 -43210 80010 -43000
rect 78850 -43220 80010 -43210
rect 77120 -43260 78030 -43250
rect 79980 -43290 80010 -43220
rect 80360 -43290 82120 -42910
rect 82490 -43290 82520 -42910
rect 59600 -43600 73200 -43400
rect 76910 -43310 77070 -43300
rect 76910 -43450 76920 -43310
rect 77060 -43450 77070 -43310
rect 79980 -43320 82520 -43290
rect 82790 -43310 82820 -42740
rect 91410 -43310 91440 -42740
rect 82790 -43340 91440 -43310
rect 76910 -43460 77070 -43450
rect 85310 -43450 90770 -43440
rect 85310 -43540 85320 -43450
rect 85390 -43540 85590 -43450
rect 86480 -43540 87040 -43450
rect 87920 -43540 88510 -43450
rect 89390 -43540 89980 -43450
rect 90760 -43540 90770 -43450
rect 85310 -43550 90770 -43540
rect 75210 -43620 78040 -43610
rect 75210 -43680 75220 -43620
rect 75340 -43680 77970 -43620
rect 78030 -43680 78040 -43620
rect 75210 -43690 78040 -43680
rect 73960 -43760 77510 -43750
rect 73960 -43830 73970 -43760
rect 74090 -43830 77430 -43760
rect 77500 -43830 77510 -43760
rect 73960 -43840 77510 -43830
rect 79400 -43860 79690 -43850
rect 79400 -44100 79410 -43860
rect 79680 -44100 79690 -43860
rect 82630 -43890 83110 -43880
rect 82630 -44000 82640 -43890
rect 82720 -44000 83040 -43890
rect 83100 -44000 83110 -43890
rect 82630 -44010 83110 -44000
rect 79400 -44110 79690 -44100
rect 91750 -44080 92160 -44050
rect 91750 -44220 91780 -44080
rect 86790 -44230 91780 -44220
rect 76480 -44250 77490 -44240
rect 76480 -44310 76490 -44250
rect 76610 -44290 77490 -44250
rect 76610 -44310 78040 -44290
rect 76480 -44320 76620 -44310
rect 77410 -44350 78040 -44310
rect 86790 -44310 86800 -44230
rect 86870 -44310 88270 -44230
rect 88340 -44310 89750 -44230
rect 89810 -44310 91210 -44230
rect 91280 -44310 91780 -44230
rect 86790 -44320 91780 -44310
rect 73460 -44380 73610 -44370
rect 73460 -44440 73470 -44380
rect 73590 -44410 77340 -44380
rect 73590 -44420 77830 -44410
rect 73590 -44440 77760 -44420
rect 73460 -44450 77760 -44440
rect 73460 -44460 73610 -44450
rect 77150 -44480 77760 -44450
rect 77820 -44480 77830 -44420
rect 77960 -44470 77970 -44350
rect 78030 -44470 78040 -44350
rect 77960 -44480 78040 -44470
rect 82790 -44440 91440 -44410
rect 77150 -44490 77830 -44480
rect 76910 -44520 77070 -44510
rect 58946 -44670 59146 -44650
rect 58946 -44830 58966 -44670
rect 59126 -44830 59146 -44670
rect 58946 -44850 59146 -44830
rect 59316 -44710 59426 -44650
rect 59316 -44850 59336 -44710
rect 59416 -44850 59426 -44710
rect 58956 -44930 59136 -44850
rect 58956 -45040 58996 -44930
rect 59106 -45040 59136 -44930
rect 58396 -45130 58896 -45040
rect 58956 -45100 59136 -45040
rect 59316 -45080 59426 -44850
rect 59946 -44720 60386 -44600
rect 76910 -44610 76920 -44520
rect 77060 -44610 77070 -44520
rect 76910 -44620 77070 -44610
rect 59946 -44840 60046 -44720
rect 60126 -44840 60386 -44720
rect 73960 -44740 77830 -44730
rect 73960 -44800 73970 -44740
rect 74090 -44800 77760 -44740
rect 77820 -44800 77830 -44740
rect 73960 -44810 77830 -44800
rect 78770 -44770 78930 -44760
rect 59946 -44890 60386 -44840
rect 77950 -44850 78030 -44840
rect 77950 -44870 77960 -44850
rect 76480 -44880 77960 -44870
rect 58396 -45490 58486 -45130
rect 58816 -45490 58896 -45130
rect 58996 -45400 59086 -45100
rect 58996 -45460 59006 -45400
rect 59066 -45460 59086 -45400
rect 58996 -45470 59086 -45460
rect 59266 -45130 59426 -45080
rect 59506 -44940 59796 -44900
rect 59506 -45040 59516 -44940
rect 59616 -45040 59796 -44940
rect 59506 -45100 59796 -45040
rect 59266 -45330 59366 -45130
rect 59266 -45390 59286 -45330
rect 59346 -45390 59366 -45330
rect 58396 -45600 58896 -45490
rect 59066 -45640 59176 -45630
rect 59066 -45710 59076 -45640
rect 59166 -45710 59176 -45640
rect 56470 -46238 56555 -46228
rect 56470 -46328 56480 -46238
rect 56550 -46328 56555 -46238
rect 56470 -46338 56555 -46328
rect 56470 -46718 56550 -46338
rect 57760 -46340 57800 -46220
rect 58240 -46340 58280 -46220
rect 57093 -46674 57373 -46664
rect 56470 -46728 56555 -46718
rect 56470 -46778 56480 -46728
rect 56475 -46788 56480 -46778
rect 56550 -46788 56555 -46728
rect 56475 -46798 56555 -46788
rect 57093 -46814 57098 -46674
rect 57368 -46814 57373 -46674
rect 57093 -46824 57373 -46814
rect 55870 -47278 55980 -46838
rect 55870 -47318 55880 -47278
rect 55875 -47358 55880 -47318
rect 55970 -47318 55980 -47278
rect 56060 -47268 56220 -47258
rect 55970 -47358 55975 -47318
rect 55875 -47368 55975 -47358
rect 55590 -47478 55620 -47388
rect 55710 -47478 55720 -47388
rect 56060 -47438 56220 -47428
rect 56060 -47448 56200 -47438
rect 55590 -47488 55720 -47478
rect 56015 -47458 56200 -47448
rect 56015 -47608 56020 -47458
rect 56080 -47608 56200 -47458
rect 56644 -47468 57008 -47463
rect 55215 -47618 55325 -47608
rect 56015 -47618 56085 -47608
rect 55215 -47718 55220 -47618
rect 55320 -47718 55325 -47618
rect 56644 -47686 56654 -47468
rect 56998 -47686 57008 -47468
rect 56644 -47691 57008 -47686
rect 55215 -47728 55325 -47718
rect 55315 -47928 55475 -47918
rect 55315 -48068 55320 -47928
rect 55470 -48068 55475 -47928
rect 55315 -48078 55475 -48068
rect 14000 -50000 25000 -49000
rect 43700 -48400 44400 -48300
rect 43700 -49000 43800 -48400
rect 44300 -48500 56200 -48400
rect 44300 -48900 55500 -48500
rect 56100 -48900 56200 -48500
rect 44300 -49000 56200 -48900
rect 43700 -49100 44400 -49000
rect 51400 -49480 55800 -49400
rect 51400 -49500 55460 -49480
rect 51400 -49700 51500 -49500
rect 52500 -49700 55460 -49500
rect 51400 -49760 55460 -49700
rect 55720 -49760 55800 -49480
rect 51400 -49800 55800 -49760
rect 55380 -49840 55800 -49800
rect 47720 -49980 48100 -49960
rect 47720 -50480 47740 -49980
rect 48080 -50120 48100 -49980
rect 48080 -50140 53800 -50120
rect 48080 -50340 53460 -50140
rect 53780 -50340 53800 -50140
rect 56496 -50180 57026 -50175
rect 48080 -50360 53800 -50340
rect 55955 -50338 56045 -50328
rect 48080 -50480 48100 -50360
rect 53515 -50458 53645 -50448
rect 47720 -50500 48100 -50480
rect 53510 -50568 53520 -50458
rect 53640 -50568 53645 -50458
rect 55955 -50488 55960 -50338
rect 56040 -50488 56200 -50338
rect 56496 -50430 56506 -50180
rect 57016 -50430 57026 -50180
rect 56496 -50435 57026 -50430
rect 55955 -50498 56200 -50488
rect 53510 -50578 53645 -50568
rect 55275 -50518 55490 -50508
rect 53045 -50758 53255 -50748
rect 53045 -52508 53050 -50758
rect 53250 -52508 53255 -50758
rect 53045 -52518 53255 -52508
rect 53510 -52718 53630 -50578
rect 55275 -50608 55280 -50518
rect 55400 -50608 55490 -50518
rect 56060 -50538 56200 -50498
rect 56060 -50548 56220 -50538
rect 55275 -50618 55490 -50608
rect 55220 -50858 55325 -50848
rect 55220 -51028 55230 -50858
rect 55320 -51028 55325 -50858
rect 55220 -51038 55325 -51028
rect 55015 -51648 55125 -51638
rect 55015 -51728 55020 -51648
rect 55120 -51728 55125 -51648
rect 55015 -51738 55125 -51728
rect 55220 -52338 55310 -51038
rect 55215 -52348 55315 -52338
rect 55215 -52518 55220 -52348
rect 55310 -52438 55315 -52348
rect 55400 -52348 55490 -50618
rect 55875 -50618 55990 -50608
rect 55875 -50658 55880 -50618
rect 55870 -50698 55880 -50658
rect 55970 -50698 55990 -50618
rect 55870 -50778 55990 -50698
rect 56060 -50718 56220 -50708
rect 55590 -50868 55720 -50858
rect 55590 -50998 55600 -50868
rect 55710 -50998 55720 -50868
rect 55400 -52358 55510 -52348
rect 55310 -52518 55320 -52438
rect 55400 -52518 55410 -52358
rect 55215 -52528 55320 -52518
rect 53505 -52728 53635 -52718
rect 53505 -52848 53510 -52728
rect 53630 -52848 53635 -52728
rect 53505 -52858 53635 -52848
rect 55220 -53008 55320 -52528
rect 55405 -52528 55410 -52518
rect 55500 -52528 55510 -52358
rect 55405 -52538 55510 -52528
rect 55590 -52788 55720 -50998
rect 55870 -51158 55980 -50778
rect 57093 -51164 57373 -51154
rect 56475 -51188 56555 -51178
rect 56470 -51248 56480 -51188
rect 56550 -51248 56555 -51188
rect 56470 -51258 56555 -51248
rect 55870 -51638 55980 -51268
rect 55870 -51728 55880 -51638
rect 55970 -51728 55980 -51638
rect 55870 -52128 55980 -51728
rect 56470 -51628 56550 -51258
rect 57093 -51304 57098 -51164
rect 57368 -51304 57373 -51164
rect 57093 -51314 57373 -51304
rect 57760 -51620 58280 -46340
rect 58516 -46260 58796 -46190
rect 58516 -46460 58556 -46260
rect 58756 -46460 58796 -46260
rect 59066 -46210 59176 -45710
rect 59266 -45820 59366 -45390
rect 59536 -45290 59616 -45100
rect 59536 -45350 59546 -45290
rect 59606 -45350 59616 -45290
rect 59536 -45410 59616 -45350
rect 59536 -45470 59546 -45410
rect 59606 -45470 59616 -45410
rect 59536 -45480 59616 -45470
rect 59266 -45830 59376 -45820
rect 59266 -45920 59286 -45830
rect 59366 -45920 59376 -45830
rect 59736 -45850 59796 -45100
rect 59856 -45340 59976 -45330
rect 59856 -45430 59866 -45340
rect 59966 -45430 59976 -45340
rect 59856 -45440 59976 -45430
rect 60036 -45520 60136 -44890
rect 61026 -44920 61136 -44910
rect 61026 -45050 61056 -44920
rect 61126 -45050 61136 -44920
rect 76480 -44950 76490 -44880
rect 76610 -44920 77960 -44880
rect 78020 -44920 78030 -44850
rect 78770 -44890 78780 -44770
rect 78920 -44800 79170 -44770
rect 78920 -44870 79070 -44800
rect 79140 -44870 79170 -44800
rect 78920 -44890 79170 -44870
rect 78770 -44900 78930 -44890
rect 76610 -44930 78030 -44920
rect 76610 -44950 77530 -44930
rect 76480 -44960 77530 -44950
rect 82790 -45010 82820 -44440
rect 91410 -45010 91440 -44440
rect 91750 -44460 91780 -44320
rect 92130 -44460 92160 -44080
rect 91750 -44490 92160 -44460
rect 82790 -45040 91440 -45010
rect 60436 -45320 60536 -45310
rect 60436 -45420 60446 -45320
rect 60526 -45420 60536 -45320
rect 60436 -45430 60536 -45420
rect 60036 -45600 60046 -45520
rect 60126 -45600 60136 -45520
rect 60036 -45610 60136 -45600
rect 60546 -45610 60636 -45600
rect 60386 -45690 60556 -45610
rect 60626 -45690 60636 -45610
rect 59966 -45700 60326 -45690
rect 59966 -45770 59976 -45700
rect 60316 -45770 60326 -45700
rect 60546 -45710 60636 -45690
rect 59966 -45780 60326 -45770
rect 59566 -45870 59796 -45850
rect 59566 -45880 59576 -45870
rect 59266 -45930 59376 -45920
rect 59516 -45930 59576 -45880
rect 59636 -45930 59796 -45870
rect 59266 -46040 59366 -45930
rect 59266 -46130 59286 -46040
rect 59356 -46130 59366 -46040
rect 59266 -46160 59366 -46130
rect 59516 -45940 59796 -45930
rect 59066 -46280 59076 -46210
rect 59166 -46280 59176 -46210
rect 59066 -46290 59176 -46280
rect 59306 -46230 59386 -46220
rect 59306 -46290 59316 -46230
rect 59376 -46290 59386 -46230
rect 59516 -46270 59596 -45940
rect 60286 -45950 60476 -45940
rect 59906 -45980 60016 -45970
rect 59906 -46160 59916 -45980
rect 60006 -46160 60016 -45980
rect 59906 -46170 60016 -46160
rect 60286 -46090 60306 -45950
rect 60456 -46090 60476 -45950
rect 60286 -46100 60476 -46090
rect 58516 -46540 58796 -46460
rect 59066 -46370 59176 -46360
rect 59066 -46440 59076 -46370
rect 59166 -46440 59176 -46370
rect 59066 -46940 59176 -46440
rect 59306 -46490 59386 -46290
rect 60076 -46280 60196 -46240
rect 60076 -46440 60096 -46280
rect 60176 -46440 60196 -46280
rect 60076 -46480 60196 -46440
rect 59066 -47000 59076 -46940
rect 59166 -47000 59176 -46940
rect 59066 -47010 59176 -47000
rect 59236 -46520 59386 -46490
rect 59236 -46610 59266 -46520
rect 59366 -46610 59386 -46520
rect 59236 -46630 59386 -46610
rect 59906 -46490 60016 -46480
rect 59236 -46760 59376 -46630
rect 59906 -46680 59916 -46490
rect 60006 -46680 60016 -46490
rect 59906 -46690 60016 -46680
rect 60286 -46510 60376 -46100
rect 60556 -46500 60626 -45710
rect 61026 -46020 61136 -45050
rect 79400 -45120 79690 -45110
rect 79400 -45360 79410 -45120
rect 79680 -45360 79690 -45120
rect 79400 -45370 79690 -45360
rect 79980 -45430 81960 -45400
rect 74460 -45480 77280 -45470
rect 74460 -45560 74470 -45480
rect 74590 -45560 77280 -45480
rect 79980 -45540 80010 -45430
rect 74460 -45570 77280 -45560
rect 77150 -45600 77280 -45570
rect 79060 -45560 80010 -45540
rect 77150 -45610 77720 -45600
rect 76910 -45640 77070 -45630
rect 61196 -45720 61356 -45710
rect 61196 -45900 61206 -45720
rect 61346 -45900 61356 -45720
rect 76910 -45740 76920 -45640
rect 77060 -45740 77070 -45640
rect 77150 -45680 77600 -45610
rect 77710 -45680 77720 -45610
rect 77150 -45690 77720 -45680
rect 79060 -45680 79080 -45560
rect 79190 -45680 80010 -45560
rect 79060 -45700 80010 -45680
rect 76910 -45750 77070 -45740
rect 79980 -45810 80010 -45700
rect 80360 -45810 81510 -45430
rect 81930 -45810 81960 -45430
rect 79980 -45840 81960 -45810
rect 61196 -45910 61356 -45900
rect 75210 -45890 78150 -45880
rect 75210 -45950 75220 -45890
rect 75340 -45950 78070 -45890
rect 78140 -45950 78150 -45890
rect 75210 -45960 78150 -45950
rect 61026 -46130 61036 -46020
rect 61126 -46130 61136 -46020
rect 61026 -46140 61136 -46130
rect 75380 -46190 79920 -46180
rect 61246 -46250 61366 -46240
rect 61246 -46260 61276 -46250
rect 61246 -46460 61256 -46260
rect 61356 -46460 61366 -46250
rect 75380 -46310 75390 -46190
rect 75550 -46310 78770 -46190
rect 78890 -46310 79740 -46190
rect 79910 -46310 79920 -46190
rect 75380 -46320 79920 -46310
rect 76900 -46440 77080 -46430
rect 61246 -46470 61366 -46460
rect 75200 -46467 75380 -46450
rect 60466 -46510 60626 -46500
rect 60286 -46570 60406 -46510
rect 60466 -46570 60476 -46510
rect 60536 -46570 60626 -46510
rect 75200 -46532 75231 -46467
rect 75322 -46480 75380 -46467
rect 76635 -46480 76739 -46467
rect 75322 -46532 76648 -46480
rect 59236 -46850 59266 -46760
rect 59366 -46850 59376 -46760
rect 59236 -46900 59376 -46850
rect 59506 -46710 59606 -46700
rect 59506 -46780 59516 -46710
rect 59596 -46780 59606 -46710
rect 59506 -46790 59606 -46780
rect 59236 -46920 59386 -46900
rect 59236 -46980 59316 -46920
rect 59376 -46980 59386 -46920
rect 58396 -47550 58896 -47050
rect 59236 -47230 59386 -46980
rect 59006 -47300 59086 -47280
rect 59236 -47290 59256 -47230
rect 59366 -47290 59386 -47230
rect 59236 -47300 59386 -47290
rect 59506 -47180 59596 -46790
rect 59986 -46920 60116 -46910
rect 59986 -46980 59996 -46920
rect 60106 -46980 60116 -46920
rect 59506 -47190 59616 -47180
rect 59506 -47260 59546 -47190
rect 59606 -47260 59616 -47190
rect 59006 -47360 59016 -47300
rect 59076 -47360 59086 -47300
rect 59006 -47550 59086 -47360
rect 59506 -47310 59616 -47260
rect 59506 -47370 59546 -47310
rect 59606 -47370 59616 -47310
rect 59796 -47210 59926 -47200
rect 59796 -47320 59806 -47210
rect 59916 -47320 59926 -47210
rect 59796 -47330 59926 -47320
rect 59006 -47640 59126 -47550
rect 59006 -47710 59016 -47640
rect 59076 -47710 59126 -47640
rect 59006 -47790 59126 -47710
rect 59506 -47640 59616 -47370
rect 59506 -47710 59546 -47640
rect 59606 -47710 59616 -47640
rect 59506 -47720 59616 -47710
rect 59986 -47790 60116 -46980
rect 60286 -47470 60376 -46570
rect 60466 -46580 60626 -46570
rect 61486 -46570 61726 -46540
rect 75200 -46545 76648 -46532
rect 76726 -46545 76739 -46480
rect 75200 -46550 76739 -46545
rect 76635 -46558 76739 -46550
rect 61486 -46620 61496 -46570
rect 61326 -46630 61496 -46620
rect 61326 -46750 61336 -46630
rect 61196 -46760 61336 -46750
rect 61456 -46740 61496 -46630
rect 61696 -46740 61726 -46570
rect 76900 -46580 76910 -46440
rect 77070 -46580 77080 -46440
rect 76900 -46590 77080 -46580
rect 74451 -46610 74620 -46597
rect 74451 -46714 74477 -46610
rect 74594 -46623 76193 -46610
rect 74594 -46701 76102 -46623
rect 76180 -46701 76193 -46623
rect 74594 -46714 76193 -46701
rect 76770 -46670 78360 -46660
rect 74451 -46727 74620 -46714
rect 61456 -46760 61726 -46740
rect 76770 -46740 76780 -46670
rect 76860 -46740 78280 -46670
rect 78350 -46740 78360 -46670
rect 76770 -46750 78360 -46740
rect 61196 -46770 61726 -46760
rect 76362 -46766 76453 -46753
rect 61196 -46940 61426 -46770
rect 76362 -46779 76375 -46766
rect 74711 -46792 76375 -46779
rect 74711 -46870 74724 -46792
rect 74841 -46844 76375 -46792
rect 76440 -46844 76453 -46766
rect 74841 -46857 76453 -46844
rect 77160 -46830 77440 -46820
rect 74841 -46870 74854 -46857
rect 74711 -46883 74854 -46870
rect 72810 -46900 73050 -46890
rect 72810 -47080 72820 -46900
rect 73040 -46910 73050 -46900
rect 73040 -47070 73370 -46910
rect 73040 -47080 73050 -47070
rect 72810 -47090 73050 -47080
rect 73210 -47080 75350 -47070
rect 62400 -47200 63000 -47100
rect 73210 -47180 75220 -47080
rect 75340 -47180 75350 -47080
rect 77160 -47080 77170 -46830
rect 77430 -47080 77440 -46830
rect 77160 -47090 77440 -47080
rect 82794 -46878 91444 -46848
rect 73210 -47190 75350 -47180
rect 63203 -47200 73103 -47199
rect 60436 -47230 60536 -47210
rect 60436 -47350 60446 -47230
rect 60526 -47350 60536 -47230
rect 60436 -47360 60536 -47350
rect 60256 -47600 60416 -47470
rect 62400 -47500 62500 -47200
rect 62900 -47230 73103 -47200
rect 62900 -47410 72820 -47230
rect 73040 -47250 73103 -47230
rect 73040 -47260 75100 -47250
rect 73040 -47380 74970 -47260
rect 75090 -47380 75100 -47260
rect 80050 -47310 80460 -47280
rect 80050 -47370 80080 -47310
rect 73040 -47390 75100 -47380
rect 79060 -47390 80080 -47370
rect 73040 -47410 73103 -47390
rect 62900 -47499 73103 -47410
rect 73960 -47470 77330 -47460
rect 62900 -47500 63600 -47499
rect 62400 -47600 63000 -47500
rect 73960 -47530 73970 -47470
rect 74090 -47480 77330 -47470
rect 74090 -47530 77230 -47480
rect 73960 -47540 77230 -47530
rect 77310 -47540 77330 -47480
rect 77200 -47560 77330 -47540
rect 79060 -47550 79080 -47390
rect 79250 -47550 80080 -47390
rect 79060 -47560 80080 -47550
rect 60256 -47730 60266 -47600
rect 60406 -47730 60416 -47600
rect 60256 -47750 60416 -47730
rect 64100 -47700 73100 -47600
rect 58956 -47800 59156 -47790
rect 58956 -47980 58966 -47800
rect 59146 -47980 59156 -47800
rect 59986 -47900 59996 -47790
rect 60106 -47900 60116 -47790
rect 64100 -47900 64200 -47700
rect 64500 -47720 73100 -47700
rect 64500 -47900 72820 -47720
rect 73040 -47730 73100 -47720
rect 76910 -47610 77070 -47600
rect 73040 -47740 74850 -47730
rect 73040 -47880 74720 -47740
rect 74840 -47880 74850 -47740
rect 76910 -47760 76920 -47610
rect 77060 -47760 77070 -47610
rect 80050 -47620 80080 -47560
rect 80430 -47620 80460 -47310
rect 82794 -47448 82824 -46878
rect 91414 -47448 91444 -46878
rect 82794 -47478 91444 -47448
rect 80050 -47630 80460 -47620
rect 85314 -47588 90774 -47578
rect 85314 -47678 85324 -47588
rect 85394 -47678 85594 -47588
rect 86484 -47678 87044 -47588
rect 87924 -47678 88514 -47588
rect 89394 -47678 89984 -47588
rect 90764 -47678 90774 -47588
rect 85314 -47688 90774 -47678
rect 76910 -47770 77070 -47760
rect 80050 -47720 80460 -47690
rect 73040 -47890 74850 -47880
rect 74960 -47820 76620 -47810
rect 74960 -47890 74980 -47820
rect 75080 -47830 76620 -47820
rect 77130 -47820 77270 -47810
rect 77130 -47830 77170 -47820
rect 75080 -47890 77170 -47830
rect 77260 -47890 77270 -47820
rect 80050 -47860 80080 -47720
rect 73040 -47900 73100 -47890
rect 74960 -47900 77270 -47890
rect 78570 -47880 80080 -47860
rect 58956 -47990 59156 -47980
rect 59600 -48000 63000 -47900
rect 64100 -48000 64600 -47900
rect 72810 -47910 73050 -47900
rect 78570 -47940 78580 -47880
rect 78640 -47940 80080 -47880
rect 78570 -47960 80080 -47940
rect 72810 -48000 73050 -47990
rect 59600 -48400 59700 -48000
rect 60400 -48400 62500 -48000
rect 62900 -48400 63000 -48000
rect 65000 -48100 72820 -48000
rect 65000 -48300 65100 -48100
rect 65400 -48180 72820 -48100
rect 73040 -48010 73100 -48000
rect 73040 -48140 74600 -48010
rect 80050 -48100 80080 -47960
rect 80430 -48100 80460 -47720
rect 80050 -48130 80460 -48100
rect 82210 -48020 83110 -48010
rect 82210 -48140 82220 -48020
rect 82340 -48140 83040 -48020
rect 83100 -48140 83110 -48020
rect 73040 -48150 77490 -48140
rect 82210 -48150 83110 -48140
rect 73040 -48170 74470 -48150
rect 73040 -48180 73100 -48170
rect 65400 -48300 73100 -48180
rect 74380 -48220 74470 -48170
rect 74590 -48220 77410 -48150
rect 77480 -48220 77490 -48150
rect 74380 -48230 77490 -48220
rect 79400 -48190 79690 -48180
rect 65000 -48400 65500 -48300
rect 59600 -48500 63000 -48400
rect 66000 -48460 73100 -48400
rect 66000 -48500 72820 -48460
rect 66000 -48700 66100 -48500
rect 66400 -48640 72820 -48500
rect 73040 -48470 73100 -48460
rect 74210 -48430 77850 -48420
rect 74210 -48470 74220 -48430
rect 73040 -48490 74220 -48470
rect 74340 -48490 77780 -48430
rect 77840 -48490 77850 -48430
rect 79400 -48430 79410 -48190
rect 79680 -48430 79690 -48190
rect 91750 -48240 92160 -48210
rect 91750 -48358 91780 -48240
rect 79400 -48440 79690 -48430
rect 86794 -48368 91780 -48358
rect 86794 -48448 86804 -48368
rect 86874 -48448 88274 -48368
rect 88344 -48448 89754 -48368
rect 89814 -48448 91214 -48368
rect 91284 -48448 91780 -48368
rect 86794 -48458 91780 -48448
rect 73040 -48500 77850 -48490
rect 73040 -48630 74350 -48500
rect 75210 -48580 77530 -48570
rect 73040 -48640 73100 -48630
rect 66400 -48700 73100 -48640
rect 75210 -48650 75220 -48580
rect 75340 -48650 77450 -48580
rect 77520 -48650 77530 -48580
rect 75210 -48660 77530 -48650
rect 82794 -48578 91444 -48548
rect 66000 -48800 66500 -48700
rect 67000 -48820 73100 -48800
rect 67000 -48900 72820 -48820
rect 67000 -49100 67100 -48900
rect 67400 -49000 72820 -48900
rect 73040 -48830 73100 -48820
rect 73040 -48840 74100 -48830
rect 73040 -48980 73970 -48840
rect 74090 -48980 74100 -48840
rect 73040 -48990 74100 -48980
rect 76910 -48860 77070 -48850
rect 73040 -49000 73100 -48990
rect 67400 -49100 73100 -49000
rect 76910 -49000 76920 -48860
rect 77060 -49000 77070 -48860
rect 76910 -49010 77070 -49000
rect 80050 -48950 82640 -48920
rect 80050 -49060 80080 -48950
rect 78660 -49070 80080 -49060
rect 67000 -49200 67500 -49100
rect 75210 -49200 77540 -49190
rect 67900 -49220 73100 -49200
rect 67900 -49300 72820 -49220
rect 67900 -49500 68000 -49300
rect 68300 -49400 72820 -49300
rect 73040 -49230 73100 -49220
rect 73040 -49240 73850 -49230
rect 73040 -49380 73720 -49240
rect 73840 -49380 73850 -49240
rect 75210 -49280 75220 -49200
rect 75340 -49280 77450 -49200
rect 77530 -49280 77540 -49200
rect 78660 -49220 78670 -49070
rect 78780 -49220 80080 -49070
rect 78660 -49230 80080 -49220
rect 75210 -49290 77540 -49280
rect 80050 -49330 80080 -49230
rect 80430 -49330 82450 -48950
rect 82610 -49330 82640 -48950
rect 82794 -49148 82824 -48578
rect 91414 -49148 91444 -48578
rect 91750 -48620 91780 -48458
rect 92130 -48620 92160 -48240
rect 91750 -48650 92160 -48620
rect 82794 -49178 91444 -49148
rect 73040 -49390 73850 -49380
rect 74460 -49360 77850 -49350
rect 80050 -49360 82640 -49330
rect 73040 -49400 73100 -49390
rect 68300 -49500 73100 -49400
rect 74460 -49420 74470 -49360
rect 74590 -49420 77780 -49360
rect 77840 -49420 77850 -49360
rect 74460 -49430 77850 -49420
rect 79400 -49420 79690 -49410
rect 67900 -49600 68400 -49500
rect 68900 -49670 73100 -49600
rect 79400 -49660 79410 -49420
rect 79680 -49660 79690 -49420
rect 68900 -49700 72820 -49670
rect 68900 -49900 69000 -49700
rect 69300 -49850 72820 -49700
rect 73040 -49680 73100 -49670
rect 74710 -49670 77850 -49660
rect 79400 -49670 79690 -49660
rect 73040 -49690 73600 -49680
rect 73040 -49830 73470 -49690
rect 73590 -49830 73600 -49690
rect 74710 -49730 74720 -49670
rect 74840 -49730 77780 -49670
rect 77840 -49730 77850 -49670
rect 74710 -49740 77850 -49730
rect 73040 -49840 73600 -49830
rect 75210 -49810 77590 -49800
rect 73040 -49850 73100 -49840
rect 69300 -49900 73100 -49850
rect 75210 -49900 75220 -49810
rect 75340 -49900 77490 -49810
rect 77580 -49900 77590 -49810
rect 68900 -50000 69400 -49900
rect 75210 -49910 77590 -49900
rect 58946 -50070 59146 -50050
rect 58946 -50230 58966 -50070
rect 59126 -50230 59146 -50070
rect 58946 -50250 59146 -50230
rect 59316 -50110 59426 -50050
rect 59316 -50250 59336 -50110
rect 59416 -50250 59426 -50110
rect 58956 -50330 59136 -50250
rect 58956 -50440 58996 -50330
rect 59106 -50440 59136 -50330
rect 58396 -50530 58896 -50440
rect 58956 -50500 59136 -50440
rect 59316 -50480 59426 -50250
rect 59946 -50120 60386 -50000
rect 59946 -50240 60046 -50120
rect 60126 -50240 60386 -50120
rect 59946 -50290 60386 -50240
rect 69900 -50040 73100 -50000
rect 69900 -50100 72820 -50040
rect 58396 -50890 58486 -50530
rect 58816 -50890 58896 -50530
rect 58996 -50800 59086 -50500
rect 58996 -50860 59006 -50800
rect 59066 -50860 59086 -50800
rect 58996 -50870 59086 -50860
rect 59266 -50530 59426 -50480
rect 59506 -50340 59796 -50300
rect 59506 -50440 59516 -50340
rect 59616 -50440 59796 -50340
rect 59506 -50500 59796 -50440
rect 59266 -50730 59366 -50530
rect 59266 -50790 59286 -50730
rect 59346 -50790 59366 -50730
rect 58396 -51000 58896 -50890
rect 59066 -51040 59176 -51030
rect 59066 -51110 59076 -51040
rect 59166 -51110 59176 -51040
rect 56470 -51638 56555 -51628
rect 56470 -51728 56480 -51638
rect 56550 -51728 56555 -51638
rect 56470 -51738 56555 -51728
rect 56470 -52118 56550 -51738
rect 57760 -51740 57800 -51620
rect 58240 -51740 58280 -51620
rect 57093 -52074 57373 -52064
rect 56470 -52128 56555 -52118
rect 56470 -52178 56480 -52128
rect 56475 -52188 56480 -52178
rect 56550 -52188 56555 -52128
rect 56475 -52198 56555 -52188
rect 57093 -52214 57098 -52074
rect 57368 -52214 57373 -52074
rect 57093 -52224 57373 -52214
rect 55870 -52678 55980 -52238
rect 55870 -52718 55880 -52678
rect 55875 -52758 55880 -52718
rect 55970 -52718 55980 -52678
rect 56060 -52668 56220 -52658
rect 55970 -52758 55975 -52718
rect 55875 -52768 55975 -52758
rect 55590 -52878 55620 -52788
rect 55710 -52878 55720 -52788
rect 56060 -52838 56220 -52828
rect 56060 -52848 56200 -52838
rect 55590 -52888 55720 -52878
rect 56015 -52858 56200 -52848
rect 56015 -53008 56020 -52858
rect 56080 -53008 56200 -52858
rect 56644 -52868 57008 -52863
rect 55215 -53018 55325 -53008
rect 56015 -53018 56085 -53008
rect 55215 -53118 55220 -53018
rect 55320 -53118 55325 -53018
rect 56644 -53086 56654 -52868
rect 56998 -53086 57008 -52868
rect 56644 -53091 57008 -53086
rect 55215 -53128 55325 -53118
rect 55315 -53328 55475 -53318
rect 55315 -53468 55320 -53328
rect 55470 -53468 55475 -53328
rect 55315 -53478 55475 -53468
rect 42800 -53800 43500 -53700
rect 42800 -54400 42900 -53800
rect 43400 -53900 56200 -53800
rect 43400 -54300 55400 -53900
rect 56100 -54300 56200 -53900
rect 43400 -54400 56200 -54300
rect 42800 -54500 43500 -54400
rect 51400 -54880 55800 -54800
rect 51400 -54900 55460 -54880
rect 51400 -55100 51500 -54900
rect 52500 -55100 55460 -54900
rect 51400 -55160 55460 -55100
rect 55720 -55160 55800 -54880
rect 51400 -55200 55800 -55160
rect 55380 -55240 55800 -55200
rect 47800 -55460 48100 -55440
rect 47800 -55820 47820 -55460
rect 48080 -55520 48100 -55460
rect 48080 -55540 53800 -55520
rect 48080 -55740 53480 -55540
rect 53780 -55740 53800 -55540
rect 56496 -55580 57026 -55575
rect 48080 -55760 53800 -55740
rect 55955 -55738 56045 -55728
rect 48080 -55820 48100 -55760
rect 47800 -55840 48100 -55820
rect 53515 -55858 53645 -55848
rect 53510 -55968 53520 -55858
rect 53640 -55968 53645 -55858
rect 55955 -55888 55960 -55738
rect 56040 -55888 56200 -55738
rect 56496 -55830 56506 -55580
rect 57016 -55830 57026 -55580
rect 56496 -55835 57026 -55830
rect 55955 -55898 56200 -55888
rect 53510 -55978 53645 -55968
rect 55275 -55918 55490 -55908
rect 53045 -56158 53255 -56148
rect 53045 -57908 53050 -56158
rect 53250 -57908 53255 -56158
rect 53045 -57918 53255 -57908
rect 53510 -58118 53630 -55978
rect 55275 -56008 55280 -55918
rect 55400 -56008 55490 -55918
rect 56060 -55938 56200 -55898
rect 56060 -55948 56220 -55938
rect 55275 -56018 55490 -56008
rect 55220 -56258 55325 -56248
rect 55220 -56428 55230 -56258
rect 55320 -56428 55325 -56258
rect 55220 -56438 55325 -56428
rect 55015 -57048 55125 -57038
rect 55015 -57128 55020 -57048
rect 55120 -57128 55125 -57048
rect 55015 -57138 55125 -57128
rect 55220 -57738 55310 -56438
rect 55215 -57748 55315 -57738
rect 55215 -57918 55220 -57748
rect 55310 -57838 55315 -57748
rect 55400 -57748 55490 -56018
rect 55875 -56018 55990 -56008
rect 55875 -56058 55880 -56018
rect 55870 -56098 55880 -56058
rect 55970 -56098 55990 -56018
rect 55870 -56178 55990 -56098
rect 56060 -56118 56220 -56108
rect 55590 -56268 55720 -56258
rect 55590 -56398 55600 -56268
rect 55710 -56398 55720 -56268
rect 55400 -57758 55510 -57748
rect 55310 -57918 55320 -57838
rect 55400 -57918 55410 -57758
rect 55215 -57928 55320 -57918
rect 53505 -58128 53635 -58118
rect 24400 -58800 36000 -58200
rect 53505 -58248 53510 -58128
rect 53630 -58248 53635 -58128
rect 53505 -58258 53635 -58248
rect 55220 -58408 55320 -57928
rect 55405 -57928 55410 -57918
rect 55500 -57928 55510 -57758
rect 55405 -57938 55510 -57928
rect 55590 -58188 55720 -56398
rect 55870 -56558 55980 -56178
rect 57093 -56564 57373 -56554
rect 56475 -56588 56555 -56578
rect 56470 -56648 56480 -56588
rect 56550 -56648 56555 -56588
rect 56470 -56658 56555 -56648
rect 55870 -57038 55980 -56668
rect 55870 -57128 55880 -57038
rect 55970 -57128 55980 -57038
rect 55870 -57528 55980 -57128
rect 56470 -57028 56550 -56658
rect 57093 -56704 57098 -56564
rect 57368 -56704 57373 -56564
rect 57093 -56714 57373 -56704
rect 57760 -57020 58280 -51740
rect 58516 -51660 58796 -51590
rect 58516 -51860 58556 -51660
rect 58756 -51860 58796 -51660
rect 59066 -51610 59176 -51110
rect 59266 -51220 59366 -50790
rect 59536 -50690 59616 -50500
rect 59536 -50750 59546 -50690
rect 59606 -50750 59616 -50690
rect 59536 -50810 59616 -50750
rect 59536 -50870 59546 -50810
rect 59606 -50870 59616 -50810
rect 59536 -50880 59616 -50870
rect 59266 -51230 59376 -51220
rect 59266 -51320 59286 -51230
rect 59366 -51320 59376 -51230
rect 59736 -51250 59796 -50500
rect 59856 -50740 59976 -50730
rect 59856 -50830 59866 -50740
rect 59966 -50830 59976 -50740
rect 59856 -50840 59976 -50830
rect 60036 -50920 60136 -50290
rect 69900 -50300 70000 -50100
rect 70300 -50220 72820 -50100
rect 73040 -50050 73100 -50040
rect 73040 -50060 73350 -50050
rect 73040 -50200 73220 -50060
rect 73340 -50200 73350 -50060
rect 73040 -50210 73350 -50200
rect 76910 -50100 77070 -50090
rect 73040 -50220 73100 -50210
rect 70300 -50300 73100 -50220
rect 76910 -50260 76920 -50100
rect 77060 -50260 77070 -50100
rect 61026 -50320 61136 -50310
rect 61026 -50450 61056 -50320
rect 61126 -50450 61136 -50320
rect 69900 -50400 70400 -50300
rect 74960 -50310 76850 -50300
rect 74960 -50370 74970 -50310
rect 75090 -50320 76850 -50310
rect 77130 -50310 77850 -50300
rect 77130 -50320 77780 -50310
rect 75090 -50370 77780 -50320
rect 77840 -50370 77850 -50310
rect 74960 -50380 77850 -50370
rect 76850 -50390 77130 -50380
rect 78130 -50400 79170 -50380
rect 78130 -50410 79050 -50400
rect 60436 -50720 60536 -50710
rect 60436 -50820 60446 -50720
rect 60526 -50820 60536 -50720
rect 60436 -50830 60536 -50820
rect 60036 -51000 60046 -50920
rect 60126 -51000 60136 -50920
rect 60036 -51010 60136 -51000
rect 60546 -51010 60636 -51000
rect 60386 -51090 60556 -51010
rect 60626 -51090 60636 -51010
rect 59966 -51100 60326 -51090
rect 59966 -51170 59976 -51100
rect 60316 -51170 60326 -51100
rect 60546 -51110 60636 -51090
rect 59966 -51180 60326 -51170
rect 59566 -51270 59796 -51250
rect 59566 -51280 59576 -51270
rect 59266 -51330 59376 -51320
rect 59516 -51330 59576 -51280
rect 59636 -51330 59796 -51270
rect 59266 -51440 59366 -51330
rect 59266 -51530 59286 -51440
rect 59356 -51530 59366 -51440
rect 59266 -51560 59366 -51530
rect 59516 -51340 59796 -51330
rect 59066 -51680 59076 -51610
rect 59166 -51680 59176 -51610
rect 59066 -51690 59176 -51680
rect 59306 -51630 59386 -51620
rect 59306 -51690 59316 -51630
rect 59376 -51690 59386 -51630
rect 59516 -51670 59596 -51340
rect 60286 -51350 60476 -51340
rect 59906 -51380 60016 -51370
rect 59906 -51560 59916 -51380
rect 60006 -51560 60016 -51380
rect 59906 -51570 60016 -51560
rect 60286 -51490 60306 -51350
rect 60456 -51490 60476 -51350
rect 60286 -51500 60476 -51490
rect 58516 -51940 58796 -51860
rect 59066 -51770 59176 -51760
rect 59066 -51840 59076 -51770
rect 59166 -51840 59176 -51770
rect 59066 -52340 59176 -51840
rect 59306 -51890 59386 -51690
rect 60076 -51680 60196 -51640
rect 60076 -51840 60096 -51680
rect 60176 -51840 60196 -51680
rect 60076 -51880 60196 -51840
rect 59066 -52400 59076 -52340
rect 59166 -52400 59176 -52340
rect 59066 -52410 59176 -52400
rect 59236 -51920 59386 -51890
rect 59236 -52010 59266 -51920
rect 59366 -52010 59386 -51920
rect 59236 -52030 59386 -52010
rect 59906 -51890 60016 -51880
rect 59236 -52160 59376 -52030
rect 59906 -52080 59916 -51890
rect 60006 -52080 60016 -51890
rect 59906 -52090 60016 -52080
rect 60286 -51910 60376 -51500
rect 60556 -51900 60626 -51110
rect 61026 -51420 61136 -50450
rect 75210 -50450 76790 -50440
rect 77190 -50450 77570 -50440
rect 75210 -50540 75220 -50450
rect 75340 -50540 77470 -50450
rect 77560 -50540 77570 -50450
rect 78130 -50510 78160 -50410
rect 78260 -50510 79050 -50410
rect 79150 -50510 79170 -50400
rect 78130 -50530 79170 -50510
rect 82790 -50530 91440 -50500
rect 75210 -50550 77570 -50540
rect 79400 -50680 79690 -50670
rect 79400 -50920 79410 -50680
rect 79680 -50920 79690 -50680
rect 79400 -50930 79690 -50920
rect 78850 -50960 79000 -50940
rect 73710 -50970 77550 -50960
rect 73710 -51040 73720 -50970
rect 73840 -51030 77470 -50970
rect 77540 -51030 77550 -50970
rect 73840 -51040 77550 -51030
rect 73710 -51050 73850 -51040
rect 77740 -51090 77930 -51080
rect 77740 -51100 77860 -51090
rect 76200 -51110 77860 -51100
rect 61196 -51120 61356 -51110
rect 61196 -51300 61206 -51120
rect 61346 -51300 61356 -51120
rect 76200 -51170 76210 -51110
rect 76340 -51150 77860 -51110
rect 77920 -51150 77930 -51090
rect 76340 -51160 77930 -51150
rect 76340 -51170 76350 -51160
rect 76200 -51180 76350 -51170
rect 75210 -51230 76140 -51220
rect 75210 -51290 75220 -51230
rect 75340 -51240 76140 -51230
rect 76410 -51230 78030 -51220
rect 76410 -51240 77960 -51230
rect 75340 -51280 77960 -51240
rect 75340 -51290 76840 -51280
rect 75210 -51300 76840 -51290
rect 77120 -51290 77960 -51280
rect 78020 -51290 78030 -51230
rect 78850 -51250 78860 -50960
rect 78980 -51040 79000 -50960
rect 79980 -50950 82080 -50920
rect 79980 -51040 80010 -50950
rect 78980 -51250 80010 -51040
rect 78850 -51260 80010 -51250
rect 77120 -51300 78030 -51290
rect 61196 -51310 61356 -51300
rect 79980 -51330 80010 -51260
rect 80360 -51140 82080 -50950
rect 82790 -51100 82820 -50530
rect 91410 -51100 91440 -50530
rect 82790 -51130 91440 -51100
rect 80360 -51330 81950 -51140
rect 61026 -51530 61036 -51420
rect 61126 -51530 61136 -51420
rect 76910 -51350 77070 -51340
rect 76910 -51490 76920 -51350
rect 77060 -51490 77070 -51350
rect 79980 -51350 81950 -51330
rect 82070 -51350 82080 -51140
rect 85310 -51240 90770 -51230
rect 85310 -51330 85320 -51240
rect 85390 -51330 85590 -51240
rect 86480 -51330 87040 -51240
rect 87920 -51330 88510 -51240
rect 89390 -51330 89980 -51240
rect 90760 -51330 90770 -51240
rect 85310 -51340 90770 -51330
rect 79980 -51360 82080 -51350
rect 76910 -51500 77070 -51490
rect 61026 -51540 61136 -51530
rect 61246 -51650 61366 -51640
rect 61246 -51660 61276 -51650
rect 61246 -51860 61256 -51660
rect 61356 -51860 61366 -51650
rect 75210 -51660 78040 -51650
rect 75210 -51720 75220 -51660
rect 75340 -51720 77970 -51660
rect 78030 -51720 78040 -51660
rect 75210 -51730 78040 -51720
rect 81630 -51680 83110 -51670
rect 81630 -51790 81640 -51680
rect 81760 -51790 83030 -51680
rect 83100 -51790 83110 -51680
rect 61246 -51870 61366 -51860
rect 73960 -51800 77510 -51790
rect 81630 -51800 83110 -51790
rect 73960 -51870 73970 -51800
rect 74090 -51870 77430 -51800
rect 77500 -51870 77510 -51800
rect 73960 -51880 77510 -51870
rect 91750 -51870 92160 -51840
rect 60466 -51910 60626 -51900
rect 60286 -51970 60406 -51910
rect 60466 -51970 60476 -51910
rect 60536 -51970 60626 -51910
rect 79400 -51900 79690 -51890
rect 59236 -52250 59266 -52160
rect 59366 -52250 59376 -52160
rect 59236 -52300 59376 -52250
rect 59506 -52110 59606 -52100
rect 59506 -52180 59516 -52110
rect 59596 -52180 59606 -52110
rect 59506 -52190 59606 -52180
rect 59236 -52320 59386 -52300
rect 59236 -52380 59316 -52320
rect 59376 -52380 59386 -52320
rect 58396 -52950 58896 -52450
rect 59236 -52630 59386 -52380
rect 59006 -52700 59086 -52680
rect 59236 -52690 59256 -52630
rect 59366 -52690 59386 -52630
rect 59236 -52700 59386 -52690
rect 59506 -52580 59596 -52190
rect 59986 -52320 60116 -52310
rect 59986 -52380 59996 -52320
rect 60106 -52380 60116 -52320
rect 59506 -52590 59616 -52580
rect 59506 -52660 59546 -52590
rect 59606 -52660 59616 -52590
rect 59006 -52760 59016 -52700
rect 59076 -52760 59086 -52700
rect 59006 -52950 59086 -52760
rect 59506 -52710 59616 -52660
rect 59506 -52770 59546 -52710
rect 59606 -52770 59616 -52710
rect 59796 -52610 59926 -52600
rect 59796 -52720 59806 -52610
rect 59916 -52720 59926 -52610
rect 59796 -52730 59926 -52720
rect 59006 -53040 59126 -52950
rect 59006 -53110 59016 -53040
rect 59076 -53110 59126 -53040
rect 59006 -53190 59126 -53110
rect 59506 -53040 59616 -52770
rect 59506 -53110 59546 -53040
rect 59606 -53110 59616 -53040
rect 59506 -53120 59616 -53110
rect 59986 -53190 60116 -52380
rect 60286 -52870 60376 -51970
rect 60466 -51980 60626 -51970
rect 61486 -51970 61726 -51940
rect 61486 -52020 61496 -51970
rect 61326 -52030 61496 -52020
rect 61326 -52150 61336 -52030
rect 61196 -52160 61336 -52150
rect 61456 -52140 61496 -52030
rect 61696 -52140 61726 -51970
rect 61456 -52160 61726 -52140
rect 79400 -52140 79410 -51900
rect 79680 -52140 79690 -51900
rect 91750 -52010 91780 -51870
rect 86790 -52020 91780 -52010
rect 86790 -52100 86800 -52020
rect 86870 -52100 88270 -52020
rect 88340 -52100 89750 -52020
rect 89810 -52100 91210 -52020
rect 91280 -52100 91780 -52020
rect 86790 -52110 91780 -52100
rect 79400 -52150 79690 -52140
rect 61196 -52170 61726 -52160
rect 61196 -52340 61426 -52170
rect 82790 -52230 91440 -52200
rect 76480 -52290 77490 -52280
rect 76480 -52350 76490 -52290
rect 76610 -52330 77490 -52290
rect 76610 -52350 78040 -52330
rect 76480 -52360 76620 -52350
rect 77410 -52390 78040 -52350
rect 73460 -52420 73610 -52410
rect 73460 -52480 73470 -52420
rect 73590 -52450 77340 -52420
rect 73590 -52460 77830 -52450
rect 73590 -52480 77760 -52460
rect 73460 -52490 77760 -52480
rect 73460 -52500 73610 -52490
rect 77150 -52520 77760 -52490
rect 77820 -52520 77830 -52460
rect 77960 -52510 77970 -52390
rect 78030 -52510 78040 -52390
rect 77960 -52520 78040 -52510
rect 77150 -52530 77830 -52520
rect 76910 -52560 77070 -52550
rect 60436 -52630 60536 -52610
rect 60436 -52750 60446 -52630
rect 60526 -52750 60536 -52630
rect 76910 -52650 76920 -52560
rect 77060 -52650 77070 -52560
rect 76910 -52660 77070 -52650
rect 60436 -52760 60536 -52750
rect 73960 -52780 77830 -52770
rect 73960 -52840 73970 -52780
rect 74090 -52840 77760 -52780
rect 77820 -52840 77830 -52780
rect 82790 -52800 82820 -52230
rect 91410 -52800 91440 -52230
rect 91750 -52250 91780 -52110
rect 92130 -52250 92160 -51870
rect 91750 -52280 92160 -52250
rect 73960 -52850 77830 -52840
rect 78770 -52810 78930 -52800
rect 60256 -53000 60416 -52870
rect 77950 -52890 78030 -52880
rect 77950 -52910 77960 -52890
rect 76480 -52920 77960 -52910
rect 76480 -52990 76490 -52920
rect 76610 -52960 77960 -52920
rect 78020 -52960 78030 -52890
rect 78770 -52930 78780 -52810
rect 78920 -52840 79170 -52810
rect 82790 -52830 91440 -52800
rect 78920 -52910 79070 -52840
rect 79140 -52910 79170 -52840
rect 78920 -52930 79170 -52910
rect 78770 -52940 78930 -52930
rect 76610 -52970 78030 -52960
rect 76610 -52990 77530 -52970
rect 76480 -53000 77530 -52990
rect 60256 -53130 60266 -53000
rect 60406 -53130 60416 -53000
rect 60256 -53150 60416 -53130
rect 58956 -53200 59156 -53190
rect 58956 -53380 58966 -53200
rect 59146 -53380 59156 -53200
rect 59986 -53300 59996 -53190
rect 60106 -53300 60116 -53190
rect 79400 -53160 79690 -53150
rect 58956 -53390 59156 -53380
rect 59600 -53400 64600 -53300
rect 59600 -53800 59700 -53400
rect 60400 -53800 64200 -53400
rect 64500 -53800 64600 -53400
rect 79400 -53400 79410 -53160
rect 79680 -53400 79690 -53160
rect 79400 -53410 79690 -53400
rect 79980 -53470 82780 -53440
rect 74460 -53520 77280 -53510
rect 74460 -53600 74470 -53520
rect 74590 -53600 77280 -53520
rect 79980 -53580 80010 -53470
rect 74460 -53610 77280 -53600
rect 77150 -53640 77280 -53610
rect 79060 -53600 80010 -53580
rect 77150 -53650 77720 -53640
rect 76910 -53680 77070 -53670
rect 76910 -53780 76920 -53680
rect 77060 -53780 77070 -53680
rect 77150 -53720 77600 -53650
rect 77710 -53720 77720 -53650
rect 77150 -53730 77720 -53720
rect 79060 -53720 79080 -53600
rect 79190 -53720 80010 -53600
rect 79060 -53740 80010 -53720
rect 76910 -53790 77070 -53780
rect 59600 -53900 64600 -53800
rect 79980 -53850 80010 -53740
rect 80360 -53850 82140 -53470
rect 82750 -53850 82780 -53470
rect 79980 -53880 82780 -53850
rect 75210 -53930 78150 -53920
rect 75210 -53990 75220 -53930
rect 75340 -53990 78070 -53930
rect 78140 -53990 78150 -53930
rect 75210 -54000 78150 -53990
rect 58946 -55470 59146 -55450
rect 58946 -55630 58966 -55470
rect 59126 -55630 59146 -55470
rect 58946 -55650 59146 -55630
rect 59316 -55510 59426 -55450
rect 59316 -55650 59336 -55510
rect 59416 -55650 59426 -55510
rect 58956 -55730 59136 -55650
rect 58956 -55840 58996 -55730
rect 59106 -55840 59136 -55730
rect 58396 -55930 58896 -55840
rect 58956 -55900 59136 -55840
rect 59316 -55880 59426 -55650
rect 59946 -55520 60386 -55400
rect 59946 -55640 60046 -55520
rect 60126 -55640 60386 -55520
rect 59946 -55690 60386 -55640
rect 58396 -56290 58486 -55930
rect 58816 -56290 58896 -55930
rect 58996 -56200 59086 -55900
rect 58996 -56260 59006 -56200
rect 59066 -56260 59086 -56200
rect 58996 -56270 59086 -56260
rect 59266 -55930 59426 -55880
rect 59506 -55740 59796 -55700
rect 59506 -55840 59516 -55740
rect 59616 -55840 59796 -55740
rect 59506 -55900 59796 -55840
rect 59266 -56130 59366 -55930
rect 59266 -56190 59286 -56130
rect 59346 -56190 59366 -56130
rect 58396 -56400 58896 -56290
rect 59066 -56440 59176 -56430
rect 59066 -56510 59076 -56440
rect 59166 -56510 59176 -56440
rect 56470 -57038 56555 -57028
rect 56470 -57128 56480 -57038
rect 56550 -57128 56555 -57038
rect 56470 -57138 56555 -57128
rect 56470 -57518 56550 -57138
rect 57760 -57140 57800 -57020
rect 58240 -57140 58280 -57020
rect 57093 -57474 57373 -57464
rect 56470 -57528 56555 -57518
rect 56470 -57578 56480 -57528
rect 56475 -57588 56480 -57578
rect 56550 -57588 56555 -57528
rect 56475 -57598 56555 -57588
rect 57093 -57614 57098 -57474
rect 57368 -57614 57373 -57474
rect 57093 -57624 57373 -57614
rect 55870 -58078 55980 -57638
rect 55870 -58118 55880 -58078
rect 55875 -58158 55880 -58118
rect 55970 -58118 55980 -58078
rect 56060 -58068 56220 -58058
rect 55970 -58158 55975 -58118
rect 55875 -58168 55975 -58158
rect 55590 -58278 55620 -58188
rect 55710 -58278 55720 -58188
rect 56060 -58238 56220 -58228
rect 56060 -58248 56200 -58238
rect 55590 -58288 55720 -58278
rect 56015 -58258 56200 -58248
rect 56015 -58408 56020 -58258
rect 56080 -58408 56200 -58258
rect 56644 -58268 57008 -58263
rect 55215 -58418 55325 -58408
rect 56015 -58418 56085 -58408
rect 55215 -58518 55220 -58418
rect 55320 -58518 55325 -58418
rect 56644 -58486 56654 -58268
rect 56998 -58486 57008 -58268
rect 56644 -58491 57008 -58486
rect 55215 -58528 55325 -58518
rect 24400 -59400 25000 -58800
rect 14600 -60000 25000 -59400
rect 14600 -64800 15200 -60000
rect 19600 -64800 25000 -60000
rect 35400 -64800 36000 -58800
rect 55315 -58728 55475 -58718
rect 55315 -58868 55320 -58728
rect 55470 -58868 55475 -58728
rect 55315 -58878 55475 -58868
rect 41900 -59200 42600 -59100
rect 41900 -59800 42000 -59200
rect 42500 -59300 56200 -59200
rect 42500 -59700 55500 -59300
rect 56100 -59700 56200 -59300
rect 42500 -59800 56200 -59700
rect 41900 -59900 42600 -59800
rect 51400 -60280 55800 -60200
rect 51400 -60300 55460 -60280
rect 51400 -60500 51500 -60300
rect 52500 -60500 55460 -60300
rect 51400 -60560 55460 -60500
rect 55720 -60560 55800 -60280
rect 51400 -60600 55800 -60560
rect 55380 -60640 55800 -60600
rect 47660 -60760 48100 -60740
rect 47660 -61300 47680 -60760
rect 48080 -60920 48100 -60760
rect 48080 -60940 53800 -60920
rect 48080 -61140 53480 -60940
rect 53780 -61140 53800 -60940
rect 56496 -60980 57026 -60975
rect 48080 -61160 53800 -61140
rect 55955 -61138 56045 -61128
rect 48080 -61300 48100 -61160
rect 53515 -61258 53645 -61248
rect 47660 -61320 48100 -61300
rect 53510 -61368 53520 -61258
rect 53640 -61368 53645 -61258
rect 55955 -61288 55960 -61138
rect 56040 -61288 56200 -61138
rect 56496 -61230 56506 -60980
rect 57016 -61230 57026 -60980
rect 56496 -61235 57026 -61230
rect 55955 -61298 56200 -61288
rect 53510 -61378 53645 -61368
rect 55275 -61318 55490 -61308
rect 53045 -61558 53255 -61548
rect 53045 -63308 53050 -61558
rect 53250 -63308 53255 -61558
rect 53045 -63318 53255 -63308
rect 53510 -63518 53630 -61378
rect 55275 -61408 55280 -61318
rect 55400 -61408 55490 -61318
rect 56060 -61338 56200 -61298
rect 56060 -61348 56220 -61338
rect 55275 -61418 55490 -61408
rect 55220 -61658 55325 -61648
rect 55220 -61828 55230 -61658
rect 55320 -61828 55325 -61658
rect 55220 -61838 55325 -61828
rect 55015 -62448 55125 -62438
rect 55015 -62528 55020 -62448
rect 55120 -62528 55125 -62448
rect 55015 -62538 55125 -62528
rect 55220 -63138 55310 -61838
rect 55215 -63148 55315 -63138
rect 55215 -63318 55220 -63148
rect 55310 -63238 55315 -63148
rect 55400 -63148 55490 -61418
rect 55875 -61418 55990 -61408
rect 55875 -61458 55880 -61418
rect 55870 -61498 55880 -61458
rect 55970 -61498 55990 -61418
rect 55870 -61578 55990 -61498
rect 56060 -61518 56220 -61508
rect 55590 -61668 55720 -61658
rect 55590 -61798 55600 -61668
rect 55710 -61798 55720 -61668
rect 55400 -63158 55510 -63148
rect 55310 -63318 55320 -63238
rect 55400 -63318 55410 -63158
rect 55215 -63328 55320 -63318
rect 53505 -63528 53635 -63518
rect 53505 -63648 53510 -63528
rect 53630 -63648 53635 -63528
rect 53505 -63658 53635 -63648
rect 55220 -63808 55320 -63328
rect 55405 -63328 55410 -63318
rect 55500 -63328 55510 -63158
rect 55405 -63338 55510 -63328
rect 55590 -63588 55720 -61798
rect 55870 -61958 55980 -61578
rect 57093 -61964 57373 -61954
rect 56475 -61988 56555 -61978
rect 56470 -62048 56480 -61988
rect 56550 -62048 56555 -61988
rect 56470 -62058 56555 -62048
rect 55870 -62438 55980 -62068
rect 55870 -62528 55880 -62438
rect 55970 -62528 55980 -62438
rect 55870 -62928 55980 -62528
rect 56470 -62428 56550 -62058
rect 57093 -62104 57098 -61964
rect 57368 -62104 57373 -61964
rect 57093 -62114 57373 -62104
rect 57760 -62420 58280 -57140
rect 58516 -57060 58796 -56990
rect 58516 -57260 58556 -57060
rect 58756 -57260 58796 -57060
rect 59066 -57010 59176 -56510
rect 59266 -56620 59366 -56190
rect 59536 -56090 59616 -55900
rect 59536 -56150 59546 -56090
rect 59606 -56150 59616 -56090
rect 59536 -56210 59616 -56150
rect 59536 -56270 59546 -56210
rect 59606 -56270 59616 -56210
rect 59536 -56280 59616 -56270
rect 59266 -56630 59376 -56620
rect 59266 -56720 59286 -56630
rect 59366 -56720 59376 -56630
rect 59736 -56650 59796 -55900
rect 59856 -56140 59976 -56130
rect 59856 -56230 59866 -56140
rect 59966 -56230 59976 -56140
rect 59856 -56240 59976 -56230
rect 60036 -56320 60136 -55690
rect 61026 -55720 61136 -55710
rect 61026 -55850 61056 -55720
rect 61126 -55850 61136 -55720
rect 60436 -56120 60536 -56110
rect 60436 -56220 60446 -56120
rect 60526 -56220 60536 -56120
rect 60436 -56230 60536 -56220
rect 60036 -56400 60046 -56320
rect 60126 -56400 60136 -56320
rect 60036 -56410 60136 -56400
rect 60546 -56410 60636 -56400
rect 60386 -56490 60556 -56410
rect 60626 -56490 60636 -56410
rect 59966 -56500 60326 -56490
rect 59966 -56570 59976 -56500
rect 60316 -56570 60326 -56500
rect 60546 -56510 60636 -56490
rect 59966 -56580 60326 -56570
rect 59566 -56670 59796 -56650
rect 59566 -56680 59576 -56670
rect 59266 -56730 59376 -56720
rect 59516 -56730 59576 -56680
rect 59636 -56730 59796 -56670
rect 59266 -56840 59366 -56730
rect 59266 -56930 59286 -56840
rect 59356 -56930 59366 -56840
rect 59266 -56960 59366 -56930
rect 59516 -56740 59796 -56730
rect 59066 -57080 59076 -57010
rect 59166 -57080 59176 -57010
rect 59066 -57090 59176 -57080
rect 59306 -57030 59386 -57020
rect 59306 -57090 59316 -57030
rect 59376 -57090 59386 -57030
rect 59516 -57070 59596 -56740
rect 60286 -56750 60476 -56740
rect 59906 -56780 60016 -56770
rect 59906 -56960 59916 -56780
rect 60006 -56960 60016 -56780
rect 59906 -56970 60016 -56960
rect 60286 -56890 60306 -56750
rect 60456 -56890 60476 -56750
rect 60286 -56900 60476 -56890
rect 58516 -57340 58796 -57260
rect 59066 -57170 59176 -57160
rect 59066 -57240 59076 -57170
rect 59166 -57240 59176 -57170
rect 59066 -57740 59176 -57240
rect 59306 -57290 59386 -57090
rect 60076 -57080 60196 -57040
rect 60076 -57240 60096 -57080
rect 60176 -57240 60196 -57080
rect 60076 -57280 60196 -57240
rect 59066 -57800 59076 -57740
rect 59166 -57800 59176 -57740
rect 59066 -57810 59176 -57800
rect 59236 -57320 59386 -57290
rect 59236 -57410 59266 -57320
rect 59366 -57410 59386 -57320
rect 59236 -57430 59386 -57410
rect 59906 -57290 60016 -57280
rect 59236 -57560 59376 -57430
rect 59906 -57480 59916 -57290
rect 60006 -57480 60016 -57290
rect 59906 -57490 60016 -57480
rect 60286 -57310 60376 -56900
rect 60556 -57300 60626 -56510
rect 61026 -56820 61136 -55850
rect 61196 -56520 61356 -56510
rect 61196 -56700 61206 -56520
rect 61346 -56700 61356 -56520
rect 61196 -56710 61356 -56700
rect 61026 -56930 61036 -56820
rect 61126 -56930 61136 -56820
rect 61026 -56940 61136 -56930
rect 61246 -57050 61366 -57040
rect 61246 -57060 61276 -57050
rect 61246 -57260 61256 -57060
rect 61356 -57260 61366 -57050
rect 61246 -57270 61366 -57260
rect 60466 -57310 60626 -57300
rect 60286 -57370 60406 -57310
rect 60466 -57370 60476 -57310
rect 60536 -57370 60626 -57310
rect 59236 -57650 59266 -57560
rect 59366 -57650 59376 -57560
rect 59236 -57700 59376 -57650
rect 59506 -57510 59606 -57500
rect 59506 -57580 59516 -57510
rect 59596 -57580 59606 -57510
rect 59506 -57590 59606 -57580
rect 59236 -57720 59386 -57700
rect 59236 -57780 59316 -57720
rect 59376 -57780 59386 -57720
rect 58396 -58350 58896 -57850
rect 59236 -58030 59386 -57780
rect 59006 -58100 59086 -58080
rect 59236 -58090 59256 -58030
rect 59366 -58090 59386 -58030
rect 59236 -58100 59386 -58090
rect 59506 -57980 59596 -57590
rect 59986 -57720 60116 -57710
rect 59986 -57780 59996 -57720
rect 60106 -57780 60116 -57720
rect 59506 -57990 59616 -57980
rect 59506 -58060 59546 -57990
rect 59606 -58060 59616 -57990
rect 59006 -58160 59016 -58100
rect 59076 -58160 59086 -58100
rect 59006 -58350 59086 -58160
rect 59506 -58110 59616 -58060
rect 59506 -58170 59546 -58110
rect 59606 -58170 59616 -58110
rect 59796 -58010 59926 -58000
rect 59796 -58120 59806 -58010
rect 59916 -58120 59926 -58010
rect 59796 -58130 59926 -58120
rect 59006 -58440 59126 -58350
rect 59006 -58510 59016 -58440
rect 59076 -58510 59126 -58440
rect 59006 -58590 59126 -58510
rect 59506 -58440 59616 -58170
rect 59506 -58510 59546 -58440
rect 59606 -58510 59616 -58440
rect 59506 -58520 59616 -58510
rect 59986 -58590 60116 -57780
rect 60286 -58270 60376 -57370
rect 60466 -57380 60626 -57370
rect 61486 -57370 61726 -57340
rect 61486 -57420 61496 -57370
rect 61326 -57430 61496 -57420
rect 61326 -57550 61336 -57430
rect 61196 -57560 61336 -57550
rect 61456 -57540 61496 -57430
rect 61696 -57540 61726 -57370
rect 61456 -57560 61726 -57540
rect 61196 -57570 61726 -57560
rect 61196 -57740 61426 -57570
rect 60436 -58030 60536 -58010
rect 60436 -58150 60446 -58030
rect 60526 -58150 60536 -58030
rect 60436 -58160 60536 -58150
rect 60256 -58400 60416 -58270
rect 60256 -58530 60266 -58400
rect 60406 -58530 60416 -58400
rect 60256 -58550 60416 -58530
rect 58956 -58600 59156 -58590
rect 58956 -58780 58966 -58600
rect 59146 -58780 59156 -58600
rect 59986 -58700 59996 -58590
rect 60106 -58700 60116 -58590
rect 58956 -58790 59156 -58780
rect 59600 -58800 65500 -58700
rect 59600 -59200 59700 -58800
rect 60400 -59200 65100 -58800
rect 65400 -59200 65500 -58800
rect 59600 -59300 65500 -59200
rect 58946 -60870 59146 -60850
rect 58946 -61030 58966 -60870
rect 59126 -61030 59146 -60870
rect 58946 -61050 59146 -61030
rect 59316 -60910 59426 -60850
rect 59316 -61050 59336 -60910
rect 59416 -61050 59426 -60910
rect 58956 -61130 59136 -61050
rect 58956 -61240 58996 -61130
rect 59106 -61240 59136 -61130
rect 58396 -61330 58896 -61240
rect 58956 -61300 59136 -61240
rect 59316 -61280 59426 -61050
rect 59946 -60920 60386 -60800
rect 59946 -61040 60046 -60920
rect 60126 -61040 60386 -60920
rect 59946 -61090 60386 -61040
rect 58396 -61690 58486 -61330
rect 58816 -61690 58896 -61330
rect 58996 -61600 59086 -61300
rect 58996 -61660 59006 -61600
rect 59066 -61660 59086 -61600
rect 58996 -61670 59086 -61660
rect 59266 -61330 59426 -61280
rect 59506 -61140 59796 -61100
rect 59506 -61240 59516 -61140
rect 59616 -61240 59796 -61140
rect 59506 -61300 59796 -61240
rect 59266 -61530 59366 -61330
rect 59266 -61590 59286 -61530
rect 59346 -61590 59366 -61530
rect 58396 -61800 58896 -61690
rect 59066 -61840 59176 -61830
rect 59066 -61910 59076 -61840
rect 59166 -61910 59176 -61840
rect 56470 -62438 56555 -62428
rect 56470 -62528 56480 -62438
rect 56550 -62528 56555 -62438
rect 56470 -62538 56555 -62528
rect 56470 -62918 56550 -62538
rect 57760 -62540 57800 -62420
rect 58240 -62540 58280 -62420
rect 57093 -62874 57373 -62864
rect 56470 -62928 56555 -62918
rect 56470 -62978 56480 -62928
rect 56475 -62988 56480 -62978
rect 56550 -62988 56555 -62928
rect 56475 -62998 56555 -62988
rect 57093 -63014 57098 -62874
rect 57368 -63014 57373 -62874
rect 57093 -63024 57373 -63014
rect 55870 -63478 55980 -63038
rect 55870 -63518 55880 -63478
rect 55875 -63558 55880 -63518
rect 55970 -63518 55980 -63478
rect 56060 -63468 56220 -63458
rect 55970 -63558 55975 -63518
rect 55875 -63568 55975 -63558
rect 55590 -63678 55620 -63588
rect 55710 -63678 55720 -63588
rect 56060 -63638 56220 -63628
rect 56060 -63648 56200 -63638
rect 55590 -63688 55720 -63678
rect 56015 -63658 56200 -63648
rect 56015 -63808 56020 -63658
rect 56080 -63808 56200 -63658
rect 56644 -63668 57008 -63663
rect 55215 -63818 55325 -63808
rect 56015 -63818 56085 -63808
rect 55215 -63918 55220 -63818
rect 55320 -63918 55325 -63818
rect 56644 -63886 56654 -63668
rect 56998 -63886 57008 -63668
rect 56644 -63891 57008 -63886
rect 55215 -63928 55325 -63918
rect 55315 -64128 55475 -64118
rect 55315 -64268 55320 -64128
rect 55470 -64268 55475 -64128
rect 55315 -64278 55475 -64268
rect 14600 -65400 36000 -64800
rect 41000 -64600 41700 -64500
rect 41000 -65200 41100 -64600
rect 41600 -64700 56200 -64600
rect 41600 -65100 55500 -64700
rect 56100 -65100 56200 -64700
rect 41600 -65200 56200 -65100
rect 41000 -65300 41700 -65200
rect 51400 -65680 55800 -65600
rect 51400 -65700 55440 -65680
rect 51400 -65900 51500 -65700
rect 52500 -65900 55440 -65700
rect 51400 -65960 55440 -65900
rect 55720 -65960 55800 -65680
rect 51400 -66000 55800 -65960
rect 55360 -66040 55800 -66000
rect 47840 -66220 48100 -66200
rect 47840 -66660 47860 -66220
rect 48080 -66320 48100 -66220
rect 48080 -66340 53800 -66320
rect 48080 -66540 53480 -66340
rect 53780 -66540 53800 -66340
rect 56496 -66380 57026 -66375
rect 48080 -66560 53800 -66540
rect 55955 -66538 56045 -66528
rect 48080 -66660 48100 -66560
rect 53515 -66658 53645 -66648
rect 47840 -66680 48100 -66660
rect 53510 -66768 53520 -66658
rect 53640 -66768 53645 -66658
rect 55955 -66688 55960 -66538
rect 56040 -66688 56200 -66538
rect 56496 -66630 56506 -66380
rect 57016 -66630 57026 -66380
rect 56496 -66635 57026 -66630
rect 55955 -66698 56200 -66688
rect 53510 -66778 53645 -66768
rect 55275 -66718 55490 -66708
rect 53045 -66958 53255 -66948
rect 53045 -68708 53050 -66958
rect 53250 -68708 53255 -66958
rect 53045 -68718 53255 -68708
rect 53510 -68918 53630 -66778
rect 55275 -66808 55280 -66718
rect 55400 -66808 55490 -66718
rect 56060 -66738 56200 -66698
rect 56060 -66748 56220 -66738
rect 55275 -66818 55490 -66808
rect 55220 -67058 55325 -67048
rect 55220 -67228 55230 -67058
rect 55320 -67228 55325 -67058
rect 55220 -67238 55325 -67228
rect 55015 -67848 55125 -67838
rect 55015 -67928 55020 -67848
rect 55120 -67928 55125 -67848
rect 55015 -67938 55125 -67928
rect 55220 -68538 55310 -67238
rect 55215 -68548 55315 -68538
rect 55215 -68718 55220 -68548
rect 55310 -68638 55315 -68548
rect 55400 -68548 55490 -66818
rect 55875 -66818 55990 -66808
rect 55875 -66858 55880 -66818
rect 55870 -66898 55880 -66858
rect 55970 -66898 55990 -66818
rect 55870 -66978 55990 -66898
rect 56060 -66918 56220 -66908
rect 55590 -67068 55720 -67058
rect 55590 -67198 55600 -67068
rect 55710 -67198 55720 -67068
rect 55400 -68558 55510 -68548
rect 55310 -68718 55320 -68638
rect 55400 -68718 55410 -68558
rect 55215 -68728 55320 -68718
rect 53505 -68928 53635 -68918
rect 53505 -69048 53510 -68928
rect 53630 -69048 53635 -68928
rect 53505 -69058 53635 -69048
rect 55220 -69208 55320 -68728
rect 55405 -68728 55410 -68718
rect 55500 -68728 55510 -68558
rect 55405 -68738 55510 -68728
rect 55590 -68988 55720 -67198
rect 55870 -67358 55980 -66978
rect 57093 -67364 57373 -67354
rect 56475 -67388 56555 -67378
rect 56470 -67448 56480 -67388
rect 56550 -67448 56555 -67388
rect 56470 -67458 56555 -67448
rect 55870 -67838 55980 -67468
rect 55870 -67928 55880 -67838
rect 55970 -67928 55980 -67838
rect 55870 -68328 55980 -67928
rect 56470 -67828 56550 -67458
rect 57093 -67504 57098 -67364
rect 57368 -67504 57373 -67364
rect 57093 -67514 57373 -67504
rect 57760 -67820 58280 -62540
rect 58516 -62460 58796 -62390
rect 58516 -62660 58556 -62460
rect 58756 -62660 58796 -62460
rect 59066 -62410 59176 -61910
rect 59266 -62020 59366 -61590
rect 59536 -61490 59616 -61300
rect 59536 -61550 59546 -61490
rect 59606 -61550 59616 -61490
rect 59536 -61610 59616 -61550
rect 59536 -61670 59546 -61610
rect 59606 -61670 59616 -61610
rect 59536 -61680 59616 -61670
rect 59266 -62030 59376 -62020
rect 59266 -62120 59286 -62030
rect 59366 -62120 59376 -62030
rect 59736 -62050 59796 -61300
rect 59856 -61540 59976 -61530
rect 59856 -61630 59866 -61540
rect 59966 -61630 59976 -61540
rect 59856 -61640 59976 -61630
rect 60036 -61720 60136 -61090
rect 61026 -61120 61136 -61110
rect 61026 -61250 61056 -61120
rect 61126 -61250 61136 -61120
rect 60436 -61520 60536 -61510
rect 60436 -61620 60446 -61520
rect 60526 -61620 60536 -61520
rect 60436 -61630 60536 -61620
rect 60036 -61800 60046 -61720
rect 60126 -61800 60136 -61720
rect 60036 -61810 60136 -61800
rect 60546 -61810 60636 -61800
rect 60386 -61890 60556 -61810
rect 60626 -61890 60636 -61810
rect 59966 -61900 60326 -61890
rect 59966 -61970 59976 -61900
rect 60316 -61970 60326 -61900
rect 60546 -61910 60636 -61890
rect 59966 -61980 60326 -61970
rect 59566 -62070 59796 -62050
rect 59566 -62080 59576 -62070
rect 59266 -62130 59376 -62120
rect 59516 -62130 59576 -62080
rect 59636 -62130 59796 -62070
rect 59266 -62240 59366 -62130
rect 59266 -62330 59286 -62240
rect 59356 -62330 59366 -62240
rect 59266 -62360 59366 -62330
rect 59516 -62140 59796 -62130
rect 59066 -62480 59076 -62410
rect 59166 -62480 59176 -62410
rect 59066 -62490 59176 -62480
rect 59306 -62430 59386 -62420
rect 59306 -62490 59316 -62430
rect 59376 -62490 59386 -62430
rect 59516 -62470 59596 -62140
rect 60286 -62150 60476 -62140
rect 59906 -62180 60016 -62170
rect 59906 -62360 59916 -62180
rect 60006 -62360 60016 -62180
rect 59906 -62370 60016 -62360
rect 60286 -62290 60306 -62150
rect 60456 -62290 60476 -62150
rect 60286 -62300 60476 -62290
rect 58516 -62740 58796 -62660
rect 59066 -62570 59176 -62560
rect 59066 -62640 59076 -62570
rect 59166 -62640 59176 -62570
rect 59066 -63140 59176 -62640
rect 59306 -62690 59386 -62490
rect 60076 -62480 60196 -62440
rect 60076 -62640 60096 -62480
rect 60176 -62640 60196 -62480
rect 60076 -62680 60196 -62640
rect 59066 -63200 59076 -63140
rect 59166 -63200 59176 -63140
rect 59066 -63210 59176 -63200
rect 59236 -62720 59386 -62690
rect 59236 -62810 59266 -62720
rect 59366 -62810 59386 -62720
rect 59236 -62830 59386 -62810
rect 59906 -62690 60016 -62680
rect 59236 -62960 59376 -62830
rect 59906 -62880 59916 -62690
rect 60006 -62880 60016 -62690
rect 59906 -62890 60016 -62880
rect 60286 -62710 60376 -62300
rect 60556 -62700 60626 -61910
rect 61026 -62220 61136 -61250
rect 61196 -61920 61356 -61910
rect 61196 -62100 61206 -61920
rect 61346 -62100 61356 -61920
rect 61196 -62110 61356 -62100
rect 61026 -62330 61036 -62220
rect 61126 -62330 61136 -62220
rect 61026 -62340 61136 -62330
rect 61246 -62450 61366 -62440
rect 61246 -62460 61276 -62450
rect 61246 -62660 61256 -62460
rect 61356 -62660 61366 -62450
rect 61246 -62670 61366 -62660
rect 60466 -62710 60626 -62700
rect 60286 -62770 60406 -62710
rect 60466 -62770 60476 -62710
rect 60536 -62770 60626 -62710
rect 59236 -63050 59266 -62960
rect 59366 -63050 59376 -62960
rect 59236 -63100 59376 -63050
rect 59506 -62910 59606 -62900
rect 59506 -62980 59516 -62910
rect 59596 -62980 59606 -62910
rect 59506 -62990 59606 -62980
rect 59236 -63120 59386 -63100
rect 59236 -63180 59316 -63120
rect 59376 -63180 59386 -63120
rect 58396 -63750 58896 -63250
rect 59236 -63430 59386 -63180
rect 59006 -63500 59086 -63480
rect 59236 -63490 59256 -63430
rect 59366 -63490 59386 -63430
rect 59236 -63500 59386 -63490
rect 59506 -63380 59596 -62990
rect 59986 -63120 60116 -63110
rect 59986 -63180 59996 -63120
rect 60106 -63180 60116 -63120
rect 59506 -63390 59616 -63380
rect 59506 -63460 59546 -63390
rect 59606 -63460 59616 -63390
rect 59006 -63560 59016 -63500
rect 59076 -63560 59086 -63500
rect 59006 -63750 59086 -63560
rect 59506 -63510 59616 -63460
rect 59506 -63570 59546 -63510
rect 59606 -63570 59616 -63510
rect 59796 -63410 59926 -63400
rect 59796 -63520 59806 -63410
rect 59916 -63520 59926 -63410
rect 59796 -63530 59926 -63520
rect 59006 -63840 59126 -63750
rect 59006 -63910 59016 -63840
rect 59076 -63910 59126 -63840
rect 59006 -63990 59126 -63910
rect 59506 -63840 59616 -63570
rect 59506 -63910 59546 -63840
rect 59606 -63910 59616 -63840
rect 59506 -63920 59616 -63910
rect 59986 -63990 60116 -63180
rect 60286 -63670 60376 -62770
rect 60466 -62780 60626 -62770
rect 61486 -62770 61726 -62740
rect 61486 -62820 61496 -62770
rect 61326 -62830 61496 -62820
rect 61326 -62950 61336 -62830
rect 61196 -62960 61336 -62950
rect 61456 -62940 61496 -62830
rect 61696 -62940 61726 -62770
rect 61456 -62960 61726 -62940
rect 61196 -62970 61726 -62960
rect 61196 -63140 61426 -62970
rect 60436 -63430 60536 -63410
rect 60436 -63550 60446 -63430
rect 60526 -63550 60536 -63430
rect 60436 -63560 60536 -63550
rect 60256 -63800 60416 -63670
rect 60256 -63930 60266 -63800
rect 60406 -63930 60416 -63800
rect 60256 -63950 60416 -63930
rect 58956 -64000 59156 -63990
rect 58956 -64180 58966 -64000
rect 59146 -64180 59156 -64000
rect 59986 -64100 59996 -63990
rect 60106 -64100 60116 -63990
rect 58956 -64190 59156 -64180
rect 59600 -64200 66500 -64100
rect 59600 -64600 59700 -64200
rect 60400 -64600 66100 -64200
rect 66400 -64600 66500 -64200
rect 59600 -64700 66500 -64600
rect 58946 -66270 59146 -66250
rect 58946 -66430 58966 -66270
rect 59126 -66430 59146 -66270
rect 58946 -66450 59146 -66430
rect 59316 -66310 59426 -66250
rect 59316 -66450 59336 -66310
rect 59416 -66450 59426 -66310
rect 58956 -66530 59136 -66450
rect 58956 -66640 58996 -66530
rect 59106 -66640 59136 -66530
rect 58396 -66730 58896 -66640
rect 58956 -66700 59136 -66640
rect 59316 -66680 59426 -66450
rect 59946 -66320 60386 -66200
rect 59946 -66440 60046 -66320
rect 60126 -66440 60386 -66320
rect 59946 -66490 60386 -66440
rect 58396 -67090 58486 -66730
rect 58816 -67090 58896 -66730
rect 58996 -67000 59086 -66700
rect 58996 -67060 59006 -67000
rect 59066 -67060 59086 -67000
rect 58996 -67070 59086 -67060
rect 59266 -66730 59426 -66680
rect 59506 -66540 59796 -66500
rect 59506 -66640 59516 -66540
rect 59616 -66640 59796 -66540
rect 59506 -66700 59796 -66640
rect 59266 -66930 59366 -66730
rect 59266 -66990 59286 -66930
rect 59346 -66990 59366 -66930
rect 58396 -67200 58896 -67090
rect 59066 -67240 59176 -67230
rect 59066 -67310 59076 -67240
rect 59166 -67310 59176 -67240
rect 56470 -67838 56555 -67828
rect 56470 -67928 56480 -67838
rect 56550 -67928 56555 -67838
rect 56470 -67938 56555 -67928
rect 56470 -68318 56550 -67938
rect 57760 -67940 57800 -67820
rect 58240 -67940 58280 -67820
rect 57093 -68274 57373 -68264
rect 56470 -68328 56555 -68318
rect 56470 -68378 56480 -68328
rect 56475 -68388 56480 -68378
rect 56550 -68388 56555 -68328
rect 56475 -68398 56555 -68388
rect 57093 -68414 57098 -68274
rect 57368 -68414 57373 -68274
rect 57093 -68424 57373 -68414
rect 55870 -68878 55980 -68438
rect 55870 -68918 55880 -68878
rect 55875 -68958 55880 -68918
rect 55970 -68918 55980 -68878
rect 56060 -68868 56220 -68858
rect 55970 -68958 55975 -68918
rect 55875 -68968 55975 -68958
rect 55590 -69078 55620 -68988
rect 55710 -69078 55720 -68988
rect 56060 -69038 56220 -69028
rect 56060 -69048 56200 -69038
rect 55590 -69088 55720 -69078
rect 56015 -69058 56200 -69048
rect 56015 -69208 56020 -69058
rect 56080 -69208 56200 -69058
rect 56644 -69068 57008 -69063
rect 55215 -69218 55325 -69208
rect 56015 -69218 56085 -69208
rect 55215 -69318 55220 -69218
rect 55320 -69318 55325 -69218
rect 56644 -69286 56654 -69068
rect 56998 -69286 57008 -69068
rect 56644 -69291 57008 -69286
rect 55215 -69328 55325 -69318
rect 55315 -69528 55475 -69518
rect 55315 -69668 55320 -69528
rect 55470 -69668 55475 -69528
rect 55315 -69678 55475 -69668
rect 40100 -70000 40800 -69900
rect 40100 -70600 40200 -70000
rect 40700 -70100 56200 -70000
rect 40700 -70500 55500 -70100
rect 56100 -70500 56200 -70100
rect 40700 -70600 56200 -70500
rect 40100 -70700 40800 -70600
rect 51400 -71080 55800 -71000
rect 51400 -71100 55460 -71080
rect 51400 -71300 51500 -71100
rect 52500 -71300 55460 -71100
rect 51400 -71360 55460 -71300
rect 55720 -71360 55800 -71080
rect 51400 -71400 55800 -71360
rect 55380 -71440 55800 -71400
rect 47700 -71600 48100 -71580
rect 47700 -72060 47720 -71600
rect 48080 -71720 48100 -71600
rect 48080 -71740 53800 -71720
rect 48080 -71940 53480 -71740
rect 53780 -71940 53800 -71740
rect 56496 -71780 57026 -71775
rect 48080 -71960 53800 -71940
rect 55955 -71938 56045 -71928
rect 48080 -72060 48100 -71960
rect 53515 -72058 53645 -72048
rect 47700 -72080 48100 -72060
rect 53510 -72168 53520 -72058
rect 53640 -72168 53645 -72058
rect 55955 -72088 55960 -71938
rect 56040 -72088 56200 -71938
rect 56496 -72030 56506 -71780
rect 57016 -72030 57026 -71780
rect 56496 -72035 57026 -72030
rect 55955 -72098 56200 -72088
rect 53510 -72178 53645 -72168
rect 55275 -72118 55490 -72108
rect 53045 -72358 53255 -72348
rect 53045 -74108 53050 -72358
rect 53250 -74108 53255 -72358
rect 53045 -74118 53255 -74108
rect 53510 -74318 53630 -72178
rect 55275 -72208 55280 -72118
rect 55400 -72208 55490 -72118
rect 56060 -72138 56200 -72098
rect 56060 -72148 56220 -72138
rect 55275 -72218 55490 -72208
rect 55220 -72458 55325 -72448
rect 55220 -72628 55230 -72458
rect 55320 -72628 55325 -72458
rect 55220 -72638 55325 -72628
rect 55015 -73248 55125 -73238
rect 55015 -73328 55020 -73248
rect 55120 -73328 55125 -73248
rect 55015 -73338 55125 -73328
rect 55220 -73938 55310 -72638
rect 55215 -73948 55315 -73938
rect 55215 -74118 55220 -73948
rect 55310 -74038 55315 -73948
rect 55400 -73948 55490 -72218
rect 55875 -72218 55990 -72208
rect 55875 -72258 55880 -72218
rect 55870 -72298 55880 -72258
rect 55970 -72298 55990 -72218
rect 55870 -72378 55990 -72298
rect 56060 -72318 56220 -72308
rect 55590 -72468 55720 -72458
rect 55590 -72598 55600 -72468
rect 55710 -72598 55720 -72468
rect 55400 -73958 55510 -73948
rect 55310 -74118 55320 -74038
rect 55400 -74118 55410 -73958
rect 55215 -74128 55320 -74118
rect 53505 -74328 53635 -74318
rect 53505 -74448 53510 -74328
rect 53630 -74448 53635 -74328
rect 53505 -74458 53635 -74448
rect 55220 -74608 55320 -74128
rect 55405 -74128 55410 -74118
rect 55500 -74128 55510 -73958
rect 55405 -74138 55510 -74128
rect 55590 -74388 55720 -72598
rect 55870 -72758 55980 -72378
rect 57093 -72764 57373 -72754
rect 56475 -72788 56555 -72778
rect 56470 -72848 56480 -72788
rect 56550 -72848 56555 -72788
rect 56470 -72858 56555 -72848
rect 55870 -73238 55980 -72868
rect 55870 -73328 55880 -73238
rect 55970 -73328 55980 -73238
rect 55870 -73728 55980 -73328
rect 56470 -73228 56550 -72858
rect 57093 -72904 57098 -72764
rect 57368 -72904 57373 -72764
rect 57093 -72914 57373 -72904
rect 57760 -73220 58280 -67940
rect 58516 -67860 58796 -67790
rect 58516 -68060 58556 -67860
rect 58756 -68060 58796 -67860
rect 59066 -67810 59176 -67310
rect 59266 -67420 59366 -66990
rect 59536 -66890 59616 -66700
rect 59536 -66950 59546 -66890
rect 59606 -66950 59616 -66890
rect 59536 -67010 59616 -66950
rect 59536 -67070 59546 -67010
rect 59606 -67070 59616 -67010
rect 59536 -67080 59616 -67070
rect 59266 -67430 59376 -67420
rect 59266 -67520 59286 -67430
rect 59366 -67520 59376 -67430
rect 59736 -67450 59796 -66700
rect 59856 -66940 59976 -66930
rect 59856 -67030 59866 -66940
rect 59966 -67030 59976 -66940
rect 59856 -67040 59976 -67030
rect 60036 -67120 60136 -66490
rect 61026 -66520 61136 -66510
rect 61026 -66650 61056 -66520
rect 61126 -66650 61136 -66520
rect 60436 -66920 60536 -66910
rect 60436 -67020 60446 -66920
rect 60526 -67020 60536 -66920
rect 60436 -67030 60536 -67020
rect 60036 -67200 60046 -67120
rect 60126 -67200 60136 -67120
rect 60036 -67210 60136 -67200
rect 60546 -67210 60636 -67200
rect 60386 -67290 60556 -67210
rect 60626 -67290 60636 -67210
rect 59966 -67300 60326 -67290
rect 59966 -67370 59976 -67300
rect 60316 -67370 60326 -67300
rect 60546 -67310 60636 -67290
rect 59966 -67380 60326 -67370
rect 59566 -67470 59796 -67450
rect 59566 -67480 59576 -67470
rect 59266 -67530 59376 -67520
rect 59516 -67530 59576 -67480
rect 59636 -67530 59796 -67470
rect 59266 -67640 59366 -67530
rect 59266 -67730 59286 -67640
rect 59356 -67730 59366 -67640
rect 59266 -67760 59366 -67730
rect 59516 -67540 59796 -67530
rect 59066 -67880 59076 -67810
rect 59166 -67880 59176 -67810
rect 59066 -67890 59176 -67880
rect 59306 -67830 59386 -67820
rect 59306 -67890 59316 -67830
rect 59376 -67890 59386 -67830
rect 59516 -67870 59596 -67540
rect 60286 -67550 60476 -67540
rect 59906 -67580 60016 -67570
rect 59906 -67760 59916 -67580
rect 60006 -67760 60016 -67580
rect 59906 -67770 60016 -67760
rect 60286 -67690 60306 -67550
rect 60456 -67690 60476 -67550
rect 60286 -67700 60476 -67690
rect 58516 -68140 58796 -68060
rect 59066 -67970 59176 -67960
rect 59066 -68040 59076 -67970
rect 59166 -68040 59176 -67970
rect 59066 -68540 59176 -68040
rect 59306 -68090 59386 -67890
rect 60076 -67880 60196 -67840
rect 60076 -68040 60096 -67880
rect 60176 -68040 60196 -67880
rect 60076 -68080 60196 -68040
rect 59066 -68600 59076 -68540
rect 59166 -68600 59176 -68540
rect 59066 -68610 59176 -68600
rect 59236 -68120 59386 -68090
rect 59236 -68210 59266 -68120
rect 59366 -68210 59386 -68120
rect 59236 -68230 59386 -68210
rect 59906 -68090 60016 -68080
rect 59236 -68360 59376 -68230
rect 59906 -68280 59916 -68090
rect 60006 -68280 60016 -68090
rect 59906 -68290 60016 -68280
rect 60286 -68110 60376 -67700
rect 60556 -68100 60626 -67310
rect 61026 -67620 61136 -66650
rect 61196 -67320 61356 -67310
rect 61196 -67500 61206 -67320
rect 61346 -67500 61356 -67320
rect 61196 -67510 61356 -67500
rect 61026 -67730 61036 -67620
rect 61126 -67730 61136 -67620
rect 61026 -67740 61136 -67730
rect 61246 -67850 61366 -67840
rect 61246 -67860 61276 -67850
rect 61246 -68060 61256 -67860
rect 61356 -68060 61366 -67850
rect 61246 -68070 61366 -68060
rect 60466 -68110 60626 -68100
rect 60286 -68170 60406 -68110
rect 60466 -68170 60476 -68110
rect 60536 -68170 60626 -68110
rect 59236 -68450 59266 -68360
rect 59366 -68450 59376 -68360
rect 59236 -68500 59376 -68450
rect 59506 -68310 59606 -68300
rect 59506 -68380 59516 -68310
rect 59596 -68380 59606 -68310
rect 59506 -68390 59606 -68380
rect 59236 -68520 59386 -68500
rect 59236 -68580 59316 -68520
rect 59376 -68580 59386 -68520
rect 58396 -69150 58896 -68650
rect 59236 -68830 59386 -68580
rect 59006 -68900 59086 -68880
rect 59236 -68890 59256 -68830
rect 59366 -68890 59386 -68830
rect 59236 -68900 59386 -68890
rect 59506 -68780 59596 -68390
rect 59986 -68520 60116 -68510
rect 59986 -68580 59996 -68520
rect 60106 -68580 60116 -68520
rect 59506 -68790 59616 -68780
rect 59506 -68860 59546 -68790
rect 59606 -68860 59616 -68790
rect 59006 -68960 59016 -68900
rect 59076 -68960 59086 -68900
rect 59006 -69150 59086 -68960
rect 59506 -68910 59616 -68860
rect 59506 -68970 59546 -68910
rect 59606 -68970 59616 -68910
rect 59796 -68810 59926 -68800
rect 59796 -68920 59806 -68810
rect 59916 -68920 59926 -68810
rect 59796 -68930 59926 -68920
rect 59006 -69240 59126 -69150
rect 59006 -69310 59016 -69240
rect 59076 -69310 59126 -69240
rect 59006 -69390 59126 -69310
rect 59506 -69240 59616 -68970
rect 59506 -69310 59546 -69240
rect 59606 -69310 59616 -69240
rect 59506 -69320 59616 -69310
rect 59986 -69390 60116 -68580
rect 60286 -69070 60376 -68170
rect 60466 -68180 60626 -68170
rect 61486 -68170 61726 -68140
rect 61486 -68220 61496 -68170
rect 61326 -68230 61496 -68220
rect 61326 -68350 61336 -68230
rect 61196 -68360 61336 -68350
rect 61456 -68340 61496 -68230
rect 61696 -68340 61726 -68170
rect 61456 -68360 61726 -68340
rect 61196 -68370 61726 -68360
rect 61196 -68540 61426 -68370
rect 60436 -68830 60536 -68810
rect 60436 -68950 60446 -68830
rect 60526 -68950 60536 -68830
rect 60436 -68960 60536 -68950
rect 60256 -69200 60416 -69070
rect 60256 -69330 60266 -69200
rect 60406 -69330 60416 -69200
rect 60256 -69350 60416 -69330
rect 58956 -69400 59156 -69390
rect 58956 -69580 58966 -69400
rect 59146 -69580 59156 -69400
rect 59986 -69500 59996 -69390
rect 60106 -69500 60116 -69390
rect 58956 -69590 59156 -69580
rect 59600 -69600 67500 -69500
rect 59600 -70000 59700 -69600
rect 60400 -70000 67100 -69600
rect 67400 -70000 67500 -69600
rect 59600 -70100 67500 -70000
rect 58946 -71670 59146 -71650
rect 58946 -71830 58966 -71670
rect 59126 -71830 59146 -71670
rect 58946 -71850 59146 -71830
rect 59316 -71710 59426 -71650
rect 59316 -71850 59336 -71710
rect 59416 -71850 59426 -71710
rect 58956 -71930 59136 -71850
rect 58956 -72040 58996 -71930
rect 59106 -72040 59136 -71930
rect 58396 -72130 58896 -72040
rect 58956 -72100 59136 -72040
rect 59316 -72080 59426 -71850
rect 59946 -71720 60386 -71600
rect 59946 -71840 60046 -71720
rect 60126 -71840 60386 -71720
rect 59946 -71890 60386 -71840
rect 58396 -72490 58486 -72130
rect 58816 -72490 58896 -72130
rect 58996 -72400 59086 -72100
rect 58996 -72460 59006 -72400
rect 59066 -72460 59086 -72400
rect 58996 -72470 59086 -72460
rect 59266 -72130 59426 -72080
rect 59506 -71940 59796 -71900
rect 59506 -72040 59516 -71940
rect 59616 -72040 59796 -71940
rect 59506 -72100 59796 -72040
rect 59266 -72330 59366 -72130
rect 59266 -72390 59286 -72330
rect 59346 -72390 59366 -72330
rect 58396 -72600 58896 -72490
rect 59066 -72640 59176 -72630
rect 59066 -72710 59076 -72640
rect 59166 -72710 59176 -72640
rect 56470 -73238 56555 -73228
rect 56470 -73328 56480 -73238
rect 56550 -73328 56555 -73238
rect 56470 -73338 56555 -73328
rect 56470 -73718 56550 -73338
rect 57760 -73340 57800 -73220
rect 58240 -73340 58280 -73220
rect 57093 -73674 57373 -73664
rect 56470 -73728 56555 -73718
rect 56470 -73778 56480 -73728
rect 56475 -73788 56480 -73778
rect 56550 -73788 56555 -73728
rect 56475 -73798 56555 -73788
rect 57093 -73814 57098 -73674
rect 57368 -73814 57373 -73674
rect 57093 -73824 57373 -73814
rect 55870 -74278 55980 -73838
rect 55870 -74318 55880 -74278
rect 55875 -74358 55880 -74318
rect 55970 -74318 55980 -74278
rect 56060 -74268 56220 -74258
rect 55970 -74358 55975 -74318
rect 55875 -74368 55975 -74358
rect 55590 -74478 55620 -74388
rect 55710 -74478 55720 -74388
rect 56060 -74438 56220 -74428
rect 56060 -74448 56200 -74438
rect 55590 -74488 55720 -74478
rect 56015 -74458 56200 -74448
rect 56015 -74608 56020 -74458
rect 56080 -74608 56200 -74458
rect 56644 -74468 57008 -74463
rect 55215 -74618 55325 -74608
rect 56015 -74618 56085 -74608
rect 55215 -74718 55220 -74618
rect 55320 -74718 55325 -74618
rect 56644 -74686 56654 -74468
rect 56998 -74686 57008 -74468
rect 56644 -74691 57008 -74686
rect 55215 -74728 55325 -74718
rect 55315 -74928 55475 -74918
rect 55315 -75068 55320 -74928
rect 55470 -75068 55475 -74928
rect 55315 -75078 55475 -75068
rect 39200 -75400 39900 -75300
rect 39200 -76000 39300 -75400
rect 39800 -75500 56200 -75400
rect 39800 -75900 55500 -75500
rect 56100 -75900 56200 -75500
rect 39800 -76000 56200 -75900
rect 39200 -76100 39900 -76000
rect 51400 -76480 55800 -76400
rect 51400 -76500 55400 -76480
rect 51400 -76700 51500 -76500
rect 52500 -76700 55400 -76500
rect 51400 -76760 55400 -76700
rect 55720 -76760 55800 -76480
rect 51400 -76800 55800 -76760
rect 55320 -76840 55800 -76800
rect 47760 -76940 48100 -76920
rect 47760 -77500 47780 -76940
rect 48080 -77120 48100 -76940
rect 48080 -77140 53800 -77120
rect 48080 -77340 53480 -77140
rect 53780 -77340 53800 -77140
rect 56496 -77180 57026 -77175
rect 48080 -77360 53800 -77340
rect 55955 -77338 56045 -77328
rect 48080 -77500 48100 -77360
rect 53515 -77458 53645 -77448
rect 47760 -77520 48100 -77500
rect 53510 -77568 53520 -77458
rect 53640 -77568 53645 -77458
rect 55955 -77488 55960 -77338
rect 56040 -77488 56200 -77338
rect 56496 -77430 56506 -77180
rect 57016 -77430 57026 -77180
rect 56496 -77435 57026 -77430
rect 55955 -77498 56200 -77488
rect 53510 -77578 53645 -77568
rect 55275 -77518 55490 -77508
rect 53045 -77758 53255 -77748
rect 53045 -79508 53050 -77758
rect 53250 -79508 53255 -77758
rect 53045 -79518 53255 -79508
rect 53510 -79718 53630 -77578
rect 55275 -77608 55280 -77518
rect 55400 -77608 55490 -77518
rect 56060 -77538 56200 -77498
rect 56060 -77548 56220 -77538
rect 55275 -77618 55490 -77608
rect 55220 -77858 55325 -77848
rect 55220 -78028 55230 -77858
rect 55320 -78028 55325 -77858
rect 55220 -78038 55325 -78028
rect 55015 -78648 55125 -78638
rect 55015 -78728 55020 -78648
rect 55120 -78728 55125 -78648
rect 55015 -78738 55125 -78728
rect 55220 -79338 55310 -78038
rect 55215 -79348 55315 -79338
rect 55215 -79518 55220 -79348
rect 55310 -79438 55315 -79348
rect 55400 -79348 55490 -77618
rect 55875 -77618 55990 -77608
rect 55875 -77658 55880 -77618
rect 55870 -77698 55880 -77658
rect 55970 -77698 55990 -77618
rect 55870 -77778 55990 -77698
rect 56060 -77718 56220 -77708
rect 55590 -77868 55720 -77858
rect 55590 -77998 55600 -77868
rect 55710 -77998 55720 -77868
rect 55400 -79358 55510 -79348
rect 55310 -79518 55320 -79438
rect 55400 -79518 55410 -79358
rect 55215 -79528 55320 -79518
rect 53505 -79728 53635 -79718
rect 53505 -79848 53510 -79728
rect 53630 -79848 53635 -79728
rect 53505 -79858 53635 -79848
rect 55220 -80008 55320 -79528
rect 55405 -79528 55410 -79518
rect 55500 -79528 55510 -79358
rect 55405 -79538 55510 -79528
rect 55590 -79788 55720 -77998
rect 55870 -78158 55980 -77778
rect 57093 -78164 57373 -78154
rect 56475 -78188 56555 -78178
rect 56470 -78248 56480 -78188
rect 56550 -78248 56555 -78188
rect 56470 -78258 56555 -78248
rect 55870 -78638 55980 -78268
rect 55870 -78728 55880 -78638
rect 55970 -78728 55980 -78638
rect 55870 -79128 55980 -78728
rect 56470 -78628 56550 -78258
rect 57093 -78304 57098 -78164
rect 57368 -78304 57373 -78164
rect 57093 -78314 57373 -78304
rect 57760 -78620 58280 -73340
rect 58516 -73260 58796 -73190
rect 58516 -73460 58556 -73260
rect 58756 -73460 58796 -73260
rect 59066 -73210 59176 -72710
rect 59266 -72820 59366 -72390
rect 59536 -72290 59616 -72100
rect 59536 -72350 59546 -72290
rect 59606 -72350 59616 -72290
rect 59536 -72410 59616 -72350
rect 59536 -72470 59546 -72410
rect 59606 -72470 59616 -72410
rect 59536 -72480 59616 -72470
rect 59266 -72830 59376 -72820
rect 59266 -72920 59286 -72830
rect 59366 -72920 59376 -72830
rect 59736 -72850 59796 -72100
rect 59856 -72340 59976 -72330
rect 59856 -72430 59866 -72340
rect 59966 -72430 59976 -72340
rect 59856 -72440 59976 -72430
rect 60036 -72520 60136 -71890
rect 61026 -71920 61136 -71910
rect 61026 -72050 61056 -71920
rect 61126 -72050 61136 -71920
rect 60436 -72320 60536 -72310
rect 60436 -72420 60446 -72320
rect 60526 -72420 60536 -72320
rect 60436 -72430 60536 -72420
rect 60036 -72600 60046 -72520
rect 60126 -72600 60136 -72520
rect 60036 -72610 60136 -72600
rect 60546 -72610 60636 -72600
rect 60386 -72690 60556 -72610
rect 60626 -72690 60636 -72610
rect 59966 -72700 60326 -72690
rect 59966 -72770 59976 -72700
rect 60316 -72770 60326 -72700
rect 60546 -72710 60636 -72690
rect 59966 -72780 60326 -72770
rect 59566 -72870 59796 -72850
rect 59566 -72880 59576 -72870
rect 59266 -72930 59376 -72920
rect 59516 -72930 59576 -72880
rect 59636 -72930 59796 -72870
rect 59266 -73040 59366 -72930
rect 59266 -73130 59286 -73040
rect 59356 -73130 59366 -73040
rect 59266 -73160 59366 -73130
rect 59516 -72940 59796 -72930
rect 59066 -73280 59076 -73210
rect 59166 -73280 59176 -73210
rect 59066 -73290 59176 -73280
rect 59306 -73230 59386 -73220
rect 59306 -73290 59316 -73230
rect 59376 -73290 59386 -73230
rect 59516 -73270 59596 -72940
rect 60286 -72950 60476 -72940
rect 59906 -72980 60016 -72970
rect 59906 -73160 59916 -72980
rect 60006 -73160 60016 -72980
rect 59906 -73170 60016 -73160
rect 60286 -73090 60306 -72950
rect 60456 -73090 60476 -72950
rect 60286 -73100 60476 -73090
rect 58516 -73540 58796 -73460
rect 59066 -73370 59176 -73360
rect 59066 -73440 59076 -73370
rect 59166 -73440 59176 -73370
rect 59066 -73940 59176 -73440
rect 59306 -73490 59386 -73290
rect 60076 -73280 60196 -73240
rect 60076 -73440 60096 -73280
rect 60176 -73440 60196 -73280
rect 60076 -73480 60196 -73440
rect 59066 -74000 59076 -73940
rect 59166 -74000 59176 -73940
rect 59066 -74010 59176 -74000
rect 59236 -73520 59386 -73490
rect 59236 -73610 59266 -73520
rect 59366 -73610 59386 -73520
rect 59236 -73630 59386 -73610
rect 59906 -73490 60016 -73480
rect 59236 -73760 59376 -73630
rect 59906 -73680 59916 -73490
rect 60006 -73680 60016 -73490
rect 59906 -73690 60016 -73680
rect 60286 -73510 60376 -73100
rect 60556 -73500 60626 -72710
rect 61026 -73020 61136 -72050
rect 61196 -72720 61356 -72710
rect 61196 -72900 61206 -72720
rect 61346 -72900 61356 -72720
rect 61196 -72910 61356 -72900
rect 61026 -73130 61036 -73020
rect 61126 -73130 61136 -73020
rect 61026 -73140 61136 -73130
rect 61246 -73250 61366 -73240
rect 61246 -73260 61276 -73250
rect 61246 -73460 61256 -73260
rect 61356 -73460 61366 -73250
rect 61246 -73470 61366 -73460
rect 60466 -73510 60626 -73500
rect 60286 -73570 60406 -73510
rect 60466 -73570 60476 -73510
rect 60536 -73570 60626 -73510
rect 59236 -73850 59266 -73760
rect 59366 -73850 59376 -73760
rect 59236 -73900 59376 -73850
rect 59506 -73710 59606 -73700
rect 59506 -73780 59516 -73710
rect 59596 -73780 59606 -73710
rect 59506 -73790 59606 -73780
rect 59236 -73920 59386 -73900
rect 59236 -73980 59316 -73920
rect 59376 -73980 59386 -73920
rect 58396 -74550 58896 -74050
rect 59236 -74230 59386 -73980
rect 59006 -74300 59086 -74280
rect 59236 -74290 59256 -74230
rect 59366 -74290 59386 -74230
rect 59236 -74300 59386 -74290
rect 59506 -74180 59596 -73790
rect 59986 -73920 60116 -73910
rect 59986 -73980 59996 -73920
rect 60106 -73980 60116 -73920
rect 59506 -74190 59616 -74180
rect 59506 -74260 59546 -74190
rect 59606 -74260 59616 -74190
rect 59006 -74360 59016 -74300
rect 59076 -74360 59086 -74300
rect 59006 -74550 59086 -74360
rect 59506 -74310 59616 -74260
rect 59506 -74370 59546 -74310
rect 59606 -74370 59616 -74310
rect 59796 -74210 59926 -74200
rect 59796 -74320 59806 -74210
rect 59916 -74320 59926 -74210
rect 59796 -74330 59926 -74320
rect 59006 -74640 59126 -74550
rect 59006 -74710 59016 -74640
rect 59076 -74710 59126 -74640
rect 59006 -74790 59126 -74710
rect 59506 -74640 59616 -74370
rect 59506 -74710 59546 -74640
rect 59606 -74710 59616 -74640
rect 59506 -74720 59616 -74710
rect 59986 -74790 60116 -73980
rect 60286 -74470 60376 -73570
rect 60466 -73580 60626 -73570
rect 61486 -73570 61726 -73540
rect 61486 -73620 61496 -73570
rect 61326 -73630 61496 -73620
rect 61326 -73750 61336 -73630
rect 61196 -73760 61336 -73750
rect 61456 -73740 61496 -73630
rect 61696 -73740 61726 -73570
rect 61456 -73760 61726 -73740
rect 61196 -73770 61726 -73760
rect 61196 -73940 61426 -73770
rect 60436 -74230 60536 -74210
rect 60436 -74350 60446 -74230
rect 60526 -74350 60536 -74230
rect 60436 -74360 60536 -74350
rect 60256 -74600 60416 -74470
rect 60256 -74730 60266 -74600
rect 60406 -74730 60416 -74600
rect 60256 -74750 60416 -74730
rect 58956 -74800 59156 -74790
rect 58956 -74980 58966 -74800
rect 59146 -74980 59156 -74800
rect 59986 -74900 59996 -74790
rect 60106 -74900 60116 -74790
rect 58956 -74990 59156 -74980
rect 59600 -75000 68400 -74900
rect 59600 -75400 59700 -75000
rect 60400 -75400 68000 -75000
rect 68300 -75400 68400 -75000
rect 59600 -75500 68400 -75400
rect 58946 -77070 59146 -77050
rect 58946 -77230 58966 -77070
rect 59126 -77230 59146 -77070
rect 58946 -77250 59146 -77230
rect 59316 -77110 59426 -77050
rect 59316 -77250 59336 -77110
rect 59416 -77250 59426 -77110
rect 58956 -77330 59136 -77250
rect 58956 -77440 58996 -77330
rect 59106 -77440 59136 -77330
rect 58396 -77530 58896 -77440
rect 58956 -77500 59136 -77440
rect 59316 -77480 59426 -77250
rect 59946 -77120 60386 -77000
rect 59946 -77240 60046 -77120
rect 60126 -77240 60386 -77120
rect 59946 -77290 60386 -77240
rect 58396 -77890 58486 -77530
rect 58816 -77890 58896 -77530
rect 58996 -77800 59086 -77500
rect 58996 -77860 59006 -77800
rect 59066 -77860 59086 -77800
rect 58996 -77870 59086 -77860
rect 59266 -77530 59426 -77480
rect 59506 -77340 59796 -77300
rect 59506 -77440 59516 -77340
rect 59616 -77440 59796 -77340
rect 59506 -77500 59796 -77440
rect 59266 -77730 59366 -77530
rect 59266 -77790 59286 -77730
rect 59346 -77790 59366 -77730
rect 58396 -78000 58896 -77890
rect 59066 -78040 59176 -78030
rect 59066 -78110 59076 -78040
rect 59166 -78110 59176 -78040
rect 56470 -78638 56555 -78628
rect 56470 -78728 56480 -78638
rect 56550 -78728 56555 -78638
rect 56470 -78738 56555 -78728
rect 56470 -79118 56550 -78738
rect 57760 -78740 57800 -78620
rect 58240 -78740 58280 -78620
rect 57093 -79074 57373 -79064
rect 56470 -79128 56555 -79118
rect 56470 -79178 56480 -79128
rect 56475 -79188 56480 -79178
rect 56550 -79188 56555 -79128
rect 56475 -79198 56555 -79188
rect 57093 -79214 57098 -79074
rect 57368 -79214 57373 -79074
rect 57093 -79224 57373 -79214
rect 55870 -79678 55980 -79238
rect 55870 -79718 55880 -79678
rect 55875 -79758 55880 -79718
rect 55970 -79718 55980 -79678
rect 56060 -79668 56220 -79658
rect 55970 -79758 55975 -79718
rect 55875 -79768 55975 -79758
rect 55590 -79878 55620 -79788
rect 55710 -79878 55720 -79788
rect 56060 -79838 56220 -79828
rect 56060 -79848 56200 -79838
rect 55590 -79888 55720 -79878
rect 56015 -79858 56200 -79848
rect 56015 -80008 56020 -79858
rect 56080 -80008 56200 -79858
rect 56644 -79868 57008 -79863
rect 55215 -80018 55325 -80008
rect 56015 -80018 56085 -80008
rect 55215 -80118 55220 -80018
rect 55320 -80118 55325 -80018
rect 56644 -80086 56654 -79868
rect 56998 -80086 57008 -79868
rect 56644 -80091 57008 -80086
rect 55215 -80128 55325 -80118
rect 55315 -80328 55475 -80318
rect 55315 -80468 55320 -80328
rect 55470 -80468 55475 -80328
rect 55315 -80478 55475 -80468
rect 38200 -80800 38900 -80700
rect 38200 -81400 38300 -80800
rect 38800 -80900 56300 -80800
rect 38800 -81300 55500 -80900
rect 56200 -81300 56300 -80900
rect 38800 -81400 56300 -81300
rect 38200 -81500 38900 -81400
rect 51400 -81880 55800 -81800
rect 51400 -81900 55440 -81880
rect 51400 -82100 51500 -81900
rect 52500 -82100 55440 -81900
rect 51400 -82160 55440 -82100
rect 55720 -82160 55800 -81880
rect 51400 -82200 55800 -82160
rect 55360 -82240 55800 -82200
rect 47780 -82380 48100 -82360
rect 47780 -82860 47800 -82380
rect 48080 -82520 48100 -82380
rect 48080 -82540 53800 -82520
rect 48080 -82740 53480 -82540
rect 53780 -82740 53800 -82540
rect 56496 -82580 57026 -82575
rect 48080 -82760 53800 -82740
rect 55955 -82738 56045 -82728
rect 48080 -82860 48100 -82760
rect 53515 -82858 53645 -82848
rect 47780 -82880 48100 -82860
rect 53510 -82968 53520 -82858
rect 53640 -82968 53645 -82858
rect 55955 -82888 55960 -82738
rect 56040 -82888 56200 -82738
rect 56496 -82830 56506 -82580
rect 57016 -82830 57026 -82580
rect 56496 -82835 57026 -82830
rect 55955 -82898 56200 -82888
rect 53510 -82978 53645 -82968
rect 55275 -82918 55490 -82908
rect 53045 -83158 53255 -83148
rect 53045 -84908 53050 -83158
rect 53250 -84908 53255 -83158
rect 53045 -84918 53255 -84908
rect 53510 -85118 53630 -82978
rect 55275 -83008 55280 -82918
rect 55400 -83008 55490 -82918
rect 56060 -82938 56200 -82898
rect 56060 -82948 56220 -82938
rect 55275 -83018 55490 -83008
rect 55220 -83258 55325 -83248
rect 55220 -83428 55230 -83258
rect 55320 -83428 55325 -83258
rect 55220 -83438 55325 -83428
rect 55015 -84048 55125 -84038
rect 55015 -84128 55020 -84048
rect 55120 -84128 55125 -84048
rect 55015 -84138 55125 -84128
rect 55220 -84738 55310 -83438
rect 55215 -84748 55315 -84738
rect 55215 -84918 55220 -84748
rect 55310 -84838 55315 -84748
rect 55400 -84748 55490 -83018
rect 55875 -83018 55990 -83008
rect 55875 -83058 55880 -83018
rect 55870 -83098 55880 -83058
rect 55970 -83098 55990 -83018
rect 55870 -83178 55990 -83098
rect 56060 -83118 56220 -83108
rect 55590 -83268 55720 -83258
rect 55590 -83398 55600 -83268
rect 55710 -83398 55720 -83268
rect 55400 -84758 55510 -84748
rect 55310 -84918 55320 -84838
rect 55400 -84918 55410 -84758
rect 55215 -84928 55320 -84918
rect 53505 -85128 53635 -85118
rect 53505 -85248 53510 -85128
rect 53630 -85248 53635 -85128
rect 53505 -85258 53635 -85248
rect 55220 -85408 55320 -84928
rect 55405 -84928 55410 -84918
rect 55500 -84928 55510 -84758
rect 55405 -84938 55510 -84928
rect 55590 -85188 55720 -83398
rect 55870 -83558 55980 -83178
rect 57093 -83564 57373 -83554
rect 56475 -83588 56555 -83578
rect 56470 -83648 56480 -83588
rect 56550 -83648 56555 -83588
rect 56470 -83658 56555 -83648
rect 55870 -84038 55980 -83668
rect 55870 -84128 55880 -84038
rect 55970 -84128 55980 -84038
rect 55870 -84528 55980 -84128
rect 56470 -84028 56550 -83658
rect 57093 -83704 57098 -83564
rect 57368 -83704 57373 -83564
rect 57093 -83714 57373 -83704
rect 57760 -84020 58280 -78740
rect 58516 -78660 58796 -78590
rect 58516 -78860 58556 -78660
rect 58756 -78860 58796 -78660
rect 59066 -78610 59176 -78110
rect 59266 -78220 59366 -77790
rect 59536 -77690 59616 -77500
rect 59536 -77750 59546 -77690
rect 59606 -77750 59616 -77690
rect 59536 -77810 59616 -77750
rect 59536 -77870 59546 -77810
rect 59606 -77870 59616 -77810
rect 59536 -77880 59616 -77870
rect 59266 -78230 59376 -78220
rect 59266 -78320 59286 -78230
rect 59366 -78320 59376 -78230
rect 59736 -78250 59796 -77500
rect 59856 -77740 59976 -77730
rect 59856 -77830 59866 -77740
rect 59966 -77830 59976 -77740
rect 59856 -77840 59976 -77830
rect 60036 -77920 60136 -77290
rect 61026 -77320 61136 -77310
rect 61026 -77450 61056 -77320
rect 61126 -77450 61136 -77320
rect 60436 -77720 60536 -77710
rect 60436 -77820 60446 -77720
rect 60526 -77820 60536 -77720
rect 60436 -77830 60536 -77820
rect 60036 -78000 60046 -77920
rect 60126 -78000 60136 -77920
rect 60036 -78010 60136 -78000
rect 60546 -78010 60636 -78000
rect 60386 -78090 60556 -78010
rect 60626 -78090 60636 -78010
rect 59966 -78100 60326 -78090
rect 59966 -78170 59976 -78100
rect 60316 -78170 60326 -78100
rect 60546 -78110 60636 -78090
rect 59966 -78180 60326 -78170
rect 59566 -78270 59796 -78250
rect 59566 -78280 59576 -78270
rect 59266 -78330 59376 -78320
rect 59516 -78330 59576 -78280
rect 59636 -78330 59796 -78270
rect 59266 -78440 59366 -78330
rect 59266 -78530 59286 -78440
rect 59356 -78530 59366 -78440
rect 59266 -78560 59366 -78530
rect 59516 -78340 59796 -78330
rect 59066 -78680 59076 -78610
rect 59166 -78680 59176 -78610
rect 59066 -78690 59176 -78680
rect 59306 -78630 59386 -78620
rect 59306 -78690 59316 -78630
rect 59376 -78690 59386 -78630
rect 59516 -78670 59596 -78340
rect 60286 -78350 60476 -78340
rect 59906 -78380 60016 -78370
rect 59906 -78560 59916 -78380
rect 60006 -78560 60016 -78380
rect 59906 -78570 60016 -78560
rect 60286 -78490 60306 -78350
rect 60456 -78490 60476 -78350
rect 60286 -78500 60476 -78490
rect 58516 -78940 58796 -78860
rect 59066 -78770 59176 -78760
rect 59066 -78840 59076 -78770
rect 59166 -78840 59176 -78770
rect 59066 -79340 59176 -78840
rect 59306 -78890 59386 -78690
rect 60076 -78680 60196 -78640
rect 60076 -78840 60096 -78680
rect 60176 -78840 60196 -78680
rect 60076 -78880 60196 -78840
rect 59066 -79400 59076 -79340
rect 59166 -79400 59176 -79340
rect 59066 -79410 59176 -79400
rect 59236 -78920 59386 -78890
rect 59236 -79010 59266 -78920
rect 59366 -79010 59386 -78920
rect 59236 -79030 59386 -79010
rect 59906 -78890 60016 -78880
rect 59236 -79160 59376 -79030
rect 59906 -79080 59916 -78890
rect 60006 -79080 60016 -78890
rect 59906 -79090 60016 -79080
rect 60286 -78910 60376 -78500
rect 60556 -78900 60626 -78110
rect 61026 -78420 61136 -77450
rect 61196 -78120 61356 -78110
rect 61196 -78300 61206 -78120
rect 61346 -78300 61356 -78120
rect 61196 -78310 61356 -78300
rect 61026 -78530 61036 -78420
rect 61126 -78530 61136 -78420
rect 61026 -78540 61136 -78530
rect 61246 -78650 61366 -78640
rect 61246 -78660 61276 -78650
rect 61246 -78860 61256 -78660
rect 61356 -78860 61366 -78650
rect 61246 -78870 61366 -78860
rect 60466 -78910 60626 -78900
rect 60286 -78970 60406 -78910
rect 60466 -78970 60476 -78910
rect 60536 -78970 60626 -78910
rect 59236 -79250 59266 -79160
rect 59366 -79250 59376 -79160
rect 59236 -79300 59376 -79250
rect 59506 -79110 59606 -79100
rect 59506 -79180 59516 -79110
rect 59596 -79180 59606 -79110
rect 59506 -79190 59606 -79180
rect 59236 -79320 59386 -79300
rect 59236 -79380 59316 -79320
rect 59376 -79380 59386 -79320
rect 58396 -79950 58896 -79450
rect 59236 -79630 59386 -79380
rect 59006 -79700 59086 -79680
rect 59236 -79690 59256 -79630
rect 59366 -79690 59386 -79630
rect 59236 -79700 59386 -79690
rect 59506 -79580 59596 -79190
rect 59986 -79320 60116 -79310
rect 59986 -79380 59996 -79320
rect 60106 -79380 60116 -79320
rect 59506 -79590 59616 -79580
rect 59506 -79660 59546 -79590
rect 59606 -79660 59616 -79590
rect 59006 -79760 59016 -79700
rect 59076 -79760 59086 -79700
rect 59006 -79950 59086 -79760
rect 59506 -79710 59616 -79660
rect 59506 -79770 59546 -79710
rect 59606 -79770 59616 -79710
rect 59796 -79610 59926 -79600
rect 59796 -79720 59806 -79610
rect 59916 -79720 59926 -79610
rect 59796 -79730 59926 -79720
rect 59006 -80040 59126 -79950
rect 59006 -80110 59016 -80040
rect 59076 -80110 59126 -80040
rect 59006 -80190 59126 -80110
rect 59506 -80040 59616 -79770
rect 59506 -80110 59546 -80040
rect 59606 -80110 59616 -80040
rect 59506 -80120 59616 -80110
rect 59986 -80190 60116 -79380
rect 60286 -79870 60376 -78970
rect 60466 -78980 60626 -78970
rect 61486 -78970 61726 -78940
rect 61486 -79020 61496 -78970
rect 61326 -79030 61496 -79020
rect 61326 -79150 61336 -79030
rect 61196 -79160 61336 -79150
rect 61456 -79140 61496 -79030
rect 61696 -79140 61726 -78970
rect 61456 -79160 61726 -79140
rect 61196 -79170 61726 -79160
rect 61196 -79340 61426 -79170
rect 60436 -79630 60536 -79610
rect 60436 -79750 60446 -79630
rect 60526 -79750 60536 -79630
rect 60436 -79760 60536 -79750
rect 60256 -80000 60416 -79870
rect 60256 -80130 60266 -80000
rect 60406 -80130 60416 -80000
rect 60256 -80150 60416 -80130
rect 58956 -80200 59156 -80190
rect 58956 -80380 58966 -80200
rect 59146 -80380 59156 -80200
rect 59986 -80300 59996 -80190
rect 60106 -80300 60116 -80190
rect 58956 -80390 59156 -80380
rect 59600 -80400 69400 -80300
rect 59600 -80800 59700 -80400
rect 60400 -80800 69000 -80400
rect 69300 -80800 69400 -80400
rect 59600 -80900 69400 -80800
rect 58946 -82470 59146 -82450
rect 58946 -82630 58966 -82470
rect 59126 -82630 59146 -82470
rect 58946 -82650 59146 -82630
rect 59316 -82510 59426 -82450
rect 59316 -82650 59336 -82510
rect 59416 -82650 59426 -82510
rect 58956 -82730 59136 -82650
rect 58956 -82840 58996 -82730
rect 59106 -82840 59136 -82730
rect 58396 -82930 58896 -82840
rect 58956 -82900 59136 -82840
rect 59316 -82880 59426 -82650
rect 59946 -82520 60386 -82400
rect 59946 -82640 60046 -82520
rect 60126 -82640 60386 -82520
rect 59946 -82690 60386 -82640
rect 58396 -83290 58486 -82930
rect 58816 -83290 58896 -82930
rect 58996 -83200 59086 -82900
rect 58996 -83260 59006 -83200
rect 59066 -83260 59086 -83200
rect 58996 -83270 59086 -83260
rect 59266 -82930 59426 -82880
rect 59506 -82740 59796 -82700
rect 59506 -82840 59516 -82740
rect 59616 -82840 59796 -82740
rect 59506 -82900 59796 -82840
rect 59266 -83130 59366 -82930
rect 59266 -83190 59286 -83130
rect 59346 -83190 59366 -83130
rect 58396 -83400 58896 -83290
rect 59066 -83440 59176 -83430
rect 59066 -83510 59076 -83440
rect 59166 -83510 59176 -83440
rect 56470 -84038 56555 -84028
rect 56470 -84128 56480 -84038
rect 56550 -84128 56555 -84038
rect 56470 -84138 56555 -84128
rect 56470 -84518 56550 -84138
rect 57760 -84140 57800 -84020
rect 58240 -84140 58280 -84020
rect 58516 -84060 58796 -83990
rect 57790 -84145 58250 -84140
rect 58516 -84260 58556 -84060
rect 58756 -84260 58796 -84060
rect 59066 -84010 59176 -83510
rect 59266 -83620 59366 -83190
rect 59536 -83090 59616 -82900
rect 59536 -83150 59546 -83090
rect 59606 -83150 59616 -83090
rect 59536 -83210 59616 -83150
rect 59536 -83270 59546 -83210
rect 59606 -83270 59616 -83210
rect 59536 -83280 59616 -83270
rect 59266 -83630 59376 -83620
rect 59266 -83720 59286 -83630
rect 59366 -83720 59376 -83630
rect 59736 -83650 59796 -82900
rect 59856 -83140 59976 -83130
rect 59856 -83230 59866 -83140
rect 59966 -83230 59976 -83140
rect 59856 -83240 59976 -83230
rect 60036 -83320 60136 -82690
rect 61026 -82720 61136 -82710
rect 61026 -82850 61056 -82720
rect 61126 -82850 61136 -82720
rect 60436 -83120 60536 -83110
rect 60436 -83220 60446 -83120
rect 60526 -83220 60536 -83120
rect 60436 -83230 60536 -83220
rect 60036 -83400 60046 -83320
rect 60126 -83400 60136 -83320
rect 60036 -83410 60136 -83400
rect 60546 -83410 60636 -83400
rect 60386 -83490 60556 -83410
rect 60626 -83490 60636 -83410
rect 59966 -83500 60326 -83490
rect 59966 -83570 59976 -83500
rect 60316 -83570 60326 -83500
rect 60546 -83510 60636 -83490
rect 59966 -83580 60326 -83570
rect 59566 -83670 59796 -83650
rect 59566 -83680 59576 -83670
rect 59266 -83730 59376 -83720
rect 59516 -83730 59576 -83680
rect 59636 -83730 59796 -83670
rect 59266 -83840 59366 -83730
rect 59266 -83930 59286 -83840
rect 59356 -83930 59366 -83840
rect 59266 -83960 59366 -83930
rect 59516 -83740 59796 -83730
rect 59066 -84080 59076 -84010
rect 59166 -84080 59176 -84010
rect 59066 -84090 59176 -84080
rect 59306 -84030 59386 -84020
rect 59306 -84090 59316 -84030
rect 59376 -84090 59386 -84030
rect 59516 -84070 59596 -83740
rect 60286 -83750 60476 -83740
rect 59906 -83780 60016 -83770
rect 59906 -83960 59916 -83780
rect 60006 -83960 60016 -83780
rect 59906 -83970 60016 -83960
rect 60286 -83890 60306 -83750
rect 60456 -83890 60476 -83750
rect 60286 -83900 60476 -83890
rect 58516 -84340 58796 -84260
rect 59066 -84170 59176 -84160
rect 59066 -84240 59076 -84170
rect 59166 -84240 59176 -84170
rect 57093 -84474 57373 -84464
rect 56470 -84528 56555 -84518
rect 56470 -84578 56480 -84528
rect 56475 -84588 56480 -84578
rect 56550 -84588 56555 -84528
rect 56475 -84598 56555 -84588
rect 57093 -84614 57098 -84474
rect 57368 -84614 57373 -84474
rect 57093 -84624 57373 -84614
rect 55870 -85078 55980 -84638
rect 59066 -84740 59176 -84240
rect 59306 -84290 59386 -84090
rect 60076 -84080 60196 -84040
rect 60076 -84240 60096 -84080
rect 60176 -84240 60196 -84080
rect 60076 -84280 60196 -84240
rect 59066 -84800 59076 -84740
rect 59166 -84800 59176 -84740
rect 59066 -84810 59176 -84800
rect 59236 -84320 59386 -84290
rect 59236 -84410 59266 -84320
rect 59366 -84410 59386 -84320
rect 59236 -84430 59386 -84410
rect 59906 -84290 60016 -84280
rect 59236 -84560 59376 -84430
rect 59906 -84480 59916 -84290
rect 60006 -84480 60016 -84290
rect 59906 -84490 60016 -84480
rect 60286 -84310 60376 -83900
rect 60556 -84300 60626 -83510
rect 61026 -83820 61136 -82850
rect 61196 -83520 61356 -83510
rect 61196 -83700 61206 -83520
rect 61346 -83700 61356 -83520
rect 61196 -83710 61356 -83700
rect 61026 -83930 61036 -83820
rect 61126 -83930 61136 -83820
rect 61026 -83940 61136 -83930
rect 61246 -84050 61366 -84040
rect 61246 -84060 61276 -84050
rect 61246 -84260 61256 -84060
rect 61356 -84260 61366 -84050
rect 61246 -84270 61366 -84260
rect 60466 -84310 60626 -84300
rect 60286 -84370 60406 -84310
rect 60466 -84370 60476 -84310
rect 60536 -84370 60626 -84310
rect 59236 -84650 59266 -84560
rect 59366 -84650 59376 -84560
rect 59236 -84700 59376 -84650
rect 59506 -84510 59606 -84500
rect 59506 -84580 59516 -84510
rect 59596 -84580 59606 -84510
rect 59506 -84590 59606 -84580
rect 59236 -84720 59386 -84700
rect 59236 -84780 59316 -84720
rect 59376 -84780 59386 -84720
rect 55870 -85118 55880 -85078
rect 55875 -85158 55880 -85118
rect 55970 -85118 55980 -85078
rect 56060 -85068 56220 -85058
rect 55970 -85158 55975 -85118
rect 55875 -85168 55975 -85158
rect 55590 -85278 55620 -85188
rect 55710 -85278 55720 -85188
rect 56060 -85238 56220 -85228
rect 56060 -85248 56200 -85238
rect 55590 -85288 55720 -85278
rect 56015 -85258 56200 -85248
rect 56015 -85408 56020 -85258
rect 56080 -85408 56200 -85258
rect 56644 -85268 57008 -85263
rect 55215 -85418 55325 -85408
rect 56015 -85418 56085 -85408
rect 55215 -85518 55220 -85418
rect 55320 -85518 55325 -85418
rect 56644 -85486 56654 -85268
rect 56998 -85486 57008 -85268
rect 58396 -85350 58896 -84850
rect 59236 -85030 59386 -84780
rect 59006 -85100 59086 -85080
rect 59236 -85090 59256 -85030
rect 59366 -85090 59386 -85030
rect 59236 -85100 59386 -85090
rect 59506 -84980 59596 -84590
rect 59986 -84720 60116 -84710
rect 59986 -84780 59996 -84720
rect 60106 -84780 60116 -84720
rect 59506 -84990 59616 -84980
rect 59506 -85060 59546 -84990
rect 59606 -85060 59616 -84990
rect 59006 -85160 59016 -85100
rect 59076 -85160 59086 -85100
rect 59006 -85350 59086 -85160
rect 59506 -85110 59616 -85060
rect 59506 -85170 59546 -85110
rect 59606 -85170 59616 -85110
rect 59796 -85010 59926 -85000
rect 59796 -85120 59806 -85010
rect 59916 -85120 59926 -85010
rect 59796 -85130 59926 -85120
rect 56644 -85491 57008 -85486
rect 59006 -85440 59126 -85350
rect 55215 -85528 55325 -85518
rect 59006 -85510 59016 -85440
rect 59076 -85510 59126 -85440
rect 59006 -85590 59126 -85510
rect 59506 -85440 59616 -85170
rect 59506 -85510 59546 -85440
rect 59606 -85510 59616 -85440
rect 59506 -85520 59616 -85510
rect 59986 -85590 60116 -84780
rect 60286 -85270 60376 -84370
rect 60466 -84380 60626 -84370
rect 61486 -84370 61726 -84340
rect 61486 -84420 61496 -84370
rect 61326 -84430 61496 -84420
rect 61326 -84550 61336 -84430
rect 61196 -84560 61336 -84550
rect 61456 -84540 61496 -84430
rect 61696 -84540 61726 -84370
rect 61456 -84560 61726 -84540
rect 61196 -84570 61726 -84560
rect 61196 -84740 61426 -84570
rect 60436 -85030 60536 -85010
rect 60436 -85150 60446 -85030
rect 60526 -85150 60536 -85030
rect 60436 -85160 60536 -85150
rect 60256 -85400 60416 -85270
rect 60256 -85530 60266 -85400
rect 60406 -85530 60416 -85400
rect 60256 -85550 60416 -85530
rect 58956 -85600 59156 -85590
rect 55315 -85728 55475 -85718
rect 55315 -85868 55320 -85728
rect 55470 -85868 55475 -85728
rect 58956 -85780 58966 -85600
rect 59146 -85780 59156 -85600
rect 59986 -85700 59996 -85590
rect 60106 -85700 60116 -85590
rect 58956 -85790 59156 -85780
rect 55315 -85878 55475 -85868
rect 59600 -85800 70400 -85700
rect 37100 -86200 37800 -86100
rect 59600 -86200 59700 -85800
rect 60400 -86200 70000 -85800
rect 70300 -86200 70400 -85800
rect 37100 -86700 37200 -86200
rect 37700 -86300 56200 -86200
rect 59600 -86300 70400 -86200
rect 37700 -86600 55500 -86300
rect 56100 -86600 56200 -86300
rect 37700 -86700 56200 -86600
rect 37100 -86800 37800 -86700
<< via3 >>
rect 38000 1400 41400 2800
rect 43000 1000 46400 2400
rect 37900 -3600 41500 -400
rect 43000 -1400 46400 0
rect 56506 -1830 57016 -1580
rect 53050 -3908 53250 -2158
rect 55020 -3128 55120 -3048
rect 56060 -2108 56220 -1948
rect 57098 -2704 57368 -2564
rect 58486 -2290 58816 -1930
rect 57098 -3614 57368 -3474
rect 56060 -4228 56220 -4068
rect 56654 -4486 56998 -4268
rect 55320 -4868 55470 -4728
rect 21000 -7400 22000 -6600
rect 56506 -7230 57016 -6980
rect 53050 -9308 53250 -7558
rect 55020 -8528 55120 -8448
rect 56060 -7508 56220 -7348
rect 57098 -8104 57368 -7964
rect 58556 -3260 58756 -3060
rect 59866 -2230 59966 -2140
rect 60446 -2220 60526 -2120
rect 59976 -2560 60316 -2500
rect 59976 -2570 60316 -2560
rect 59916 -2960 60006 -2780
rect 60096 -3240 60176 -3080
rect 59916 -3480 60006 -3290
rect 61206 -2700 61346 -2520
rect 61256 -3260 61276 -3060
rect 61276 -3260 61326 -3060
rect 59806 -4120 59916 -4010
rect 61496 -3540 61696 -3370
rect 60446 -4150 60526 -4030
rect 58486 -7690 58816 -7330
rect 57098 -9014 57368 -8874
rect 56060 -9628 56220 -9468
rect 56654 -9886 56998 -9668
rect 55320 -10268 55470 -10128
rect 27200 -13000 34400 -10600
rect 56506 -12630 57016 -12380
rect 53050 -14708 53250 -12958
rect 55020 -13928 55120 -13848
rect 56060 -12908 56220 -12748
rect 57098 -13504 57368 -13364
rect 58556 -8660 58756 -8460
rect 59866 -7630 59966 -7540
rect 60446 -7620 60526 -7520
rect 59976 -7960 60316 -7900
rect 59976 -7970 60316 -7960
rect 59916 -8360 60006 -8180
rect 60096 -8640 60176 -8480
rect 59916 -8880 60006 -8690
rect 61206 -8100 61346 -7920
rect 61256 -8660 61276 -8460
rect 61276 -8660 61326 -8460
rect 59806 -9520 59916 -9410
rect 61496 -8940 61696 -8770
rect 60446 -9550 60526 -9430
rect 58486 -13090 58816 -12730
rect 57098 -14414 57368 -14274
rect 56060 -15028 56220 -14868
rect 56654 -15286 56998 -15068
rect 55320 -15668 55470 -15528
rect 56506 -18030 57016 -17780
rect 53050 -20108 53250 -18358
rect 55020 -19328 55120 -19248
rect 56060 -18308 56220 -18148
rect 57098 -18904 57368 -18764
rect 58556 -14060 58756 -13860
rect 59866 -13030 59966 -12940
rect 60446 -13020 60526 -12920
rect 59976 -13360 60316 -13300
rect 59976 -13370 60316 -13360
rect 59916 -13760 60006 -13580
rect 60096 -14040 60176 -13880
rect 59916 -14280 60006 -14090
rect 61206 -13500 61346 -13320
rect 61256 -14060 61276 -13860
rect 61276 -14060 61326 -13860
rect 59806 -14920 59916 -14810
rect 61496 -14340 61696 -14170
rect 60446 -14950 60526 -14830
rect 58486 -18490 58816 -18130
rect 57098 -19814 57368 -19674
rect 56060 -20428 56220 -20268
rect 56654 -20686 56998 -20468
rect 55320 -21068 55470 -20928
rect 56506 -23430 57016 -23180
rect 53050 -25508 53250 -23758
rect 55020 -24728 55120 -24648
rect 56060 -23708 56220 -23548
rect 57098 -24304 57368 -24164
rect 58556 -19460 58756 -19260
rect 59866 -18430 59966 -18340
rect 60446 -18420 60526 -18320
rect 59976 -18760 60316 -18700
rect 59976 -18770 60316 -18760
rect 59916 -19160 60006 -18980
rect 60096 -19440 60176 -19280
rect 59916 -19680 60006 -19490
rect 61206 -18900 61346 -18720
rect 61256 -19460 61276 -19260
rect 61276 -19460 61326 -19260
rect 59806 -20320 59916 -20210
rect 61496 -19740 61696 -19570
rect 60446 -20350 60526 -20230
rect 58486 -23890 58816 -23530
rect 57098 -25214 57368 -25074
rect 56060 -25828 56220 -25668
rect 56654 -26086 56998 -25868
rect 55320 -26468 55470 -26328
rect 56506 -28830 57016 -28580
rect 53050 -30908 53250 -29158
rect 55020 -30128 55120 -30048
rect 56060 -29108 56220 -28948
rect 57098 -29704 57368 -29564
rect 58556 -24860 58756 -24660
rect 59866 -23830 59966 -23740
rect 60446 -23820 60526 -23720
rect 59976 -24160 60316 -24100
rect 59976 -24170 60316 -24160
rect 59916 -24560 60006 -24380
rect 60096 -24840 60176 -24680
rect 59916 -25080 60006 -24890
rect 61206 -24300 61346 -24120
rect 61256 -24860 61276 -24660
rect 61276 -24860 61326 -24660
rect 59806 -25720 59916 -25610
rect 61496 -25140 61696 -24970
rect 60446 -25750 60526 -25630
rect 58486 -29290 58816 -28930
rect 57098 -30614 57368 -30474
rect 56060 -31228 56220 -31068
rect 56654 -31486 56998 -31268
rect 55320 -31868 55470 -31728
rect 56506 -34230 57016 -33980
rect 53050 -36308 53250 -34558
rect 55020 -35528 55120 -35448
rect 56060 -34508 56220 -34348
rect 57098 -35104 57368 -34964
rect 58556 -30260 58756 -30060
rect 59866 -29230 59966 -29140
rect 60446 -29220 60526 -29120
rect 59976 -29560 60316 -29500
rect 59976 -29570 60316 -29560
rect 59916 -29960 60006 -29780
rect 60096 -30240 60176 -30080
rect 59916 -30480 60006 -30290
rect 61206 -29700 61346 -29520
rect 61256 -30260 61276 -30060
rect 61276 -30260 61326 -30060
rect 59806 -31120 59916 -31010
rect 61496 -30540 61696 -30370
rect 60446 -31150 60526 -31030
rect 58486 -34690 58816 -34330
rect 57098 -36014 57368 -35874
rect 56060 -36628 56220 -36468
rect 56654 -36886 56998 -36668
rect 55320 -37268 55470 -37128
rect 15000 -49000 24000 -38000
rect 56506 -39630 57016 -39380
rect 53050 -41708 53250 -39958
rect 55020 -40928 55120 -40848
rect 56060 -39908 56220 -39748
rect 57098 -40504 57368 -40364
rect 58556 -35660 58756 -35460
rect 59866 -34630 59966 -34540
rect 60446 -34620 60526 -34520
rect 59976 -34960 60316 -34900
rect 59976 -34970 60316 -34960
rect 59916 -35360 60006 -35180
rect 60096 -35640 60176 -35480
rect 59916 -35880 60006 -35690
rect 61206 -35100 61346 -34920
rect 61256 -35660 61276 -35460
rect 61276 -35660 61326 -35460
rect 72000 -35500 74000 -34100
rect 59806 -36520 59916 -36410
rect 61496 -35940 61696 -35770
rect 60446 -36550 60526 -36430
rect 76910 -38410 77070 -38400
rect 76910 -38530 76920 -38410
rect 76920 -38530 77060 -38410
rect 77060 -38530 77070 -38410
rect 76910 -38540 77070 -38530
rect 84960 -38480 85400 -38050
rect 77170 -39040 77430 -38790
rect 88150 -38820 88590 -38390
rect 58486 -40090 58816 -39730
rect 57098 -41414 57368 -41274
rect 56060 -42028 56220 -41868
rect 56654 -42286 56998 -42068
rect 55320 -42668 55470 -42528
rect 56506 -45030 57016 -44780
rect 53050 -47108 53250 -45358
rect 55020 -46328 55120 -46248
rect 56060 -45308 56220 -45148
rect 57098 -45904 57368 -45764
rect 58556 -41060 58756 -40860
rect 59866 -40030 59966 -39940
rect 60446 -40020 60526 -39920
rect 59976 -40360 60316 -40300
rect 59976 -40370 60316 -40360
rect 59916 -40760 60006 -40580
rect 60096 -41040 60176 -40880
rect 59916 -41280 60006 -41090
rect 76920 -39720 77060 -39570
rect 61206 -40500 61346 -40320
rect 79410 -40390 79680 -40150
rect 83150 -40180 83510 -39830
rect 81140 -40510 81570 -40250
rect 87830 -40590 88190 -40240
rect 61256 -41060 61276 -40860
rect 61276 -41060 61326 -40860
rect 76920 -40960 77060 -40820
rect 59806 -41920 59916 -41810
rect 61496 -41340 61696 -41170
rect 79410 -41620 79680 -41380
rect 60446 -41950 60526 -41830
rect 76920 -42210 77060 -42060
rect 76920 -42220 77060 -42210
rect 79410 -42880 79680 -42640
rect 76920 -43450 77060 -43310
rect 82820 -43310 91410 -42740
rect 79410 -44100 79680 -43860
rect 76920 -44610 77060 -44520
rect 58486 -45490 58816 -45130
rect 57098 -46814 57368 -46674
rect 56060 -47428 56220 -47268
rect 56654 -47686 56998 -47468
rect 55320 -48068 55470 -47928
rect 56506 -50430 57016 -50180
rect 53050 -52508 53250 -50758
rect 55020 -51728 55120 -51648
rect 56060 -50708 56220 -50548
rect 57098 -51304 57368 -51164
rect 58556 -46460 58756 -46260
rect 59866 -45430 59966 -45340
rect 82820 -45010 91410 -44440
rect 60446 -45420 60526 -45320
rect 59976 -45760 60316 -45700
rect 59976 -45770 60316 -45760
rect 59916 -46160 60006 -45980
rect 60096 -46440 60176 -46280
rect 59916 -46680 60006 -46490
rect 79410 -45360 79680 -45120
rect 61206 -45900 61346 -45720
rect 76920 -45740 77060 -45640
rect 61256 -46460 61276 -46260
rect 61276 -46460 61326 -46260
rect 59806 -47320 59916 -47210
rect 61496 -46740 61696 -46570
rect 76910 -46450 77070 -46440
rect 76910 -46570 76920 -46450
rect 76920 -46570 77060 -46450
rect 77060 -46570 77070 -46450
rect 76910 -46580 77070 -46570
rect 77170 -47080 77430 -46830
rect 60446 -47350 60526 -47230
rect 76920 -47760 77060 -47610
rect 82824 -47448 91414 -46878
rect 79410 -48430 79680 -48190
rect 76920 -49000 77060 -48860
rect 82824 -49148 91414 -48578
rect 79410 -49660 79680 -49420
rect 58486 -50890 58816 -50530
rect 57098 -52214 57368 -52074
rect 56060 -52828 56220 -52668
rect 56654 -53086 56998 -52868
rect 55320 -53468 55470 -53328
rect 56506 -55830 57016 -55580
rect 53050 -57908 53250 -56158
rect 55020 -57128 55120 -57048
rect 56060 -56108 56220 -55948
rect 57098 -56704 57368 -56564
rect 58556 -51860 58756 -51660
rect 59866 -50830 59966 -50740
rect 76920 -50250 77060 -50100
rect 76920 -50260 77060 -50250
rect 60446 -50820 60526 -50720
rect 59976 -51160 60316 -51100
rect 59976 -51170 60316 -51160
rect 59916 -51560 60006 -51380
rect 60096 -51840 60176 -51680
rect 59916 -52080 60006 -51890
rect 79410 -50920 79680 -50680
rect 61206 -51300 61346 -51120
rect 82820 -51100 91410 -50530
rect 76920 -51490 77060 -51350
rect 61256 -51860 61276 -51660
rect 61276 -51860 61326 -51660
rect 59806 -52720 59916 -52610
rect 61496 -52140 61696 -51970
rect 79410 -52140 79680 -51900
rect 60446 -52750 60526 -52630
rect 76920 -52650 77060 -52560
rect 82820 -52800 91410 -52230
rect 79410 -53400 79680 -53160
rect 76920 -53780 77060 -53680
rect 58486 -56290 58816 -55930
rect 57098 -57614 57368 -57474
rect 56060 -58228 56220 -58068
rect 56654 -58486 56998 -58268
rect 55320 -58868 55470 -58728
rect 56506 -61230 57016 -60980
rect 53050 -63308 53250 -61558
rect 55020 -62528 55120 -62448
rect 56060 -61508 56220 -61348
rect 57098 -62104 57368 -61964
rect 58556 -57260 58756 -57060
rect 59866 -56230 59966 -56140
rect 60446 -56220 60526 -56120
rect 59976 -56560 60316 -56500
rect 59976 -56570 60316 -56560
rect 59916 -56960 60006 -56780
rect 60096 -57240 60176 -57080
rect 59916 -57480 60006 -57290
rect 61206 -56700 61346 -56520
rect 61256 -57260 61276 -57060
rect 61276 -57260 61326 -57060
rect 59806 -58120 59916 -58010
rect 61496 -57540 61696 -57370
rect 60446 -58150 60526 -58030
rect 58486 -61690 58816 -61330
rect 57098 -63014 57368 -62874
rect 56060 -63628 56220 -63468
rect 56654 -63886 56998 -63668
rect 55320 -64268 55470 -64128
rect 56506 -66630 57016 -66380
rect 53050 -68708 53250 -66958
rect 55020 -67928 55120 -67848
rect 56060 -66908 56220 -66748
rect 57098 -67504 57368 -67364
rect 58556 -62660 58756 -62460
rect 59866 -61630 59966 -61540
rect 60446 -61620 60526 -61520
rect 59976 -61960 60316 -61900
rect 59976 -61970 60316 -61960
rect 59916 -62360 60006 -62180
rect 60096 -62640 60176 -62480
rect 59916 -62880 60006 -62690
rect 61206 -62100 61346 -61920
rect 61256 -62660 61276 -62460
rect 61276 -62660 61326 -62460
rect 59806 -63520 59916 -63410
rect 61496 -62940 61696 -62770
rect 60446 -63550 60526 -63430
rect 58486 -67090 58816 -66730
rect 57098 -68414 57368 -68274
rect 56060 -69028 56220 -68868
rect 56654 -69286 56998 -69068
rect 55320 -69668 55470 -69528
rect 56506 -72030 57016 -71780
rect 53050 -74108 53250 -72358
rect 55020 -73328 55120 -73248
rect 56060 -72308 56220 -72148
rect 57098 -72904 57368 -72764
rect 58556 -68060 58756 -67860
rect 59866 -67030 59966 -66940
rect 60446 -67020 60526 -66920
rect 59976 -67360 60316 -67300
rect 59976 -67370 60316 -67360
rect 59916 -67760 60006 -67580
rect 60096 -68040 60176 -67880
rect 59916 -68280 60006 -68090
rect 61206 -67500 61346 -67320
rect 61256 -68060 61276 -67860
rect 61276 -68060 61326 -67860
rect 59806 -68920 59916 -68810
rect 61496 -68340 61696 -68170
rect 60446 -68950 60526 -68830
rect 58486 -72490 58816 -72130
rect 57098 -73814 57368 -73674
rect 56060 -74428 56220 -74268
rect 56654 -74686 56998 -74468
rect 55320 -75068 55470 -74928
rect 56506 -77430 57016 -77180
rect 53050 -79508 53250 -77758
rect 55020 -78728 55120 -78648
rect 56060 -77708 56220 -77548
rect 57098 -78304 57368 -78164
rect 58556 -73460 58756 -73260
rect 59866 -72430 59966 -72340
rect 60446 -72420 60526 -72320
rect 59976 -72760 60316 -72700
rect 59976 -72770 60316 -72760
rect 59916 -73160 60006 -72980
rect 60096 -73440 60176 -73280
rect 59916 -73680 60006 -73490
rect 61206 -72900 61346 -72720
rect 61256 -73460 61276 -73260
rect 61276 -73460 61326 -73260
rect 59806 -74320 59916 -74210
rect 61496 -73740 61696 -73570
rect 60446 -74350 60526 -74230
rect 58486 -77890 58816 -77530
rect 57098 -79214 57368 -79074
rect 56060 -79828 56220 -79668
rect 56654 -80086 56998 -79868
rect 55320 -80468 55470 -80328
rect 56506 -82830 57016 -82580
rect 53050 -84908 53250 -83158
rect 55020 -84128 55120 -84048
rect 56060 -83108 56220 -82948
rect 57098 -83704 57368 -83564
rect 58556 -78860 58756 -78660
rect 59866 -77830 59966 -77740
rect 60446 -77820 60526 -77720
rect 59976 -78160 60316 -78100
rect 59976 -78170 60316 -78160
rect 59916 -78560 60006 -78380
rect 60096 -78840 60176 -78680
rect 59916 -79080 60006 -78890
rect 61206 -78300 61346 -78120
rect 61256 -78860 61276 -78660
rect 61276 -78860 61326 -78660
rect 59806 -79720 59916 -79610
rect 61496 -79140 61696 -78970
rect 60446 -79750 60526 -79630
rect 58486 -83290 58816 -82930
rect 58556 -84260 58756 -84060
rect 59866 -83230 59966 -83140
rect 60446 -83220 60526 -83120
rect 59976 -83560 60316 -83500
rect 59976 -83570 60316 -83560
rect 59916 -83960 60006 -83780
rect 57098 -84614 57368 -84474
rect 60096 -84240 60176 -84080
rect 59916 -84480 60006 -84290
rect 61206 -83700 61346 -83520
rect 61256 -84260 61276 -84060
rect 61276 -84260 61326 -84060
rect 56060 -85228 56220 -85068
rect 56654 -85486 56998 -85268
rect 59806 -85120 59916 -85010
rect 61496 -84540 61696 -84370
rect 60446 -85150 60526 -85030
rect 55320 -85868 55470 -85728
<< metal4 >>
rect 37800 3000 69400 5000
rect 37800 2800 41600 3000
rect 37800 1400 38000 2800
rect 41400 1400 41600 2800
rect 37800 1200 41600 1400
rect 42800 2400 46600 2600
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 800 46600 1000
rect 42800 0 46600 200
rect 37800 -400 41600 -300
rect 37800 -3600 37900 -400
rect 41500 -2000 41600 -400
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 42800 -1600 46600 -1400
rect 56505 -1580 57017 -1579
rect 56505 -1830 56506 -1580
rect 57016 -1830 57017 -1580
rect 56505 -1831 57017 -1830
rect 58396 -1930 58896 -1840
rect 56059 -1948 56221 -1947
rect 56059 -2000 56060 -1948
rect 41500 -2108 56060 -2000
rect 56220 -2108 56221 -1948
rect 41500 -2109 56221 -2108
rect 41500 -2158 56220 -2109
rect 41500 -3600 53050 -2158
rect 37800 -3908 53050 -3600
rect 53250 -2554 56220 -2158
rect 58396 -2290 58486 -1930
rect 58816 -2290 58896 -1930
rect 60436 -2120 60536 -2110
rect 58396 -2400 58896 -2290
rect 59826 -2140 59976 -2130
rect 59826 -2230 59866 -2140
rect 59966 -2230 59976 -2140
rect 59826 -2240 59976 -2230
rect 60436 -2220 60446 -2120
rect 60526 -2220 60536 -2120
rect 59826 -2470 59946 -2240
rect 60436 -2470 60536 -2220
rect 59666 -2500 60536 -2470
rect 53250 -2564 57378 -2554
rect 53250 -2704 57098 -2564
rect 57368 -2704 57378 -2564
rect 59666 -2570 59976 -2500
rect 60316 -2570 60536 -2500
rect 61820 -2510 69400 3000
rect 59666 -2590 60536 -2570
rect 61186 -2520 69400 -2510
rect 59666 -2640 59776 -2590
rect 53250 -2714 57378 -2704
rect 53250 -3048 56220 -2714
rect 53250 -3128 55020 -3048
rect 55120 -3128 56220 -3048
rect 53250 -3464 56220 -3128
rect 59656 -3040 59776 -2640
rect 61186 -2700 61206 -2520
rect 61346 -2700 69400 -2520
rect 61186 -2720 69400 -2700
rect 59906 -2780 60026 -2750
rect 59906 -2960 59916 -2780
rect 60006 -2960 60026 -2780
rect 59906 -3040 60026 -2960
rect 61186 -3040 61366 -2720
rect 59656 -3060 61366 -3040
rect 59656 -3080 61256 -3060
rect 59656 -3240 60096 -3080
rect 60176 -3240 61256 -3080
rect 59656 -3260 61256 -3240
rect 61326 -3260 61366 -3060
rect 59656 -3280 61366 -3260
rect 53250 -3474 57378 -3464
rect 53250 -3614 57098 -3474
rect 57368 -3614 57378 -3474
rect 53250 -3624 57378 -3614
rect 53250 -3908 56220 -3624
rect 59656 -3650 59776 -3280
rect 59906 -3290 60026 -3280
rect 59906 -3480 59916 -3290
rect 60006 -3480 60026 -3290
rect 61256 -3390 61366 -3280
rect 59906 -3490 60026 -3480
rect 61426 -3500 61446 -3260
rect 61686 -3370 61726 -3260
rect 61426 -3540 61496 -3500
rect 61696 -3540 61726 -3370
rect 61426 -3570 61726 -3540
rect 59656 -3770 60536 -3650
rect 37800 -4067 56220 -3908
rect 58396 -3930 58896 -3850
rect 37800 -4068 56221 -4067
rect 37800 -4228 56060 -4068
rect 56220 -4228 56221 -4068
rect 37800 -4229 56221 -4228
rect 37800 -4690 56200 -4229
rect 58396 -4290 58486 -3930
rect 58816 -4290 58896 -3930
rect 59796 -4010 59926 -3770
rect 59796 -4120 59806 -4010
rect 59916 -4120 59926 -4010
rect 59796 -4130 59926 -4120
rect 60436 -4030 60536 -3770
rect 60436 -4150 60446 -4030
rect 60526 -4150 60536 -4030
rect 60436 -4160 60536 -4150
rect 58396 -4350 58896 -4290
rect 61820 -4690 69400 -2720
rect 37800 -4728 69400 -4690
rect 37800 -4868 55320 -4728
rect 55470 -4868 69400 -4728
rect 37800 -4940 69400 -4868
rect 20800 -6600 22200 -6400
rect 20800 -7400 21000 -6600
rect 22000 -7400 22200 -6600
rect 20800 -7600 22200 -7400
rect 37800 -7347 56200 -4940
rect 56505 -6980 57017 -6979
rect 56505 -7230 56506 -6980
rect 57016 -7230 57017 -6980
rect 56505 -7231 57017 -7230
rect 58396 -7330 58896 -7240
rect 37800 -7348 56221 -7347
rect 37800 -7508 56060 -7348
rect 56220 -7508 56221 -7348
rect 37800 -7509 56221 -7508
rect 37800 -7558 56220 -7509
rect 37800 -9308 53050 -7558
rect 53250 -7954 56220 -7558
rect 58396 -7690 58486 -7330
rect 58816 -7690 58896 -7330
rect 60436 -7520 60536 -7510
rect 58396 -7800 58896 -7690
rect 59826 -7540 59976 -7530
rect 59826 -7630 59866 -7540
rect 59966 -7630 59976 -7540
rect 59826 -7640 59976 -7630
rect 60436 -7620 60446 -7520
rect 60526 -7620 60536 -7520
rect 59826 -7870 59946 -7640
rect 60436 -7870 60536 -7620
rect 59666 -7900 60536 -7870
rect 53250 -7964 57378 -7954
rect 53250 -8104 57098 -7964
rect 57368 -8104 57378 -7964
rect 59666 -7970 59976 -7900
rect 60316 -7970 60536 -7900
rect 61820 -7910 69400 -4940
rect 59666 -7990 60536 -7970
rect 61186 -7920 69400 -7910
rect 59666 -8040 59776 -7990
rect 53250 -8114 57378 -8104
rect 53250 -8448 56220 -8114
rect 53250 -8528 55020 -8448
rect 55120 -8528 56220 -8448
rect 53250 -8864 56220 -8528
rect 59656 -8440 59776 -8040
rect 61186 -8100 61206 -7920
rect 61346 -8100 69400 -7920
rect 61186 -8120 69400 -8100
rect 59906 -8180 60026 -8150
rect 59906 -8360 59916 -8180
rect 60006 -8360 60026 -8180
rect 59906 -8440 60026 -8360
rect 61186 -8440 61366 -8120
rect 59656 -8460 61366 -8440
rect 59656 -8480 61256 -8460
rect 59656 -8640 60096 -8480
rect 60176 -8640 61256 -8480
rect 59656 -8660 61256 -8640
rect 61326 -8660 61366 -8460
rect 59656 -8680 61366 -8660
rect 53250 -8874 57378 -8864
rect 53250 -9014 57098 -8874
rect 57368 -9014 57378 -8874
rect 53250 -9024 57378 -9014
rect 53250 -9308 56220 -9024
rect 59656 -9050 59776 -8680
rect 59906 -8690 60026 -8680
rect 59906 -8880 59916 -8690
rect 60006 -8880 60026 -8690
rect 61256 -8790 61366 -8680
rect 59906 -8890 60026 -8880
rect 61426 -8900 61446 -8660
rect 61686 -8770 61726 -8660
rect 61426 -8940 61496 -8900
rect 61696 -8940 61726 -8770
rect 61426 -8970 61726 -8940
rect 59656 -9170 60536 -9050
rect 37800 -9467 56220 -9308
rect 58396 -9330 58896 -9250
rect 37800 -9468 56221 -9467
rect 37800 -9628 56060 -9468
rect 56220 -9628 56221 -9468
rect 37800 -9629 56221 -9628
rect 37800 -10090 56200 -9629
rect 58396 -9690 58486 -9330
rect 58816 -9690 58896 -9330
rect 59796 -9410 59926 -9170
rect 59796 -9520 59806 -9410
rect 59916 -9520 59926 -9410
rect 59796 -9530 59926 -9520
rect 60436 -9430 60536 -9170
rect 60436 -9550 60446 -9430
rect 60526 -9550 60536 -9430
rect 60436 -9560 60536 -9550
rect 58396 -9750 58896 -9690
rect 61820 -10090 69400 -8120
rect 37800 -10128 69400 -10090
rect 37800 -10268 55320 -10128
rect 55470 -10268 69400 -10128
rect 37800 -10340 69400 -10268
rect 37800 -10400 56200 -10340
rect 27000 -10600 56200 -10400
rect 27000 -13000 27200 -10600
rect 34400 -12747 56200 -10600
rect 56505 -12380 57017 -12379
rect 56505 -12630 56506 -12380
rect 57016 -12630 57017 -12380
rect 56505 -12631 57017 -12630
rect 58396 -12730 58896 -12640
rect 34400 -12748 56221 -12747
rect 34400 -12908 56060 -12748
rect 56220 -12908 56221 -12748
rect 34400 -12909 56221 -12908
rect 34400 -12958 56220 -12909
rect 34400 -13000 53050 -12958
rect 27000 -13200 53050 -13000
rect 37800 -14708 53050 -13200
rect 53250 -13354 56220 -12958
rect 58396 -13090 58486 -12730
rect 58816 -13090 58896 -12730
rect 60436 -12920 60536 -12910
rect 58396 -13200 58896 -13090
rect 59826 -12940 59976 -12930
rect 59826 -13030 59866 -12940
rect 59966 -13030 59976 -12940
rect 59826 -13040 59976 -13030
rect 60436 -13020 60446 -12920
rect 60526 -13020 60536 -12920
rect 59826 -13270 59946 -13040
rect 60436 -13270 60536 -13020
rect 59666 -13300 60536 -13270
rect 53250 -13364 57378 -13354
rect 53250 -13504 57098 -13364
rect 57368 -13504 57378 -13364
rect 59666 -13370 59976 -13300
rect 60316 -13370 60536 -13300
rect 61820 -13310 69400 -10340
rect 59666 -13390 60536 -13370
rect 61186 -13320 69400 -13310
rect 59666 -13440 59776 -13390
rect 53250 -13514 57378 -13504
rect 53250 -13848 56220 -13514
rect 53250 -13928 55020 -13848
rect 55120 -13928 56220 -13848
rect 53250 -14264 56220 -13928
rect 59656 -13840 59776 -13440
rect 61186 -13500 61206 -13320
rect 61346 -13500 69400 -13320
rect 61186 -13520 69400 -13500
rect 59906 -13580 60026 -13550
rect 59906 -13760 59916 -13580
rect 60006 -13760 60026 -13580
rect 59906 -13840 60026 -13760
rect 61186 -13840 61366 -13520
rect 59656 -13860 61366 -13840
rect 59656 -13880 61256 -13860
rect 59656 -14040 60096 -13880
rect 60176 -14040 61256 -13880
rect 59656 -14060 61256 -14040
rect 61326 -14060 61366 -13860
rect 59656 -14080 61366 -14060
rect 53250 -14274 57378 -14264
rect 53250 -14414 57098 -14274
rect 57368 -14414 57378 -14274
rect 53250 -14424 57378 -14414
rect 53250 -14708 56220 -14424
rect 59656 -14450 59776 -14080
rect 59906 -14090 60026 -14080
rect 59906 -14280 59916 -14090
rect 60006 -14280 60026 -14090
rect 61256 -14190 61366 -14080
rect 59906 -14290 60026 -14280
rect 61426 -14300 61446 -14060
rect 61686 -14170 61726 -14060
rect 61426 -14340 61496 -14300
rect 61696 -14340 61726 -14170
rect 61426 -14370 61726 -14340
rect 59656 -14570 60536 -14450
rect 37800 -14867 56220 -14708
rect 58396 -14730 58896 -14650
rect 37800 -14868 56221 -14867
rect 37800 -15028 56060 -14868
rect 56220 -15028 56221 -14868
rect 37800 -15029 56221 -15028
rect 37800 -15490 56200 -15029
rect 58396 -15090 58486 -14730
rect 58816 -15090 58896 -14730
rect 59796 -14810 59926 -14570
rect 59796 -14920 59806 -14810
rect 59916 -14920 59926 -14810
rect 59796 -14930 59926 -14920
rect 60436 -14830 60536 -14570
rect 60436 -14950 60446 -14830
rect 60526 -14950 60536 -14830
rect 60436 -14960 60536 -14950
rect 58396 -15150 58896 -15090
rect 61820 -15490 69400 -13520
rect 37800 -15528 69400 -15490
rect 37800 -15668 55320 -15528
rect 55470 -15668 69400 -15528
rect 37800 -15740 69400 -15668
rect 37800 -18147 56200 -15740
rect 56505 -17780 57017 -17779
rect 56505 -18030 56506 -17780
rect 57016 -18030 57017 -17780
rect 56505 -18031 57017 -18030
rect 58396 -18130 58896 -18040
rect 37800 -18148 56221 -18147
rect 37800 -18308 56060 -18148
rect 56220 -18308 56221 -18148
rect 37800 -18309 56221 -18308
rect 37800 -18358 56220 -18309
rect 37800 -20108 53050 -18358
rect 53250 -18754 56220 -18358
rect 58396 -18490 58486 -18130
rect 58816 -18490 58896 -18130
rect 60436 -18320 60536 -18310
rect 58396 -18600 58896 -18490
rect 59826 -18340 59976 -18330
rect 59826 -18430 59866 -18340
rect 59966 -18430 59976 -18340
rect 59826 -18440 59976 -18430
rect 60436 -18420 60446 -18320
rect 60526 -18420 60536 -18320
rect 59826 -18670 59946 -18440
rect 60436 -18670 60536 -18420
rect 59666 -18700 60536 -18670
rect 53250 -18764 57378 -18754
rect 53250 -18904 57098 -18764
rect 57368 -18904 57378 -18764
rect 59666 -18770 59976 -18700
rect 60316 -18770 60536 -18700
rect 61820 -18710 69400 -15740
rect 59666 -18790 60536 -18770
rect 61186 -18720 69400 -18710
rect 59666 -18840 59776 -18790
rect 53250 -18914 57378 -18904
rect 53250 -19248 56220 -18914
rect 53250 -19328 55020 -19248
rect 55120 -19328 56220 -19248
rect 53250 -19664 56220 -19328
rect 59656 -19240 59776 -18840
rect 61186 -18900 61206 -18720
rect 61346 -18900 69400 -18720
rect 61186 -18920 69400 -18900
rect 59906 -18980 60026 -18950
rect 59906 -19160 59916 -18980
rect 60006 -19160 60026 -18980
rect 59906 -19240 60026 -19160
rect 61186 -19240 61366 -18920
rect 59656 -19260 61366 -19240
rect 59656 -19280 61256 -19260
rect 59656 -19440 60096 -19280
rect 60176 -19440 61256 -19280
rect 59656 -19460 61256 -19440
rect 61326 -19460 61366 -19260
rect 59656 -19480 61366 -19460
rect 53250 -19674 57378 -19664
rect 53250 -19814 57098 -19674
rect 57368 -19814 57378 -19674
rect 53250 -19824 57378 -19814
rect 53250 -20108 56220 -19824
rect 59656 -19850 59776 -19480
rect 59906 -19490 60026 -19480
rect 59906 -19680 59916 -19490
rect 60006 -19680 60026 -19490
rect 61256 -19590 61366 -19480
rect 59906 -19690 60026 -19680
rect 61426 -19700 61446 -19460
rect 61686 -19570 61726 -19460
rect 61426 -19740 61496 -19700
rect 61696 -19740 61726 -19570
rect 61426 -19770 61726 -19740
rect 59656 -19970 60536 -19850
rect 37800 -20267 56220 -20108
rect 58396 -20130 58896 -20050
rect 37800 -20268 56221 -20267
rect 37800 -20428 56060 -20268
rect 56220 -20428 56221 -20268
rect 37800 -20429 56221 -20428
rect 37800 -20890 56200 -20429
rect 58396 -20490 58486 -20130
rect 58816 -20490 58896 -20130
rect 59796 -20210 59926 -19970
rect 59796 -20320 59806 -20210
rect 59916 -20320 59926 -20210
rect 59796 -20330 59926 -20320
rect 60436 -20230 60536 -19970
rect 60436 -20350 60446 -20230
rect 60526 -20350 60536 -20230
rect 60436 -20360 60536 -20350
rect 58396 -20550 58896 -20490
rect 61820 -20890 69400 -18920
rect 37800 -20928 69400 -20890
rect 37800 -21068 55320 -20928
rect 55470 -21068 69400 -20928
rect 37800 -21140 69400 -21068
rect 37800 -23547 56200 -21140
rect 56505 -23180 57017 -23179
rect 56505 -23430 56506 -23180
rect 57016 -23430 57017 -23180
rect 56505 -23431 57017 -23430
rect 58396 -23530 58896 -23440
rect 37800 -23548 56221 -23547
rect 37800 -23708 56060 -23548
rect 56220 -23708 56221 -23548
rect 37800 -23709 56221 -23708
rect 37800 -23758 56220 -23709
rect 37800 -25508 53050 -23758
rect 53250 -24154 56220 -23758
rect 58396 -23890 58486 -23530
rect 58816 -23890 58896 -23530
rect 60436 -23720 60536 -23710
rect 58396 -24000 58896 -23890
rect 59826 -23740 59976 -23730
rect 59826 -23830 59866 -23740
rect 59966 -23830 59976 -23740
rect 59826 -23840 59976 -23830
rect 60436 -23820 60446 -23720
rect 60526 -23820 60536 -23720
rect 59826 -24070 59946 -23840
rect 60436 -24070 60536 -23820
rect 59666 -24100 60536 -24070
rect 53250 -24164 57378 -24154
rect 53250 -24304 57098 -24164
rect 57368 -24304 57378 -24164
rect 59666 -24170 59976 -24100
rect 60316 -24170 60536 -24100
rect 61820 -24110 69400 -21140
rect 59666 -24190 60536 -24170
rect 61186 -24120 69400 -24110
rect 59666 -24240 59776 -24190
rect 53250 -24314 57378 -24304
rect 53250 -24648 56220 -24314
rect 53250 -24728 55020 -24648
rect 55120 -24728 56220 -24648
rect 53250 -25064 56220 -24728
rect 59656 -24640 59776 -24240
rect 61186 -24300 61206 -24120
rect 61346 -24300 69400 -24120
rect 61186 -24320 69400 -24300
rect 59906 -24380 60026 -24350
rect 59906 -24560 59916 -24380
rect 60006 -24560 60026 -24380
rect 59906 -24640 60026 -24560
rect 61186 -24640 61366 -24320
rect 59656 -24660 61366 -24640
rect 59656 -24680 61256 -24660
rect 59656 -24840 60096 -24680
rect 60176 -24840 61256 -24680
rect 59656 -24860 61256 -24840
rect 61326 -24860 61366 -24660
rect 59656 -24880 61366 -24860
rect 53250 -25074 57378 -25064
rect 53250 -25214 57098 -25074
rect 57368 -25214 57378 -25074
rect 53250 -25224 57378 -25214
rect 53250 -25508 56220 -25224
rect 59656 -25250 59776 -24880
rect 59906 -24890 60026 -24880
rect 59906 -25080 59916 -24890
rect 60006 -25080 60026 -24890
rect 61256 -24990 61366 -24880
rect 59906 -25090 60026 -25080
rect 61426 -25100 61446 -24860
rect 61686 -24970 61726 -24860
rect 61426 -25140 61496 -25100
rect 61696 -25140 61726 -24970
rect 61426 -25170 61726 -25140
rect 59656 -25370 60536 -25250
rect 37800 -25667 56220 -25508
rect 58396 -25530 58896 -25450
rect 37800 -25668 56221 -25667
rect 37800 -25828 56060 -25668
rect 56220 -25828 56221 -25668
rect 37800 -25829 56221 -25828
rect 37800 -26290 56200 -25829
rect 58396 -25890 58486 -25530
rect 58816 -25890 58896 -25530
rect 59796 -25610 59926 -25370
rect 59796 -25720 59806 -25610
rect 59916 -25720 59926 -25610
rect 59796 -25730 59926 -25720
rect 60436 -25630 60536 -25370
rect 60436 -25750 60446 -25630
rect 60526 -25750 60536 -25630
rect 60436 -25760 60536 -25750
rect 58396 -25950 58896 -25890
rect 61820 -26290 69400 -24320
rect 37800 -26328 69400 -26290
rect 37800 -26468 55320 -26328
rect 55470 -26468 69400 -26328
rect 37800 -26540 69400 -26468
rect 37800 -28947 56200 -26540
rect 56505 -28580 57017 -28579
rect 56505 -28830 56506 -28580
rect 57016 -28830 57017 -28580
rect 56505 -28831 57017 -28830
rect 58396 -28930 58896 -28840
rect 37800 -28948 56221 -28947
rect 37800 -29108 56060 -28948
rect 56220 -29108 56221 -28948
rect 37800 -29109 56221 -29108
rect 37800 -29158 56220 -29109
rect 37800 -30908 53050 -29158
rect 53250 -29554 56220 -29158
rect 58396 -29290 58486 -28930
rect 58816 -29290 58896 -28930
rect 60436 -29120 60536 -29110
rect 58396 -29400 58896 -29290
rect 59826 -29140 59976 -29130
rect 59826 -29230 59866 -29140
rect 59966 -29230 59976 -29140
rect 59826 -29240 59976 -29230
rect 60436 -29220 60446 -29120
rect 60526 -29220 60536 -29120
rect 59826 -29470 59946 -29240
rect 60436 -29470 60536 -29220
rect 59666 -29500 60536 -29470
rect 53250 -29564 57378 -29554
rect 53250 -29704 57098 -29564
rect 57368 -29704 57378 -29564
rect 59666 -29570 59976 -29500
rect 60316 -29570 60536 -29500
rect 61820 -29510 69400 -26540
rect 59666 -29590 60536 -29570
rect 61186 -29520 69400 -29510
rect 59666 -29640 59776 -29590
rect 53250 -29714 57378 -29704
rect 53250 -30048 56220 -29714
rect 53250 -30128 55020 -30048
rect 55120 -30128 56220 -30048
rect 53250 -30464 56220 -30128
rect 59656 -30040 59776 -29640
rect 61186 -29700 61206 -29520
rect 61346 -29700 69400 -29520
rect 61186 -29720 69400 -29700
rect 59906 -29780 60026 -29750
rect 59906 -29960 59916 -29780
rect 60006 -29960 60026 -29780
rect 59906 -30040 60026 -29960
rect 61186 -30040 61366 -29720
rect 59656 -30060 61366 -30040
rect 59656 -30080 61256 -30060
rect 59656 -30240 60096 -30080
rect 60176 -30240 61256 -30080
rect 59656 -30260 61256 -30240
rect 61326 -30260 61366 -30060
rect 59656 -30280 61366 -30260
rect 53250 -30474 57378 -30464
rect 53250 -30614 57098 -30474
rect 57368 -30614 57378 -30474
rect 53250 -30624 57378 -30614
rect 53250 -30908 56220 -30624
rect 59656 -30650 59776 -30280
rect 59906 -30290 60026 -30280
rect 59906 -30480 59916 -30290
rect 60006 -30480 60026 -30290
rect 61256 -30390 61366 -30280
rect 59906 -30490 60026 -30480
rect 61426 -30500 61446 -30260
rect 61686 -30370 61726 -30260
rect 61426 -30540 61496 -30500
rect 61696 -30540 61726 -30370
rect 61426 -30570 61726 -30540
rect 59656 -30770 60536 -30650
rect 37800 -31067 56220 -30908
rect 58396 -30930 58896 -30850
rect 37800 -31068 56221 -31067
rect 37800 -31228 56060 -31068
rect 56220 -31228 56221 -31068
rect 37800 -31229 56221 -31228
rect 37800 -31690 56200 -31229
rect 58396 -31290 58486 -30930
rect 58816 -31290 58896 -30930
rect 59796 -31010 59926 -30770
rect 59796 -31120 59806 -31010
rect 59916 -31120 59926 -31010
rect 59796 -31130 59926 -31120
rect 60436 -31030 60536 -30770
rect 60436 -31150 60446 -31030
rect 60526 -31150 60536 -31030
rect 60436 -31160 60536 -31150
rect 58396 -31350 58896 -31290
rect 61820 -31690 69400 -29720
rect 37800 -31728 69400 -31690
rect 37800 -31868 55320 -31728
rect 55470 -31868 69400 -31728
rect 37800 -31940 69400 -31868
rect 37800 -34347 56200 -31940
rect 56505 -33980 57017 -33979
rect 56505 -34230 56506 -33980
rect 57016 -34230 57017 -33980
rect 56505 -34231 57017 -34230
rect 58396 -34330 58896 -34240
rect 37800 -34348 56221 -34347
rect 37800 -34508 56060 -34348
rect 56220 -34508 56221 -34348
rect 37800 -34509 56221 -34508
rect 37800 -34558 56220 -34509
rect 37800 -36308 53050 -34558
rect 53250 -34954 56220 -34558
rect 58396 -34690 58486 -34330
rect 58816 -34690 58896 -34330
rect 60436 -34520 60536 -34510
rect 58396 -34800 58896 -34690
rect 59826 -34540 59976 -34530
rect 59826 -34630 59866 -34540
rect 59966 -34630 59976 -34540
rect 59826 -34640 59976 -34630
rect 60436 -34620 60446 -34520
rect 60526 -34620 60536 -34520
rect 59826 -34870 59946 -34640
rect 60436 -34870 60536 -34620
rect 59666 -34900 60536 -34870
rect 53250 -34964 57378 -34954
rect 53250 -35104 57098 -34964
rect 57368 -35104 57378 -34964
rect 59666 -34970 59976 -34900
rect 60316 -34970 60536 -34900
rect 61820 -34910 69400 -31940
rect 59666 -34990 60536 -34970
rect 61186 -34920 69400 -34910
rect 59666 -35040 59776 -34990
rect 53250 -35114 57378 -35104
rect 53250 -35448 56220 -35114
rect 53250 -35528 55020 -35448
rect 55120 -35528 56220 -35448
rect 53250 -35864 56220 -35528
rect 59656 -35440 59776 -35040
rect 61186 -35100 61206 -34920
rect 61346 -35100 69400 -34920
rect 61186 -35120 69400 -35100
rect 59906 -35180 60026 -35150
rect 59906 -35360 59916 -35180
rect 60006 -35360 60026 -35180
rect 59906 -35440 60026 -35360
rect 61186 -35440 61366 -35120
rect 59656 -35460 61366 -35440
rect 59656 -35480 61256 -35460
rect 59656 -35640 60096 -35480
rect 60176 -35640 61256 -35480
rect 59656 -35660 61256 -35640
rect 61326 -35660 61366 -35460
rect 59656 -35680 61366 -35660
rect 53250 -35874 57378 -35864
rect 53250 -36014 57098 -35874
rect 57368 -36014 57378 -35874
rect 53250 -36024 57378 -36014
rect 53250 -36308 56220 -36024
rect 59656 -36050 59776 -35680
rect 59906 -35690 60026 -35680
rect 59906 -35880 59916 -35690
rect 60006 -35880 60026 -35690
rect 61256 -35790 61366 -35680
rect 59906 -35890 60026 -35880
rect 61426 -35900 61446 -35660
rect 61686 -35770 61726 -35660
rect 61426 -35940 61496 -35900
rect 61696 -35940 61726 -35770
rect 61426 -35970 61726 -35940
rect 59656 -36170 60536 -36050
rect 37800 -36467 56220 -36308
rect 58396 -36330 58896 -36250
rect 37800 -36468 56221 -36467
rect 37800 -36628 56060 -36468
rect 56220 -36628 56221 -36468
rect 37800 -36629 56221 -36628
rect 37800 -37000 56200 -36629
rect 58396 -36690 58486 -36330
rect 58816 -36690 58896 -36330
rect 59796 -36410 59926 -36170
rect 59796 -36520 59806 -36410
rect 59916 -36520 59926 -36410
rect 59796 -36530 59926 -36520
rect 60436 -36430 60536 -36170
rect 60436 -36550 60446 -36430
rect 60526 -36550 60536 -36430
rect 60436 -36560 60536 -36550
rect 58396 -36750 58896 -36690
rect 61820 -36800 69400 -35120
rect 71900 -34100 74100 -34000
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 14000 -37090 56200 -37000
rect 61820 -37090 80600 -36800
rect 14000 -37128 80600 -37090
rect 14000 -37268 55320 -37128
rect 55470 -37268 80600 -37128
rect 14000 -37340 80600 -37268
rect 14000 -38000 56200 -37340
rect 14000 -49000 15000 -38000
rect 24000 -39747 56200 -38000
rect 61820 -38000 80600 -37340
rect 56505 -39380 57017 -39379
rect 56505 -39630 56506 -39380
rect 57016 -39630 57017 -39380
rect 56505 -39631 57017 -39630
rect 58396 -39730 58896 -39640
rect 24000 -39748 56221 -39747
rect 24000 -39908 56060 -39748
rect 56220 -39908 56221 -39748
rect 24000 -39909 56221 -39908
rect 24000 -39958 56220 -39909
rect 24000 -41708 53050 -39958
rect 53250 -40354 56220 -39958
rect 58396 -40090 58486 -39730
rect 58816 -40090 58896 -39730
rect 60436 -39920 60536 -39910
rect 58396 -40200 58896 -40090
rect 59826 -39940 59976 -39930
rect 59826 -40030 59866 -39940
rect 59966 -40030 59976 -39940
rect 59826 -40040 59976 -40030
rect 60436 -40020 60446 -39920
rect 60526 -40020 60536 -39920
rect 59826 -40270 59946 -40040
rect 60436 -40270 60536 -40020
rect 59666 -40300 60536 -40270
rect 53250 -40364 57378 -40354
rect 53250 -40504 57098 -40364
rect 57368 -40504 57378 -40364
rect 59666 -40370 59976 -40300
rect 60316 -40370 60536 -40300
rect 61820 -40310 69400 -38000
rect 59666 -40390 60536 -40370
rect 61186 -40320 69400 -40310
rect 59666 -40440 59776 -40390
rect 53250 -40514 57378 -40504
rect 53250 -40848 56220 -40514
rect 53250 -40928 55020 -40848
rect 55120 -40928 56220 -40848
rect 53250 -41264 56220 -40928
rect 59656 -40840 59776 -40440
rect 61186 -40500 61206 -40320
rect 61346 -40500 69400 -40320
rect 61186 -40520 69400 -40500
rect 59906 -40580 60026 -40550
rect 59906 -40760 59916 -40580
rect 60006 -40760 60026 -40580
rect 59906 -40840 60026 -40760
rect 61186 -40840 61366 -40520
rect 59656 -40860 61366 -40840
rect 59656 -40880 61256 -40860
rect 59656 -41040 60096 -40880
rect 60176 -41040 61256 -40880
rect 59656 -41060 61256 -41040
rect 61326 -41060 61366 -40860
rect 59656 -41080 61366 -41060
rect 53250 -41274 57378 -41264
rect 53250 -41414 57098 -41274
rect 57368 -41414 57378 -41274
rect 53250 -41424 57378 -41414
rect 53250 -41708 56220 -41424
rect 59656 -41450 59776 -41080
rect 59906 -41090 60026 -41080
rect 59906 -41280 59916 -41090
rect 60006 -41280 60026 -41090
rect 61256 -41190 61366 -41080
rect 59906 -41290 60026 -41280
rect 61426 -41300 61446 -41060
rect 61686 -41170 61726 -41060
rect 61426 -41340 61496 -41300
rect 61696 -41340 61726 -41170
rect 61426 -41370 61726 -41340
rect 59656 -41570 60536 -41450
rect 24000 -41867 56220 -41708
rect 58396 -41730 58896 -41650
rect 24000 -41868 56221 -41867
rect 24000 -42028 56060 -41868
rect 56220 -42028 56221 -41868
rect 24000 -42029 56221 -42028
rect 24000 -42490 56200 -42029
rect 58396 -42090 58486 -41730
rect 58816 -42090 58896 -41730
rect 59796 -41810 59926 -41570
rect 59796 -41920 59806 -41810
rect 59916 -41920 59926 -41810
rect 59796 -41930 59926 -41920
rect 60436 -41830 60536 -41570
rect 60436 -41950 60446 -41830
rect 60526 -41950 60536 -41830
rect 60436 -41960 60536 -41950
rect 58396 -42150 58896 -42090
rect 61820 -42490 69400 -40520
rect 24000 -42528 69400 -42490
rect 24000 -42668 55320 -42528
rect 55470 -42668 69400 -42528
rect 24000 -42740 69400 -42668
rect 24000 -45147 56200 -42740
rect 56505 -44780 57017 -44779
rect 56505 -45030 56506 -44780
rect 57016 -45030 57017 -44780
rect 56505 -45031 57017 -45030
rect 58396 -45130 58896 -45040
rect 24000 -45148 56221 -45147
rect 24000 -45308 56060 -45148
rect 56220 -45308 56221 -45148
rect 24000 -45309 56221 -45308
rect 24000 -45358 56220 -45309
rect 24000 -47108 53050 -45358
rect 53250 -45754 56220 -45358
rect 58396 -45490 58486 -45130
rect 58816 -45490 58896 -45130
rect 60436 -45320 60536 -45310
rect 58396 -45600 58896 -45490
rect 59826 -45340 59976 -45330
rect 59826 -45430 59866 -45340
rect 59966 -45430 59976 -45340
rect 59826 -45440 59976 -45430
rect 60436 -45420 60446 -45320
rect 60526 -45420 60536 -45320
rect 59826 -45670 59946 -45440
rect 60436 -45670 60536 -45420
rect 59666 -45700 60536 -45670
rect 53250 -45764 57378 -45754
rect 53250 -45904 57098 -45764
rect 57368 -45904 57378 -45764
rect 59666 -45770 59976 -45700
rect 60316 -45770 60536 -45700
rect 61820 -45710 69400 -42740
rect 59666 -45790 60536 -45770
rect 61186 -45720 69400 -45710
rect 59666 -45840 59776 -45790
rect 53250 -45914 57378 -45904
rect 53250 -46248 56220 -45914
rect 53250 -46328 55020 -46248
rect 55120 -46328 56220 -46248
rect 53250 -46664 56220 -46328
rect 59656 -46240 59776 -45840
rect 61186 -45900 61206 -45720
rect 61346 -45900 69400 -45720
rect 61186 -45920 69400 -45900
rect 59906 -45980 60026 -45950
rect 59906 -46160 59916 -45980
rect 60006 -46160 60026 -45980
rect 59906 -46240 60026 -46160
rect 61186 -46240 61366 -45920
rect 59656 -46260 61366 -46240
rect 59656 -46280 61256 -46260
rect 59656 -46440 60096 -46280
rect 60176 -46440 61256 -46280
rect 59656 -46460 61256 -46440
rect 61326 -46460 61366 -46260
rect 59656 -46480 61366 -46460
rect 53250 -46674 57378 -46664
rect 53250 -46814 57098 -46674
rect 57368 -46814 57378 -46674
rect 53250 -46824 57378 -46814
rect 53250 -47108 56220 -46824
rect 59656 -46850 59776 -46480
rect 59906 -46490 60026 -46480
rect 59906 -46680 59916 -46490
rect 60006 -46680 60026 -46490
rect 61256 -46590 61366 -46480
rect 59906 -46690 60026 -46680
rect 61426 -46700 61446 -46460
rect 61686 -46570 61726 -46460
rect 61426 -46740 61496 -46700
rect 61696 -46740 61726 -46570
rect 61426 -46770 61726 -46740
rect 59656 -46970 60536 -46850
rect 24000 -47267 56220 -47108
rect 58396 -47130 58896 -47050
rect 24000 -47268 56221 -47267
rect 24000 -47428 56060 -47268
rect 56220 -47428 56221 -47268
rect 24000 -47429 56221 -47428
rect 24000 -47890 56200 -47429
rect 58396 -47490 58486 -47130
rect 58816 -47490 58896 -47130
rect 59796 -47210 59926 -46970
rect 59796 -47320 59806 -47210
rect 59916 -47320 59926 -47210
rect 59796 -47330 59926 -47320
rect 60436 -47230 60536 -46970
rect 60436 -47350 60446 -47230
rect 60526 -47350 60536 -47230
rect 60436 -47360 60536 -47350
rect 58396 -47550 58896 -47490
rect 61820 -47890 69400 -45920
rect 24000 -47928 69400 -47890
rect 24000 -48068 55320 -47928
rect 55470 -48068 69400 -47928
rect 24000 -48140 69400 -48068
rect 24000 -49000 56200 -48140
rect 14000 -50000 56200 -49000
rect 37800 -50547 56200 -50000
rect 56505 -50180 57017 -50179
rect 56505 -50430 56506 -50180
rect 57016 -50430 57017 -50180
rect 56505 -50431 57017 -50430
rect 58396 -50530 58896 -50440
rect 37800 -50548 56221 -50547
rect 37800 -50708 56060 -50548
rect 56220 -50708 56221 -50548
rect 37800 -50709 56221 -50708
rect 37800 -50758 56220 -50709
rect 37800 -52508 53050 -50758
rect 53250 -51154 56220 -50758
rect 58396 -50890 58486 -50530
rect 58816 -50890 58896 -50530
rect 60436 -50720 60536 -50710
rect 58396 -51000 58896 -50890
rect 59826 -50740 59976 -50730
rect 59826 -50830 59866 -50740
rect 59966 -50830 59976 -50740
rect 59826 -50840 59976 -50830
rect 60436 -50820 60446 -50720
rect 60526 -50820 60536 -50720
rect 59826 -51070 59946 -50840
rect 60436 -51070 60536 -50820
rect 59666 -51100 60536 -51070
rect 53250 -51164 57378 -51154
rect 53250 -51304 57098 -51164
rect 57368 -51304 57378 -51164
rect 59666 -51170 59976 -51100
rect 60316 -51170 60536 -51100
rect 61820 -51110 69400 -48140
rect 59666 -51190 60536 -51170
rect 61186 -51120 69400 -51110
rect 59666 -51240 59776 -51190
rect 53250 -51314 57378 -51304
rect 53250 -51648 56220 -51314
rect 53250 -51728 55020 -51648
rect 55120 -51728 56220 -51648
rect 53250 -52064 56220 -51728
rect 59656 -51640 59776 -51240
rect 61186 -51300 61206 -51120
rect 61346 -51300 69400 -51120
rect 61186 -51320 69400 -51300
rect 59906 -51380 60026 -51350
rect 59906 -51560 59916 -51380
rect 60006 -51560 60026 -51380
rect 59906 -51640 60026 -51560
rect 61186 -51640 61366 -51320
rect 59656 -51660 61366 -51640
rect 59656 -51680 61256 -51660
rect 59656 -51840 60096 -51680
rect 60176 -51840 61256 -51680
rect 59656 -51860 61256 -51840
rect 61326 -51860 61366 -51660
rect 59656 -51880 61366 -51860
rect 53250 -52074 57378 -52064
rect 53250 -52214 57098 -52074
rect 57368 -52214 57378 -52074
rect 53250 -52224 57378 -52214
rect 53250 -52508 56220 -52224
rect 59656 -52250 59776 -51880
rect 59906 -51890 60026 -51880
rect 59906 -52080 59916 -51890
rect 60006 -52080 60026 -51890
rect 61256 -51990 61366 -51880
rect 59906 -52090 60026 -52080
rect 61426 -52100 61446 -51860
rect 61686 -51970 61726 -51860
rect 61426 -52140 61496 -52100
rect 61696 -52140 61726 -51970
rect 61426 -52170 61726 -52140
rect 59656 -52370 60536 -52250
rect 37800 -52667 56220 -52508
rect 58396 -52530 58896 -52450
rect 37800 -52668 56221 -52667
rect 37800 -52828 56060 -52668
rect 56220 -52828 56221 -52668
rect 37800 -52829 56221 -52828
rect 37800 -53290 56200 -52829
rect 58396 -52890 58486 -52530
rect 58816 -52890 58896 -52530
rect 59796 -52610 59926 -52370
rect 59796 -52720 59806 -52610
rect 59916 -52720 59926 -52610
rect 59796 -52730 59926 -52720
rect 60436 -52630 60536 -52370
rect 60436 -52750 60446 -52630
rect 60526 -52750 60536 -52630
rect 60436 -52760 60536 -52750
rect 58396 -52950 58896 -52890
rect 61820 -53290 69400 -51320
rect 37800 -53328 69400 -53290
rect 37800 -53468 55320 -53328
rect 55470 -53468 69400 -53328
rect 37800 -53540 69400 -53468
rect 37800 -55947 56200 -53540
rect 61820 -54400 69400 -53540
rect 76270 -38400 80600 -38000
rect 76270 -38540 76910 -38400
rect 77070 -38540 80600 -38400
rect 76270 -38630 80600 -38540
rect 76270 -39570 77080 -38630
rect 77160 -38790 77440 -38780
rect 77160 -39040 77170 -38790
rect 77430 -39040 77440 -38790
rect 77160 -39050 77440 -39040
rect 76270 -39720 76920 -39570
rect 77060 -39720 77080 -39570
rect 76270 -40820 77080 -39720
rect 79910 -39600 80600 -38630
rect 84700 -38050 85660 -37780
rect 84700 -38480 84960 -38050
rect 85400 -38480 85660 -38050
rect 84700 -38690 85660 -38480
rect 87880 -38390 88840 -38140
rect 87880 -38820 88150 -38390
rect 88590 -38820 88840 -38390
rect 87880 -39050 88840 -38820
rect 79910 -39830 88480 -39600
rect 79910 -39980 83150 -39830
rect 79400 -40150 79690 -40140
rect 79400 -40390 79410 -40150
rect 79680 -40390 79690 -40150
rect 79400 -40400 79690 -40390
rect 76270 -40960 76920 -40820
rect 77060 -40960 77080 -40820
rect 76270 -42060 77080 -40960
rect 79400 -41380 79690 -41370
rect 79400 -41620 79410 -41380
rect 79680 -41620 79690 -41380
rect 79400 -41630 79690 -41620
rect 76270 -42220 76920 -42060
rect 77060 -42220 77080 -42060
rect 76270 -43310 77080 -42220
rect 79400 -42640 79690 -42630
rect 79400 -42880 79410 -42640
rect 79680 -42880 79690 -42640
rect 79400 -42890 79690 -42880
rect 76270 -43450 76920 -43310
rect 77060 -43450 77080 -43310
rect 76270 -44520 77080 -43450
rect 79400 -43860 79690 -43850
rect 79400 -44100 79410 -43860
rect 79680 -44100 79690 -43860
rect 79400 -44110 79690 -44100
rect 76270 -44610 76920 -44520
rect 77060 -44610 77080 -44520
rect 76270 -45640 77080 -44610
rect 79910 -44410 80600 -39980
rect 83000 -40180 83150 -39980
rect 83510 -39980 88480 -39830
rect 83510 -40180 83640 -39980
rect 81110 -40250 81600 -40220
rect 81110 -40510 81140 -40250
rect 81570 -40510 81600 -40250
rect 83000 -40290 83640 -40180
rect 87520 -40240 88480 -39980
rect 81110 -40540 81600 -40510
rect 87520 -40590 87830 -40240
rect 88190 -40590 88480 -40240
rect 87520 -40890 88480 -40590
rect 82790 -42740 91440 -42710
rect 82790 -43310 82820 -42740
rect 91410 -43310 91440 -42740
rect 82790 -43340 91440 -43310
rect 79910 -44440 91440 -44410
rect 79910 -45010 82820 -44440
rect 91410 -45010 91440 -44440
rect 79910 -45040 91440 -45010
rect 79400 -45120 79690 -45110
rect 79400 -45360 79410 -45120
rect 79680 -45360 79690 -45120
rect 79400 -45370 79690 -45360
rect 76270 -45740 76920 -45640
rect 77060 -45740 77080 -45640
rect 76270 -46440 77080 -45740
rect 76270 -46580 76910 -46440
rect 77070 -46580 77080 -46440
rect 76270 -47610 77080 -46580
rect 77160 -46830 77440 -46820
rect 77160 -47080 77170 -46830
rect 77430 -47080 77440 -46830
rect 77160 -47090 77440 -47080
rect 76270 -47760 76920 -47610
rect 77060 -47760 77080 -47610
rect 76270 -48860 77080 -47760
rect 79400 -48190 79690 -48180
rect 79400 -48430 79410 -48190
rect 79680 -48430 79690 -48190
rect 79400 -48440 79690 -48430
rect 76270 -49000 76920 -48860
rect 77060 -49000 77080 -48860
rect 76270 -50100 77080 -49000
rect 79910 -48540 80600 -45040
rect 82794 -46878 91444 -46848
rect 82794 -47448 82824 -46878
rect 91414 -47448 91444 -46878
rect 82794 -47478 91444 -47448
rect 79910 -48578 91450 -48540
rect 79910 -49148 82824 -48578
rect 91414 -49148 91450 -48578
rect 79910 -49180 91450 -49148
rect 79400 -49420 79690 -49410
rect 79400 -49660 79410 -49420
rect 79680 -49660 79690 -49420
rect 79400 -49670 79690 -49660
rect 76270 -50260 76920 -50100
rect 77060 -50260 77080 -50100
rect 76270 -51350 77080 -50260
rect 79400 -50680 79690 -50670
rect 79400 -50920 79410 -50680
rect 79680 -50920 79690 -50680
rect 79400 -50930 79690 -50920
rect 76270 -51490 76920 -51350
rect 77060 -51490 77080 -51350
rect 76270 -52560 77080 -51490
rect 79400 -51900 79690 -51890
rect 79400 -52140 79410 -51900
rect 79680 -52140 79690 -51900
rect 79400 -52150 79690 -52140
rect 76270 -52650 76920 -52560
rect 77060 -52650 77080 -52560
rect 76270 -53680 77080 -52650
rect 79910 -52200 80600 -49180
rect 82790 -50530 91440 -50500
rect 82790 -51100 82820 -50530
rect 91410 -51100 91440 -50530
rect 82790 -51130 91440 -51100
rect 79910 -52230 91440 -52200
rect 79910 -52800 82820 -52230
rect 91410 -52800 91440 -52230
rect 79910 -52830 91440 -52800
rect 79400 -53160 79690 -53150
rect 79400 -53400 79410 -53160
rect 79680 -53400 79690 -53160
rect 79400 -53410 79690 -53400
rect 76270 -53780 76920 -53680
rect 77060 -53780 77080 -53680
rect 76270 -53800 77080 -53780
rect 81400 -54400 91400 -52830
rect 56505 -55580 57017 -55579
rect 56505 -55830 56506 -55580
rect 57016 -55830 57017 -55580
rect 56505 -55831 57017 -55830
rect 58396 -55930 58896 -55840
rect 37800 -55948 56221 -55947
rect 37800 -56108 56060 -55948
rect 56220 -56108 56221 -55948
rect 37800 -56109 56221 -56108
rect 37800 -56158 56220 -56109
rect 37800 -57908 53050 -56158
rect 53250 -56554 56220 -56158
rect 58396 -56290 58486 -55930
rect 58816 -56290 58896 -55930
rect 61820 -56000 91400 -54400
rect 60436 -56120 60536 -56110
rect 58396 -56400 58896 -56290
rect 59826 -56140 59976 -56130
rect 59826 -56230 59866 -56140
rect 59966 -56230 59976 -56140
rect 59826 -56240 59976 -56230
rect 60436 -56220 60446 -56120
rect 60526 -56220 60536 -56120
rect 59826 -56470 59946 -56240
rect 60436 -56470 60536 -56220
rect 59666 -56500 60536 -56470
rect 53250 -56564 57378 -56554
rect 53250 -56704 57098 -56564
rect 57368 -56704 57378 -56564
rect 59666 -56570 59976 -56500
rect 60316 -56570 60536 -56500
rect 61820 -56510 69300 -56000
rect 59666 -56590 60536 -56570
rect 61186 -56520 69300 -56510
rect 59666 -56640 59776 -56590
rect 53250 -56714 57378 -56704
rect 53250 -57048 56220 -56714
rect 53250 -57128 55020 -57048
rect 55120 -57128 56220 -57048
rect 53250 -57464 56220 -57128
rect 59656 -57040 59776 -56640
rect 61186 -56700 61206 -56520
rect 61346 -56700 69300 -56520
rect 61186 -56720 69300 -56700
rect 59906 -56780 60026 -56750
rect 59906 -56960 59916 -56780
rect 60006 -56960 60026 -56780
rect 59906 -57040 60026 -56960
rect 61186 -57040 61366 -56720
rect 59656 -57060 61366 -57040
rect 59656 -57080 61256 -57060
rect 59656 -57240 60096 -57080
rect 60176 -57240 61256 -57080
rect 59656 -57260 61256 -57240
rect 61326 -57260 61366 -57060
rect 59656 -57280 61366 -57260
rect 53250 -57474 57378 -57464
rect 53250 -57614 57098 -57474
rect 57368 -57614 57378 -57474
rect 53250 -57624 57378 -57614
rect 53250 -57908 56220 -57624
rect 59656 -57650 59776 -57280
rect 59906 -57290 60026 -57280
rect 59906 -57480 59916 -57290
rect 60006 -57480 60026 -57290
rect 61256 -57390 61366 -57280
rect 59906 -57490 60026 -57480
rect 61426 -57500 61446 -57260
rect 61686 -57370 61726 -57260
rect 61426 -57540 61496 -57500
rect 61696 -57540 61726 -57370
rect 61426 -57570 61726 -57540
rect 59656 -57770 60536 -57650
rect 37800 -58067 56220 -57908
rect 58396 -57930 58896 -57850
rect 37800 -58068 56221 -58067
rect 37800 -58228 56060 -58068
rect 56220 -58228 56221 -58068
rect 37800 -58229 56221 -58228
rect 37800 -58690 56200 -58229
rect 58396 -58290 58486 -57930
rect 58816 -58290 58896 -57930
rect 59796 -58010 59926 -57770
rect 59796 -58120 59806 -58010
rect 59916 -58120 59926 -58010
rect 59796 -58130 59926 -58120
rect 60436 -58030 60536 -57770
rect 60436 -58150 60446 -58030
rect 60526 -58150 60536 -58030
rect 60436 -58160 60536 -58150
rect 58396 -58350 58896 -58290
rect 61820 -58690 69300 -56720
rect 37800 -58728 69300 -58690
rect 37800 -58868 55320 -58728
rect 55470 -58868 69300 -58728
rect 37800 -58940 69300 -58868
rect 37800 -61347 56200 -58940
rect 56505 -60980 57017 -60979
rect 56505 -61230 56506 -60980
rect 57016 -61230 57017 -60980
rect 56505 -61231 57017 -61230
rect 58396 -61330 58896 -61240
rect 37800 -61348 56221 -61347
rect 37800 -61508 56060 -61348
rect 56220 -61508 56221 -61348
rect 37800 -61509 56221 -61508
rect 37800 -61558 56220 -61509
rect 37800 -63308 53050 -61558
rect 53250 -61954 56220 -61558
rect 58396 -61690 58486 -61330
rect 58816 -61690 58896 -61330
rect 60436 -61520 60536 -61510
rect 58396 -61800 58896 -61690
rect 59826 -61540 59976 -61530
rect 59826 -61630 59866 -61540
rect 59966 -61630 59976 -61540
rect 59826 -61640 59976 -61630
rect 60436 -61620 60446 -61520
rect 60526 -61620 60536 -61520
rect 59826 -61870 59946 -61640
rect 60436 -61870 60536 -61620
rect 59666 -61900 60536 -61870
rect 53250 -61964 57378 -61954
rect 53250 -62104 57098 -61964
rect 57368 -62104 57378 -61964
rect 59666 -61970 59976 -61900
rect 60316 -61970 60536 -61900
rect 61820 -61910 69300 -58940
rect 59666 -61990 60536 -61970
rect 61186 -61920 69300 -61910
rect 59666 -62040 59776 -61990
rect 53250 -62114 57378 -62104
rect 53250 -62448 56220 -62114
rect 53250 -62528 55020 -62448
rect 55120 -62528 56220 -62448
rect 53250 -62864 56220 -62528
rect 59656 -62440 59776 -62040
rect 61186 -62100 61206 -61920
rect 61346 -62100 69300 -61920
rect 61186 -62120 69300 -62100
rect 59906 -62180 60026 -62150
rect 59906 -62360 59916 -62180
rect 60006 -62360 60026 -62180
rect 59906 -62440 60026 -62360
rect 61186 -62440 61366 -62120
rect 59656 -62460 61366 -62440
rect 59656 -62480 61256 -62460
rect 59656 -62640 60096 -62480
rect 60176 -62640 61256 -62480
rect 59656 -62660 61256 -62640
rect 61326 -62660 61366 -62460
rect 59656 -62680 61366 -62660
rect 53250 -62874 57378 -62864
rect 53250 -63014 57098 -62874
rect 57368 -63014 57378 -62874
rect 53250 -63024 57378 -63014
rect 53250 -63308 56220 -63024
rect 59656 -63050 59776 -62680
rect 59906 -62690 60026 -62680
rect 59906 -62880 59916 -62690
rect 60006 -62880 60026 -62690
rect 61256 -62790 61366 -62680
rect 59906 -62890 60026 -62880
rect 61426 -62900 61446 -62660
rect 61686 -62770 61726 -62660
rect 61426 -62940 61496 -62900
rect 61696 -62940 61726 -62770
rect 61426 -62970 61726 -62940
rect 59656 -63170 60536 -63050
rect 37800 -63467 56220 -63308
rect 58396 -63330 58896 -63250
rect 37800 -63468 56221 -63467
rect 37800 -63628 56060 -63468
rect 56220 -63628 56221 -63468
rect 37800 -63629 56221 -63628
rect 37800 -64090 56200 -63629
rect 58396 -63690 58486 -63330
rect 58816 -63690 58896 -63330
rect 59796 -63410 59926 -63170
rect 59796 -63520 59806 -63410
rect 59916 -63520 59926 -63410
rect 59796 -63530 59926 -63520
rect 60436 -63430 60536 -63170
rect 60436 -63550 60446 -63430
rect 60526 -63550 60536 -63430
rect 60436 -63560 60536 -63550
rect 58396 -63750 58896 -63690
rect 61820 -64090 69300 -62120
rect 37800 -64128 69300 -64090
rect 37800 -64268 55320 -64128
rect 55470 -64268 69300 -64128
rect 37800 -64340 69300 -64268
rect 37800 -66747 56200 -64340
rect 56505 -66380 57017 -66379
rect 56505 -66630 56506 -66380
rect 57016 -66630 57017 -66380
rect 56505 -66631 57017 -66630
rect 58396 -66730 58896 -66640
rect 37800 -66748 56221 -66747
rect 37800 -66908 56060 -66748
rect 56220 -66908 56221 -66748
rect 37800 -66909 56221 -66908
rect 37800 -66958 56220 -66909
rect 37800 -68708 53050 -66958
rect 53250 -67354 56220 -66958
rect 58396 -67090 58486 -66730
rect 58816 -67090 58896 -66730
rect 60436 -66920 60536 -66910
rect 58396 -67200 58896 -67090
rect 59826 -66940 59976 -66930
rect 59826 -67030 59866 -66940
rect 59966 -67030 59976 -66940
rect 59826 -67040 59976 -67030
rect 60436 -67020 60446 -66920
rect 60526 -67020 60536 -66920
rect 59826 -67270 59946 -67040
rect 60436 -67270 60536 -67020
rect 59666 -67300 60536 -67270
rect 53250 -67364 57378 -67354
rect 53250 -67504 57098 -67364
rect 57368 -67504 57378 -67364
rect 59666 -67370 59976 -67300
rect 60316 -67370 60536 -67300
rect 61820 -67310 69300 -64340
rect 59666 -67390 60536 -67370
rect 61186 -67320 69300 -67310
rect 59666 -67440 59776 -67390
rect 53250 -67514 57378 -67504
rect 53250 -67848 56220 -67514
rect 53250 -67928 55020 -67848
rect 55120 -67928 56220 -67848
rect 53250 -68264 56220 -67928
rect 59656 -67840 59776 -67440
rect 61186 -67500 61206 -67320
rect 61346 -67500 69300 -67320
rect 61186 -67520 69300 -67500
rect 59906 -67580 60026 -67550
rect 59906 -67760 59916 -67580
rect 60006 -67760 60026 -67580
rect 59906 -67840 60026 -67760
rect 61186 -67840 61366 -67520
rect 59656 -67860 61366 -67840
rect 59656 -67880 61256 -67860
rect 59656 -68040 60096 -67880
rect 60176 -68040 61256 -67880
rect 59656 -68060 61256 -68040
rect 61326 -68060 61366 -67860
rect 59656 -68080 61366 -68060
rect 53250 -68274 57378 -68264
rect 53250 -68414 57098 -68274
rect 57368 -68414 57378 -68274
rect 53250 -68424 57378 -68414
rect 53250 -68708 56220 -68424
rect 59656 -68450 59776 -68080
rect 59906 -68090 60026 -68080
rect 59906 -68280 59916 -68090
rect 60006 -68280 60026 -68090
rect 61256 -68190 61366 -68080
rect 59906 -68290 60026 -68280
rect 61426 -68300 61446 -68060
rect 61686 -68170 61726 -68060
rect 61426 -68340 61496 -68300
rect 61696 -68340 61726 -68170
rect 61426 -68370 61726 -68340
rect 59656 -68570 60536 -68450
rect 37800 -68867 56220 -68708
rect 58396 -68730 58896 -68650
rect 37800 -68868 56221 -68867
rect 37800 -69028 56060 -68868
rect 56220 -69028 56221 -68868
rect 37800 -69029 56221 -69028
rect 37800 -69490 56200 -69029
rect 58396 -69090 58486 -68730
rect 58816 -69090 58896 -68730
rect 59796 -68810 59926 -68570
rect 59796 -68920 59806 -68810
rect 59916 -68920 59926 -68810
rect 59796 -68930 59926 -68920
rect 60436 -68830 60536 -68570
rect 60436 -68950 60446 -68830
rect 60526 -68950 60536 -68830
rect 60436 -68960 60536 -68950
rect 58396 -69150 58896 -69090
rect 61820 -69490 69300 -67520
rect 37800 -69528 69300 -69490
rect 37800 -69668 55320 -69528
rect 55470 -69668 69300 -69528
rect 37800 -69740 69300 -69668
rect 37800 -72147 56200 -69740
rect 56505 -71780 57017 -71779
rect 56505 -72030 56506 -71780
rect 57016 -72030 57017 -71780
rect 56505 -72031 57017 -72030
rect 58396 -72130 58896 -72040
rect 37800 -72148 56221 -72147
rect 37800 -72308 56060 -72148
rect 56220 -72308 56221 -72148
rect 37800 -72309 56221 -72308
rect 37800 -72358 56220 -72309
rect 37800 -74108 53050 -72358
rect 53250 -72754 56220 -72358
rect 58396 -72490 58486 -72130
rect 58816 -72490 58896 -72130
rect 60436 -72320 60536 -72310
rect 58396 -72600 58896 -72490
rect 59826 -72340 59976 -72330
rect 59826 -72430 59866 -72340
rect 59966 -72430 59976 -72340
rect 59826 -72440 59976 -72430
rect 60436 -72420 60446 -72320
rect 60526 -72420 60536 -72320
rect 59826 -72670 59946 -72440
rect 60436 -72670 60536 -72420
rect 59666 -72700 60536 -72670
rect 53250 -72764 57378 -72754
rect 53250 -72904 57098 -72764
rect 57368 -72904 57378 -72764
rect 59666 -72770 59976 -72700
rect 60316 -72770 60536 -72700
rect 61820 -72710 69300 -69740
rect 59666 -72790 60536 -72770
rect 61186 -72720 69300 -72710
rect 59666 -72840 59776 -72790
rect 53250 -72914 57378 -72904
rect 53250 -73248 56220 -72914
rect 53250 -73328 55020 -73248
rect 55120 -73328 56220 -73248
rect 53250 -73664 56220 -73328
rect 59656 -73240 59776 -72840
rect 61186 -72900 61206 -72720
rect 61346 -72900 69300 -72720
rect 61186 -72920 69300 -72900
rect 59906 -72980 60026 -72950
rect 59906 -73160 59916 -72980
rect 60006 -73160 60026 -72980
rect 59906 -73240 60026 -73160
rect 61186 -73240 61366 -72920
rect 59656 -73260 61366 -73240
rect 59656 -73280 61256 -73260
rect 59656 -73440 60096 -73280
rect 60176 -73440 61256 -73280
rect 59656 -73460 61256 -73440
rect 61326 -73460 61366 -73260
rect 59656 -73480 61366 -73460
rect 53250 -73674 57378 -73664
rect 53250 -73814 57098 -73674
rect 57368 -73814 57378 -73674
rect 53250 -73824 57378 -73814
rect 53250 -74108 56220 -73824
rect 59656 -73850 59776 -73480
rect 59906 -73490 60026 -73480
rect 59906 -73680 59916 -73490
rect 60006 -73680 60026 -73490
rect 61256 -73590 61366 -73480
rect 59906 -73690 60026 -73680
rect 61426 -73700 61446 -73460
rect 61686 -73570 61726 -73460
rect 61426 -73740 61496 -73700
rect 61696 -73740 61726 -73570
rect 61426 -73770 61726 -73740
rect 59656 -73970 60536 -73850
rect 37800 -74267 56220 -74108
rect 58396 -74130 58896 -74050
rect 37800 -74268 56221 -74267
rect 37800 -74428 56060 -74268
rect 56220 -74428 56221 -74268
rect 37800 -74429 56221 -74428
rect 37800 -74890 56200 -74429
rect 58396 -74490 58486 -74130
rect 58816 -74490 58896 -74130
rect 59796 -74210 59926 -73970
rect 59796 -74320 59806 -74210
rect 59916 -74320 59926 -74210
rect 59796 -74330 59926 -74320
rect 60436 -74230 60536 -73970
rect 60436 -74350 60446 -74230
rect 60526 -74350 60536 -74230
rect 60436 -74360 60536 -74350
rect 58396 -74550 58896 -74490
rect 61820 -74890 69300 -72920
rect 37800 -74928 69300 -74890
rect 37800 -75068 55320 -74928
rect 55470 -75068 69300 -74928
rect 37800 -75140 69300 -75068
rect 37800 -77547 56200 -75140
rect 56505 -77180 57017 -77179
rect 56505 -77430 56506 -77180
rect 57016 -77430 57017 -77180
rect 56505 -77431 57017 -77430
rect 58396 -77530 58896 -77440
rect 37800 -77548 56221 -77547
rect 37800 -77708 56060 -77548
rect 56220 -77708 56221 -77548
rect 37800 -77709 56221 -77708
rect 37800 -77758 56220 -77709
rect 37800 -79508 53050 -77758
rect 53250 -78154 56220 -77758
rect 58396 -77890 58486 -77530
rect 58816 -77890 58896 -77530
rect 60436 -77720 60536 -77710
rect 58396 -78000 58896 -77890
rect 59826 -77740 59976 -77730
rect 59826 -77830 59866 -77740
rect 59966 -77830 59976 -77740
rect 59826 -77840 59976 -77830
rect 60436 -77820 60446 -77720
rect 60526 -77820 60536 -77720
rect 59826 -78070 59946 -77840
rect 60436 -78070 60536 -77820
rect 59666 -78100 60536 -78070
rect 53250 -78164 57378 -78154
rect 53250 -78304 57098 -78164
rect 57368 -78304 57378 -78164
rect 59666 -78170 59976 -78100
rect 60316 -78170 60536 -78100
rect 61820 -78110 69300 -75140
rect 59666 -78190 60536 -78170
rect 61186 -78120 69300 -78110
rect 59666 -78240 59776 -78190
rect 53250 -78314 57378 -78304
rect 53250 -78648 56220 -78314
rect 53250 -78728 55020 -78648
rect 55120 -78728 56220 -78648
rect 53250 -79064 56220 -78728
rect 59656 -78640 59776 -78240
rect 61186 -78300 61206 -78120
rect 61346 -78300 69300 -78120
rect 61186 -78320 69300 -78300
rect 59906 -78380 60026 -78350
rect 59906 -78560 59916 -78380
rect 60006 -78560 60026 -78380
rect 59906 -78640 60026 -78560
rect 61186 -78640 61366 -78320
rect 59656 -78660 61366 -78640
rect 59656 -78680 61256 -78660
rect 59656 -78840 60096 -78680
rect 60176 -78840 61256 -78680
rect 59656 -78860 61256 -78840
rect 61326 -78860 61366 -78660
rect 59656 -78880 61366 -78860
rect 53250 -79074 57378 -79064
rect 53250 -79214 57098 -79074
rect 57368 -79214 57378 -79074
rect 53250 -79224 57378 -79214
rect 53250 -79508 56220 -79224
rect 59656 -79250 59776 -78880
rect 59906 -78890 60026 -78880
rect 59906 -79080 59916 -78890
rect 60006 -79080 60026 -78890
rect 61256 -78990 61366 -78880
rect 59906 -79090 60026 -79080
rect 61426 -79100 61446 -78860
rect 61686 -78970 61726 -78860
rect 61426 -79140 61496 -79100
rect 61696 -79140 61726 -78970
rect 61426 -79170 61726 -79140
rect 59656 -79370 60536 -79250
rect 37800 -79667 56220 -79508
rect 58396 -79530 58896 -79450
rect 37800 -79668 56221 -79667
rect 37800 -79828 56060 -79668
rect 56220 -79828 56221 -79668
rect 37800 -79829 56221 -79828
rect 37800 -80290 56200 -79829
rect 58396 -79890 58486 -79530
rect 58816 -79890 58896 -79530
rect 59796 -79610 59926 -79370
rect 59796 -79720 59806 -79610
rect 59916 -79720 59926 -79610
rect 59796 -79730 59926 -79720
rect 60436 -79630 60536 -79370
rect 60436 -79750 60446 -79630
rect 60526 -79750 60536 -79630
rect 60436 -79760 60536 -79750
rect 58396 -79950 58896 -79890
rect 61820 -80290 69300 -78320
rect 37800 -80328 69300 -80290
rect 37800 -80468 55320 -80328
rect 55470 -80468 69300 -80328
rect 37800 -80540 69300 -80468
rect 37800 -82947 56200 -80540
rect 56505 -82580 57017 -82579
rect 56505 -82830 56506 -82580
rect 57016 -82830 57017 -82580
rect 56505 -82831 57017 -82830
rect 58396 -82930 58896 -82840
rect 37800 -82948 56221 -82947
rect 37800 -83108 56060 -82948
rect 56220 -83108 56221 -82948
rect 37800 -83109 56221 -83108
rect 37800 -83158 56220 -83109
rect 37800 -84908 53050 -83158
rect 53250 -83554 56220 -83158
rect 58396 -83290 58486 -82930
rect 58816 -83290 58896 -82930
rect 60436 -83120 60536 -83110
rect 58396 -83400 58896 -83290
rect 59826 -83140 59976 -83130
rect 59826 -83230 59866 -83140
rect 59966 -83230 59976 -83140
rect 59826 -83240 59976 -83230
rect 60436 -83220 60446 -83120
rect 60526 -83220 60536 -83120
rect 59826 -83470 59946 -83240
rect 60436 -83470 60536 -83220
rect 59666 -83500 60536 -83470
rect 53250 -83564 57378 -83554
rect 53250 -83704 57098 -83564
rect 57368 -83704 57378 -83564
rect 59666 -83570 59976 -83500
rect 60316 -83570 60536 -83500
rect 61820 -83510 69300 -80540
rect 59666 -83590 60536 -83570
rect 61186 -83520 69300 -83510
rect 59666 -83640 59776 -83590
rect 53250 -83714 57378 -83704
rect 53250 -84048 56220 -83714
rect 53250 -84128 55020 -84048
rect 55120 -84128 56220 -84048
rect 53250 -84464 56220 -84128
rect 59656 -84040 59776 -83640
rect 61186 -83700 61206 -83520
rect 61346 -83700 69300 -83520
rect 61186 -83720 69300 -83700
rect 59906 -83780 60026 -83750
rect 59906 -83960 59916 -83780
rect 60006 -83960 60026 -83780
rect 59906 -84040 60026 -83960
rect 61186 -84040 61366 -83720
rect 59656 -84060 61366 -84040
rect 59656 -84080 61256 -84060
rect 59656 -84240 60096 -84080
rect 60176 -84240 61256 -84080
rect 59656 -84260 61256 -84240
rect 61326 -84260 61366 -84060
rect 59656 -84280 61366 -84260
rect 53250 -84474 57378 -84464
rect 53250 -84614 57098 -84474
rect 57368 -84614 57378 -84474
rect 53250 -84624 57378 -84614
rect 53250 -84908 56220 -84624
rect 59656 -84650 59776 -84280
rect 59906 -84290 60026 -84280
rect 59906 -84480 59916 -84290
rect 60006 -84480 60026 -84290
rect 61256 -84390 61366 -84280
rect 59906 -84490 60026 -84480
rect 61426 -84500 61446 -84260
rect 61686 -84370 61726 -84260
rect 61426 -84540 61496 -84500
rect 61696 -84540 61726 -84370
rect 61426 -84570 61726 -84540
rect 59656 -84770 60536 -84650
rect 37800 -85067 56220 -84908
rect 58396 -84930 58896 -84850
rect 37800 -85068 56221 -85067
rect 37800 -85228 56060 -85068
rect 56220 -85228 56221 -85068
rect 37800 -85229 56221 -85228
rect 37800 -85690 56200 -85229
rect 58396 -85290 58486 -84930
rect 58816 -85290 58896 -84930
rect 59796 -85010 59926 -84770
rect 59796 -85120 59806 -85010
rect 59916 -85120 59926 -85010
rect 59796 -85130 59926 -85120
rect 60436 -85030 60536 -84770
rect 60436 -85150 60446 -85030
rect 60526 -85150 60536 -85030
rect 60436 -85160 60536 -85150
rect 58396 -85350 58896 -85290
rect 61820 -85690 69300 -83720
rect 37800 -85728 69300 -85690
rect 37800 -85868 55320 -85728
rect 55470 -85868 69300 -85728
rect 37800 -85940 69300 -85868
rect 37800 -86700 56200 -85940
rect 53200 -86800 56200 -86700
<< via4 >>
rect 43000 1000 46400 2400
rect 43000 -1400 46400 0
rect 56506 -1830 57016 -1580
rect 58486 -2290 58816 -1930
rect 58516 -3060 58796 -2990
rect 58516 -3260 58556 -3060
rect 58556 -3260 58756 -3060
rect 58756 -3260 58796 -3060
rect 58516 -3340 58796 -3260
rect 61446 -3370 61686 -3260
rect 61446 -3500 61496 -3370
rect 61496 -3500 61686 -3370
rect 56628 -4268 57026 -4222
rect 56628 -4486 56654 -4268
rect 56654 -4486 56998 -4268
rect 56998 -4486 57026 -4268
rect 58486 -4290 58816 -3930
rect 56628 -4526 57026 -4486
rect 21000 -7400 22000 -6600
rect 56506 -7230 57016 -6980
rect 58486 -7690 58816 -7330
rect 58516 -8460 58796 -8390
rect 58516 -8660 58556 -8460
rect 58556 -8660 58756 -8460
rect 58756 -8660 58796 -8460
rect 58516 -8740 58796 -8660
rect 61446 -8770 61686 -8660
rect 61446 -8900 61496 -8770
rect 61496 -8900 61686 -8770
rect 56628 -9668 57026 -9622
rect 56628 -9886 56654 -9668
rect 56654 -9886 56998 -9668
rect 56998 -9886 57026 -9668
rect 58486 -9690 58816 -9330
rect 56628 -9926 57026 -9886
rect 56506 -12630 57016 -12380
rect 58486 -13090 58816 -12730
rect 58516 -13860 58796 -13790
rect 58516 -14060 58556 -13860
rect 58556 -14060 58756 -13860
rect 58756 -14060 58796 -13860
rect 58516 -14140 58796 -14060
rect 61446 -14170 61686 -14060
rect 61446 -14300 61496 -14170
rect 61496 -14300 61686 -14170
rect 56628 -15068 57026 -15022
rect 56628 -15286 56654 -15068
rect 56654 -15286 56998 -15068
rect 56998 -15286 57026 -15068
rect 58486 -15090 58816 -14730
rect 56628 -15326 57026 -15286
rect 56506 -18030 57016 -17780
rect 58486 -18490 58816 -18130
rect 58516 -19260 58796 -19190
rect 58516 -19460 58556 -19260
rect 58556 -19460 58756 -19260
rect 58756 -19460 58796 -19260
rect 58516 -19540 58796 -19460
rect 61446 -19570 61686 -19460
rect 61446 -19700 61496 -19570
rect 61496 -19700 61686 -19570
rect 56628 -20468 57026 -20422
rect 56628 -20686 56654 -20468
rect 56654 -20686 56998 -20468
rect 56998 -20686 57026 -20468
rect 58486 -20490 58816 -20130
rect 56628 -20726 57026 -20686
rect 56506 -23430 57016 -23180
rect 58486 -23890 58816 -23530
rect 58516 -24660 58796 -24590
rect 58516 -24860 58556 -24660
rect 58556 -24860 58756 -24660
rect 58756 -24860 58796 -24660
rect 58516 -24940 58796 -24860
rect 61446 -24970 61686 -24860
rect 61446 -25100 61496 -24970
rect 61496 -25100 61686 -24970
rect 56628 -25868 57026 -25822
rect 56628 -26086 56654 -25868
rect 56654 -26086 56998 -25868
rect 56998 -26086 57026 -25868
rect 58486 -25890 58816 -25530
rect 56628 -26126 57026 -26086
rect 56506 -28830 57016 -28580
rect 58486 -29290 58816 -28930
rect 58516 -30060 58796 -29990
rect 58516 -30260 58556 -30060
rect 58556 -30260 58756 -30060
rect 58756 -30260 58796 -30060
rect 58516 -30340 58796 -30260
rect 61446 -30370 61686 -30260
rect 61446 -30500 61496 -30370
rect 61496 -30500 61686 -30370
rect 56628 -31268 57026 -31222
rect 56628 -31486 56654 -31268
rect 56654 -31486 56998 -31268
rect 56998 -31486 57026 -31268
rect 58486 -31290 58816 -30930
rect 56628 -31526 57026 -31486
rect 56506 -34230 57016 -33980
rect 58486 -34690 58816 -34330
rect 58516 -35460 58796 -35390
rect 58516 -35660 58556 -35460
rect 58556 -35660 58756 -35460
rect 58756 -35660 58796 -35460
rect 58516 -35740 58796 -35660
rect 61446 -35770 61686 -35660
rect 61446 -35900 61496 -35770
rect 61496 -35900 61686 -35770
rect 56628 -36668 57026 -36622
rect 56628 -36886 56654 -36668
rect 56654 -36886 56998 -36668
rect 56998 -36886 57026 -36668
rect 58486 -36690 58816 -36330
rect 56628 -36926 57026 -36886
rect 72000 -35500 74000 -34100
rect 56506 -39630 57016 -39380
rect 58486 -40090 58816 -39730
rect 58516 -40860 58796 -40790
rect 58516 -41060 58556 -40860
rect 58556 -41060 58756 -40860
rect 58756 -41060 58796 -40860
rect 58516 -41140 58796 -41060
rect 61446 -41170 61686 -41060
rect 61446 -41300 61496 -41170
rect 61496 -41300 61686 -41170
rect 56628 -42068 57026 -42022
rect 56628 -42286 56654 -42068
rect 56654 -42286 56998 -42068
rect 56998 -42286 57026 -42068
rect 58486 -42090 58816 -41730
rect 56628 -42326 57026 -42286
rect 56506 -45030 57016 -44780
rect 58486 -45490 58816 -45130
rect 58516 -46260 58796 -46190
rect 58516 -46460 58556 -46260
rect 58556 -46460 58756 -46260
rect 58756 -46460 58796 -46260
rect 58516 -46540 58796 -46460
rect 61446 -46570 61686 -46460
rect 61446 -46700 61496 -46570
rect 61496 -46700 61686 -46570
rect 56628 -47468 57026 -47422
rect 56628 -47686 56654 -47468
rect 56654 -47686 56998 -47468
rect 56998 -47686 57026 -47468
rect 58486 -47490 58816 -47130
rect 56628 -47726 57026 -47686
rect 56506 -50430 57016 -50180
rect 58486 -50890 58816 -50530
rect 58516 -51660 58796 -51590
rect 58516 -51860 58556 -51660
rect 58556 -51860 58756 -51660
rect 58756 -51860 58796 -51660
rect 58516 -51940 58796 -51860
rect 61446 -51970 61686 -51860
rect 61446 -52100 61496 -51970
rect 61496 -52100 61686 -51970
rect 56628 -52868 57026 -52822
rect 56628 -53086 56654 -52868
rect 56654 -53086 56998 -52868
rect 56998 -53086 57026 -52868
rect 58486 -52890 58816 -52530
rect 56628 -53126 57026 -53086
rect 77170 -39040 77430 -38790
rect 84960 -38480 85400 -38050
rect 88150 -38820 88590 -38390
rect 79410 -40390 79680 -40150
rect 79410 -41620 79680 -41380
rect 79410 -42880 79680 -42640
rect 79410 -44100 79680 -43860
rect 81140 -40510 81570 -40250
rect 82820 -43310 91410 -42740
rect 79410 -45360 79680 -45120
rect 77170 -47080 77430 -46830
rect 79410 -48430 79680 -48190
rect 82824 -47448 91414 -46878
rect 79410 -49660 79680 -49420
rect 79410 -50920 79680 -50680
rect 79410 -52140 79680 -51900
rect 82820 -51100 91410 -50530
rect 79410 -53400 79680 -53160
rect 56506 -55830 57016 -55580
rect 58486 -56290 58816 -55930
rect 58516 -57060 58796 -56990
rect 58516 -57260 58556 -57060
rect 58556 -57260 58756 -57060
rect 58756 -57260 58796 -57060
rect 58516 -57340 58796 -57260
rect 61446 -57370 61686 -57260
rect 61446 -57500 61496 -57370
rect 61496 -57500 61686 -57370
rect 56628 -58268 57026 -58222
rect 56628 -58486 56654 -58268
rect 56654 -58486 56998 -58268
rect 56998 -58486 57026 -58268
rect 58486 -58290 58816 -57930
rect 56628 -58526 57026 -58486
rect 56506 -61230 57016 -60980
rect 58486 -61690 58816 -61330
rect 58516 -62460 58796 -62390
rect 58516 -62660 58556 -62460
rect 58556 -62660 58756 -62460
rect 58756 -62660 58796 -62460
rect 58516 -62740 58796 -62660
rect 61446 -62770 61686 -62660
rect 61446 -62900 61496 -62770
rect 61496 -62900 61686 -62770
rect 56628 -63668 57026 -63622
rect 56628 -63886 56654 -63668
rect 56654 -63886 56998 -63668
rect 56998 -63886 57026 -63668
rect 58486 -63690 58816 -63330
rect 56628 -63926 57026 -63886
rect 56506 -66630 57016 -66380
rect 58486 -67090 58816 -66730
rect 58516 -67860 58796 -67790
rect 58516 -68060 58556 -67860
rect 58556 -68060 58756 -67860
rect 58756 -68060 58796 -67860
rect 58516 -68140 58796 -68060
rect 61446 -68170 61686 -68060
rect 61446 -68300 61496 -68170
rect 61496 -68300 61686 -68170
rect 56628 -69068 57026 -69022
rect 56628 -69286 56654 -69068
rect 56654 -69286 56998 -69068
rect 56998 -69286 57026 -69068
rect 58486 -69090 58816 -68730
rect 56628 -69326 57026 -69286
rect 56506 -72030 57016 -71780
rect 58486 -72490 58816 -72130
rect 58516 -73260 58796 -73190
rect 58516 -73460 58556 -73260
rect 58556 -73460 58756 -73260
rect 58756 -73460 58796 -73260
rect 58516 -73540 58796 -73460
rect 61446 -73570 61686 -73460
rect 61446 -73700 61496 -73570
rect 61496 -73700 61686 -73570
rect 56628 -74468 57026 -74422
rect 56628 -74686 56654 -74468
rect 56654 -74686 56998 -74468
rect 56998 -74686 57026 -74468
rect 58486 -74490 58816 -74130
rect 56628 -74726 57026 -74686
rect 56506 -77430 57016 -77180
rect 58486 -77890 58816 -77530
rect 58516 -78660 58796 -78590
rect 58516 -78860 58556 -78660
rect 58556 -78860 58756 -78660
rect 58756 -78860 58796 -78660
rect 58516 -78940 58796 -78860
rect 61446 -78970 61686 -78860
rect 61446 -79100 61496 -78970
rect 61496 -79100 61686 -78970
rect 56628 -79868 57026 -79822
rect 56628 -80086 56654 -79868
rect 56654 -80086 56998 -79868
rect 56998 -80086 57026 -79868
rect 58486 -79890 58816 -79530
rect 56628 -80126 57026 -80086
rect 56506 -82830 57016 -82580
rect 58486 -83290 58816 -82930
rect 58516 -84060 58796 -83990
rect 58516 -84260 58556 -84060
rect 58556 -84260 58756 -84060
rect 58756 -84260 58796 -84060
rect 58516 -84340 58796 -84260
rect 61446 -84370 61686 -84260
rect 61446 -84500 61496 -84370
rect 61496 -84500 61686 -84370
rect 56628 -85268 57026 -85222
rect 56628 -85486 56654 -85268
rect 56654 -85486 56998 -85268
rect 56998 -85486 57026 -85268
rect 58486 -85290 58816 -84930
rect 56628 -85526 57026 -85486
<< metal5 >>
rect 42800 2400 65600 2600
rect 42800 1000 43000 2400
rect 46400 1000 65600 2400
rect 42800 800 65600 1000
rect 42800 0 46600 200
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 42800 -1500 46600 -1400
rect 56476 -1500 58896 -1470
rect 42800 -1580 58900 -1500
rect 42800 -1830 56506 -1580
rect 57016 -1830 58900 -1580
rect 42800 -1930 58900 -1830
rect 42800 -2290 58486 -1930
rect 58816 -2290 58900 -1930
rect 42800 -2890 58900 -2290
rect 42800 -2990 61726 -2890
rect 42800 -3340 58516 -2990
rect 58796 -3260 61726 -2990
rect 58796 -3340 61446 -3260
rect 42800 -3500 61446 -3340
rect 61686 -3500 61726 -3260
rect 42800 -3580 61726 -3500
rect 42800 -3930 58900 -3580
rect 42800 -4222 58486 -3930
rect 42800 -4526 56628 -4222
rect 57026 -4290 58486 -4222
rect 58816 -4290 58900 -3930
rect 57026 -4526 58900 -4290
rect 42800 -4600 58900 -4526
rect 42800 -6400 53300 -4600
rect 56486 -4610 58886 -4600
rect 20800 -6600 53300 -6400
rect 20800 -7400 21000 -6600
rect 22000 -6900 53300 -6600
rect 56476 -6900 58896 -6870
rect 22000 -6980 58896 -6900
rect 22000 -7230 56506 -6980
rect 57016 -7230 58896 -6980
rect 22000 -7330 58896 -7230
rect 22000 -7400 58486 -7330
rect 20800 -7600 58486 -7400
rect 42700 -7690 58486 -7600
rect 58816 -7690 58896 -7330
rect 42700 -8290 58896 -7690
rect 42700 -8390 61726 -8290
rect 42700 -8740 58516 -8390
rect 58796 -8660 61726 -8390
rect 58796 -8740 61446 -8660
rect 42700 -8900 61446 -8740
rect 61686 -8900 61726 -8660
rect 42700 -8980 61726 -8900
rect 42700 -9330 58896 -8980
rect 42700 -9622 58486 -9330
rect 42700 -9926 56628 -9622
rect 57026 -9690 58486 -9622
rect 58816 -9690 58896 -9330
rect 57026 -9750 58896 -9690
rect 57026 -9926 58886 -9750
rect 42700 -10000 58886 -9926
rect 42800 -12300 53300 -10000
rect 56486 -10010 58886 -10000
rect 56476 -12300 58896 -12270
rect 42800 -12380 58900 -12300
rect 42800 -12630 56506 -12380
rect 57016 -12630 58900 -12380
rect 42800 -12730 58900 -12630
rect 42800 -13090 58486 -12730
rect 58816 -13090 58900 -12730
rect 42800 -13690 58900 -13090
rect 42800 -13790 61726 -13690
rect 42800 -14140 58516 -13790
rect 58796 -14060 61726 -13790
rect 58796 -14140 61446 -14060
rect 42800 -14300 61446 -14140
rect 61686 -14300 61726 -14060
rect 42800 -14380 61726 -14300
rect 42800 -14730 58900 -14380
rect 42800 -15022 58486 -14730
rect 42800 -15326 56628 -15022
rect 57026 -15090 58486 -15022
rect 58816 -15090 58900 -14730
rect 57026 -15326 58900 -15090
rect 42800 -15400 58900 -15326
rect 42800 -17700 53300 -15400
rect 56486 -15410 58886 -15400
rect 56476 -17700 58896 -17670
rect 42800 -17780 58900 -17700
rect 42800 -18030 56506 -17780
rect 57016 -18030 58900 -17780
rect 42800 -18130 58900 -18030
rect 42800 -18490 58486 -18130
rect 58816 -18490 58900 -18130
rect 42800 -19090 58900 -18490
rect 42800 -19190 61726 -19090
rect 42800 -19540 58516 -19190
rect 58796 -19460 61726 -19190
rect 58796 -19540 61446 -19460
rect 42800 -19700 61446 -19540
rect 61686 -19700 61726 -19460
rect 42800 -19780 61726 -19700
rect 42800 -20130 58900 -19780
rect 42800 -20422 58486 -20130
rect 42800 -20726 56628 -20422
rect 57026 -20490 58486 -20422
rect 58816 -20490 58900 -20130
rect 57026 -20726 58900 -20490
rect 42800 -20800 58900 -20726
rect 42800 -23100 53300 -20800
rect 56486 -20810 58886 -20800
rect 56476 -23100 58896 -23070
rect 42800 -23180 58900 -23100
rect 42800 -23430 56506 -23180
rect 57016 -23430 58900 -23180
rect 42800 -23530 58900 -23430
rect 42800 -23890 58486 -23530
rect 58816 -23890 58900 -23530
rect 42800 -24490 58900 -23890
rect 42800 -24590 61726 -24490
rect 42800 -24940 58516 -24590
rect 58796 -24860 61726 -24590
rect 58796 -24940 61446 -24860
rect 42800 -25100 61446 -24940
rect 61686 -25100 61726 -24860
rect 42800 -25180 61726 -25100
rect 42800 -25530 58900 -25180
rect 42800 -25822 58486 -25530
rect 42800 -26126 56628 -25822
rect 57026 -25890 58486 -25822
rect 58816 -25890 58900 -25530
rect 57026 -26126 58900 -25890
rect 42800 -26200 58900 -26126
rect 42800 -28500 53300 -26200
rect 56486 -26210 58886 -26200
rect 56476 -28500 58896 -28470
rect 42800 -28580 58900 -28500
rect 42800 -28830 56506 -28580
rect 57016 -28830 58900 -28580
rect 42800 -28930 58900 -28830
rect 42800 -29290 58486 -28930
rect 58816 -29290 58900 -28930
rect 42800 -29890 58900 -29290
rect 42800 -29990 61726 -29890
rect 42800 -30340 58516 -29990
rect 58796 -30260 61726 -29990
rect 58796 -30340 61446 -30260
rect 42800 -30500 61446 -30340
rect 61686 -30500 61726 -30260
rect 42800 -30580 61726 -30500
rect 42800 -30930 58900 -30580
rect 42800 -31222 58486 -30930
rect 42800 -31526 56628 -31222
rect 57026 -31290 58486 -31222
rect 58816 -31290 58900 -30930
rect 57026 -31526 58900 -31290
rect 42800 -31600 58900 -31526
rect 42800 -33900 53300 -31600
rect 56486 -31610 58886 -31600
rect 56476 -33900 58896 -33870
rect 42800 -33980 58900 -33900
rect 42800 -34230 56506 -33980
rect 57016 -34230 58900 -33980
rect 42800 -34330 58900 -34230
rect 42800 -34690 58486 -34330
rect 58816 -34690 58900 -34330
rect 42800 -35290 58900 -34690
rect 63200 -34000 65600 800
rect 63200 -34100 89600 -34000
rect 42800 -35390 61726 -35290
rect 42800 -35740 58516 -35390
rect 58796 -35660 61726 -35390
rect 58796 -35740 61446 -35660
rect 42800 -35900 61446 -35740
rect 61686 -35900 61726 -35660
rect 42800 -35980 61726 -35900
rect 63200 -35500 72000 -34100
rect 74000 -35500 89600 -34100
rect 63200 -35600 89600 -35500
rect 42800 -36330 58900 -35980
rect 42800 -36622 58486 -36330
rect 42800 -36926 56628 -36622
rect 57026 -36690 58486 -36622
rect 58816 -36690 58900 -36330
rect 57026 -36926 58900 -36690
rect 42800 -37000 58900 -36926
rect 42800 -39300 53300 -37000
rect 56486 -37010 58886 -37000
rect 56476 -39300 58896 -39270
rect 42800 -39380 58900 -39300
rect 42800 -39630 56506 -39380
rect 57016 -39630 58900 -39380
rect 42800 -39730 58900 -39630
rect 42800 -40090 58486 -39730
rect 58816 -40090 58900 -39730
rect 42800 -40690 58900 -40090
rect 42800 -40790 61726 -40690
rect 42800 -41140 58516 -40790
rect 58796 -41060 61726 -40790
rect 58796 -41140 61446 -41060
rect 42800 -41300 61446 -41140
rect 61686 -41300 61726 -41060
rect 42800 -41380 61726 -41300
rect 63200 -41000 65600 -35600
rect 79200 -38050 89600 -35600
rect 79200 -38480 84960 -38050
rect 85400 -38390 89600 -38050
rect 85400 -38480 88150 -38390
rect 79200 -38760 88150 -38480
rect 75500 -38790 88150 -38760
rect 75500 -39040 77170 -38790
rect 77430 -38820 88150 -38790
rect 88590 -38800 89600 -38390
rect 88590 -38820 89440 -38800
rect 77430 -39040 89440 -38820
rect 75500 -39080 89440 -39040
rect 79290 -39260 89440 -39080
rect 79290 -39890 80530 -39260
rect 79290 -40150 81600 -39890
rect 79290 -40390 79410 -40150
rect 79680 -40250 81600 -40150
rect 79680 -40390 81140 -40250
rect 79290 -40510 81140 -40390
rect 81570 -40510 81600 -40250
rect 79290 -40540 81600 -40510
rect 79290 -41000 80530 -40540
rect 42800 -41730 58900 -41380
rect 42800 -42022 58486 -41730
rect 42800 -42326 56628 -42022
rect 57026 -42090 58486 -42022
rect 58816 -42090 58900 -41730
rect 57026 -42326 58900 -42090
rect 42800 -42400 58900 -42326
rect 63200 -41792 69418 -41000
rect 72648 -41380 91400 -41000
rect 72648 -41620 79410 -41380
rect 79680 -41620 91400 -41380
rect 72648 -41792 91400 -41620
rect 42800 -44700 53300 -42400
rect 56486 -42410 58886 -42400
rect 63200 -42640 91400 -41792
rect 63200 -42800 79410 -42640
rect 56476 -44700 58896 -44670
rect 42800 -44780 58900 -44700
rect 42800 -45030 56506 -44780
rect 57016 -45030 58900 -44780
rect 42800 -45130 58900 -45030
rect 42800 -45490 58486 -45130
rect 58816 -45490 58900 -45130
rect 42800 -46090 58900 -45490
rect 63200 -45600 65600 -42800
rect 79290 -42880 79410 -42800
rect 79680 -42710 91400 -42640
rect 79680 -42740 91440 -42710
rect 79680 -42880 82820 -42740
rect 79290 -43310 82820 -42880
rect 91410 -43310 91440 -42740
rect 79290 -43340 91440 -43310
rect 79290 -43860 80530 -43340
rect 79290 -44100 79410 -43860
rect 79680 -44100 80530 -43860
rect 79290 -45120 80530 -44100
rect 79290 -45360 79410 -45120
rect 79680 -45360 80530 -45120
rect 79290 -45600 80530 -45360
rect 42800 -46190 61726 -46090
rect 42800 -46540 58516 -46190
rect 58796 -46460 61726 -46190
rect 58796 -46540 61446 -46460
rect 42800 -46700 61446 -46540
rect 61686 -46700 61726 -46460
rect 42800 -46780 61726 -46700
rect 42800 -47130 58900 -46780
rect 42800 -47422 58486 -47130
rect 42800 -47726 56628 -47422
rect 57026 -47490 58486 -47422
rect 58816 -47490 58900 -47130
rect 57026 -47726 58900 -47490
rect 42800 -47800 58900 -47726
rect 63200 -46830 91400 -45600
rect 63200 -47080 77170 -46830
rect 77430 -46840 91400 -46830
rect 77430 -46878 91450 -46840
rect 77430 -47080 82824 -46878
rect 63200 -47400 82824 -47080
rect 42800 -50100 53300 -47800
rect 56486 -47810 58886 -47800
rect 63200 -49600 65600 -47400
rect 79290 -47448 82824 -47400
rect 91414 -47448 91450 -46878
rect 79290 -47480 91450 -47448
rect 79290 -48190 80530 -47480
rect 79290 -48430 79410 -48190
rect 79680 -48430 80530 -48190
rect 79290 -49420 80530 -48430
rect 79290 -49600 79410 -49420
rect 56476 -50100 58896 -50070
rect 42800 -50180 58900 -50100
rect 42800 -50430 56506 -50180
rect 57016 -50430 58900 -50180
rect 42800 -50530 58900 -50430
rect 42800 -50890 58486 -50530
rect 58816 -50890 58900 -50530
rect 42800 -51490 58900 -50890
rect 63200 -50492 69234 -49600
rect 73098 -49660 79410 -49600
rect 79680 -49600 80530 -49420
rect 79680 -49660 91400 -49600
rect 73098 -50492 91400 -49660
rect 63200 -50500 91400 -50492
rect 63200 -50530 91440 -50500
rect 63200 -50680 82820 -50530
rect 63200 -50920 79410 -50680
rect 79680 -50920 82820 -50680
rect 63200 -51100 82820 -50920
rect 91410 -51100 91440 -50530
rect 63200 -51130 91440 -51100
rect 63200 -51400 91400 -51130
rect 42800 -51590 61726 -51490
rect 42800 -51940 58516 -51590
rect 58796 -51860 61726 -51590
rect 58796 -51940 61446 -51860
rect 42800 -52100 61446 -51940
rect 61686 -52100 61726 -51860
rect 42800 -52180 61726 -52100
rect 79290 -51900 80530 -51400
rect 79290 -52140 79410 -51900
rect 79680 -52140 80530 -51900
rect 42800 -52530 58900 -52180
rect 42800 -52822 58486 -52530
rect 42800 -53126 56628 -52822
rect 57026 -52890 58486 -52822
rect 58816 -52890 58900 -52530
rect 57026 -53126 58900 -52890
rect 42800 -53200 58900 -53126
rect 79290 -53160 80530 -52140
rect 42800 -55500 53300 -53200
rect 56486 -53210 58886 -53200
rect 79290 -53400 79410 -53160
rect 79680 -53400 80530 -53160
rect 79290 -53430 80530 -53400
rect 56476 -55500 58896 -55470
rect 42800 -55580 58900 -55500
rect 42800 -55830 56506 -55580
rect 57016 -55830 58900 -55580
rect 42800 -55930 58900 -55830
rect 42800 -56290 58486 -55930
rect 58816 -56290 58900 -55930
rect 42800 -56890 58900 -56290
rect 42800 -56990 61726 -56890
rect 42800 -57340 58516 -56990
rect 58796 -57260 61726 -56990
rect 58796 -57340 61446 -57260
rect 42800 -57500 61446 -57340
rect 61686 -57500 61726 -57260
rect 42800 -57580 61726 -57500
rect 42800 -57930 58900 -57580
rect 42800 -58222 58486 -57930
rect 42800 -58526 56628 -58222
rect 57026 -58290 58486 -58222
rect 58816 -58290 58900 -57930
rect 57026 -58526 58900 -58290
rect 42800 -58600 58900 -58526
rect 42800 -60900 53300 -58600
rect 56486 -58610 58886 -58600
rect 56476 -60900 58896 -60870
rect 42800 -60980 58900 -60900
rect 42800 -61230 56506 -60980
rect 57016 -61230 58900 -60980
rect 42800 -61330 58900 -61230
rect 42800 -61690 58486 -61330
rect 58816 -61690 58900 -61330
rect 42800 -62290 58900 -61690
rect 42800 -62390 61726 -62290
rect 42800 -62740 58516 -62390
rect 58796 -62660 61726 -62390
rect 58796 -62740 61446 -62660
rect 42800 -62900 61446 -62740
rect 61686 -62900 61726 -62660
rect 42800 -62980 61726 -62900
rect 42800 -63330 58900 -62980
rect 42800 -63622 58486 -63330
rect 42800 -63926 56628 -63622
rect 57026 -63690 58486 -63622
rect 58816 -63690 58900 -63330
rect 57026 -63926 58900 -63690
rect 42800 -64000 58900 -63926
rect 42800 -66300 53300 -64000
rect 56486 -64010 58886 -64000
rect 56476 -66300 58896 -66270
rect 42800 -66380 58900 -66300
rect 42800 -66630 56506 -66380
rect 57016 -66630 58900 -66380
rect 42800 -66730 58900 -66630
rect 42800 -67090 58486 -66730
rect 58816 -67090 58900 -66730
rect 42800 -67690 58900 -67090
rect 42800 -67790 61726 -67690
rect 42800 -68140 58516 -67790
rect 58796 -68060 61726 -67790
rect 58796 -68140 61446 -68060
rect 42800 -68300 61446 -68140
rect 61686 -68300 61726 -68060
rect 42800 -68380 61726 -68300
rect 42800 -68730 58900 -68380
rect 42800 -69022 58486 -68730
rect 42800 -69326 56628 -69022
rect 57026 -69090 58486 -69022
rect 58816 -69090 58900 -68730
rect 57026 -69326 58900 -69090
rect 42800 -69400 58900 -69326
rect 42800 -71700 53300 -69400
rect 56486 -69410 58886 -69400
rect 56476 -71700 58896 -71670
rect 42800 -71780 58900 -71700
rect 42800 -72030 56506 -71780
rect 57016 -72030 58900 -71780
rect 42800 -72130 58900 -72030
rect 42800 -72490 58486 -72130
rect 58816 -72490 58900 -72130
rect 42800 -73090 58900 -72490
rect 42800 -73190 61726 -73090
rect 42800 -73540 58516 -73190
rect 58796 -73460 61726 -73190
rect 58796 -73540 61446 -73460
rect 42800 -73700 61446 -73540
rect 61686 -73700 61726 -73460
rect 42800 -73780 61726 -73700
rect 42800 -74130 58900 -73780
rect 42800 -74422 58486 -74130
rect 42800 -74726 56628 -74422
rect 57026 -74490 58486 -74422
rect 58816 -74490 58900 -74130
rect 57026 -74726 58900 -74490
rect 42800 -74800 58900 -74726
rect 42800 -77100 53300 -74800
rect 56486 -74810 58886 -74800
rect 56476 -77100 58896 -77070
rect 42800 -77180 58900 -77100
rect 42800 -77430 56506 -77180
rect 57016 -77430 58900 -77180
rect 42800 -77520 58900 -77430
rect 42800 -78230 56224 -77520
rect 57194 -77530 58900 -77520
rect 57194 -77890 58486 -77530
rect 58816 -77890 58900 -77530
rect 57194 -78230 58900 -77890
rect 42800 -78490 58900 -78230
rect 42800 -78590 61726 -78490
rect 42800 -78940 58516 -78590
rect 58796 -78860 61726 -78590
rect 58796 -78940 61446 -78860
rect 42800 -79100 61446 -78940
rect 61686 -79100 61726 -78860
rect 42800 -79106 61726 -79100
rect 42800 -79798 56126 -79106
rect 57196 -79180 61726 -79106
rect 57196 -79530 58900 -79180
rect 57196 -79680 58486 -79530
rect 56486 -79798 58486 -79680
rect 42800 -79822 58486 -79798
rect 42800 -80126 56628 -79822
rect 57026 -79890 58486 -79822
rect 58816 -79890 58900 -79530
rect 57026 -80126 58900 -79890
rect 42800 -80200 58900 -80126
rect 42800 -82500 53300 -80200
rect 56486 -80210 58886 -80200
rect 56476 -82500 58896 -82470
rect 42800 -82580 58900 -82500
rect 42800 -82830 56506 -82580
rect 57016 -82830 58900 -82580
rect 42800 -82930 58900 -82830
rect 42800 -83000 58486 -82930
rect 42800 -83540 56342 -83000
rect 57110 -83290 58486 -83000
rect 58816 -83290 58900 -82930
rect 57110 -83540 58900 -83290
rect 42800 -83890 58900 -83540
rect 42800 -83990 61726 -83890
rect 42800 -84340 58516 -83990
rect 58796 -84260 61726 -83990
rect 58796 -84340 61446 -84260
rect 42800 -84500 61446 -84340
rect 61686 -84500 61726 -84260
rect 42800 -84580 61726 -84500
rect 42800 -84586 58900 -84580
rect 42800 -85078 56350 -84586
rect 57054 -84930 58900 -84586
rect 57054 -85078 58486 -84930
rect 42800 -85222 58486 -85078
rect 42800 -85526 56628 -85222
rect 57026 -85290 58486 -85222
rect 58816 -85290 58900 -84930
rect 57026 -85526 58900 -85290
rect 42800 -85600 58900 -85526
rect 56486 -85610 58886 -85600
<< labels >>
flabel metal1 12400 -29200 12600 -29000 0 FreeSans 256 0 0 0 VFS
port 0 nsew
flabel metal1 12400 -62800 12600 -62600 0 FreeSans 256 0 0 0 VL
port 9 nsew
flabel metal1 39700 600 39900 800 0 FreeSans 256 0 0 0 GND
port 8 nsew
flabel metal1 44600 400 44800 600 0 FreeSans 256 0 0 0 VDD
port 5 nsew
flabel metal1 52000 1100 52200 1300 0 FreeSans 256 0 0 0 VIN
port 6 nsew
flabel metal1 94000 -39800 94200 -39600 0 FreeSans 256 0 0 0 OUT3
port 1 nsew
flabel metal1 93800 -44400 94000 -44200 0 FreeSans 256 0 0 0 OUT2
port 2 nsew
flabel metal1 93800 -48400 94000 -48200 0 FreeSans 256 0 0 0 OUT1
port 3 nsew
flabel metal1 93800 -52200 94000 -52000 0 FreeSans 256 0 0 0 OUT0
port 4 nsew
flabel metal1 57920 1100 58120 1300 0 FreeSans 256 0 0 0 CLK
port 7 nsew
rlabel metal3 37700 -86700 55500 -86200 1 VV1
port 10 n
rlabel metal3 38800 -81400 55500 -80800 1 VV2
port 11 n
rlabel metal3 39800 -76000 55500 -75400 1 VV3
port 12 n
rlabel metal3 40700 -70600 55500 -70000 1 VV4
port 13 n
rlabel metal3 41600 -65200 55500 -64600 1 VV5
port 14 n
rlabel metal3 42500 -59800 55500 -59200 1 VV6
port 15 n
rlabel metal3 43400 -54400 55400 -53800 1 VV7
port 16 n
rlabel metal3 44300 -49000 55500 -48400 1 VV8
port 17 n
rlabel metal3 44300 -43600 55500 -43000 1 VV9
port 18 n
rlabel metal3 43100 -38200 55400 -37600 1 VV10
port 19 n
rlabel metal3 42100 -32800 55500 -32200 1 VV11
port 20 n
rlabel metal3 41000 -27400 55500 -26800 1 VV12
port 21 n
rlabel metal3 40000 -22000 55500 -21400 1 VV13
port 22 n
rlabel metal3 39000 -16600 55500 -16000 1 VV14
port 23 n
rlabel metal3 38100 -11200 55500 -10600 1 VV15
port 24 n
rlabel metal3 37000 -5700 55600 -5200 1 VV16
port 25 n
rlabel metal1 56374 -85082 57010 -84958 1 R0
port 26 n
flabel metal1 56592 -83258 57024 -83024 0 FreeSans 192 0 0 0 S0
port 27 n
rlabel metal1 56362 -79722 57006 -79558 1 R1
port 28 n
rlabel metal1 56580 -77892 57066 -77610 1 S1
port 29 n
rlabel metal3 68600 -39240 73080 -39060 1 I15
port 30 n
rlabel metal3 67400 -39740 73200 -39560 1 I14
port 31 n
rlabel metal3 66600 -40020 72399 -39839 1 I13
port 32 n
rlabel metal3 65400 -40480 73200 -40300 1 I12
port 33 n
rlabel metal3 64160 -40840 73200 -40660 1 I11
port 34 n
rlabel metal3 63300 -41300 73200 -41000 1 I10
port 35 n
rlabel metal3 62500 -41700 73100 -41500 1 I9
port 36 n
rlabel metal3 60400 -43600 73200 -42600 1 I8
port 37 n
rlabel metal3 63203 -47499 73103 -47199 1 I7
port 38 n
rlabel metal3 64500 -47900 73100 -47600 1 I6
port 39 n
rlabel metal3 65400 -48300 73100 -48000 1 I5
port 40 n
rlabel metal3 66400 -48700 73100 -48400 1 I4
port 41 n
rlabel metal3 67400 -49100 73100 -48800 1 I3
port 42 n
rlabel metal3 68300 -49500 73100 -49200 1 I2
port 43 n
rlabel metal3 69300 -49900 73100 -49600 1 I1
port 44 n
rlabel metal3 70300 -50300 73100 -50000 1 I0
port 45 n
flabel metal1 36000 -56720 36200 -56520 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V1
flabel metal1 35990 -55110 36190 -54910 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V2
flabel metal1 36030 -53490 36230 -53290 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V3
flabel metal1 36050 -51920 36250 -51720 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V4
flabel metal1 36050 -50320 36250 -50120 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V5
flabel metal1 36010 -48740 36210 -48540 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V6
flabel metal1 36030 -47120 36230 -46920 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V7
flabel metal1 36020 -45540 36220 -45340 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V8
flabel metal1 36040 -43930 36240 -43730 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V9
flabel metal1 36060 -42330 36260 -42130 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V10
flabel metal1 36060 -40700 36260 -40500 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V11
flabel metal1 36030 -39130 36230 -38930 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V12
flabel metal1 36010 -37550 36210 -37350 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V13
flabel metal1 36040 -35920 36240 -35720 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V14
flabel metal1 36020 -34410 36220 -34210 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V15
flabel metal1 36060 -32740 36260 -32540 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.V16
flabel metal1 30740 -58750 30940 -58550 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.VL
flabel metal1 30820 -30870 31020 -30670 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.VFS
flabel metal1 25040 -44680 25240 -44480 0 FreeSans 256 0 0 0 resistorDivider_v0p0p1_0.GND
flabel metal1 57096 -55760 57296 -55560 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.VDD
flabel metal1 53056 -57750 53256 -57550 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.GND
flabel metal1 53586 -55740 53786 -55540 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.IB
flabel metal1 55576 -55240 55776 -55040 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.VIN
flabel metal1 55706 -59400 55906 -59200 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.VN
flabel metal1 57036 -57190 57236 -56990 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.CLK
flabel metal1 59956 -58910 60156 -58710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.Q
flabel metal1 56510 -55938 56710 -55738 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.VDD
flabel metal4 53070 -57188 53270 -56988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.VSS
flabel metal1 55580 -55238 55780 -55038 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.VIP
flabel metal1 56800 -56468 57000 -56268 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.VOP
flabel metal1 56800 -57958 57000 -57758 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.VON
flabel metal1 56860 -57188 57060 -56988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.CLK
flabel metal1 55710 -59398 55910 -59198 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.VIN
flabel metal1 53590 -55718 53790 -55518 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.class_AB_v3_sym_0.IB
flabel metal1 57127 -56623 57161 -56589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.VGND
flabel metal1 57125 -56079 57159 -56045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.VPWR
flabel locali 57125 -56079 57159 -56045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.VPWR
flabel locali 57127 -56623 57161 -56589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.VGND
flabel locali 57307 -56521 57341 -56487 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.X
flabel locali 57307 -56249 57341 -56215 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.X
flabel locali 57307 -56181 57341 -56147 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.X
flabel locali 57125 -56385 57159 -56351 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.A
flabel nwell 57125 -56079 57159 -56045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.VPB
flabel pwell 57127 -56623 57161 -56589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x65.VNB
rlabel comment 57096 -56606 57096 -56606 4 frontAnalog_v0p0p1_10.x65.buf_1
rlabel metal1 57096 -56654 57372 -56558 1 frontAnalog_v0p0p1_10.x65.VGND
rlabel metal1 57096 -56110 57372 -56014 1 frontAnalog_v0p0p1_10.x65.VPWR
flabel metal1 57127 -57599 57161 -57565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.VGND
flabel metal1 57125 -58143 57159 -58109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.VPWR
flabel locali 57125 -58143 57159 -58109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.VPWR
flabel locali 57127 -57599 57161 -57565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.VGND
flabel locali 57307 -57701 57341 -57667 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.X
flabel locali 57307 -57973 57341 -57939 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.X
flabel locali 57307 -58041 57341 -58007 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.X
flabel locali 57125 -57837 57159 -57803 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.A
flabel nwell 57125 -58143 57159 -58109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.VPB
flabel pwell 57127 -57599 57161 -57565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.x63.VNB
rlabel comment 57096 -57582 57096 -57582 2 frontAnalog_v0p0p1_10.x63.buf_1
rlabel metal1 57096 -57630 57372 -57534 5 frontAnalog_v0p0p1_10.x63.VGND
rlabel metal1 57096 -58174 57372 -58078 5 frontAnalog_v0p0p1_10.x63.VPWR
flabel metal1 58556 -57260 58756 -57060 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.VDD
flabel metal1 61166 -56710 61366 -56510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.GND
flabel metal1 58956 -58790 59156 -58590 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.R
flabel metal1 58946 -55650 59146 -55450 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.S
flabel metal1 59956 -58910 60156 -58710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.Q
flabel metal1 60186 -55680 60386 -55480 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.QN
flabel locali 60297 -57359 60331 -57325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y
flabel locali 60365 -57359 60399 -57325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y
flabel locali 60433 -57359 60467 -57325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y
flabel locali 60365 -56991 60399 -56957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.A
flabel locali 60365 -57083 60399 -57049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.A
flabel locali 60365 -57175 60399 -57141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.A
flabel locali 60365 -57267 60399 -57233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.A
flabel nwell 60671 -56991 60705 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.VPB
flabel pwell 60127 -56991 60161 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.VNB
flabel metal1 60671 -56991 60705 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.VPWR
flabel metal1 60127 -56991 60161 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.VGND
rlabel comment 60144 -56928 60144 -56928 6 frontAnalog_v0p0p1_10.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -57388 60192 -56928 3 frontAnalog_v0p0p1_10.RSfetsym_0.x1.VGND
rlabel metal1 60640 -57388 60736 -56928 3 frontAnalog_v0p0p1_10.RSfetsym_0.x1.VPWR
flabel locali 61121 -57359 61155 -57325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y
flabel locali 61053 -57359 61087 -57325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y
flabel locali 60985 -57359 61019 -57325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y
flabel locali 61053 -56991 61087 -56957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.A
flabel locali 61053 -57083 61087 -57049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.A
flabel locali 61053 -57175 61087 -57141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.A
flabel locali 61053 -57267 61087 -57233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.A
flabel nwell 60747 -56991 60781 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.VPB
flabel pwell 61291 -56991 61325 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.VNB
flabel metal1 60747 -56991 60781 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.VPWR
flabel metal1 61291 -56991 61325 -56957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.VGND
rlabel comment 61308 -56928 61308 -56928 4 frontAnalog_v0p0p1_10.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -57388 61356 -56928 7 frontAnalog_v0p0p1_10.RSfetsym_0.x2.VGND
rlabel metal1 60716 -57388 60812 -56928 7 frontAnalog_v0p0p1_10.RSfetsym_0.x2.VPWR
flabel metal1 57096 -61160 57296 -60960 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.VDD
flabel metal1 53056 -63150 53256 -62950 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.GND
flabel metal1 53586 -61140 53786 -60940 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.IB
flabel metal1 55576 -60640 55776 -60440 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.VIN
flabel metal1 55706 -64800 55906 -64600 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.VN
flabel metal1 57036 -62590 57236 -62390 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.CLK
flabel metal1 59956 -64310 60156 -64110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.Q
flabel metal1 56510 -61338 56710 -61138 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.VDD
flabel metal4 53070 -62588 53270 -62388 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.VSS
flabel metal1 55580 -60638 55780 -60438 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.VIP
flabel metal1 56800 -61868 57000 -61668 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.VOP
flabel metal1 56800 -63358 57000 -63158 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.VON
flabel metal1 56860 -62588 57060 -62388 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.CLK
flabel metal1 55710 -64798 55910 -64598 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.VIN
flabel metal1 53590 -61118 53790 -60918 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.class_AB_v3_sym_0.IB
flabel metal1 57127 -62023 57161 -61989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.VGND
flabel metal1 57125 -61479 57159 -61445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.VPWR
flabel locali 57125 -61479 57159 -61445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.VPWR
flabel locali 57127 -62023 57161 -61989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.VGND
flabel locali 57307 -61921 57341 -61887 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.X
flabel locali 57307 -61649 57341 -61615 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.X
flabel locali 57307 -61581 57341 -61547 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.X
flabel locali 57125 -61785 57159 -61751 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.A
flabel nwell 57125 -61479 57159 -61445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.VPB
flabel pwell 57127 -62023 57161 -61989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x65.VNB
rlabel comment 57096 -62006 57096 -62006 4 frontAnalog_v0p0p1_11.x65.buf_1
rlabel metal1 57096 -62054 57372 -61958 1 frontAnalog_v0p0p1_11.x65.VGND
rlabel metal1 57096 -61510 57372 -61414 1 frontAnalog_v0p0p1_11.x65.VPWR
flabel metal1 57127 -62999 57161 -62965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.VGND
flabel metal1 57125 -63543 57159 -63509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.VPWR
flabel locali 57125 -63543 57159 -63509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.VPWR
flabel locali 57127 -62999 57161 -62965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.VGND
flabel locali 57307 -63101 57341 -63067 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.X
flabel locali 57307 -63373 57341 -63339 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.X
flabel locali 57307 -63441 57341 -63407 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.X
flabel locali 57125 -63237 57159 -63203 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.A
flabel nwell 57125 -63543 57159 -63509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.VPB
flabel pwell 57127 -62999 57161 -62965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.x63.VNB
rlabel comment 57096 -62982 57096 -62982 2 frontAnalog_v0p0p1_11.x63.buf_1
rlabel metal1 57096 -63030 57372 -62934 5 frontAnalog_v0p0p1_11.x63.VGND
rlabel metal1 57096 -63574 57372 -63478 5 frontAnalog_v0p0p1_11.x63.VPWR
flabel metal1 58556 -62660 58756 -62460 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.VDD
flabel metal1 61166 -62110 61366 -61910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.GND
flabel metal1 58956 -64190 59156 -63990 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.R
flabel metal1 58946 -61050 59146 -60850 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.S
flabel metal1 59956 -64310 60156 -64110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.Q
flabel metal1 60186 -61080 60386 -60880 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.QN
flabel locali 60297 -62759 60331 -62725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y
flabel locali 60365 -62759 60399 -62725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y
flabel locali 60433 -62759 60467 -62725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y
flabel locali 60365 -62391 60399 -62357 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.A
flabel locali 60365 -62483 60399 -62449 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.A
flabel locali 60365 -62575 60399 -62541 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.A
flabel locali 60365 -62667 60399 -62633 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.A
flabel nwell 60671 -62391 60705 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.VPB
flabel pwell 60127 -62391 60161 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.VNB
flabel metal1 60671 -62391 60705 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.VPWR
flabel metal1 60127 -62391 60161 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.VGND
rlabel comment 60144 -62328 60144 -62328 6 frontAnalog_v0p0p1_11.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -62788 60192 -62328 3 frontAnalog_v0p0p1_11.RSfetsym_0.x1.VGND
rlabel metal1 60640 -62788 60736 -62328 3 frontAnalog_v0p0p1_11.RSfetsym_0.x1.VPWR
flabel locali 61121 -62759 61155 -62725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y
flabel locali 61053 -62759 61087 -62725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y
flabel locali 60985 -62759 61019 -62725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y
flabel locali 61053 -62391 61087 -62357 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.A
flabel locali 61053 -62483 61087 -62449 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.A
flabel locali 61053 -62575 61087 -62541 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.A
flabel locali 61053 -62667 61087 -62633 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.A
flabel nwell 60747 -62391 60781 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.VPB
flabel pwell 61291 -62391 61325 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.VNB
flabel metal1 60747 -62391 60781 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.VPWR
flabel metal1 61291 -62391 61325 -62357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.VGND
rlabel comment 61308 -62328 61308 -62328 4 frontAnalog_v0p0p1_11.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -62788 61356 -62328 7 frontAnalog_v0p0p1_11.RSfetsym_0.x2.VGND
rlabel metal1 60716 -62788 60812 -62328 7 frontAnalog_v0p0p1_11.RSfetsym_0.x2.VPWR
flabel metal1 57096 -71960 57296 -71760 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.VDD
flabel metal1 53056 -73950 53256 -73750 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.GND
flabel metal1 53586 -71940 53786 -71740 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.IB
flabel metal1 55576 -71440 55776 -71240 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.VIN
flabel metal1 55706 -75600 55906 -75400 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.VN
flabel metal1 57036 -73390 57236 -73190 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.CLK
flabel metal1 59956 -75110 60156 -74910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.Q
flabel metal1 56510 -72138 56710 -71938 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.VDD
flabel metal4 53070 -73388 53270 -73188 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.VSS
flabel metal1 55580 -71438 55780 -71238 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.VIP
flabel metal1 56800 -72668 57000 -72468 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.VOP
flabel metal1 56800 -74158 57000 -73958 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.VON
flabel metal1 56860 -73388 57060 -73188 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.CLK
flabel metal1 55710 -75598 55910 -75398 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.VIN
flabel metal1 53590 -71918 53790 -71718 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.class_AB_v3_sym_0.IB
flabel metal1 57127 -72823 57161 -72789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.VGND
flabel metal1 57125 -72279 57159 -72245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.VPWR
flabel locali 57125 -72279 57159 -72245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.VPWR
flabel locali 57127 -72823 57161 -72789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.VGND
flabel locali 57307 -72721 57341 -72687 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.X
flabel locali 57307 -72449 57341 -72415 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.X
flabel locali 57307 -72381 57341 -72347 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.X
flabel locali 57125 -72585 57159 -72551 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.A
flabel nwell 57125 -72279 57159 -72245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.VPB
flabel pwell 57127 -72823 57161 -72789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x65.VNB
rlabel comment 57096 -72806 57096 -72806 4 frontAnalog_v0p0p1_12.x65.buf_1
rlabel metal1 57096 -72854 57372 -72758 1 frontAnalog_v0p0p1_12.x65.VGND
rlabel metal1 57096 -72310 57372 -72214 1 frontAnalog_v0p0p1_12.x65.VPWR
flabel metal1 57127 -73799 57161 -73765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.VGND
flabel metal1 57125 -74343 57159 -74309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.VPWR
flabel locali 57125 -74343 57159 -74309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.VPWR
flabel locali 57127 -73799 57161 -73765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.VGND
flabel locali 57307 -73901 57341 -73867 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.X
flabel locali 57307 -74173 57341 -74139 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.X
flabel locali 57307 -74241 57341 -74207 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.X
flabel locali 57125 -74037 57159 -74003 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.A
flabel nwell 57125 -74343 57159 -74309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.VPB
flabel pwell 57127 -73799 57161 -73765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.x63.VNB
rlabel comment 57096 -73782 57096 -73782 2 frontAnalog_v0p0p1_12.x63.buf_1
rlabel metal1 57096 -73830 57372 -73734 5 frontAnalog_v0p0p1_12.x63.VGND
rlabel metal1 57096 -74374 57372 -74278 5 frontAnalog_v0p0p1_12.x63.VPWR
flabel metal1 58556 -73460 58756 -73260 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.VDD
flabel metal1 61166 -72910 61366 -72710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.GND
flabel metal1 58956 -74990 59156 -74790 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.R
flabel metal1 58946 -71850 59146 -71650 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.S
flabel metal1 59956 -75110 60156 -74910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.Q
flabel metal1 60186 -71880 60386 -71680 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.QN
flabel locali 60297 -73559 60331 -73525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y
flabel locali 60365 -73559 60399 -73525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y
flabel locali 60433 -73559 60467 -73525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y
flabel locali 60365 -73191 60399 -73157 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.A
flabel locali 60365 -73283 60399 -73249 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.A
flabel locali 60365 -73375 60399 -73341 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.A
flabel locali 60365 -73467 60399 -73433 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.A
flabel nwell 60671 -73191 60705 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.VPB
flabel pwell 60127 -73191 60161 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.VNB
flabel metal1 60671 -73191 60705 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.VPWR
flabel metal1 60127 -73191 60161 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x1.VGND
rlabel comment 60144 -73128 60144 -73128 6 frontAnalog_v0p0p1_12.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -73588 60192 -73128 3 frontAnalog_v0p0p1_12.RSfetsym_0.x1.VGND
rlabel metal1 60640 -73588 60736 -73128 3 frontAnalog_v0p0p1_12.RSfetsym_0.x1.VPWR
flabel locali 61121 -73559 61155 -73525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y
flabel locali 61053 -73559 61087 -73525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y
flabel locali 60985 -73559 61019 -73525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y
flabel locali 61053 -73191 61087 -73157 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.A
flabel locali 61053 -73283 61087 -73249 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.A
flabel locali 61053 -73375 61087 -73341 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.A
flabel locali 61053 -73467 61087 -73433 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.A
flabel nwell 60747 -73191 60781 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.VPB
flabel pwell 61291 -73191 61325 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.VNB
flabel metal1 60747 -73191 60781 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.VPWR
flabel metal1 61291 -73191 61325 -73157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_12.RSfetsym_0.x2.VGND
rlabel comment 61308 -73128 61308 -73128 4 frontAnalog_v0p0p1_12.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -73588 61356 -73128 7 frontAnalog_v0p0p1_12.RSfetsym_0.x2.VGND
rlabel metal1 60716 -73588 60812 -73128 7 frontAnalog_v0p0p1_12.RSfetsym_0.x2.VPWR
flabel metal1 57096 -66560 57296 -66360 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.VDD
flabel metal1 53056 -68550 53256 -68350 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.GND
flabel metal1 53586 -66540 53786 -66340 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.IB
flabel metal1 55576 -66040 55776 -65840 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.VIN
flabel metal1 55706 -70200 55906 -70000 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.VN
flabel metal1 57036 -67990 57236 -67790 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.CLK
flabel metal1 59956 -69710 60156 -69510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.Q
flabel metal1 56510 -66738 56710 -66538 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.VDD
flabel metal4 53070 -67988 53270 -67788 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.VSS
flabel metal1 55580 -66038 55780 -65838 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.VIP
flabel metal1 56800 -67268 57000 -67068 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.VOP
flabel metal1 56800 -68758 57000 -68558 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.VON
flabel metal1 56860 -67988 57060 -67788 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.CLK
flabel metal1 55710 -70198 55910 -69998 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.VIN
flabel metal1 53590 -66518 53790 -66318 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.class_AB_v3_sym_0.IB
flabel metal1 57127 -67423 57161 -67389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.VGND
flabel metal1 57125 -66879 57159 -66845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.VPWR
flabel locali 57125 -66879 57159 -66845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.VPWR
flabel locali 57127 -67423 57161 -67389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.VGND
flabel locali 57307 -67321 57341 -67287 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.X
flabel locali 57307 -67049 57341 -67015 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.X
flabel locali 57307 -66981 57341 -66947 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.X
flabel locali 57125 -67185 57159 -67151 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.A
flabel nwell 57125 -66879 57159 -66845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.VPB
flabel pwell 57127 -67423 57161 -67389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x65.VNB
rlabel comment 57096 -67406 57096 -67406 4 frontAnalog_v0p0p1_13.x65.buf_1
rlabel metal1 57096 -67454 57372 -67358 1 frontAnalog_v0p0p1_13.x65.VGND
rlabel metal1 57096 -66910 57372 -66814 1 frontAnalog_v0p0p1_13.x65.VPWR
flabel metal1 57127 -68399 57161 -68365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.VGND
flabel metal1 57125 -68943 57159 -68909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.VPWR
flabel locali 57125 -68943 57159 -68909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.VPWR
flabel locali 57127 -68399 57161 -68365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.VGND
flabel locali 57307 -68501 57341 -68467 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.X
flabel locali 57307 -68773 57341 -68739 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.X
flabel locali 57307 -68841 57341 -68807 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.X
flabel locali 57125 -68637 57159 -68603 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.A
flabel nwell 57125 -68943 57159 -68909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.VPB
flabel pwell 57127 -68399 57161 -68365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.x63.VNB
rlabel comment 57096 -68382 57096 -68382 2 frontAnalog_v0p0p1_13.x63.buf_1
rlabel metal1 57096 -68430 57372 -68334 5 frontAnalog_v0p0p1_13.x63.VGND
rlabel metal1 57096 -68974 57372 -68878 5 frontAnalog_v0p0p1_13.x63.VPWR
flabel metal1 58556 -68060 58756 -67860 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.VDD
flabel metal1 61166 -67510 61366 -67310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.GND
flabel metal1 58956 -69590 59156 -69390 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.R
flabel metal1 58946 -66450 59146 -66250 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.S
flabel metal1 59956 -69710 60156 -69510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.Q
flabel metal1 60186 -66480 60386 -66280 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.QN
flabel locali 60297 -68159 60331 -68125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y
flabel locali 60365 -68159 60399 -68125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y
flabel locali 60433 -68159 60467 -68125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y
flabel locali 60365 -67791 60399 -67757 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.A
flabel locali 60365 -67883 60399 -67849 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.A
flabel locali 60365 -67975 60399 -67941 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.A
flabel locali 60365 -68067 60399 -68033 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.A
flabel nwell 60671 -67791 60705 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.VPB
flabel pwell 60127 -67791 60161 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.VNB
flabel metal1 60671 -67791 60705 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.VPWR
flabel metal1 60127 -67791 60161 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.VGND
rlabel comment 60144 -67728 60144 -67728 6 frontAnalog_v0p0p1_13.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -68188 60192 -67728 3 frontAnalog_v0p0p1_13.RSfetsym_0.x1.VGND
rlabel metal1 60640 -68188 60736 -67728 3 frontAnalog_v0p0p1_13.RSfetsym_0.x1.VPWR
flabel locali 61121 -68159 61155 -68125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y
flabel locali 61053 -68159 61087 -68125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y
flabel locali 60985 -68159 61019 -68125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y
flabel locali 61053 -67791 61087 -67757 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.A
flabel locali 61053 -67883 61087 -67849 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.A
flabel locali 61053 -67975 61087 -67941 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.A
flabel locali 61053 -68067 61087 -68033 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.A
flabel nwell 60747 -67791 60781 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.VPB
flabel pwell 61291 -67791 61325 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.VNB
flabel metal1 60747 -67791 60781 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.VPWR
flabel metal1 61291 -67791 61325 -67757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.VGND
rlabel comment 61308 -67728 61308 -67728 4 frontAnalog_v0p0p1_13.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -68188 61356 -67728 7 frontAnalog_v0p0p1_13.RSfetsym_0.x2.VGND
rlabel metal1 60716 -68188 60812 -67728 7 frontAnalog_v0p0p1_13.RSfetsym_0.x2.VPWR
flabel metal1 57096 -77360 57296 -77160 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.VDD
flabel metal1 53056 -79350 53256 -79150 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.GND
flabel metal1 53586 -77340 53786 -77140 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.IB
flabel metal1 55576 -76840 55776 -76640 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.VIN
flabel metal1 55706 -81000 55906 -80800 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.VN
flabel metal1 57036 -78790 57236 -78590 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.CLK
flabel metal1 59956 -80510 60156 -80310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.Q
flabel metal1 56510 -77538 56710 -77338 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.VDD
flabel metal4 53070 -78788 53270 -78588 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.VSS
flabel metal1 55580 -76838 55780 -76638 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.VIP
flabel metal1 56800 -78068 57000 -77868 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.VOP
flabel metal1 56800 -79558 57000 -79358 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.VON
flabel metal1 56860 -78788 57060 -78588 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.CLK
flabel metal1 55710 -80998 55910 -80798 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.VIN
flabel metal1 53590 -77318 53790 -77118 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.class_AB_v3_sym_0.IB
flabel metal1 57127 -78223 57161 -78189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.VGND
flabel metal1 57125 -77679 57159 -77645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.VPWR
flabel locali 57125 -77679 57159 -77645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.VPWR
flabel locali 57127 -78223 57161 -78189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.VGND
flabel locali 57307 -78121 57341 -78087 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.X
flabel locali 57307 -77849 57341 -77815 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.X
flabel locali 57307 -77781 57341 -77747 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.X
flabel locali 57125 -77985 57159 -77951 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.A
flabel nwell 57125 -77679 57159 -77645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.VPB
flabel pwell 57127 -78223 57161 -78189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x65.VNB
rlabel comment 57096 -78206 57096 -78206 4 frontAnalog_v0p0p1_14.x65.buf_1
rlabel metal1 57096 -78254 57372 -78158 1 frontAnalog_v0p0p1_14.x65.VGND
rlabel metal1 57096 -77710 57372 -77614 1 frontAnalog_v0p0p1_14.x65.VPWR
flabel metal1 57127 -79199 57161 -79165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.VGND
flabel metal1 57125 -79743 57159 -79709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.VPWR
flabel locali 57125 -79743 57159 -79709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.VPWR
flabel locali 57127 -79199 57161 -79165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.VGND
flabel locali 57307 -79301 57341 -79267 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.X
flabel locali 57307 -79573 57341 -79539 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.X
flabel locali 57307 -79641 57341 -79607 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.X
flabel locali 57125 -79437 57159 -79403 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.A
flabel nwell 57125 -79743 57159 -79709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.VPB
flabel pwell 57127 -79199 57161 -79165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.x63.VNB
rlabel comment 57096 -79182 57096 -79182 2 frontAnalog_v0p0p1_14.x63.buf_1
rlabel metal1 57096 -79230 57372 -79134 5 frontAnalog_v0p0p1_14.x63.VGND
rlabel metal1 57096 -79774 57372 -79678 5 frontAnalog_v0p0p1_14.x63.VPWR
flabel metal1 58556 -78860 58756 -78660 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.VDD
flabel metal1 61166 -78310 61366 -78110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.GND
flabel metal1 58956 -80390 59156 -80190 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.R
flabel metal1 58946 -77250 59146 -77050 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.S
flabel metal1 59956 -80510 60156 -80310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.Q
flabel metal1 60186 -77280 60386 -77080 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.QN
flabel locali 60297 -78959 60331 -78925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y
flabel locali 60365 -78959 60399 -78925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y
flabel locali 60433 -78959 60467 -78925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y
flabel locali 60365 -78591 60399 -78557 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.A
flabel locali 60365 -78683 60399 -78649 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.A
flabel locali 60365 -78775 60399 -78741 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.A
flabel locali 60365 -78867 60399 -78833 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.A
flabel nwell 60671 -78591 60705 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.VPB
flabel pwell 60127 -78591 60161 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.VNB
flabel metal1 60671 -78591 60705 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.VPWR
flabel metal1 60127 -78591 60161 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.VGND
rlabel comment 60144 -78528 60144 -78528 6 frontAnalog_v0p0p1_14.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -78988 60192 -78528 3 frontAnalog_v0p0p1_14.RSfetsym_0.x1.VGND
rlabel metal1 60640 -78988 60736 -78528 3 frontAnalog_v0p0p1_14.RSfetsym_0.x1.VPWR
flabel locali 61121 -78959 61155 -78925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y
flabel locali 61053 -78959 61087 -78925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y
flabel locali 60985 -78959 61019 -78925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y
flabel locali 61053 -78591 61087 -78557 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.A
flabel locali 61053 -78683 61087 -78649 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.A
flabel locali 61053 -78775 61087 -78741 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.A
flabel locali 61053 -78867 61087 -78833 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.A
flabel nwell 60747 -78591 60781 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.VPB
flabel pwell 61291 -78591 61325 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.VNB
flabel metal1 60747 -78591 60781 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.VPWR
flabel metal1 61291 -78591 61325 -78557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_14.RSfetsym_0.x2.VGND
rlabel comment 61308 -78528 61308 -78528 4 frontAnalog_v0p0p1_14.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -78988 61356 -78528 7 frontAnalog_v0p0p1_14.RSfetsym_0.x2.VGND
rlabel metal1 60716 -78988 60812 -78528 7 frontAnalog_v0p0p1_14.RSfetsym_0.x2.VPWR
flabel metal1 57096 -82760 57296 -82560 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.VDD
flabel metal1 53056 -84750 53256 -84550 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.GND
flabel metal1 53586 -82740 53786 -82540 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.IB
flabel metal1 55576 -82240 55776 -82040 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.VIN
flabel metal1 55706 -86400 55906 -86200 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.VN
flabel metal1 57036 -84190 57236 -83990 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.CLK
flabel metal1 59956 -85910 60156 -85710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.Q
flabel metal1 56510 -82938 56710 -82738 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.VDD
flabel metal4 53070 -84188 53270 -83988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.VSS
flabel metal1 55580 -82238 55780 -82038 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.VIP
flabel metal1 56800 -83468 57000 -83268 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.VOP
flabel metal1 56800 -84958 57000 -84758 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.VON
flabel metal1 56860 -84188 57060 -83988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.CLK
flabel metal1 55710 -86398 55910 -86198 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.VIN
flabel metal1 53590 -82718 53790 -82518 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.class_AB_v3_sym_0.IB
flabel metal1 57127 -83623 57161 -83589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.VGND
flabel metal1 57125 -83079 57159 -83045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.VPWR
flabel locali 57125 -83079 57159 -83045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.VPWR
flabel locali 57127 -83623 57161 -83589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.VGND
flabel locali 57307 -83521 57341 -83487 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.X
flabel locali 57307 -83249 57341 -83215 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.X
flabel locali 57307 -83181 57341 -83147 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.X
flabel locali 57125 -83385 57159 -83351 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.A
flabel nwell 57125 -83079 57159 -83045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.VPB
flabel pwell 57127 -83623 57161 -83589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x65.VNB
rlabel comment 57096 -83606 57096 -83606 4 frontAnalog_v0p0p1_15.x65.buf_1
rlabel metal1 57096 -83654 57372 -83558 1 frontAnalog_v0p0p1_15.x65.VGND
rlabel metal1 57096 -83110 57372 -83014 1 frontAnalog_v0p0p1_15.x65.VPWR
flabel metal1 57127 -84599 57161 -84565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.VGND
flabel metal1 57125 -85143 57159 -85109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.VPWR
flabel locali 57125 -85143 57159 -85109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.VPWR
flabel locali 57127 -84599 57161 -84565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.VGND
flabel locali 57307 -84701 57341 -84667 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.X
flabel locali 57307 -84973 57341 -84939 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.X
flabel locali 57307 -85041 57341 -85007 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.X
flabel locali 57125 -84837 57159 -84803 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.A
flabel nwell 57125 -85143 57159 -85109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.VPB
flabel pwell 57127 -84599 57161 -84565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.x63.VNB
rlabel comment 57096 -84582 57096 -84582 2 frontAnalog_v0p0p1_15.x63.buf_1
rlabel metal1 57096 -84630 57372 -84534 5 frontAnalog_v0p0p1_15.x63.VGND
rlabel metal1 57096 -85174 57372 -85078 5 frontAnalog_v0p0p1_15.x63.VPWR
flabel metal1 58556 -84260 58756 -84060 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.VDD
flabel metal1 61166 -83710 61366 -83510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.GND
flabel metal1 58956 -85790 59156 -85590 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.R
flabel metal1 58946 -82650 59146 -82450 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.S
flabel metal1 59956 -85910 60156 -85710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.Q
flabel metal1 60186 -82680 60386 -82480 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.QN
flabel locali 60297 -84359 60331 -84325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y
flabel locali 60365 -84359 60399 -84325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y
flabel locali 60433 -84359 60467 -84325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y
flabel locali 60365 -83991 60399 -83957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.A
flabel locali 60365 -84083 60399 -84049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.A
flabel locali 60365 -84175 60399 -84141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.A
flabel locali 60365 -84267 60399 -84233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.A
flabel nwell 60671 -83991 60705 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.VPB
flabel pwell 60127 -83991 60161 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.VNB
flabel metal1 60671 -83991 60705 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.VPWR
flabel metal1 60127 -83991 60161 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.VGND
rlabel comment 60144 -83928 60144 -83928 6 frontAnalog_v0p0p1_15.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -84388 60192 -83928 3 frontAnalog_v0p0p1_15.RSfetsym_0.x1.VGND
rlabel metal1 60640 -84388 60736 -83928 3 frontAnalog_v0p0p1_15.RSfetsym_0.x1.VPWR
flabel locali 61121 -84359 61155 -84325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y
flabel locali 61053 -84359 61087 -84325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y
flabel locali 60985 -84359 61019 -84325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y
flabel locali 61053 -83991 61087 -83957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.A
flabel locali 61053 -84083 61087 -84049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.A
flabel locali 61053 -84175 61087 -84141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.A
flabel locali 61053 -84267 61087 -84233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.A
flabel nwell 60747 -83991 60781 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.VPB
flabel pwell 61291 -83991 61325 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.VNB
flabel metal1 60747 -83991 60781 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.VPWR
flabel metal1 61291 -83991 61325 -83957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_15.RSfetsym_0.x2.VGND
rlabel comment 61308 -83928 61308 -83928 4 frontAnalog_v0p0p1_15.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -84388 61356 -83928 7 frontAnalog_v0p0p1_15.RSfetsym_0.x2.VGND
rlabel metal1 60716 -84388 60812 -83928 7 frontAnalog_v0p0p1_15.RSfetsym_0.x2.VPWR
flabel metal1 57096 -39560 57296 -39360 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.VDD
flabel metal1 53056 -41550 53256 -41350 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.GND
flabel metal1 53586 -39540 53786 -39340 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.IB
flabel metal1 55576 -39040 55776 -38840 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.VIN
flabel metal1 55706 -43200 55906 -43000 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.VN
flabel metal1 57036 -40990 57236 -40790 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.CLK
flabel metal1 59956 -42710 60156 -42510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.Q
flabel metal1 56510 -39738 56710 -39538 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.VDD
flabel metal4 53070 -40988 53270 -40788 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.VSS
flabel metal1 55580 -39038 55780 -38838 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.VIP
flabel metal1 56800 -40268 57000 -40068 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.VOP
flabel metal1 56800 -41758 57000 -41558 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.VON
flabel metal1 56860 -40988 57060 -40788 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.CLK
flabel metal1 55710 -43198 55910 -42998 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.VIN
flabel metal1 53590 -39518 53790 -39318 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.class_AB_v3_sym_0.IB
flabel metal1 57127 -40423 57161 -40389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.VGND
flabel metal1 57125 -39879 57159 -39845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.VPWR
flabel locali 57125 -39879 57159 -39845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.VPWR
flabel locali 57127 -40423 57161 -40389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.VGND
flabel locali 57307 -40321 57341 -40287 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.X
flabel locali 57307 -40049 57341 -40015 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.X
flabel locali 57307 -39981 57341 -39947 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.X
flabel locali 57125 -40185 57159 -40151 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.A
flabel nwell 57125 -39879 57159 -39845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.VPB
flabel pwell 57127 -40423 57161 -40389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x65.VNB
rlabel comment 57096 -40406 57096 -40406 4 frontAnalog_v0p0p1_1.x65.buf_1
rlabel metal1 57096 -40454 57372 -40358 1 frontAnalog_v0p0p1_1.x65.VGND
rlabel metal1 57096 -39910 57372 -39814 1 frontAnalog_v0p0p1_1.x65.VPWR
flabel metal1 57127 -41399 57161 -41365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.VGND
flabel metal1 57125 -41943 57159 -41909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.VPWR
flabel locali 57125 -41943 57159 -41909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.VPWR
flabel locali 57127 -41399 57161 -41365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.VGND
flabel locali 57307 -41501 57341 -41467 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.X
flabel locali 57307 -41773 57341 -41739 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.X
flabel locali 57307 -41841 57341 -41807 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.X
flabel locali 57125 -41637 57159 -41603 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.A
flabel nwell 57125 -41943 57159 -41909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.VPB
flabel pwell 57127 -41399 57161 -41365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.x63.VNB
rlabel comment 57096 -41382 57096 -41382 2 frontAnalog_v0p0p1_1.x63.buf_1
rlabel metal1 57096 -41430 57372 -41334 5 frontAnalog_v0p0p1_1.x63.VGND
rlabel metal1 57096 -41974 57372 -41878 5 frontAnalog_v0p0p1_1.x63.VPWR
flabel metal1 58556 -41060 58756 -40860 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.VDD
flabel metal1 61166 -40510 61366 -40310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.GND
flabel metal1 58956 -42590 59156 -42390 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.R
flabel metal1 58946 -39450 59146 -39250 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.S
flabel metal1 59956 -42710 60156 -42510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.Q
flabel metal1 60186 -39480 60386 -39280 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.QN
flabel locali 60297 -41159 60331 -41125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y
flabel locali 60365 -41159 60399 -41125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y
flabel locali 60433 -41159 60467 -41125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y
flabel locali 60365 -40791 60399 -40757 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.A
flabel locali 60365 -40883 60399 -40849 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.A
flabel locali 60365 -40975 60399 -40941 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.A
flabel locali 60365 -41067 60399 -41033 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.A
flabel nwell 60671 -40791 60705 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.VPB
flabel pwell 60127 -40791 60161 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.VNB
flabel metal1 60671 -40791 60705 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.VPWR
flabel metal1 60127 -40791 60161 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.VGND
rlabel comment 60144 -40728 60144 -40728 6 frontAnalog_v0p0p1_1.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -41188 60192 -40728 3 frontAnalog_v0p0p1_1.RSfetsym_0.x1.VGND
rlabel metal1 60640 -41188 60736 -40728 3 frontAnalog_v0p0p1_1.RSfetsym_0.x1.VPWR
flabel locali 61121 -41159 61155 -41125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y
flabel locali 61053 -41159 61087 -41125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y
flabel locali 60985 -41159 61019 -41125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y
flabel locali 61053 -40791 61087 -40757 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.A
flabel locali 61053 -40883 61087 -40849 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.A
flabel locali 61053 -40975 61087 -40941 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.A
flabel locali 61053 -41067 61087 -41033 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.A
flabel nwell 60747 -40791 60781 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.VPB
flabel pwell 61291 -40791 61325 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.VNB
flabel metal1 60747 -40791 60781 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.VPWR
flabel metal1 61291 -40791 61325 -40757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.VGND
rlabel comment 61308 -40728 61308 -40728 4 frontAnalog_v0p0p1_1.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -41188 61356 -40728 7 frontAnalog_v0p0p1_1.RSfetsym_0.x2.VGND
rlabel metal1 60716 -41188 60812 -40728 7 frontAnalog_v0p0p1_1.RSfetsym_0.x2.VPWR
flabel metal1 57096 -28760 57296 -28560 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.VDD
flabel metal1 53056 -30750 53256 -30550 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.GND
flabel metal1 53586 -28740 53786 -28540 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.IB
flabel metal1 55576 -28240 55776 -28040 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.VIN
flabel metal1 55706 -32400 55906 -32200 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.VN
flabel metal1 57036 -30190 57236 -29990 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.CLK
flabel metal1 59956 -31910 60156 -31710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.Q
flabel metal1 56510 -28938 56710 -28738 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.VDD
flabel metal4 53070 -30188 53270 -29988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.VSS
flabel metal1 55580 -28238 55780 -28038 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.VIP
flabel metal1 56800 -29468 57000 -29268 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.VOP
flabel metal1 56800 -30958 57000 -30758 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.VON
flabel metal1 56860 -30188 57060 -29988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.CLK
flabel metal1 55710 -32398 55910 -32198 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.VIN
flabel metal1 53590 -28718 53790 -28518 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.class_AB_v3_sym_0.IB
flabel metal1 57127 -29623 57161 -29589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.VGND
flabel metal1 57125 -29079 57159 -29045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.VPWR
flabel locali 57125 -29079 57159 -29045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.VPWR
flabel locali 57127 -29623 57161 -29589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.VGND
flabel locali 57307 -29521 57341 -29487 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.X
flabel locali 57307 -29249 57341 -29215 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.X
flabel locali 57307 -29181 57341 -29147 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.X
flabel locali 57125 -29385 57159 -29351 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.A
flabel nwell 57125 -29079 57159 -29045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.VPB
flabel pwell 57127 -29623 57161 -29589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x65.VNB
rlabel comment 57096 -29606 57096 -29606 4 frontAnalog_v0p0p1_6.x65.buf_1
rlabel metal1 57096 -29654 57372 -29558 1 frontAnalog_v0p0p1_6.x65.VGND
rlabel metal1 57096 -29110 57372 -29014 1 frontAnalog_v0p0p1_6.x65.VPWR
flabel metal1 57127 -30599 57161 -30565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.VGND
flabel metal1 57125 -31143 57159 -31109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.VPWR
flabel locali 57125 -31143 57159 -31109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.VPWR
flabel locali 57127 -30599 57161 -30565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.VGND
flabel locali 57307 -30701 57341 -30667 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.X
flabel locali 57307 -30973 57341 -30939 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.X
flabel locali 57307 -31041 57341 -31007 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.X
flabel locali 57125 -30837 57159 -30803 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.A
flabel nwell 57125 -31143 57159 -31109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.VPB
flabel pwell 57127 -30599 57161 -30565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.x63.VNB
rlabel comment 57096 -30582 57096 -30582 2 frontAnalog_v0p0p1_6.x63.buf_1
rlabel metal1 57096 -30630 57372 -30534 5 frontAnalog_v0p0p1_6.x63.VGND
rlabel metal1 57096 -31174 57372 -31078 5 frontAnalog_v0p0p1_6.x63.VPWR
flabel metal1 58556 -30260 58756 -30060 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.VDD
flabel metal1 61166 -29710 61366 -29510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.GND
flabel metal1 58956 -31790 59156 -31590 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.R
flabel metal1 58946 -28650 59146 -28450 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.S
flabel metal1 59956 -31910 60156 -31710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.Q
flabel metal1 60186 -28680 60386 -28480 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.QN
flabel locali 60297 -30359 60331 -30325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y
flabel locali 60365 -30359 60399 -30325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y
flabel locali 60433 -30359 60467 -30325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y
flabel locali 60365 -29991 60399 -29957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.A
flabel locali 60365 -30083 60399 -30049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.A
flabel locali 60365 -30175 60399 -30141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.A
flabel locali 60365 -30267 60399 -30233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.A
flabel nwell 60671 -29991 60705 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.VPB
flabel pwell 60127 -29991 60161 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.VNB
flabel metal1 60671 -29991 60705 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.VPWR
flabel metal1 60127 -29991 60161 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x1.VGND
rlabel comment 60144 -29928 60144 -29928 6 frontAnalog_v0p0p1_6.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -30388 60192 -29928 3 frontAnalog_v0p0p1_6.RSfetsym_0.x1.VGND
rlabel metal1 60640 -30388 60736 -29928 3 frontAnalog_v0p0p1_6.RSfetsym_0.x1.VPWR
flabel locali 61121 -30359 61155 -30325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y
flabel locali 61053 -30359 61087 -30325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y
flabel locali 60985 -30359 61019 -30325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y
flabel locali 61053 -29991 61087 -29957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.A
flabel locali 61053 -30083 61087 -30049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.A
flabel locali 61053 -30175 61087 -30141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.A
flabel locali 61053 -30267 61087 -30233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.A
flabel nwell 60747 -29991 60781 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.VPB
flabel pwell 61291 -29991 61325 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.VNB
flabel metal1 60747 -29991 60781 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.VPWR
flabel metal1 61291 -29991 61325 -29957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_6.RSfetsym_0.x2.VGND
rlabel comment 61308 -29928 61308 -29928 4 frontAnalog_v0p0p1_6.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -30388 61356 -29928 7 frontAnalog_v0p0p1_6.RSfetsym_0.x2.VGND
rlabel metal1 60716 -30388 60812 -29928 7 frontAnalog_v0p0p1_6.RSfetsym_0.x2.VPWR
flabel metal1 57096 -34160 57296 -33960 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.VDD
flabel metal1 53056 -36150 53256 -35950 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.GND
flabel metal1 53586 -34140 53786 -33940 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.IB
flabel metal1 55576 -33640 55776 -33440 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.VIN
flabel metal1 55706 -37800 55906 -37600 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.VN
flabel metal1 57036 -35590 57236 -35390 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.CLK
flabel metal1 59956 -37310 60156 -37110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.Q
flabel metal1 56510 -34338 56710 -34138 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.VDD
flabel metal4 53070 -35588 53270 -35388 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.VSS
flabel metal1 55580 -33638 55780 -33438 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.VIP
flabel metal1 56800 -34868 57000 -34668 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.VOP
flabel metal1 56800 -36358 57000 -36158 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.VON
flabel metal1 56860 -35588 57060 -35388 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.CLK
flabel metal1 55710 -37798 55910 -37598 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.VIN
flabel metal1 53590 -34118 53790 -33918 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.class_AB_v3_sym_0.IB
flabel metal1 57127 -35023 57161 -34989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.VGND
flabel metal1 57125 -34479 57159 -34445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.VPWR
flabel locali 57125 -34479 57159 -34445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.VPWR
flabel locali 57127 -35023 57161 -34989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.VGND
flabel locali 57307 -34921 57341 -34887 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.X
flabel locali 57307 -34649 57341 -34615 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.X
flabel locali 57307 -34581 57341 -34547 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.X
flabel locali 57125 -34785 57159 -34751 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.A
flabel nwell 57125 -34479 57159 -34445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.VPB
flabel pwell 57127 -35023 57161 -34989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x65.VNB
rlabel comment 57096 -35006 57096 -35006 4 frontAnalog_v0p0p1_7.x65.buf_1
rlabel metal1 57096 -35054 57372 -34958 1 frontAnalog_v0p0p1_7.x65.VGND
rlabel metal1 57096 -34510 57372 -34414 1 frontAnalog_v0p0p1_7.x65.VPWR
flabel metal1 57127 -35999 57161 -35965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.VGND
flabel metal1 57125 -36543 57159 -36509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.VPWR
flabel locali 57125 -36543 57159 -36509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.VPWR
flabel locali 57127 -35999 57161 -35965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.VGND
flabel locali 57307 -36101 57341 -36067 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.X
flabel locali 57307 -36373 57341 -36339 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.X
flabel locali 57307 -36441 57341 -36407 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.X
flabel locali 57125 -36237 57159 -36203 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.A
flabel nwell 57125 -36543 57159 -36509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.VPB
flabel pwell 57127 -35999 57161 -35965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.x63.VNB
rlabel comment 57096 -35982 57096 -35982 2 frontAnalog_v0p0p1_7.x63.buf_1
rlabel metal1 57096 -36030 57372 -35934 5 frontAnalog_v0p0p1_7.x63.VGND
rlabel metal1 57096 -36574 57372 -36478 5 frontAnalog_v0p0p1_7.x63.VPWR
flabel metal1 58556 -35660 58756 -35460 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.VDD
flabel metal1 61166 -35110 61366 -34910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.GND
flabel metal1 58956 -37190 59156 -36990 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.R
flabel metal1 58946 -34050 59146 -33850 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.S
flabel metal1 59956 -37310 60156 -37110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.Q
flabel metal1 60186 -34080 60386 -33880 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.QN
flabel locali 60297 -35759 60331 -35725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y
flabel locali 60365 -35759 60399 -35725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y
flabel locali 60433 -35759 60467 -35725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y
flabel locali 60365 -35391 60399 -35357 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.A
flabel locali 60365 -35483 60399 -35449 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.A
flabel locali 60365 -35575 60399 -35541 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.A
flabel locali 60365 -35667 60399 -35633 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.A
flabel nwell 60671 -35391 60705 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.VPB
flabel pwell 60127 -35391 60161 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.VNB
flabel metal1 60671 -35391 60705 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.VPWR
flabel metal1 60127 -35391 60161 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.VGND
rlabel comment 60144 -35328 60144 -35328 6 frontAnalog_v0p0p1_7.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -35788 60192 -35328 3 frontAnalog_v0p0p1_7.RSfetsym_0.x1.VGND
rlabel metal1 60640 -35788 60736 -35328 3 frontAnalog_v0p0p1_7.RSfetsym_0.x1.VPWR
flabel locali 61121 -35759 61155 -35725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y
flabel locali 61053 -35759 61087 -35725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y
flabel locali 60985 -35759 61019 -35725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y
flabel locali 61053 -35391 61087 -35357 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.A
flabel locali 61053 -35483 61087 -35449 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.A
flabel locali 61053 -35575 61087 -35541 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.A
flabel locali 61053 -35667 61087 -35633 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.A
flabel nwell 60747 -35391 60781 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.VPB
flabel pwell 61291 -35391 61325 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.VNB
flabel metal1 60747 -35391 60781 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.VPWR
flabel metal1 61291 -35391 61325 -35357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_7.RSfetsym_0.x2.VGND
rlabel comment 61308 -35328 61308 -35328 4 frontAnalog_v0p0p1_7.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -35788 61356 -35328 7 frontAnalog_v0p0p1_7.RSfetsym_0.x2.VGND
rlabel metal1 60716 -35788 60812 -35328 7 frontAnalog_v0p0p1_7.RSfetsym_0.x2.VPWR
flabel metal1 57096 -44960 57296 -44760 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.VDD
flabel metal1 53056 -46950 53256 -46750 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.GND
flabel metal1 53586 -44940 53786 -44740 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.IB
flabel metal1 55576 -44440 55776 -44240 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.VIN
flabel metal1 55706 -48600 55906 -48400 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.VN
flabel metal1 57036 -46390 57236 -46190 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.CLK
flabel metal1 59956 -48110 60156 -47910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.Q
flabel metal1 56510 -45138 56710 -44938 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.VDD
flabel metal4 53070 -46388 53270 -46188 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.VSS
flabel metal1 55580 -44438 55780 -44238 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.VIP
flabel metal1 56800 -45668 57000 -45468 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.VOP
flabel metal1 56800 -47158 57000 -46958 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.VON
flabel metal1 56860 -46388 57060 -46188 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.CLK
flabel metal1 55710 -48598 55910 -48398 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.VIN
flabel metal1 53590 -44918 53790 -44718 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.class_AB_v3_sym_0.IB
flabel metal1 57127 -45823 57161 -45789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.VGND
flabel metal1 57125 -45279 57159 -45245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.VPWR
flabel locali 57125 -45279 57159 -45245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.VPWR
flabel locali 57127 -45823 57161 -45789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.VGND
flabel locali 57307 -45721 57341 -45687 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.X
flabel locali 57307 -45449 57341 -45415 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.X
flabel locali 57307 -45381 57341 -45347 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.X
flabel locali 57125 -45585 57159 -45551 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.A
flabel nwell 57125 -45279 57159 -45245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.VPB
flabel pwell 57127 -45823 57161 -45789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x65.VNB
rlabel comment 57096 -45806 57096 -45806 4 frontAnalog_v0p0p1_8.x65.buf_1
rlabel metal1 57096 -45854 57372 -45758 1 frontAnalog_v0p0p1_8.x65.VGND
rlabel metal1 57096 -45310 57372 -45214 1 frontAnalog_v0p0p1_8.x65.VPWR
flabel metal1 57127 -46799 57161 -46765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.VGND
flabel metal1 57125 -47343 57159 -47309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.VPWR
flabel locali 57125 -47343 57159 -47309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.VPWR
flabel locali 57127 -46799 57161 -46765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.VGND
flabel locali 57307 -46901 57341 -46867 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.X
flabel locali 57307 -47173 57341 -47139 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.X
flabel locali 57307 -47241 57341 -47207 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.X
flabel locali 57125 -47037 57159 -47003 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.A
flabel nwell 57125 -47343 57159 -47309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.VPB
flabel pwell 57127 -46799 57161 -46765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.x63.VNB
rlabel comment 57096 -46782 57096 -46782 2 frontAnalog_v0p0p1_8.x63.buf_1
rlabel metal1 57096 -46830 57372 -46734 5 frontAnalog_v0p0p1_8.x63.VGND
rlabel metal1 57096 -47374 57372 -47278 5 frontAnalog_v0p0p1_8.x63.VPWR
flabel metal1 58556 -46460 58756 -46260 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.VDD
flabel metal1 61166 -45910 61366 -45710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.GND
flabel metal1 58956 -47990 59156 -47790 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.R
flabel metal1 58946 -44850 59146 -44650 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.S
flabel metal1 59956 -48110 60156 -47910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.Q
flabel metal1 60186 -44880 60386 -44680 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.QN
flabel locali 60297 -46559 60331 -46525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y
flabel locali 60365 -46559 60399 -46525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y
flabel locali 60433 -46559 60467 -46525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y
flabel locali 60365 -46191 60399 -46157 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.A
flabel locali 60365 -46283 60399 -46249 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.A
flabel locali 60365 -46375 60399 -46341 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.A
flabel locali 60365 -46467 60399 -46433 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.A
flabel nwell 60671 -46191 60705 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.VPB
flabel pwell 60127 -46191 60161 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.VNB
flabel metal1 60671 -46191 60705 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.VPWR
flabel metal1 60127 -46191 60161 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.VGND
rlabel comment 60144 -46128 60144 -46128 6 frontAnalog_v0p0p1_8.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -46588 60192 -46128 3 frontAnalog_v0p0p1_8.RSfetsym_0.x1.VGND
rlabel metal1 60640 -46588 60736 -46128 3 frontAnalog_v0p0p1_8.RSfetsym_0.x1.VPWR
flabel locali 61121 -46559 61155 -46525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y
flabel locali 61053 -46559 61087 -46525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y
flabel locali 60985 -46559 61019 -46525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y
flabel locali 61053 -46191 61087 -46157 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.A
flabel locali 61053 -46283 61087 -46249 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.A
flabel locali 61053 -46375 61087 -46341 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.A
flabel locali 61053 -46467 61087 -46433 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.A
flabel nwell 60747 -46191 60781 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.VPB
flabel pwell 61291 -46191 61325 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.VNB
flabel metal1 60747 -46191 60781 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.VPWR
flabel metal1 61291 -46191 61325 -46157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_8.RSfetsym_0.x2.VGND
rlabel comment 61308 -46128 61308 -46128 4 frontAnalog_v0p0p1_8.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -46588 61356 -46128 7 frontAnalog_v0p0p1_8.RSfetsym_0.x2.VGND
rlabel metal1 60716 -46588 60812 -46128 7 frontAnalog_v0p0p1_8.RSfetsym_0.x2.VPWR
flabel metal1 57096 -50360 57296 -50160 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.VDD
flabel metal1 53056 -52350 53256 -52150 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.GND
flabel metal1 53586 -50340 53786 -50140 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.IB
flabel metal1 55576 -49840 55776 -49640 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.VIN
flabel metal1 55706 -54000 55906 -53800 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.VN
flabel metal1 57036 -51790 57236 -51590 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.CLK
flabel metal1 59956 -53510 60156 -53310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.Q
flabel metal1 56510 -50538 56710 -50338 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.VDD
flabel metal4 53070 -51788 53270 -51588 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.VSS
flabel metal1 55580 -49838 55780 -49638 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.VIP
flabel metal1 56800 -51068 57000 -50868 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.VOP
flabel metal1 56800 -52558 57000 -52358 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.VON
flabel metal1 56860 -51788 57060 -51588 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.CLK
flabel metal1 55710 -53998 55910 -53798 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.VIN
flabel metal1 53590 -50318 53790 -50118 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.class_AB_v3_sym_0.IB
flabel metal1 57127 -51223 57161 -51189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.VGND
flabel metal1 57125 -50679 57159 -50645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.VPWR
flabel locali 57125 -50679 57159 -50645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.VPWR
flabel locali 57127 -51223 57161 -51189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.VGND
flabel locali 57307 -51121 57341 -51087 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.X
flabel locali 57307 -50849 57341 -50815 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.X
flabel locali 57307 -50781 57341 -50747 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.X
flabel locali 57125 -50985 57159 -50951 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.A
flabel nwell 57125 -50679 57159 -50645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.VPB
flabel pwell 57127 -51223 57161 -51189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x65.VNB
rlabel comment 57096 -51206 57096 -51206 4 frontAnalog_v0p0p1_9.x65.buf_1
rlabel metal1 57096 -51254 57372 -51158 1 frontAnalog_v0p0p1_9.x65.VGND
rlabel metal1 57096 -50710 57372 -50614 1 frontAnalog_v0p0p1_9.x65.VPWR
flabel metal1 57127 -52199 57161 -52165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.VGND
flabel metal1 57125 -52743 57159 -52709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.VPWR
flabel locali 57125 -52743 57159 -52709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.VPWR
flabel locali 57127 -52199 57161 -52165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.VGND
flabel locali 57307 -52301 57341 -52267 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.X
flabel locali 57307 -52573 57341 -52539 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.X
flabel locali 57307 -52641 57341 -52607 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.X
flabel locali 57125 -52437 57159 -52403 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.A
flabel nwell 57125 -52743 57159 -52709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.VPB
flabel pwell 57127 -52199 57161 -52165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.x63.VNB
rlabel comment 57096 -52182 57096 -52182 2 frontAnalog_v0p0p1_9.x63.buf_1
rlabel metal1 57096 -52230 57372 -52134 5 frontAnalog_v0p0p1_9.x63.VGND
rlabel metal1 57096 -52774 57372 -52678 5 frontAnalog_v0p0p1_9.x63.VPWR
flabel metal1 58556 -51860 58756 -51660 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.VDD
flabel metal1 61166 -51310 61366 -51110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.GND
flabel metal1 58956 -53390 59156 -53190 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.R
flabel metal1 58946 -50250 59146 -50050 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.S
flabel metal1 59956 -53510 60156 -53310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.Q
flabel metal1 60186 -50280 60386 -50080 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.QN
flabel locali 60297 -51959 60331 -51925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y
flabel locali 60365 -51959 60399 -51925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y
flabel locali 60433 -51959 60467 -51925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y
flabel locali 60365 -51591 60399 -51557 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.A
flabel locali 60365 -51683 60399 -51649 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.A
flabel locali 60365 -51775 60399 -51741 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.A
flabel locali 60365 -51867 60399 -51833 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.A
flabel nwell 60671 -51591 60705 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.VPB
flabel pwell 60127 -51591 60161 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.VNB
flabel metal1 60671 -51591 60705 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.VPWR
flabel metal1 60127 -51591 60161 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.VGND
rlabel comment 60144 -51528 60144 -51528 6 frontAnalog_v0p0p1_9.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -51988 60192 -51528 3 frontAnalog_v0p0p1_9.RSfetsym_0.x1.VGND
rlabel metal1 60640 -51988 60736 -51528 3 frontAnalog_v0p0p1_9.RSfetsym_0.x1.VPWR
flabel locali 61121 -51959 61155 -51925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y
flabel locali 61053 -51959 61087 -51925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y
flabel locali 60985 -51959 61019 -51925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y
flabel locali 61053 -51591 61087 -51557 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.A
flabel locali 61053 -51683 61087 -51649 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.A
flabel locali 61053 -51775 61087 -51741 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.A
flabel locali 61053 -51867 61087 -51833 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.A
flabel nwell 60747 -51591 60781 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.VPB
flabel pwell 61291 -51591 61325 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.VNB
flabel metal1 60747 -51591 60781 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.VPWR
flabel metal1 61291 -51591 61325 -51557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.VGND
rlabel comment 61308 -51528 61308 -51528 4 frontAnalog_v0p0p1_9.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -51988 61356 -51528 7 frontAnalog_v0p0p1_9.RSfetsym_0.x2.VGND
rlabel metal1 60716 -51988 60812 -51528 7 frontAnalog_v0p0p1_9.RSfetsym_0.x2.VPWR
flabel metal1 72610 -39260 72810 -39060 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I15
flabel metal1 72610 -38930 72810 -38730 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.EI
flabel metal1 72610 -39750 72810 -39550 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I14
flabel metal1 72610 -40030 72810 -39830 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I13
flabel metal1 72610 -40490 72810 -40290 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I12
flabel metal1 72610 -40850 72810 -40650 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I11
flabel metal1 72610 -41250 72810 -41050 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I10
flabel metal1 72610 -41700 72810 -41500 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I9
flabel metal1 72610 -42070 72810 -41870 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I8
flabel metal1 72610 -50230 72810 -50030 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I0
flabel metal1 72600 -49860 72800 -49660 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I1
flabel metal1 72600 -49410 72800 -49210 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I2
flabel metal1 72600 -49010 72800 -48810 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I3
flabel metal1 72600 -48650 72800 -48450 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I4
flabel metal1 72600 -48190 72800 -47990 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I5
flabel metal1 72600 -47910 72800 -47710 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I6
flabel metal1 72600 -47420 72800 -47220 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.I7
flabel metal1 92160 -44390 92360 -44190 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.A2
flabel metal1 92160 -39860 92360 -39660 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.A3
flabel metal1 92160 -48540 92360 -48340 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.A1
flabel metal1 92160 -52150 92360 -51950 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.A0
flabel metal5 79290 -53430 80530 -37780 0 FreeSans 512 0 0 0 16to4_PriorityEncoder_v0p0p1_0.VDD
flabel metal4 76270 -53800 77080 -37780 1 FreeSans 512 0 0 0 16to4_PriorityEncoder_v0p0p1_0.GND
flabel metal1 73180 -46380 73380 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I0
flabel metal1 73430 -46380 73630 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I1
flabel metal1 73680 -46380 73880 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I2
flabel metal1 73930 -46380 74130 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I3
flabel metal1 74180 -46380 74380 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I4
flabel metal1 74430 -46380 74630 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I5
flabel metal1 74680 -46380 74880 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I6
flabel metal1 74930 -46380 75130 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.I7
flabel metal1 75180 -46380 75380 -46180 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.EI
flabel metal1 80460 -48020 80660 -47820 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.EO
flabel metal1 80460 -47570 80660 -47370 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.GS
flabel metal1 80460 -49240 80660 -49040 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.A2
flabel metal1 80390 -51230 80590 -51030 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.A1
flabel metal1 80390 -53770 80590 -53570 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.A0
flabel metal5 79380 -48190 79710 -46170 0 FreeSans 512 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.VDD
flabel metal4 76900 -53680 77080 -52650 0 FreeSans 512 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.GND
flabel locali 78159 -53147 78193 -53113 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X
flabel locali 77883 -52807 77917 -52773 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C
flabel locali 77883 -52875 77917 -52841 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C
flabel locali 77607 -52943 77641 -52909 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.A
flabel locali 77883 -52943 77917 -52909 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C
flabel locali 77791 -52807 77825 -52773 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.B
flabel locali 77791 -52875 77825 -52841 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.B
flabel locali 77975 -52943 78009 -52909 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D
flabel locali 78159 -52807 78193 -52773 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X
flabel locali 78159 -52875 78193 -52841 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X
flabel locali 78159 -52943 78193 -52909 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X
flabel locali 78159 -53011 78193 -52977 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X
flabel locali 78159 -53079 78193 -53045 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X
flabel metal1 77607 -52705 77641 -52671 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.VGND
flabel metal1 77607 -53249 77641 -53215 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.VPWR
flabel nwell 77607 -53249 77641 -53215 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.VPB
flabel pwell 77607 -52705 77641 -52671 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.VNB
rlabel comment 77578 -52688 77578 -52688 2 16to4_PriorityEncoder_v0p0p1_0.x3.x19.and4_1
rlabel metal1 77578 -52736 78222 -52640 5 16to4_PriorityEncoder_v0p0p1_0.x3.x19.VGND
rlabel metal1 77578 -53280 78222 -53184 5 16to4_PriorityEncoder_v0p0p1_0.x3.x19.VPWR
flabel metal1 77607 -53869 77641 -53835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.VGND
flabel metal1 77607 -53325 77641 -53291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.VPWR
flabel locali 77975 -53427 78009 -53393 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X
flabel locali 77975 -53767 78009 -53733 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X
flabel locali 77791 -53427 77825 -53393 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B
flabel locali 77607 -53699 77641 -53665 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.A
flabel locali 77813 -53699 77847 -53665 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.C
flabel nwell 77607 -53325 77641 -53291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.VPB
flabel pwell 77607 -53869 77641 -53835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.VNB
rlabel comment 77578 -53852 77578 -53852 4 16to4_PriorityEncoder_v0p0p1_0.x3.x20.and3_1
rlabel metal1 77578 -53900 78038 -53804 1 16to4_PriorityEncoder_v0p0p1_0.x3.x20.VGND
rlabel metal1 77578 -53356 78038 -53260 1 16to4_PriorityEncoder_v0p0p1_0.x3.x20.VPWR
flabel metal1 78067 -53325 78101 -53291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.VPWR
flabel metal1 78067 -53869 78101 -53835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.VGND
flabel locali 78435 -53699 78469 -53665 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X
flabel locali 78435 -53767 78469 -53733 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X
flabel locali 78435 -53631 78469 -53597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X
flabel locali 78435 -53563 78469 -53529 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X
flabel locali 78435 -53495 78469 -53461 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X
flabel locali 78435 -53427 78469 -53393 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X
flabel locali 78251 -53631 78285 -53597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B
flabel locali 78159 -53631 78193 -53597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.A
flabel locali 78067 -53631 78101 -53597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.A
flabel nwell 78067 -53325 78101 -53291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.VPB
flabel pwell 78067 -53869 78101 -53835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x21.VNB
rlabel comment 78038 -53852 78038 -53852 4 16to4_PriorityEncoder_v0p0p1_0.x3.x21.and2_1
rlabel metal1 78038 -53900 78498 -53804 1 16to4_PriorityEncoder_v0p0p1_0.x3.x21.VGND
rlabel metal1 78038 -53356 78498 -53260 1 16to4_PriorityEncoder_v0p0p1_0.x3.x21.VPWR
flabel locali 78712 -53631 78746 -53597 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C
flabel locali 78804 -53631 78838 -53597 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A
flabel locali 78988 -53495 79022 -53461 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.X
flabel locali 78620 -53631 78654 -53597 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C
flabel locali 78712 -53427 78746 -53393 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B
flabel locali 78620 -53427 78654 -53393 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B
flabel locali 78620 -53563 78654 -53529 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C
flabel locali 78528 -53427 78562 -53393 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B
flabel locali 78712 -53563 78746 -53529 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C
flabel locali 78528 -53631 78562 -53597 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D
flabel locali 78528 -53699 78562 -53665 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D
flabel metal1 78528 -53325 78562 -53291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.VPWR
flabel metal1 78528 -53869 78562 -53835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.VGND
flabel nwell 78528 -53325 78562 -53291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.VPB
flabel pwell 78528 -53869 78562 -53835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.VNB
rlabel comment 78498 -53852 78498 -53852 4 16to4_PriorityEncoder_v0p0p1_0.x3.x22.or4_1
rlabel metal1 78498 -53900 79050 -53804 1 16to4_PriorityEncoder_v0p0p1_0.x3.x22.VGND
rlabel metal1 78498 -53356 79050 -53260 1 16to4_PriorityEncoder_v0p0p1_0.x3.x22.VPWR
flabel locali 78159 -51913 78193 -51879 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X
flabel locali 77883 -51573 77917 -51539 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C
flabel locali 77883 -51641 77917 -51607 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C
flabel locali 77607 -51709 77641 -51675 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.A
flabel locali 77883 -51709 77917 -51675 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C
flabel locali 77791 -51573 77825 -51539 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.B
flabel locali 77791 -51641 77825 -51607 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.B
flabel locali 77975 -51709 78009 -51675 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.D
flabel locali 78159 -51573 78193 -51539 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X
flabel locali 78159 -51641 78193 -51607 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X
flabel locali 78159 -51709 78193 -51675 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X
flabel locali 78159 -51777 78193 -51743 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X
flabel locali 78159 -51845 78193 -51811 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X
flabel metal1 77607 -51471 77641 -51437 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.VGND
flabel metal1 77607 -52015 77641 -51981 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.VPWR
flabel nwell 77607 -52015 77641 -51981 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.VPB
flabel pwell 77607 -51471 77641 -51437 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x16.VNB
rlabel comment 77578 -51454 77578 -51454 2 16to4_PriorityEncoder_v0p0p1_0.x3.x16.and4_1
rlabel metal1 77578 -51502 78222 -51406 5 16to4_PriorityEncoder_v0p0p1_0.x3.x16.VGND
rlabel metal1 77578 -52046 78222 -51950 5 16to4_PriorityEncoder_v0p0p1_0.x3.x16.VPWR
flabel locali 78159 -52189 78193 -52155 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.X
flabel locali 77883 -52529 77917 -52495 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C
flabel locali 77883 -52461 77917 -52427 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C
flabel locali 77607 -52393 77641 -52359 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.A
flabel locali 77883 -52393 77917 -52359 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C
flabel locali 77791 -52529 77825 -52495 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.B
flabel locali 77791 -52461 77825 -52427 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.B
flabel locali 77975 -52393 78009 -52359 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.D
flabel locali 78159 -52529 78193 -52495 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.X
flabel locali 78159 -52461 78193 -52427 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.X
flabel locali 78159 -52393 78193 -52359 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.X
flabel locali 78159 -52325 78193 -52291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.X
flabel locali 78159 -52257 78193 -52223 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.X
flabel metal1 77607 -52631 77641 -52597 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.VGND
flabel metal1 77607 -52087 77641 -52053 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.VPWR
flabel nwell 77607 -52087 77641 -52053 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.VPB
flabel pwell 77607 -52631 77641 -52597 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x18.VNB
rlabel comment 77578 -52614 77578 -52614 4 16to4_PriorityEncoder_v0p0p1_0.x3.x18.and4_1
rlabel metal1 77578 -52662 78222 -52566 1 16to4_PriorityEncoder_v0p0p1_0.x3.x18.VGND
rlabel metal1 77578 -52118 78222 -52022 1 16to4_PriorityEncoder_v0p0p1_0.x3.x18.VPWR
flabel metal1 77609 -50783 77643 -50749 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.VPWR
flabel metal1 77609 -50239 77643 -50205 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.VGND
flabel locali 77977 -50409 78011 -50375 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.X
flabel locali 77977 -50341 78011 -50307 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.X
flabel locali 77977 -50477 78011 -50443 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.X
flabel locali 77977 -50545 78011 -50511 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.X
flabel locali 77977 -50613 78011 -50579 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.X
flabel locali 77977 -50681 78011 -50647 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.X
flabel locali 77793 -50477 77827 -50443 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.B
flabel locali 77701 -50477 77735 -50443 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.A
flabel locali 77609 -50477 77643 -50443 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.A
flabel nwell 77609 -50783 77643 -50749 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.VPB
flabel pwell 77609 -50239 77643 -50205 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x13.VNB
rlabel comment 77580 -50222 77580 -50222 2 16to4_PriorityEncoder_v0p0p1_0.x3.x13.and2_1
rlabel metal1 77580 -50270 78040 -50174 5 16to4_PriorityEncoder_v0p0p1_0.x3.x13.VGND
rlabel metal1 77580 -50814 78040 -50718 5 16to4_PriorityEncoder_v0p0p1_0.x3.x13.VPWR
flabel locali 78159 -50957 78193 -50923 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X
flabel locali 77883 -51297 77917 -51263 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.C
flabel locali 77883 -51229 77917 -51195 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.C
flabel locali 77607 -51161 77641 -51127 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.A
flabel locali 77883 -51161 77917 -51127 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.C
flabel locali 77791 -51297 77825 -51263 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.B
flabel locali 77791 -51229 77825 -51195 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.B
flabel locali 77975 -51161 78009 -51127 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.D
flabel locali 78159 -51297 78193 -51263 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X
flabel locali 78159 -51229 78193 -51195 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X
flabel locali 78159 -51161 78193 -51127 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X
flabel locali 78159 -51093 78193 -51059 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X
flabel locali 78159 -51025 78193 -50991 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X
flabel metal1 77607 -51399 77641 -51365 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.VGND
flabel metal1 77607 -50855 77641 -50821 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.VPWR
flabel nwell 77607 -50855 77641 -50821 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.VPB
flabel pwell 77607 -51399 77641 -51365 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x15.VNB
rlabel comment 77578 -51382 77578 -51382 4 16to4_PriorityEncoder_v0p0p1_0.x3.x15.and4_1
rlabel metal1 77578 -51430 78222 -51334 1 16to4_PriorityEncoder_v0p0p1_0.x3.x15.VGND
rlabel metal1 77578 -50886 78222 -50790 1 16to4_PriorityEncoder_v0p0p1_0.x3.x15.VPWR
flabel locali 78536 -51161 78570 -51127 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C
flabel locali 78628 -51161 78662 -51127 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A
flabel locali 78812 -51025 78846 -50991 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.X
flabel locali 78444 -51161 78478 -51127 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C
flabel locali 78536 -50957 78570 -50923 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.B
flabel locali 78444 -50957 78478 -50923 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.B
flabel locali 78444 -51093 78478 -51059 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C
flabel locali 78352 -50957 78386 -50923 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.B
flabel locali 78536 -51093 78570 -51059 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C
flabel locali 78352 -51161 78386 -51127 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D
flabel locali 78352 -51229 78386 -51195 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D
flabel metal1 78352 -50855 78386 -50821 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.VPWR
flabel metal1 78352 -51399 78386 -51365 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.VGND
flabel nwell 78352 -50855 78386 -50821 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.VPB
flabel pwell 78352 -51399 78386 -51365 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x17.VNB
rlabel comment 78322 -51382 78322 -51382 4 16to4_PriorityEncoder_v0p0p1_0.x3.x17.or4_1
rlabel metal1 78322 -51430 78874 -51334 1 16to4_PriorityEncoder_v0p0p1_0.x3.x17.VGND
rlabel metal1 78322 -50886 78874 -50790 1 16to4_PriorityEncoder_v0p0p1_0.x3.x17.VPWR
flabel metal1 77607 -49529 77641 -49495 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.VPWR
flabel metal1 77607 -48985 77641 -48951 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.VGND
flabel locali 77975 -49155 78009 -49121 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X
flabel locali 77975 -49087 78009 -49053 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X
flabel locali 77975 -49223 78009 -49189 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X
flabel locali 77975 -49291 78009 -49257 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X
flabel locali 77975 -49359 78009 -49325 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X
flabel locali 77975 -49427 78009 -49393 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X
flabel locali 77791 -49223 77825 -49189 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.B
flabel locali 77699 -49223 77733 -49189 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.A
flabel locali 77607 -49223 77641 -49189 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.A
flabel nwell 77607 -49529 77641 -49495 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.VPB
flabel pwell 77607 -48985 77641 -48951 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x11.VNB
rlabel comment 77578 -48968 77578 -48968 2 16to4_PriorityEncoder_v0p0p1_0.x3.x11.and2_1
rlabel metal1 77578 -49016 78038 -48920 5 16to4_PriorityEncoder_v0p0p1_0.x3.x11.VGND
rlabel metal1 77578 -49560 78038 -49464 5 16to4_PriorityEncoder_v0p0p1_0.x3.x11.VPWR
flabel metal1 77607 -49605 77641 -49571 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.VPWR
flabel metal1 77607 -50149 77641 -50115 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.VGND
flabel locali 77975 -49979 78009 -49945 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.X
flabel locali 77975 -50047 78009 -50013 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.X
flabel locali 77975 -49911 78009 -49877 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.X
flabel locali 77975 -49843 78009 -49809 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.X
flabel locali 77975 -49775 78009 -49741 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.X
flabel locali 77975 -49707 78009 -49673 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.X
flabel locali 77791 -49911 77825 -49877 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.B
flabel locali 77699 -49911 77733 -49877 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.A
flabel locali 77607 -49911 77641 -49877 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.A
flabel nwell 77607 -49605 77641 -49571 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.VPB
flabel pwell 77607 -50149 77641 -50115 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x12.VNB
rlabel comment 77578 -50132 77578 -50132 4 16to4_PriorityEncoder_v0p0p1_0.x3.x12.and2_1
rlabel metal1 77578 -50180 78038 -50084 1 16to4_PriorityEncoder_v0p0p1_0.x3.x12.VGND
rlabel metal1 77578 -49636 78038 -49540 1 16to4_PriorityEncoder_v0p0p1_0.x3.x12.VPWR
flabel locali 78252 -49223 78286 -49189 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.C
flabel locali 78344 -49223 78378 -49189 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A
flabel locali 78528 -49359 78562 -49325 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.X
flabel locali 78160 -49223 78194 -49189 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.C
flabel locali 78252 -49427 78286 -49393 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B
flabel locali 78160 -49427 78194 -49393 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B
flabel locali 78160 -49291 78194 -49257 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.C
flabel locali 78068 -49427 78102 -49393 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B
flabel locali 78252 -49291 78286 -49257 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.C
flabel locali 78068 -49223 78102 -49189 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.D
flabel locali 78068 -49155 78102 -49121 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.D
flabel metal1 78068 -49529 78102 -49495 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.VPWR
flabel metal1 78068 -48985 78102 -48951 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.VGND
flabel nwell 78068 -49529 78102 -49495 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.VPB
flabel pwell 78068 -48985 78102 -48951 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x14.VNB
rlabel comment 78038 -48968 78038 -48968 2 16to4_PriorityEncoder_v0p0p1_0.x3.x14.or4_1
rlabel metal1 78038 -49016 78590 -48920 5 16to4_PriorityEncoder_v0p0p1_0.x3.x14.VGND
rlabel metal1 78038 -49560 78590 -49464 5 16to4_PriorityEncoder_v0p0p1_0.x3.x14.VPWR
flabel metal1 77607 -48365 77641 -48331 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.VPWR
flabel metal1 77607 -48909 77641 -48875 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.VGND
flabel locali 77975 -48739 78009 -48705 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.X
flabel locali 77975 -48807 78009 -48773 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.X
flabel locali 77975 -48671 78009 -48637 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.X
flabel locali 77975 -48603 78009 -48569 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.X
flabel locali 77975 -48535 78009 -48501 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.X
flabel locali 77975 -48467 78009 -48433 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.X
flabel locali 77791 -48671 77825 -48637 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.B
flabel locali 77699 -48671 77733 -48637 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.A
flabel locali 77607 -48671 77641 -48637 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.A
flabel nwell 77607 -48365 77641 -48331 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.VPB
flabel pwell 77607 -48909 77641 -48875 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x10.VNB
rlabel comment 77578 -48892 77578 -48892 4 16to4_PriorityEncoder_v0p0p1_0.x3.x10.and2_1
rlabel metal1 77578 -48940 78038 -48844 1 16to4_PriorityEncoder_v0p0p1_0.x3.x10.VGND
rlabel metal1 77578 -48396 78038 -48300 1 16to4_PriorityEncoder_v0p0p1_0.x3.x10.VPWR
flabel locali 77792 -47421 77826 -47387 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.C
flabel locali 77884 -47421 77918 -47387 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.A
flabel locali 78068 -47285 78102 -47251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X
flabel locali 77700 -47421 77734 -47387 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.C
flabel locali 77792 -47217 77826 -47183 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.B
flabel locali 77700 -47217 77734 -47183 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.B
flabel locali 77700 -47353 77734 -47319 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.C
flabel locali 77608 -47217 77642 -47183 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.B
flabel locali 77792 -47353 77826 -47319 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.C
flabel locali 77608 -47421 77642 -47387 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.D
flabel locali 77608 -47489 77642 -47455 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.D
flabel metal1 77608 -47115 77642 -47081 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.VPWR
flabel metal1 77608 -47659 77642 -47625 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.VGND
flabel nwell 77608 -47115 77642 -47081 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.VPB
flabel pwell 77608 -47659 77642 -47625 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x1.VNB
rlabel comment 77578 -47642 77578 -47642 4 16to4_PriorityEncoder_v0p0p1_0.x3.x1.or4_1
rlabel metal1 77578 -47690 78130 -47594 1 16to4_PriorityEncoder_v0p0p1_0.x3.x1.VGND
rlabel metal1 77578 -47146 78130 -47050 1 16to4_PriorityEncoder_v0p0p1_0.x3.x1.VPWR
flabel locali 77792 -47983 77826 -47949 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.C
flabel locali 77884 -47983 77918 -47949 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.A
flabel locali 78068 -48119 78102 -48085 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X
flabel locali 77700 -47983 77734 -47949 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.C
flabel locali 77792 -48187 77826 -48153 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.B
flabel locali 77700 -48187 77734 -48153 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.B
flabel locali 77700 -48051 77734 -48017 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.C
flabel locali 77608 -48187 77642 -48153 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.B
flabel locali 77792 -48051 77826 -48017 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.C
flabel locali 77608 -47983 77642 -47949 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.D
flabel locali 77608 -47915 77642 -47881 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.D
flabel metal1 77608 -48289 77642 -48255 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.VPWR
flabel metal1 77608 -47745 77642 -47711 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.VGND
flabel nwell 77608 -48289 77642 -48255 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.VPB
flabel pwell 77608 -47745 77642 -47711 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x2.VNB
rlabel comment 77578 -47728 77578 -47728 2 16to4_PriorityEncoder_v0p0p1_0.x3.x2.or4_1
rlabel metal1 77578 -47776 78130 -47680 5 16to4_PriorityEncoder_v0p0p1_0.x3.x2.VGND
rlabel metal1 77578 -48320 78130 -48224 5 16to4_PriorityEncoder_v0p0p1_0.x3.x2.VPWR
flabel locali 78342 -47421 78376 -47387 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A
flabel locali 78250 -47421 78284 -47387 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A
flabel locali 78526 -47285 78560 -47251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.X
flabel locali 78250 -47353 78284 -47319 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A
flabel locali 78158 -47217 78192 -47183 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B
flabel locali 78250 -47217 78284 -47183 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B
flabel locali 78158 -47421 78192 -47387 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C
flabel metal1 78158 -47115 78192 -47081 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.VPWR
flabel metal1 78158 -47659 78192 -47625 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.VGND
flabel nwell 78158 -47115 78192 -47081 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.VPB
flabel pwell 78158 -47659 78192 -47625 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x4.VNB
rlabel comment 78130 -47642 78130 -47642 4 16to4_PriorityEncoder_v0p0p1_0.x3.x4.or3_1
rlabel metal1 78130 -47690 78590 -47594 1 16to4_PriorityEncoder_v0p0p1_0.x3.x4.VGND
rlabel metal1 78130 -47146 78590 -47050 1 16to4_PriorityEncoder_v0p0p1_0.x3.x4.VPWR
flabel metal1 78619 -47115 78653 -47081 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.VPWR
flabel metal1 78619 -47659 78653 -47625 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.VGND
flabel locali 78987 -47489 79021 -47455 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.X
flabel locali 78987 -47557 79021 -47523 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.X
flabel locali 78987 -47421 79021 -47387 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.X
flabel locali 78987 -47353 79021 -47319 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.X
flabel locali 78987 -47285 79021 -47251 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.X
flabel locali 78987 -47217 79021 -47183 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.X
flabel locali 78803 -47421 78837 -47387 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.B
flabel locali 78711 -47421 78745 -47387 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.A
flabel locali 78619 -47421 78653 -47387 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.A
flabel nwell 78619 -47115 78653 -47081 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.VPB
flabel pwell 78619 -47659 78653 -47625 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x8.VNB
rlabel comment 78590 -47642 78590 -47642 4 16to4_PriorityEncoder_v0p0p1_0.x3.x8.and2_1
rlabel metal1 78590 -47690 79050 -47594 1 16to4_PriorityEncoder_v0p0p1_0.x3.x8.VGND
rlabel metal1 78590 -47146 79050 -47050 1 16to4_PriorityEncoder_v0p0p1_0.x3.x8.VPWR
flabel locali 76496 -46751 76530 -46717 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x3.Y
flabel locali 76496 -46683 76530 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x3.Y
flabel locali 76404 -46683 76438 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x3.A
flabel nwell 76361 -46989 76395 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x3.VPB
flabel pwell 76361 -46445 76395 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x3.VNB
flabel metal1 76361 -46445 76395 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x3.VGND
flabel metal1 76361 -46989 76395 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x3.VPWR
rlabel comment 76332 -46428 76332 -46428 2 16to4_PriorityEncoder_v0p0p1_0.x3.x3.inv_1
rlabel metal1 76332 -46476 76608 -46380 5 16to4_PriorityEncoder_v0p0p1_0.x3.x3.VGND
rlabel metal1 76332 -47020 76608 -46924 5 16to4_PriorityEncoder_v0p0p1_0.x3.x3.VPWR
flabel locali 76220 -46751 76254 -46717 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x5.Y
flabel locali 76220 -46683 76254 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x5.Y
flabel locali 76128 -46683 76162 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x5.A
flabel nwell 76085 -46989 76119 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x5.VPB
flabel pwell 76085 -46445 76119 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x5.VNB
flabel metal1 76085 -46445 76119 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x5.VGND
flabel metal1 76085 -46989 76119 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x5.VPWR
rlabel comment 76056 -46428 76056 -46428 2 16to4_PriorityEncoder_v0p0p1_0.x3.x5.inv_1
rlabel metal1 76056 -46476 76332 -46380 5 16to4_PriorityEncoder_v0p0p1_0.x3.x5.VGND
rlabel metal1 76056 -47020 76332 -46924 5 16to4_PriorityEncoder_v0p0p1_0.x3.x5.VPWR
flabel locali 75946 -46751 75980 -46717 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x6.Y
flabel locali 75946 -46683 75980 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x6.Y
flabel locali 75854 -46683 75888 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x6.A
flabel nwell 75811 -46989 75845 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x6.VPB
flabel pwell 75811 -46445 75845 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x6.VNB
flabel metal1 75811 -46445 75845 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x6.VGND
flabel metal1 75811 -46989 75845 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x6.VPWR
rlabel comment 75782 -46428 75782 -46428 2 16to4_PriorityEncoder_v0p0p1_0.x3.x6.inv_1
rlabel metal1 75782 -46476 76058 -46380 5 16to4_PriorityEncoder_v0p0p1_0.x3.x6.VGND
rlabel metal1 75782 -47020 76058 -46924 5 16to4_PriorityEncoder_v0p0p1_0.x3.x6.VPWR
flabel locali 75670 -46751 75704 -46717 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x7.Y
flabel locali 75670 -46683 75704 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x7.Y
flabel locali 75578 -46683 75612 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x7.A
flabel nwell 75535 -46989 75569 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x7.VPB
flabel pwell 75535 -46445 75569 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x7.VNB
flabel metal1 75535 -46445 75569 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x7.VGND
flabel metal1 75535 -46989 75569 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x7.VPWR
rlabel comment 75506 -46428 75506 -46428 2 16to4_PriorityEncoder_v0p0p1_0.x3.x7.inv_1
rlabel metal1 75506 -46476 75782 -46380 5 16to4_PriorityEncoder_v0p0p1_0.x3.x7.VGND
rlabel metal1 75506 -47020 75782 -46924 5 16to4_PriorityEncoder_v0p0p1_0.x3.x7.VPWR
flabel locali 76772 -46751 76806 -46717 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y
flabel locali 76772 -46683 76806 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y
flabel locali 76680 -46683 76714 -46649 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x9.A
flabel nwell 76637 -46989 76671 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x9.VPB
flabel pwell 76637 -46445 76671 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x9.VNB
flabel metal1 76637 -46445 76671 -46411 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x9.VGND
flabel metal1 76637 -46989 76671 -46955 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x3.x9.VPWR
rlabel comment 76608 -46428 76608 -46428 2 16to4_PriorityEncoder_v0p0p1_0.x3.x9.inv_1
rlabel metal1 76608 -46476 76884 -46380 5 16to4_PriorityEncoder_v0p0p1_0.x3.x9.VGND
rlabel metal1 76608 -47020 76884 -46924 5 16to4_PriorityEncoder_v0p0p1_0.x3.x9.VPWR
flabel locali 83051 -51721 83085 -51687 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x2.A
flabel locali 83235 -51585 83269 -51551 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x2.X
flabel locali 82867 -51721 82901 -51687 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x2.B
flabel nwell 82867 -51415 82901 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x2.VPB
flabel pwell 82867 -51959 82901 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x2.VNB
flabel metal1 82867 -51959 82901 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x2.VGND
flabel metal1 82867 -51415 82901 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x2.VPWR
rlabel comment 82838 -51942 82838 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x2.or2_1
rlabel metal1 82838 -51990 83298 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x2.VGND
rlabel metal1 82838 -51446 83298 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x2.VPWR
flabel locali 85351 -51721 85385 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.Y
flabel locali 85351 -51789 85385 -51755 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.Y
flabel locali 84063 -51721 84097 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.A
flabel locali 84431 -51721 84465 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.A
flabel locali 84799 -51721 84833 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.A
flabel locali 84891 -51721 84925 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.A
flabel nwell 84063 -51415 84097 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.VPB
flabel pwell 84063 -51959 84097 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.VNB
flabel metal1 84063 -51959 84097 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.VGND
flabel metal1 84063 -51415 84097 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x22.VPWR
rlabel comment 84034 -51942 84034 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x22.inv_16
rlabel metal1 84034 -51990 85506 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x22.VGND
rlabel metal1 84034 -51446 85506 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x22.VPWR
flabel locali 83971 -51789 84005 -51755 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.Y
flabel locali 83971 -51721 84005 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.Y
flabel locali 83971 -51653 84005 -51619 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.Y
flabel locali 83603 -51721 83637 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.A
flabel locali 83695 -51721 83729 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.A
flabel locali 83787 -51721 83821 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.A
flabel locali 83879 -51721 83913 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.A
flabel nwell 83603 -51415 83637 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.VPB
flabel pwell 83603 -51959 83637 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.VNB
flabel metal1 83603 -51415 83637 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.VPWR
flabel metal1 83603 -51959 83637 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x21.VGND
rlabel comment 83574 -51942 83574 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x21.inv_4
rlabel metal1 83574 -51990 84034 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x21.VGND
rlabel metal1 83574 -51446 84034 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x21.VPWR
flabel locali 83462 -51653 83496 -51619 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x20.Y
flabel locali 83462 -51721 83496 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x20.Y
flabel locali 83370 -51721 83404 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x20.A
flabel nwell 83327 -51415 83361 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x20.VPB
flabel pwell 83327 -51959 83361 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x20.VNB
flabel metal1 83327 -51959 83361 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x20.VGND
flabel metal1 83327 -51415 83361 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x20.VPWR
rlabel comment 83298 -51942 83298 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x20.inv_1
rlabel metal1 83298 -51990 83574 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x20.VGND
rlabel metal1 83298 -51446 83574 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x20.VPWR
flabel locali 88295 -51721 88329 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.Y
flabel locali 88295 -51789 88329 -51755 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.Y
flabel locali 87007 -51721 87041 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.A
flabel locali 87375 -51721 87409 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.A
flabel locali 87743 -51721 87777 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.A
flabel locali 87835 -51721 87869 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.A
flabel nwell 87007 -51415 87041 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.VPB
flabel pwell 87007 -51959 87041 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.VNB
flabel metal1 87007 -51959 87041 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.VGND
flabel metal1 87007 -51415 87041 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x23.VPWR
rlabel comment 86978 -51942 86978 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x23.inv_16
rlabel metal1 86978 -51990 88450 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x23.VGND
rlabel metal1 86978 -51446 88450 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x23.VPWR
flabel locali 86823 -51721 86857 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.Y
flabel locali 86823 -51789 86857 -51755 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.Y
flabel locali 85535 -51721 85569 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.A
flabel locali 85903 -51721 85937 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.A
flabel locali 86271 -51721 86305 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.A
flabel locali 86363 -51721 86397 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.A
flabel nwell 85535 -51415 85569 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.VPB
flabel pwell 85535 -51959 85569 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.VNB
flabel metal1 85535 -51959 85569 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.VGND
flabel metal1 85535 -51415 85569 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x19.VPWR
rlabel comment 85506 -51942 85506 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x19.inv_16
rlabel metal1 85506 -51990 86978 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x19.VGND
rlabel metal1 85506 -51446 86978 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x19.VPWR
flabel locali 83051 -48071 83085 -48037 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x1.A
flabel locali 83235 -47935 83269 -47901 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x1.X
flabel locali 82867 -48071 82901 -48037 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x1.B
flabel nwell 82867 -47765 82901 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x1.VPB
flabel pwell 82867 -48309 82901 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x1.VNB
flabel metal1 82867 -48309 82901 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x1.VGND
flabel metal1 82867 -47765 82901 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x1.VPWR
rlabel comment 82838 -48292 82838 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x1.or2_1
rlabel metal1 82838 -48340 83298 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x1.VGND
rlabel metal1 82838 -47796 83298 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x1.VPWR
flabel locali 85351 -48071 85385 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.Y
flabel locali 85351 -48139 85385 -48105 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.Y
flabel locali 84063 -48071 84097 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.A
flabel locali 84431 -48071 84465 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.A
flabel locali 84799 -48071 84833 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.A
flabel locali 84891 -48071 84925 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.A
flabel nwell 84063 -47765 84097 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.VPB
flabel pwell 84063 -48309 84097 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.VNB
flabel metal1 84063 -48309 84097 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.VGND
flabel metal1 84063 -47765 84097 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x29.VPWR
rlabel comment 84034 -48292 84034 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x29.inv_16
rlabel metal1 84034 -48340 85506 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x29.VGND
rlabel metal1 84034 -47796 85506 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x29.VPWR
flabel locali 83971 -48139 84005 -48105 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.Y
flabel locali 83971 -48071 84005 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.Y
flabel locali 83971 -48003 84005 -47969 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.Y
flabel locali 83603 -48071 83637 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.A
flabel locali 83695 -48071 83729 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.A
flabel locali 83787 -48071 83821 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.A
flabel locali 83879 -48071 83913 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.A
flabel nwell 83603 -47765 83637 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.VPB
flabel pwell 83603 -48309 83637 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.VNB
flabel metal1 83603 -47765 83637 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.VPWR
flabel metal1 83603 -48309 83637 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x28.VGND
rlabel comment 83574 -48292 83574 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x28.inv_4
rlabel metal1 83574 -48340 84034 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x28.VGND
rlabel metal1 83574 -47796 84034 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x28.VPWR
flabel locali 83462 -48003 83496 -47969 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x27.Y
flabel locali 83462 -48071 83496 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x27.Y
flabel locali 83370 -48071 83404 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x27.A
flabel nwell 83327 -47765 83361 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x27.VPB
flabel pwell 83327 -48309 83361 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x27.VNB
flabel metal1 83327 -48309 83361 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x27.VGND
flabel metal1 83327 -47765 83361 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x27.VPWR
rlabel comment 83298 -48292 83298 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x27.inv_1
rlabel metal1 83298 -48340 83574 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x27.VGND
rlabel metal1 83298 -47796 83574 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x27.VPWR
flabel locali 88295 -48071 88329 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.Y
flabel locali 88295 -48139 88329 -48105 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.Y
flabel locali 87007 -48071 87041 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.A
flabel locali 87375 -48071 87409 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.A
flabel locali 87743 -48071 87777 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.A
flabel locali 87835 -48071 87869 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.A
flabel nwell 87007 -47765 87041 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.VPB
flabel pwell 87007 -48309 87041 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.VNB
flabel metal1 87007 -48309 87041 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.VGND
flabel metal1 87007 -47765 87041 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x16.VPWR
rlabel comment 86978 -48292 86978 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x16.inv_16
rlabel metal1 86978 -48340 88450 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x16.VGND
rlabel metal1 86978 -47796 88450 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x16.VPWR
flabel locali 86823 -48071 86857 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.Y
flabel locali 86823 -48139 86857 -48105 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.Y
flabel locali 85535 -48071 85569 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.A
flabel locali 85903 -48071 85937 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.A
flabel locali 86271 -48071 86305 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.A
flabel locali 86363 -48071 86397 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.A
flabel nwell 85535 -47765 85569 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.VPB
flabel pwell 85535 -48309 85569 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.VNB
flabel metal1 85535 -48309 85569 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.VGND
flabel metal1 85535 -47765 85569 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x15.VPWR
rlabel comment 85506 -48292 85506 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x15.inv_16
rlabel metal1 85506 -48340 86978 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x15.VGND
rlabel metal1 85506 -47796 86978 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x15.VPWR
flabel locali 89767 -48071 89801 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.Y
flabel locali 89767 -48139 89801 -48105 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.Y
flabel locali 88479 -48071 88513 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.A
flabel locali 88847 -48071 88881 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.A
flabel locali 89215 -48071 89249 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.A
flabel locali 89307 -48071 89341 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.A
flabel nwell 88479 -47765 88513 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.VPB
flabel pwell 88479 -48309 88513 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.VNB
flabel metal1 88479 -48309 88513 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.VGND
flabel metal1 88479 -47765 88513 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x17.VPWR
rlabel comment 88450 -48292 88450 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x17.inv_16
rlabel metal1 88450 -48340 89922 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x17.VGND
rlabel metal1 88450 -47796 89922 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x17.VPWR
flabel locali 91239 -48071 91273 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.Y
flabel locali 91239 -48139 91273 -48105 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.Y
flabel locali 89951 -48071 89985 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.A
flabel locali 90319 -48071 90353 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.A
flabel locali 90687 -48071 90721 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.A
flabel locali 90779 -48071 90813 -48037 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.A
flabel nwell 89951 -47765 89985 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.VPB
flabel pwell 89951 -48309 89985 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.VNB
flabel metal1 89951 -48309 89985 -48275 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.VGND
flabel metal1 89951 -47765 89985 -47731 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x18.VPWR
rlabel comment 89922 -48292 89922 -48292 4 16to4_PriorityEncoder_v0p0p1_0.x18.inv_16
rlabel metal1 89922 -48340 91394 -48244 1 16to4_PriorityEncoder_v0p0p1_0.x18.VGND
rlabel metal1 89922 -47796 91394 -47700 1 16to4_PriorityEncoder_v0p0p1_0.x18.VPWR
flabel locali 89767 -51721 89801 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.Y
flabel locali 89767 -51789 89801 -51755 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.Y
flabel locali 88479 -51721 88513 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.A
flabel locali 88847 -51721 88881 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.A
flabel locali 89215 -51721 89249 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.A
flabel locali 89307 -51721 89341 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.A
flabel nwell 88479 -51415 88513 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.VPB
flabel pwell 88479 -51959 88513 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.VNB
flabel metal1 88479 -51959 88513 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.VGND
flabel metal1 88479 -51415 88513 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x24.VPWR
rlabel comment 88450 -51942 88450 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x24.inv_16
rlabel metal1 88450 -51990 89922 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x24.VGND
rlabel metal1 88450 -51446 89922 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x24.VPWR
flabel locali 91239 -51721 91273 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.Y
flabel locali 91239 -51789 91273 -51755 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.Y
flabel locali 89951 -51721 89985 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.A
flabel locali 90319 -51721 90353 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.A
flabel locali 90687 -51721 90721 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.A
flabel locali 90779 -51721 90813 -51687 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.A
flabel nwell 89951 -51415 89985 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.VPB
flabel pwell 89951 -51959 89985 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.VNB
flabel metal1 89951 -51959 89985 -51925 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.VGND
flabel metal1 89951 -51415 89985 -51381 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x25.VPWR
rlabel comment 89922 -51942 89922 -51942 4 16to4_PriorityEncoder_v0p0p1_0.x25.inv_16
rlabel metal1 89922 -51990 91394 -51894 1 16to4_PriorityEncoder_v0p0p1_0.x25.VGND
rlabel metal1 89922 -51446 91394 -51350 1 16to4_PriorityEncoder_v0p0p1_0.x25.VPWR
flabel metal1 73180 -38340 73380 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I0
flabel metal1 73430 -38340 73630 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I1
flabel metal1 73680 -38340 73880 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I2
flabel metal1 73930 -38340 74130 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I3
flabel metal1 74180 -38340 74380 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I4
flabel metal1 74430 -38340 74630 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I5
flabel metal1 74680 -38340 74880 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I6
flabel metal1 74930 -38340 75130 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.I7
flabel metal1 75180 -38340 75380 -38140 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.EI
flabel metal1 80460 -39980 80660 -39780 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.EO
flabel metal1 80460 -39530 80660 -39330 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.GS
flabel metal1 80460 -41200 80660 -41000 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.A2
flabel metal1 80390 -43190 80590 -42990 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.A1
flabel metal1 80390 -45730 80590 -45530 0 FreeSans 256 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.A0
flabel metal5 79380 -40150 79710 -38130 0 FreeSans 512 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.VDD
flabel metal4 76900 -45640 77080 -44610 0 FreeSans 512 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.GND
flabel locali 78159 -45107 78193 -45073 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X
flabel locali 77883 -44767 77917 -44733 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C
flabel locali 77883 -44835 77917 -44801 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C
flabel locali 77607 -44903 77641 -44869 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.A
flabel locali 77883 -44903 77917 -44869 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C
flabel locali 77791 -44767 77825 -44733 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.B
flabel locali 77791 -44835 77825 -44801 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.B
flabel locali 77975 -44903 78009 -44869 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D
flabel locali 78159 -44767 78193 -44733 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X
flabel locali 78159 -44835 78193 -44801 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X
flabel locali 78159 -44903 78193 -44869 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X
flabel locali 78159 -44971 78193 -44937 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X
flabel locali 78159 -45039 78193 -45005 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X
flabel metal1 77607 -44665 77641 -44631 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.VGND
flabel metal1 77607 -45209 77641 -45175 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.VPWR
flabel nwell 77607 -45209 77641 -45175 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.VPB
flabel pwell 77607 -44665 77641 -44631 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x19.VNB
rlabel comment 77578 -44648 77578 -44648 2 16to4_PriorityEncoder_v0p0p1_0.x5.x19.and4_1
rlabel metal1 77578 -44696 78222 -44600 5 16to4_PriorityEncoder_v0p0p1_0.x5.x19.VGND
rlabel metal1 77578 -45240 78222 -45144 5 16to4_PriorityEncoder_v0p0p1_0.x5.x19.VPWR
flabel metal1 77607 -45829 77641 -45795 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.VGND
flabel metal1 77607 -45285 77641 -45251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.VPWR
flabel locali 77975 -45387 78009 -45353 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X
flabel locali 77975 -45727 78009 -45693 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X
flabel locali 77791 -45387 77825 -45353 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B
flabel locali 77607 -45659 77641 -45625 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.A
flabel locali 77813 -45659 77847 -45625 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.C
flabel nwell 77607 -45285 77641 -45251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.VPB
flabel pwell 77607 -45829 77641 -45795 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x20.VNB
rlabel comment 77578 -45812 77578 -45812 4 16to4_PriorityEncoder_v0p0p1_0.x5.x20.and3_1
rlabel metal1 77578 -45860 78038 -45764 1 16to4_PriorityEncoder_v0p0p1_0.x5.x20.VGND
rlabel metal1 77578 -45316 78038 -45220 1 16to4_PriorityEncoder_v0p0p1_0.x5.x20.VPWR
flabel metal1 78067 -45285 78101 -45251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.VPWR
flabel metal1 78067 -45829 78101 -45795 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.VGND
flabel locali 78435 -45659 78469 -45625 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X
flabel locali 78435 -45727 78469 -45693 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X
flabel locali 78435 -45591 78469 -45557 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X
flabel locali 78435 -45523 78469 -45489 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X
flabel locali 78435 -45455 78469 -45421 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X
flabel locali 78435 -45387 78469 -45353 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X
flabel locali 78251 -45591 78285 -45557 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B
flabel locali 78159 -45591 78193 -45557 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.A
flabel locali 78067 -45591 78101 -45557 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.A
flabel nwell 78067 -45285 78101 -45251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.VPB
flabel pwell 78067 -45829 78101 -45795 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x21.VNB
rlabel comment 78038 -45812 78038 -45812 4 16to4_PriorityEncoder_v0p0p1_0.x5.x21.and2_1
rlabel metal1 78038 -45860 78498 -45764 1 16to4_PriorityEncoder_v0p0p1_0.x5.x21.VGND
rlabel metal1 78038 -45316 78498 -45220 1 16to4_PriorityEncoder_v0p0p1_0.x5.x21.VPWR
flabel locali 78712 -45591 78746 -45557 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C
flabel locali 78804 -45591 78838 -45557 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A
flabel locali 78988 -45455 79022 -45421 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.X
flabel locali 78620 -45591 78654 -45557 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C
flabel locali 78712 -45387 78746 -45353 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B
flabel locali 78620 -45387 78654 -45353 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B
flabel locali 78620 -45523 78654 -45489 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C
flabel locali 78528 -45387 78562 -45353 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B
flabel locali 78712 -45523 78746 -45489 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C
flabel locali 78528 -45591 78562 -45557 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D
flabel locali 78528 -45659 78562 -45625 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D
flabel metal1 78528 -45285 78562 -45251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.VPWR
flabel metal1 78528 -45829 78562 -45795 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.VGND
flabel nwell 78528 -45285 78562 -45251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.VPB
flabel pwell 78528 -45829 78562 -45795 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x22.VNB
rlabel comment 78498 -45812 78498 -45812 4 16to4_PriorityEncoder_v0p0p1_0.x5.x22.or4_1
rlabel metal1 78498 -45860 79050 -45764 1 16to4_PriorityEncoder_v0p0p1_0.x5.x22.VGND
rlabel metal1 78498 -45316 79050 -45220 1 16to4_PriorityEncoder_v0p0p1_0.x5.x22.VPWR
flabel locali 78159 -43873 78193 -43839 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X
flabel locali 77883 -43533 77917 -43499 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C
flabel locali 77883 -43601 77917 -43567 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C
flabel locali 77607 -43669 77641 -43635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.A
flabel locali 77883 -43669 77917 -43635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C
flabel locali 77791 -43533 77825 -43499 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.B
flabel locali 77791 -43601 77825 -43567 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.B
flabel locali 77975 -43669 78009 -43635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.D
flabel locali 78159 -43533 78193 -43499 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X
flabel locali 78159 -43601 78193 -43567 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X
flabel locali 78159 -43669 78193 -43635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X
flabel locali 78159 -43737 78193 -43703 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X
flabel locali 78159 -43805 78193 -43771 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X
flabel metal1 77607 -43431 77641 -43397 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.VGND
flabel metal1 77607 -43975 77641 -43941 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.VPWR
flabel nwell 77607 -43975 77641 -43941 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.VPB
flabel pwell 77607 -43431 77641 -43397 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x16.VNB
rlabel comment 77578 -43414 77578 -43414 2 16to4_PriorityEncoder_v0p0p1_0.x5.x16.and4_1
rlabel metal1 77578 -43462 78222 -43366 5 16to4_PriorityEncoder_v0p0p1_0.x5.x16.VGND
rlabel metal1 77578 -44006 78222 -43910 5 16to4_PriorityEncoder_v0p0p1_0.x5.x16.VPWR
flabel locali 78159 -44149 78193 -44115 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.X
flabel locali 77883 -44489 77917 -44455 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C
flabel locali 77883 -44421 77917 -44387 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C
flabel locali 77607 -44353 77641 -44319 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.A
flabel locali 77883 -44353 77917 -44319 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C
flabel locali 77791 -44489 77825 -44455 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.B
flabel locali 77791 -44421 77825 -44387 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.B
flabel locali 77975 -44353 78009 -44319 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.D
flabel locali 78159 -44489 78193 -44455 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.X
flabel locali 78159 -44421 78193 -44387 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.X
flabel locali 78159 -44353 78193 -44319 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.X
flabel locali 78159 -44285 78193 -44251 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.X
flabel locali 78159 -44217 78193 -44183 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.X
flabel metal1 77607 -44591 77641 -44557 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.VGND
flabel metal1 77607 -44047 77641 -44013 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.VPWR
flabel nwell 77607 -44047 77641 -44013 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.VPB
flabel pwell 77607 -44591 77641 -44557 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x18.VNB
rlabel comment 77578 -44574 77578 -44574 4 16to4_PriorityEncoder_v0p0p1_0.x5.x18.and4_1
rlabel metal1 77578 -44622 78222 -44526 1 16to4_PriorityEncoder_v0p0p1_0.x5.x18.VGND
rlabel metal1 77578 -44078 78222 -43982 1 16to4_PriorityEncoder_v0p0p1_0.x5.x18.VPWR
flabel metal1 77609 -42743 77643 -42709 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.VPWR
flabel metal1 77609 -42199 77643 -42165 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.VGND
flabel locali 77977 -42369 78011 -42335 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.X
flabel locali 77977 -42301 78011 -42267 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.X
flabel locali 77977 -42437 78011 -42403 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.X
flabel locali 77977 -42505 78011 -42471 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.X
flabel locali 77977 -42573 78011 -42539 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.X
flabel locali 77977 -42641 78011 -42607 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.X
flabel locali 77793 -42437 77827 -42403 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.B
flabel locali 77701 -42437 77735 -42403 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.A
flabel locali 77609 -42437 77643 -42403 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.A
flabel nwell 77609 -42743 77643 -42709 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.VPB
flabel pwell 77609 -42199 77643 -42165 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x13.VNB
rlabel comment 77580 -42182 77580 -42182 2 16to4_PriorityEncoder_v0p0p1_0.x5.x13.and2_1
rlabel metal1 77580 -42230 78040 -42134 5 16to4_PriorityEncoder_v0p0p1_0.x5.x13.VGND
rlabel metal1 77580 -42774 78040 -42678 5 16to4_PriorityEncoder_v0p0p1_0.x5.x13.VPWR
flabel locali 78159 -42917 78193 -42883 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X
flabel locali 77883 -43257 77917 -43223 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.C
flabel locali 77883 -43189 77917 -43155 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.C
flabel locali 77607 -43121 77641 -43087 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.A
flabel locali 77883 -43121 77917 -43087 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.C
flabel locali 77791 -43257 77825 -43223 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.B
flabel locali 77791 -43189 77825 -43155 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.B
flabel locali 77975 -43121 78009 -43087 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.D
flabel locali 78159 -43257 78193 -43223 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X
flabel locali 78159 -43189 78193 -43155 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X
flabel locali 78159 -43121 78193 -43087 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X
flabel locali 78159 -43053 78193 -43019 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X
flabel locali 78159 -42985 78193 -42951 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X
flabel metal1 77607 -43359 77641 -43325 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.VGND
flabel metal1 77607 -42815 77641 -42781 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.VPWR
flabel nwell 77607 -42815 77641 -42781 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.VPB
flabel pwell 77607 -43359 77641 -43325 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x15.VNB
rlabel comment 77578 -43342 77578 -43342 4 16to4_PriorityEncoder_v0p0p1_0.x5.x15.and4_1
rlabel metal1 77578 -43390 78222 -43294 1 16to4_PriorityEncoder_v0p0p1_0.x5.x15.VGND
rlabel metal1 77578 -42846 78222 -42750 1 16to4_PriorityEncoder_v0p0p1_0.x5.x15.VPWR
flabel locali 78536 -43121 78570 -43087 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C
flabel locali 78628 -43121 78662 -43087 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A
flabel locali 78812 -42985 78846 -42951 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.X
flabel locali 78444 -43121 78478 -43087 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C
flabel locali 78536 -42917 78570 -42883 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.B
flabel locali 78444 -42917 78478 -42883 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.B
flabel locali 78444 -43053 78478 -43019 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C
flabel locali 78352 -42917 78386 -42883 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.B
flabel locali 78536 -43053 78570 -43019 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C
flabel locali 78352 -43121 78386 -43087 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D
flabel locali 78352 -43189 78386 -43155 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D
flabel metal1 78352 -42815 78386 -42781 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.VPWR
flabel metal1 78352 -43359 78386 -43325 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.VGND
flabel nwell 78352 -42815 78386 -42781 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.VPB
flabel pwell 78352 -43359 78386 -43325 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x17.VNB
rlabel comment 78322 -43342 78322 -43342 4 16to4_PriorityEncoder_v0p0p1_0.x5.x17.or4_1
rlabel metal1 78322 -43390 78874 -43294 1 16to4_PriorityEncoder_v0p0p1_0.x5.x17.VGND
rlabel metal1 78322 -42846 78874 -42750 1 16to4_PriorityEncoder_v0p0p1_0.x5.x17.VPWR
flabel metal1 77607 -41489 77641 -41455 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.VPWR
flabel metal1 77607 -40945 77641 -40911 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.VGND
flabel locali 77975 -41115 78009 -41081 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X
flabel locali 77975 -41047 78009 -41013 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X
flabel locali 77975 -41183 78009 -41149 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X
flabel locali 77975 -41251 78009 -41217 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X
flabel locali 77975 -41319 78009 -41285 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X
flabel locali 77975 -41387 78009 -41353 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X
flabel locali 77791 -41183 77825 -41149 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.B
flabel locali 77699 -41183 77733 -41149 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.A
flabel locali 77607 -41183 77641 -41149 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.A
flabel nwell 77607 -41489 77641 -41455 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.VPB
flabel pwell 77607 -40945 77641 -40911 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x11.VNB
rlabel comment 77578 -40928 77578 -40928 2 16to4_PriorityEncoder_v0p0p1_0.x5.x11.and2_1
rlabel metal1 77578 -40976 78038 -40880 5 16to4_PriorityEncoder_v0p0p1_0.x5.x11.VGND
rlabel metal1 77578 -41520 78038 -41424 5 16to4_PriorityEncoder_v0p0p1_0.x5.x11.VPWR
flabel metal1 77607 -41565 77641 -41531 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.VPWR
flabel metal1 77607 -42109 77641 -42075 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.VGND
flabel locali 77975 -41939 78009 -41905 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.X
flabel locali 77975 -42007 78009 -41973 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.X
flabel locali 77975 -41871 78009 -41837 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.X
flabel locali 77975 -41803 78009 -41769 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.X
flabel locali 77975 -41735 78009 -41701 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.X
flabel locali 77975 -41667 78009 -41633 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.X
flabel locali 77791 -41871 77825 -41837 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.B
flabel locali 77699 -41871 77733 -41837 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.A
flabel locali 77607 -41871 77641 -41837 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.A
flabel nwell 77607 -41565 77641 -41531 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.VPB
flabel pwell 77607 -42109 77641 -42075 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x12.VNB
rlabel comment 77578 -42092 77578 -42092 4 16to4_PriorityEncoder_v0p0p1_0.x5.x12.and2_1
rlabel metal1 77578 -42140 78038 -42044 1 16to4_PriorityEncoder_v0p0p1_0.x5.x12.VGND
rlabel metal1 77578 -41596 78038 -41500 1 16to4_PriorityEncoder_v0p0p1_0.x5.x12.VPWR
flabel locali 78252 -41183 78286 -41149 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.C
flabel locali 78344 -41183 78378 -41149 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A
flabel locali 78528 -41319 78562 -41285 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.X
flabel locali 78160 -41183 78194 -41149 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.C
flabel locali 78252 -41387 78286 -41353 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B
flabel locali 78160 -41387 78194 -41353 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B
flabel locali 78160 -41251 78194 -41217 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.C
flabel locali 78068 -41387 78102 -41353 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B
flabel locali 78252 -41251 78286 -41217 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.C
flabel locali 78068 -41183 78102 -41149 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.D
flabel locali 78068 -41115 78102 -41081 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.D
flabel metal1 78068 -41489 78102 -41455 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.VPWR
flabel metal1 78068 -40945 78102 -40911 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.VGND
flabel nwell 78068 -41489 78102 -41455 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.VPB
flabel pwell 78068 -40945 78102 -40911 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x14.VNB
rlabel comment 78038 -40928 78038 -40928 2 16to4_PriorityEncoder_v0p0p1_0.x5.x14.or4_1
rlabel metal1 78038 -40976 78590 -40880 5 16to4_PriorityEncoder_v0p0p1_0.x5.x14.VGND
rlabel metal1 78038 -41520 78590 -41424 5 16to4_PriorityEncoder_v0p0p1_0.x5.x14.VPWR
flabel metal1 77607 -40325 77641 -40291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.VPWR
flabel metal1 77607 -40869 77641 -40835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.VGND
flabel locali 77975 -40699 78009 -40665 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.X
flabel locali 77975 -40767 78009 -40733 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.X
flabel locali 77975 -40631 78009 -40597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.X
flabel locali 77975 -40563 78009 -40529 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.X
flabel locali 77975 -40495 78009 -40461 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.X
flabel locali 77975 -40427 78009 -40393 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.X
flabel locali 77791 -40631 77825 -40597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.B
flabel locali 77699 -40631 77733 -40597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.A
flabel locali 77607 -40631 77641 -40597 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.A
flabel nwell 77607 -40325 77641 -40291 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.VPB
flabel pwell 77607 -40869 77641 -40835 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x10.VNB
rlabel comment 77578 -40852 77578 -40852 4 16to4_PriorityEncoder_v0p0p1_0.x5.x10.and2_1
rlabel metal1 77578 -40900 78038 -40804 1 16to4_PriorityEncoder_v0p0p1_0.x5.x10.VGND
rlabel metal1 77578 -40356 78038 -40260 1 16to4_PriorityEncoder_v0p0p1_0.x5.x10.VPWR
flabel locali 77792 -39381 77826 -39347 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.C
flabel locali 77884 -39381 77918 -39347 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.A
flabel locali 78068 -39245 78102 -39211 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X
flabel locali 77700 -39381 77734 -39347 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.C
flabel locali 77792 -39177 77826 -39143 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.B
flabel locali 77700 -39177 77734 -39143 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.B
flabel locali 77700 -39313 77734 -39279 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.C
flabel locali 77608 -39177 77642 -39143 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.B
flabel locali 77792 -39313 77826 -39279 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.C
flabel locali 77608 -39381 77642 -39347 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.D
flabel locali 77608 -39449 77642 -39415 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.D
flabel metal1 77608 -39075 77642 -39041 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.VPWR
flabel metal1 77608 -39619 77642 -39585 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.VGND
flabel nwell 77608 -39075 77642 -39041 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.VPB
flabel pwell 77608 -39619 77642 -39585 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x1.VNB
rlabel comment 77578 -39602 77578 -39602 4 16to4_PriorityEncoder_v0p0p1_0.x5.x1.or4_1
rlabel metal1 77578 -39650 78130 -39554 1 16to4_PriorityEncoder_v0p0p1_0.x5.x1.VGND
rlabel metal1 77578 -39106 78130 -39010 1 16to4_PriorityEncoder_v0p0p1_0.x5.x1.VPWR
flabel locali 77792 -39943 77826 -39909 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.C
flabel locali 77884 -39943 77918 -39909 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.A
flabel locali 78068 -40079 78102 -40045 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X
flabel locali 77700 -39943 77734 -39909 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.C
flabel locali 77792 -40147 77826 -40113 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.B
flabel locali 77700 -40147 77734 -40113 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.B
flabel locali 77700 -40011 77734 -39977 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.C
flabel locali 77608 -40147 77642 -40113 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.B
flabel locali 77792 -40011 77826 -39977 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.C
flabel locali 77608 -39943 77642 -39909 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.D
flabel locali 77608 -39875 77642 -39841 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.D
flabel metal1 77608 -40249 77642 -40215 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.VPWR
flabel metal1 77608 -39705 77642 -39671 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.VGND
flabel nwell 77608 -40249 77642 -40215 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.VPB
flabel pwell 77608 -39705 77642 -39671 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x2.VNB
rlabel comment 77578 -39688 77578 -39688 2 16to4_PriorityEncoder_v0p0p1_0.x5.x2.or4_1
rlabel metal1 77578 -39736 78130 -39640 5 16to4_PriorityEncoder_v0p0p1_0.x5.x2.VGND
rlabel metal1 77578 -40280 78130 -40184 5 16to4_PriorityEncoder_v0p0p1_0.x5.x2.VPWR
flabel locali 78342 -39381 78376 -39347 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A
flabel locali 78250 -39381 78284 -39347 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A
flabel locali 78526 -39245 78560 -39211 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.X
flabel locali 78250 -39313 78284 -39279 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A
flabel locali 78158 -39177 78192 -39143 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B
flabel locali 78250 -39177 78284 -39143 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B
flabel locali 78158 -39381 78192 -39347 0 FreeSans 400 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C
flabel metal1 78158 -39075 78192 -39041 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.VPWR
flabel metal1 78158 -39619 78192 -39585 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.VGND
flabel nwell 78158 -39075 78192 -39041 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.VPB
flabel pwell 78158 -39619 78192 -39585 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x4.VNB
rlabel comment 78130 -39602 78130 -39602 4 16to4_PriorityEncoder_v0p0p1_0.x5.x4.or3_1
rlabel metal1 78130 -39650 78590 -39554 1 16to4_PriorityEncoder_v0p0p1_0.x5.x4.VGND
rlabel metal1 78130 -39106 78590 -39010 1 16to4_PriorityEncoder_v0p0p1_0.x5.x4.VPWR
flabel metal1 78619 -39075 78653 -39041 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.VPWR
flabel metal1 78619 -39619 78653 -39585 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.VGND
flabel locali 78987 -39449 79021 -39415 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.X
flabel locali 78987 -39517 79021 -39483 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.X
flabel locali 78987 -39381 79021 -39347 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.X
flabel locali 78987 -39313 79021 -39279 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.X
flabel locali 78987 -39245 79021 -39211 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.X
flabel locali 78987 -39177 79021 -39143 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.X
flabel locali 78803 -39381 78837 -39347 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.B
flabel locali 78711 -39381 78745 -39347 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.A
flabel locali 78619 -39381 78653 -39347 0 FreeSans 250 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.A
flabel nwell 78619 -39075 78653 -39041 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.VPB
flabel pwell 78619 -39619 78653 -39585 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x8.VNB
rlabel comment 78590 -39602 78590 -39602 4 16to4_PriorityEncoder_v0p0p1_0.x5.x8.and2_1
rlabel metal1 78590 -39650 79050 -39554 1 16to4_PriorityEncoder_v0p0p1_0.x5.x8.VGND
rlabel metal1 78590 -39106 79050 -39010 1 16to4_PriorityEncoder_v0p0p1_0.x5.x8.VPWR
flabel locali 76496 -38711 76530 -38677 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x3.Y
flabel locali 76496 -38643 76530 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x3.Y
flabel locali 76404 -38643 76438 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x3.A
flabel nwell 76361 -38949 76395 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x3.VPB
flabel pwell 76361 -38405 76395 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x3.VNB
flabel metal1 76361 -38405 76395 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x3.VGND
flabel metal1 76361 -38949 76395 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x3.VPWR
rlabel comment 76332 -38388 76332 -38388 2 16to4_PriorityEncoder_v0p0p1_0.x5.x3.inv_1
rlabel metal1 76332 -38436 76608 -38340 5 16to4_PriorityEncoder_v0p0p1_0.x5.x3.VGND
rlabel metal1 76332 -38980 76608 -38884 5 16to4_PriorityEncoder_v0p0p1_0.x5.x3.VPWR
flabel locali 76220 -38711 76254 -38677 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x5.Y
flabel locali 76220 -38643 76254 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x5.Y
flabel locali 76128 -38643 76162 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x5.A
flabel nwell 76085 -38949 76119 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x5.VPB
flabel pwell 76085 -38405 76119 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x5.VNB
flabel metal1 76085 -38405 76119 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x5.VGND
flabel metal1 76085 -38949 76119 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x5.VPWR
rlabel comment 76056 -38388 76056 -38388 2 16to4_PriorityEncoder_v0p0p1_0.x5.x5.inv_1
rlabel metal1 76056 -38436 76332 -38340 5 16to4_PriorityEncoder_v0p0p1_0.x5.x5.VGND
rlabel metal1 76056 -38980 76332 -38884 5 16to4_PriorityEncoder_v0p0p1_0.x5.x5.VPWR
flabel locali 75946 -38711 75980 -38677 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x6.Y
flabel locali 75946 -38643 75980 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x6.Y
flabel locali 75854 -38643 75888 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x6.A
flabel nwell 75811 -38949 75845 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x6.VPB
flabel pwell 75811 -38405 75845 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x6.VNB
flabel metal1 75811 -38405 75845 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x6.VGND
flabel metal1 75811 -38949 75845 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x6.VPWR
rlabel comment 75782 -38388 75782 -38388 2 16to4_PriorityEncoder_v0p0p1_0.x5.x6.inv_1
rlabel metal1 75782 -38436 76058 -38340 5 16to4_PriorityEncoder_v0p0p1_0.x5.x6.VGND
rlabel metal1 75782 -38980 76058 -38884 5 16to4_PriorityEncoder_v0p0p1_0.x5.x6.VPWR
flabel locali 75670 -38711 75704 -38677 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x7.Y
flabel locali 75670 -38643 75704 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x7.Y
flabel locali 75578 -38643 75612 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x7.A
flabel nwell 75535 -38949 75569 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x7.VPB
flabel pwell 75535 -38405 75569 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x7.VNB
flabel metal1 75535 -38405 75569 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x7.VGND
flabel metal1 75535 -38949 75569 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x7.VPWR
rlabel comment 75506 -38388 75506 -38388 2 16to4_PriorityEncoder_v0p0p1_0.x5.x7.inv_1
rlabel metal1 75506 -38436 75782 -38340 5 16to4_PriorityEncoder_v0p0p1_0.x5.x7.VGND
rlabel metal1 75506 -38980 75782 -38884 5 16to4_PriorityEncoder_v0p0p1_0.x5.x7.VPWR
flabel locali 76772 -38711 76806 -38677 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y
flabel locali 76772 -38643 76806 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y
flabel locali 76680 -38643 76714 -38609 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x9.A
flabel nwell 76637 -38949 76671 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x9.VPB
flabel pwell 76637 -38405 76671 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x9.VNB
flabel metal1 76637 -38405 76671 -38371 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x9.VGND
flabel metal1 76637 -38949 76671 -38915 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x5.x9.VPWR
rlabel comment 76608 -38388 76608 -38388 2 16to4_PriorityEncoder_v0p0p1_0.x5.x9.inv_1
rlabel metal1 76608 -38436 76884 -38340 5 16to4_PriorityEncoder_v0p0p1_0.x5.x9.VGND
rlabel metal1 76608 -38980 76884 -38884 5 16to4_PriorityEncoder_v0p0p1_0.x5.x9.VPWR
flabel locali 85351 -43931 85385 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.Y
flabel locali 85351 -43999 85385 -43965 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.Y
flabel locali 84063 -43931 84097 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.A
flabel locali 84431 -43931 84465 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.A
flabel locali 84799 -43931 84833 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.A
flabel locali 84891 -43931 84925 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.A
flabel nwell 84063 -43625 84097 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.VPB
flabel pwell 84063 -44169 84097 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.VNB
flabel metal1 84063 -44169 84097 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.VGND
flabel metal1 84063 -43625 84097 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x36.VPWR
rlabel comment 84034 -44152 84034 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x36.inv_16
rlabel metal1 84034 -44200 85506 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x36.VGND
rlabel metal1 84034 -43656 85506 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x36.VPWR
flabel locali 83971 -43999 84005 -43965 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.Y
flabel locali 83971 -43931 84005 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.Y
flabel locali 83971 -43863 84005 -43829 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.Y
flabel locali 83603 -43931 83637 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.A
flabel locali 83695 -43931 83729 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.A
flabel locali 83787 -43931 83821 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.A
flabel locali 83879 -43931 83913 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.A
flabel nwell 83603 -43625 83637 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.VPB
flabel pwell 83603 -44169 83637 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.VNB
flabel metal1 83603 -43625 83637 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.VPWR
flabel metal1 83603 -44169 83637 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x35.VGND
rlabel comment 83574 -44152 83574 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x35.inv_4
rlabel metal1 83574 -44200 84034 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x35.VGND
rlabel metal1 83574 -43656 84034 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x35.VPWR
flabel locali 83462 -43863 83496 -43829 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x34.Y
flabel locali 83462 -43931 83496 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x34.Y
flabel locali 83370 -43931 83404 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x34.A
flabel nwell 83327 -43625 83361 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x34.VPB
flabel pwell 83327 -44169 83361 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x34.VNB
flabel metal1 83327 -44169 83361 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x34.VGND
flabel metal1 83327 -43625 83361 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x34.VPWR
rlabel comment 83298 -44152 83298 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x34.inv_1
rlabel metal1 83298 -44200 83574 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x34.VGND
rlabel metal1 83298 -43656 83574 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x34.VPWR
flabel locali 83051 -43931 83085 -43897 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x11.A
flabel locali 83235 -43795 83269 -43761 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x11.X
flabel locali 82867 -43931 82901 -43897 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x11.B
flabel nwell 82867 -43625 82901 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x11.VPB
flabel pwell 82867 -44169 82901 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x11.VNB
flabel metal1 82867 -44169 82901 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x11.VGND
flabel metal1 82867 -43625 82901 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x11.VPWR
rlabel comment 82838 -44152 82838 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x11.or2_1
rlabel metal1 82838 -44200 83298 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x11.VGND
rlabel metal1 82838 -43656 83298 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x11.VPWR
flabel locali 86823 -43931 86857 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.Y
flabel locali 86823 -43999 86857 -43965 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.Y
flabel locali 85535 -43931 85569 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.A
flabel locali 85903 -43931 85937 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.A
flabel locali 86271 -43931 86305 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.A
flabel locali 86363 -43931 86397 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.A
flabel nwell 85535 -43625 85569 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.VPB
flabel pwell 85535 -44169 85569 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.VNB
flabel metal1 85535 -44169 85569 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.VGND
flabel metal1 85535 -43625 85569 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x10.VPWR
rlabel comment 85506 -44152 85506 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x10.inv_16
rlabel metal1 85506 -44200 86978 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x10.VGND
rlabel metal1 85506 -43656 86978 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x10.VPWR
flabel locali 88295 -43931 88329 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.Y
flabel locali 88295 -43999 88329 -43965 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.Y
flabel locali 87007 -43931 87041 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.A
flabel locali 87375 -43931 87409 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.A
flabel locali 87743 -43931 87777 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.A
flabel locali 87835 -43931 87869 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.A
flabel nwell 87007 -43625 87041 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.VPB
flabel pwell 87007 -44169 87041 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.VNB
flabel metal1 87007 -44169 87041 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.VGND
flabel metal1 87007 -43625 87041 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x12.VPWR
rlabel comment 86978 -44152 86978 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x12.inv_16
rlabel metal1 86978 -44200 88450 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x12.VGND
rlabel metal1 86978 -43656 88450 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x12.VPWR
flabel locali 80952 -40051 80986 -40017 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x7.Y
flabel locali 80952 -39983 80986 -39949 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x7.Y
flabel locali 80860 -39983 80894 -39949 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x7.A
flabel nwell 80817 -40289 80851 -40255 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x7.VPB
flabel pwell 80817 -39745 80851 -39711 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x7.VNB
flabel metal1 80817 -39745 80851 -39711 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x7.VGND
flabel metal1 80817 -40289 80851 -40255 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x7.VPWR
rlabel comment 80788 -39728 80788 -39728 2 16to4_PriorityEncoder_v0p0p1_0.x7.inv_1
rlabel metal1 80788 -39776 81064 -39680 5 16to4_PriorityEncoder_v0p0p1_0.x7.VGND
rlabel metal1 80788 -40320 81064 -40224 5 16to4_PriorityEncoder_v0p0p1_0.x7.VPWR
flabel locali 82791 -39431 82825 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.Y
flabel locali 82791 -39499 82825 -39465 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.Y
flabel locali 81503 -39431 81537 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.A
flabel locali 81871 -39431 81905 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.A
flabel locali 82239 -39431 82273 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.A
flabel locali 82331 -39431 82365 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.A
flabel nwell 81503 -39125 81537 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.VPB
flabel pwell 81503 -39669 81537 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.VNB
flabel metal1 81503 -39669 81537 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.VGND
flabel metal1 81503 -39125 81537 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x43.VPWR
rlabel comment 81474 -39652 81474 -39652 4 16to4_PriorityEncoder_v0p0p1_0.x43.inv_16
rlabel metal1 81474 -39700 82946 -39604 1 16to4_PriorityEncoder_v0p0p1_0.x43.VGND
rlabel metal1 81474 -39156 82946 -39060 1 16to4_PriorityEncoder_v0p0p1_0.x43.VPWR
flabel locali 81411 -39499 81445 -39465 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.Y
flabel locali 81411 -39431 81445 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.Y
flabel locali 81411 -39363 81445 -39329 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.Y
flabel locali 81043 -39431 81077 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.A
flabel locali 81135 -39431 81169 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.A
flabel locali 81227 -39431 81261 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.A
flabel locali 81319 -39431 81353 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.A
flabel nwell 81043 -39125 81077 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.VPB
flabel pwell 81043 -39669 81077 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.VNB
flabel metal1 81043 -39125 81077 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.VPWR
flabel metal1 81043 -39669 81077 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x42.VGND
rlabel comment 81014 -39652 81014 -39652 4 16to4_PriorityEncoder_v0p0p1_0.x42.inv_4
rlabel metal1 81014 -39700 81474 -39604 1 16to4_PriorityEncoder_v0p0p1_0.x42.VGND
rlabel metal1 81014 -39156 81474 -39060 1 16to4_PriorityEncoder_v0p0p1_0.x42.VPWR
flabel locali 80902 -39363 80936 -39329 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x41.Y
flabel locali 80902 -39431 80936 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x41.Y
flabel locali 80810 -39431 80844 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x41.A
flabel nwell 80767 -39125 80801 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x41.VPB
flabel pwell 80767 -39669 80801 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x41.VNB
flabel metal1 80767 -39669 80801 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x41.VGND
flabel metal1 80767 -39125 80801 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x41.VPWR
rlabel comment 80738 -39652 80738 -39652 4 16to4_PriorityEncoder_v0p0p1_0.x41.inv_1
rlabel metal1 80738 -39700 81014 -39604 1 16to4_PriorityEncoder_v0p0p1_0.x41.VGND
rlabel metal1 80738 -39156 81014 -39060 1 16to4_PriorityEncoder_v0p0p1_0.x41.VPWR
flabel locali 84263 -39431 84297 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.Y
flabel locali 84263 -39499 84297 -39465 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.Y
flabel locali 82975 -39431 83009 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.A
flabel locali 83343 -39431 83377 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.A
flabel locali 83711 -39431 83745 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.A
flabel locali 83803 -39431 83837 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.A
flabel nwell 82975 -39125 83009 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.VPB
flabel pwell 82975 -39669 83009 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.VNB
flabel metal1 82975 -39669 83009 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.VGND
flabel metal1 82975 -39125 83009 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x6.VPWR
rlabel comment 82946 -39652 82946 -39652 4 16to4_PriorityEncoder_v0p0p1_0.x6.inv_16
rlabel metal1 82946 -39700 84418 -39604 1 16to4_PriorityEncoder_v0p0p1_0.x6.VGND
rlabel metal1 82946 -39156 84418 -39060 1 16to4_PriorityEncoder_v0p0p1_0.x6.VPWR
flabel locali 85735 -39431 85769 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.Y
flabel locali 85735 -39499 85769 -39465 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.Y
flabel locali 84447 -39431 84481 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.A
flabel locali 84815 -39431 84849 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.A
flabel locali 85183 -39431 85217 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.A
flabel locali 85275 -39431 85309 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.A
flabel nwell 84447 -39125 84481 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.VPB
flabel pwell 84447 -39669 84481 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.VNB
flabel metal1 84447 -39669 84481 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.VGND
flabel metal1 84447 -39125 84481 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x4.VPWR
rlabel comment 84418 -39652 84418 -39652 4 16to4_PriorityEncoder_v0p0p1_0.x4.inv_16
rlabel metal1 84418 -39700 85890 -39604 1 16to4_PriorityEncoder_v0p0p1_0.x4.VGND
rlabel metal1 84418 -39156 85890 -39060 1 16to4_PriorityEncoder_v0p0p1_0.x4.VPWR
flabel locali 87207 -39431 87241 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.Y
flabel locali 87207 -39499 87241 -39465 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.Y
flabel locali 85919 -39431 85953 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.A
flabel locali 86287 -39431 86321 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.A
flabel locali 86655 -39431 86689 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.A
flabel locali 86747 -39431 86781 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.A
flabel nwell 85919 -39125 85953 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.VPB
flabel pwell 85919 -39669 85953 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.VNB
flabel metal1 85919 -39669 85953 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.VGND
flabel metal1 85919 -39125 85953 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x8.VPWR
rlabel comment 85890 -39652 85890 -39652 4 16to4_PriorityEncoder_v0p0p1_0.x8.inv_16
rlabel metal1 85890 -39700 87362 -39604 1 16to4_PriorityEncoder_v0p0p1_0.x8.VGND
rlabel metal1 85890 -39156 87362 -39060 1 16to4_PriorityEncoder_v0p0p1_0.x8.VPWR
flabel locali 88679 -39431 88713 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.Y
flabel locali 88679 -39499 88713 -39465 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.Y
flabel locali 87391 -39431 87425 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.A
flabel locali 87759 -39431 87793 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.A
flabel locali 88127 -39431 88161 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.A
flabel locali 88219 -39431 88253 -39397 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.A
flabel nwell 87391 -39125 87425 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.VPB
flabel pwell 87391 -39669 87425 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.VNB
flabel metal1 87391 -39669 87425 -39635 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.VGND
flabel metal1 87391 -39125 87425 -39091 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x9.VPWR
rlabel comment 87362 -39652 87362 -39652 4 16to4_PriorityEncoder_v0p0p1_0.x9.inv_16
rlabel metal1 87362 -39700 88834 -39604 1 16to4_PriorityEncoder_v0p0p1_0.x9.VGND
rlabel metal1 87362 -39156 88834 -39060 1 16to4_PriorityEncoder_v0p0p1_0.x9.VPWR
flabel locali 89767 -43931 89801 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.Y
flabel locali 89767 -43999 89801 -43965 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.Y
flabel locali 88479 -43931 88513 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.A
flabel locali 88847 -43931 88881 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.A
flabel locali 89215 -43931 89249 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.A
flabel locali 89307 -43931 89341 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.A
flabel nwell 88479 -43625 88513 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.VPB
flabel pwell 88479 -44169 88513 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.VNB
flabel metal1 88479 -44169 88513 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.VGND
flabel metal1 88479 -43625 88513 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x13.VPWR
rlabel comment 88450 -44152 88450 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x13.inv_16
rlabel metal1 88450 -44200 89922 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x13.VGND
rlabel metal1 88450 -43656 89922 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x13.VPWR
flabel locali 91239 -43931 91273 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.Y
flabel locali 91239 -43999 91273 -43965 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.Y
flabel locali 89951 -43931 89985 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.A
flabel locali 90319 -43931 90353 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.A
flabel locali 90687 -43931 90721 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.A
flabel locali 90779 -43931 90813 -43897 0 FreeSans 340 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.A
flabel nwell 89951 -43625 89985 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.VPB
flabel pwell 89951 -44169 89985 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.VNB
flabel metal1 89951 -44169 89985 -44135 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.VGND
flabel metal1 89951 -43625 89985 -43591 0 FreeSans 200 0 0 0 16to4_PriorityEncoder_v0p0p1_0.x14.VPWR
rlabel comment 89922 -44152 89922 -44152 4 16to4_PriorityEncoder_v0p0p1_0.x14.inv_16
rlabel metal1 89922 -44200 91394 -44104 1 16to4_PriorityEncoder_v0p0p1_0.x14.VGND
rlabel metal1 89922 -43656 91394 -43560 1 16to4_PriorityEncoder_v0p0p1_0.x14.VPWR
flabel metal1 21396 -7609 21596 -7409 0 FreeSans 256 0 0 0 PTAT_v0p0p0_mag_0.VDD
flabel metal1 25310 -11592 25510 -11392 0 FreeSans 256 0 0 0 PTAT_v0p0p0_mag_0.VOUT
flabel metal1 28410 -13092 28610 -12892 0 FreeSans 256 0 0 0 PTAT_v0p0p0_mag_0.VSS
flabel metal1 57096 -7160 57296 -6960 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.VDD
flabel metal1 53056 -9150 53256 -8950 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.GND
flabel metal1 53586 -7140 53786 -6940 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.IB
flabel metal1 55576 -6640 55776 -6440 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.VIN
flabel metal1 55706 -10800 55906 -10600 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.VN
flabel metal1 57036 -8590 57236 -8390 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.CLK
flabel metal1 59956 -10310 60156 -10110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.Q
flabel metal1 56510 -7338 56710 -7138 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.VDD
flabel metal4 53070 -8588 53270 -8388 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.VSS
flabel metal1 55580 -6638 55780 -6438 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.VIP
flabel metal1 56800 -7868 57000 -7668 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.VOP
flabel metal1 56800 -9358 57000 -9158 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.VON
flabel metal1 56860 -8588 57060 -8388 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.CLK
flabel metal1 55710 -10798 55910 -10598 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.VIN
flabel metal1 53590 -7118 53790 -6918 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.class_AB_v3_sym_0.IB
flabel metal1 57127 -8023 57161 -7989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.VGND
flabel metal1 57125 -7479 57159 -7445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.VPWR
flabel locali 57125 -7479 57159 -7445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.VPWR
flabel locali 57127 -8023 57161 -7989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.VGND
flabel locali 57307 -7921 57341 -7887 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.X
flabel locali 57307 -7649 57341 -7615 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.X
flabel locali 57307 -7581 57341 -7547 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.X
flabel locali 57125 -7785 57159 -7751 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.A
flabel nwell 57125 -7479 57159 -7445 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.VPB
flabel pwell 57127 -8023 57161 -7989 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x65.VNB
rlabel comment 57096 -8006 57096 -8006 4 frontAnalog_v0p0p1_0.x65.buf_1
rlabel metal1 57096 -8054 57372 -7958 1 frontAnalog_v0p0p1_0.x65.VGND
rlabel metal1 57096 -7510 57372 -7414 1 frontAnalog_v0p0p1_0.x65.VPWR
flabel metal1 57127 -8999 57161 -8965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.VGND
flabel metal1 57125 -9543 57159 -9509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.VPWR
flabel locali 57125 -9543 57159 -9509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.VPWR
flabel locali 57127 -8999 57161 -8965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.VGND
flabel locali 57307 -9101 57341 -9067 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.X
flabel locali 57307 -9373 57341 -9339 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.X
flabel locali 57307 -9441 57341 -9407 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.X
flabel locali 57125 -9237 57159 -9203 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.A
flabel nwell 57125 -9543 57159 -9509 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.VPB
flabel pwell 57127 -8999 57161 -8965 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.x63.VNB
rlabel comment 57096 -8982 57096 -8982 2 frontAnalog_v0p0p1_0.x63.buf_1
rlabel metal1 57096 -9030 57372 -8934 5 frontAnalog_v0p0p1_0.x63.VGND
rlabel metal1 57096 -9574 57372 -9478 5 frontAnalog_v0p0p1_0.x63.VPWR
flabel metal1 58556 -8660 58756 -8460 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.VDD
flabel metal1 61166 -8110 61366 -7910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.GND
flabel metal1 58956 -10190 59156 -9990 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.R
flabel metal1 58946 -7050 59146 -6850 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.S
flabel metal1 59956 -10310 60156 -10110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.Q
flabel metal1 60186 -7080 60386 -6880 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.QN
flabel locali 60297 -8759 60331 -8725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y
flabel locali 60365 -8759 60399 -8725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y
flabel locali 60433 -8759 60467 -8725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y
flabel locali 60365 -8391 60399 -8357 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.A
flabel locali 60365 -8483 60399 -8449 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.A
flabel locali 60365 -8575 60399 -8541 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.A
flabel locali 60365 -8667 60399 -8633 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.A
flabel nwell 60671 -8391 60705 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.VPB
flabel pwell 60127 -8391 60161 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.VNB
flabel metal1 60671 -8391 60705 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.VPWR
flabel metal1 60127 -8391 60161 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.VGND
rlabel comment 60144 -8328 60144 -8328 6 frontAnalog_v0p0p1_0.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -8788 60192 -8328 3 frontAnalog_v0p0p1_0.RSfetsym_0.x1.VGND
rlabel metal1 60640 -8788 60736 -8328 3 frontAnalog_v0p0p1_0.RSfetsym_0.x1.VPWR
flabel locali 61121 -8759 61155 -8725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y
flabel locali 61053 -8759 61087 -8725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y
flabel locali 60985 -8759 61019 -8725 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y
flabel locali 61053 -8391 61087 -8357 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.A
flabel locali 61053 -8483 61087 -8449 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.A
flabel locali 61053 -8575 61087 -8541 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.A
flabel locali 61053 -8667 61087 -8633 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.A
flabel nwell 60747 -8391 60781 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.VPB
flabel pwell 61291 -8391 61325 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.VNB
flabel metal1 60747 -8391 60781 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.VPWR
flabel metal1 61291 -8391 61325 -8357 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_0.RSfetsym_0.x2.VGND
rlabel comment 61308 -8328 61308 -8328 4 frontAnalog_v0p0p1_0.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -8788 61356 -8328 7 frontAnalog_v0p0p1_0.RSfetsym_0.x2.VGND
rlabel metal1 60716 -8788 60812 -8328 7 frontAnalog_v0p0p1_0.RSfetsym_0.x2.VPWR
flabel metal1 57096 -1760 57296 -1560 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.VDD
flabel metal1 53056 -3750 53256 -3550 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.GND
flabel metal1 53586 -1740 53786 -1540 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.IB
flabel metal1 55576 -1240 55776 -1040 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.VIN
flabel metal1 55706 -5400 55906 -5200 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.VN
flabel metal1 57036 -3190 57236 -2990 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.CLK
flabel metal1 59956 -4910 60156 -4710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.Q
flabel metal1 56510 -1938 56710 -1738 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.VDD
flabel metal4 53070 -3188 53270 -2988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.VSS
flabel metal1 55580 -1238 55780 -1038 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.VIP
flabel metal1 56800 -2468 57000 -2268 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.VOP
flabel metal1 56800 -3958 57000 -3758 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.VON
flabel metal1 56860 -3188 57060 -2988 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.CLK
flabel metal1 55710 -5398 55910 -5198 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.VIN
flabel metal1 53590 -1718 53790 -1518 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.class_AB_v3_sym_0.IB
flabel metal1 57127 -2623 57161 -2589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.VGND
flabel metal1 57125 -2079 57159 -2045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.VPWR
flabel locali 57125 -2079 57159 -2045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.VPWR
flabel locali 57127 -2623 57161 -2589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.VGND
flabel locali 57307 -2521 57341 -2487 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.X
flabel locali 57307 -2249 57341 -2215 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.X
flabel locali 57307 -2181 57341 -2147 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.X
flabel locali 57125 -2385 57159 -2351 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.A
flabel nwell 57125 -2079 57159 -2045 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.VPB
flabel pwell 57127 -2623 57161 -2589 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x65.VNB
rlabel comment 57096 -2606 57096 -2606 4 frontAnalog_v0p0p1_2.x65.buf_1
rlabel metal1 57096 -2654 57372 -2558 1 frontAnalog_v0p0p1_2.x65.VGND
rlabel metal1 57096 -2110 57372 -2014 1 frontAnalog_v0p0p1_2.x65.VPWR
flabel metal1 57127 -3599 57161 -3565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.VGND
flabel metal1 57125 -4143 57159 -4109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.VPWR
flabel locali 57125 -4143 57159 -4109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.VPWR
flabel locali 57127 -3599 57161 -3565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.VGND
flabel locali 57307 -3701 57341 -3667 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.X
flabel locali 57307 -3973 57341 -3939 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.X
flabel locali 57307 -4041 57341 -4007 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.X
flabel locali 57125 -3837 57159 -3803 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.A
flabel nwell 57125 -4143 57159 -4109 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.VPB
flabel pwell 57127 -3599 57161 -3565 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.x63.VNB
rlabel comment 57096 -3582 57096 -3582 2 frontAnalog_v0p0p1_2.x63.buf_1
rlabel metal1 57096 -3630 57372 -3534 5 frontAnalog_v0p0p1_2.x63.VGND
rlabel metal1 57096 -4174 57372 -4078 5 frontAnalog_v0p0p1_2.x63.VPWR
flabel metal1 58556 -3260 58756 -3060 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.VDD
flabel metal1 61166 -2710 61366 -2510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.GND
flabel metal1 58956 -4790 59156 -4590 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.R
flabel metal1 58946 -1650 59146 -1450 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.S
flabel metal1 59956 -4910 60156 -4710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.Q
flabel metal1 60186 -1680 60386 -1480 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.QN
flabel locali 60297 -3359 60331 -3325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y
flabel locali 60365 -3359 60399 -3325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y
flabel locali 60433 -3359 60467 -3325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y
flabel locali 60365 -2991 60399 -2957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.A
flabel locali 60365 -3083 60399 -3049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.A
flabel locali 60365 -3175 60399 -3141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.A
flabel locali 60365 -3267 60399 -3233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.A
flabel nwell 60671 -2991 60705 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.VPB
flabel pwell 60127 -2991 60161 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.VNB
flabel metal1 60671 -2991 60705 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.VPWR
flabel metal1 60127 -2991 60161 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.VGND
rlabel comment 60144 -2928 60144 -2928 6 frontAnalog_v0p0p1_2.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -3388 60192 -2928 3 frontAnalog_v0p0p1_2.RSfetsym_0.x1.VGND
rlabel metal1 60640 -3388 60736 -2928 3 frontAnalog_v0p0p1_2.RSfetsym_0.x1.VPWR
flabel locali 61121 -3359 61155 -3325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y
flabel locali 61053 -3359 61087 -3325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y
flabel locali 60985 -3359 61019 -3325 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y
flabel locali 61053 -2991 61087 -2957 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.A
flabel locali 61053 -3083 61087 -3049 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.A
flabel locali 61053 -3175 61087 -3141 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.A
flabel locali 61053 -3267 61087 -3233 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.A
flabel nwell 60747 -2991 60781 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.VPB
flabel pwell 61291 -2991 61325 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.VNB
flabel metal1 60747 -2991 60781 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.VPWR
flabel metal1 61291 -2991 61325 -2957 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_2.RSfetsym_0.x2.VGND
rlabel comment 61308 -2928 61308 -2928 4 frontAnalog_v0p0p1_2.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -3388 61356 -2928 7 frontAnalog_v0p0p1_2.RSfetsym_0.x2.VGND
rlabel metal1 60716 -3388 60812 -2928 7 frontAnalog_v0p0p1_2.RSfetsym_0.x2.VPWR
flabel metal1 57096 -12560 57296 -12360 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.VDD
flabel metal1 53056 -14550 53256 -14350 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.GND
flabel metal1 53586 -12540 53786 -12340 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.IB
flabel metal1 55576 -12040 55776 -11840 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.VIN
flabel metal1 55706 -16200 55906 -16000 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.VN
flabel metal1 57036 -13990 57236 -13790 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.CLK
flabel metal1 59956 -15710 60156 -15510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.Q
flabel metal1 56510 -12738 56710 -12538 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.VDD
flabel metal4 53070 -13988 53270 -13788 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.VSS
flabel metal1 55580 -12038 55780 -11838 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.VIP
flabel metal1 56800 -13268 57000 -13068 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.VOP
flabel metal1 56800 -14758 57000 -14558 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.VON
flabel metal1 56860 -13988 57060 -13788 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.CLK
flabel metal1 55710 -16198 55910 -15998 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.VIN
flabel metal1 53590 -12518 53790 -12318 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.class_AB_v3_sym_0.IB
flabel metal1 57127 -13423 57161 -13389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.VGND
flabel metal1 57125 -12879 57159 -12845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.VPWR
flabel locali 57125 -12879 57159 -12845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.VPWR
flabel locali 57127 -13423 57161 -13389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.VGND
flabel locali 57307 -13321 57341 -13287 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.X
flabel locali 57307 -13049 57341 -13015 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.X
flabel locali 57307 -12981 57341 -12947 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.X
flabel locali 57125 -13185 57159 -13151 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.A
flabel nwell 57125 -12879 57159 -12845 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.VPB
flabel pwell 57127 -13423 57161 -13389 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x65.VNB
rlabel comment 57096 -13406 57096 -13406 4 frontAnalog_v0p0p1_3.x65.buf_1
rlabel metal1 57096 -13454 57372 -13358 1 frontAnalog_v0p0p1_3.x65.VGND
rlabel metal1 57096 -12910 57372 -12814 1 frontAnalog_v0p0p1_3.x65.VPWR
flabel metal1 57127 -14399 57161 -14365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.VGND
flabel metal1 57125 -14943 57159 -14909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.VPWR
flabel locali 57125 -14943 57159 -14909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.VPWR
flabel locali 57127 -14399 57161 -14365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.VGND
flabel locali 57307 -14501 57341 -14467 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.X
flabel locali 57307 -14773 57341 -14739 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.X
flabel locali 57307 -14841 57341 -14807 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.X
flabel locali 57125 -14637 57159 -14603 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.A
flabel nwell 57125 -14943 57159 -14909 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.VPB
flabel pwell 57127 -14399 57161 -14365 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.x63.VNB
rlabel comment 57096 -14382 57096 -14382 2 frontAnalog_v0p0p1_3.x63.buf_1
rlabel metal1 57096 -14430 57372 -14334 5 frontAnalog_v0p0p1_3.x63.VGND
rlabel metal1 57096 -14974 57372 -14878 5 frontAnalog_v0p0p1_3.x63.VPWR
flabel metal1 58556 -14060 58756 -13860 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.VDD
flabel metal1 61166 -13510 61366 -13310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.GND
flabel metal1 58956 -15590 59156 -15390 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.R
flabel metal1 58946 -12450 59146 -12250 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.S
flabel metal1 59956 -15710 60156 -15510 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.Q
flabel metal1 60186 -12480 60386 -12280 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.QN
flabel locali 60297 -14159 60331 -14125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y
flabel locali 60365 -14159 60399 -14125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y
flabel locali 60433 -14159 60467 -14125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y
flabel locali 60365 -13791 60399 -13757 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.A
flabel locali 60365 -13883 60399 -13849 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.A
flabel locali 60365 -13975 60399 -13941 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.A
flabel locali 60365 -14067 60399 -14033 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.A
flabel nwell 60671 -13791 60705 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.VPB
flabel pwell 60127 -13791 60161 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.VNB
flabel metal1 60671 -13791 60705 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.VPWR
flabel metal1 60127 -13791 60161 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.VGND
rlabel comment 60144 -13728 60144 -13728 6 frontAnalog_v0p0p1_3.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -14188 60192 -13728 3 frontAnalog_v0p0p1_3.RSfetsym_0.x1.VGND
rlabel metal1 60640 -14188 60736 -13728 3 frontAnalog_v0p0p1_3.RSfetsym_0.x1.VPWR
flabel locali 61121 -14159 61155 -14125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y
flabel locali 61053 -14159 61087 -14125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y
flabel locali 60985 -14159 61019 -14125 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y
flabel locali 61053 -13791 61087 -13757 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.A
flabel locali 61053 -13883 61087 -13849 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.A
flabel locali 61053 -13975 61087 -13941 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.A
flabel locali 61053 -14067 61087 -14033 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.A
flabel nwell 60747 -13791 60781 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.VPB
flabel pwell 61291 -13791 61325 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.VNB
flabel metal1 60747 -13791 60781 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.VPWR
flabel metal1 61291 -13791 61325 -13757 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.VGND
rlabel comment 61308 -13728 61308 -13728 4 frontAnalog_v0p0p1_3.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -14188 61356 -13728 7 frontAnalog_v0p0p1_3.RSfetsym_0.x2.VGND
rlabel metal1 60716 -14188 60812 -13728 7 frontAnalog_v0p0p1_3.RSfetsym_0.x2.VPWR
flabel metal1 57096 -17960 57296 -17760 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.VDD
flabel metal1 53056 -19950 53256 -19750 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.GND
flabel metal1 53586 -17940 53786 -17740 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.IB
flabel metal1 55576 -17440 55776 -17240 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.VIN
flabel metal1 55706 -21600 55906 -21400 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.VN
flabel metal1 57036 -19390 57236 -19190 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.CLK
flabel metal1 59956 -21110 60156 -20910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.Q
flabel metal1 56510 -18138 56710 -17938 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.VDD
flabel metal4 53070 -19388 53270 -19188 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.VSS
flabel metal1 55580 -17438 55780 -17238 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.VIP
flabel metal1 56800 -18668 57000 -18468 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.VOP
flabel metal1 56800 -20158 57000 -19958 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.VON
flabel metal1 56860 -19388 57060 -19188 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.CLK
flabel metal1 55710 -21598 55910 -21398 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.VIN
flabel metal1 53590 -17918 53790 -17718 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.class_AB_v3_sym_0.IB
flabel metal1 57127 -18823 57161 -18789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.VGND
flabel metal1 57125 -18279 57159 -18245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.VPWR
flabel locali 57125 -18279 57159 -18245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.VPWR
flabel locali 57127 -18823 57161 -18789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.VGND
flabel locali 57307 -18721 57341 -18687 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.X
flabel locali 57307 -18449 57341 -18415 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.X
flabel locali 57307 -18381 57341 -18347 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.X
flabel locali 57125 -18585 57159 -18551 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.A
flabel nwell 57125 -18279 57159 -18245 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.VPB
flabel pwell 57127 -18823 57161 -18789 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x65.VNB
rlabel comment 57096 -18806 57096 -18806 4 frontAnalog_v0p0p1_4.x65.buf_1
rlabel metal1 57096 -18854 57372 -18758 1 frontAnalog_v0p0p1_4.x65.VGND
rlabel metal1 57096 -18310 57372 -18214 1 frontAnalog_v0p0p1_4.x65.VPWR
flabel metal1 57127 -19799 57161 -19765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.VGND
flabel metal1 57125 -20343 57159 -20309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.VPWR
flabel locali 57125 -20343 57159 -20309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.VPWR
flabel locali 57127 -19799 57161 -19765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.VGND
flabel locali 57307 -19901 57341 -19867 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.X
flabel locali 57307 -20173 57341 -20139 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.X
flabel locali 57307 -20241 57341 -20207 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.X
flabel locali 57125 -20037 57159 -20003 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.A
flabel nwell 57125 -20343 57159 -20309 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.VPB
flabel pwell 57127 -19799 57161 -19765 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.x63.VNB
rlabel comment 57096 -19782 57096 -19782 2 frontAnalog_v0p0p1_4.x63.buf_1
rlabel metal1 57096 -19830 57372 -19734 5 frontAnalog_v0p0p1_4.x63.VGND
rlabel metal1 57096 -20374 57372 -20278 5 frontAnalog_v0p0p1_4.x63.VPWR
flabel metal1 58556 -19460 58756 -19260 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.VDD
flabel metal1 61166 -18910 61366 -18710 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.GND
flabel metal1 58956 -20990 59156 -20790 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.R
flabel metal1 58946 -17850 59146 -17650 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.S
flabel metal1 59956 -21110 60156 -20910 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.Q
flabel metal1 60186 -17880 60386 -17680 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.QN
flabel locali 60297 -19559 60331 -19525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y
flabel locali 60365 -19559 60399 -19525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y
flabel locali 60433 -19559 60467 -19525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y
flabel locali 60365 -19191 60399 -19157 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.A
flabel locali 60365 -19283 60399 -19249 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.A
flabel locali 60365 -19375 60399 -19341 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.A
flabel locali 60365 -19467 60399 -19433 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.A
flabel nwell 60671 -19191 60705 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.VPB
flabel pwell 60127 -19191 60161 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.VNB
flabel metal1 60671 -19191 60705 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.VPWR
flabel metal1 60127 -19191 60161 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.VGND
rlabel comment 60144 -19128 60144 -19128 6 frontAnalog_v0p0p1_4.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -19588 60192 -19128 3 frontAnalog_v0p0p1_4.RSfetsym_0.x1.VGND
rlabel metal1 60640 -19588 60736 -19128 3 frontAnalog_v0p0p1_4.RSfetsym_0.x1.VPWR
flabel locali 61121 -19559 61155 -19525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y
flabel locali 61053 -19559 61087 -19525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y
flabel locali 60985 -19559 61019 -19525 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y
flabel locali 61053 -19191 61087 -19157 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.A
flabel locali 61053 -19283 61087 -19249 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.A
flabel locali 61053 -19375 61087 -19341 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.A
flabel locali 61053 -19467 61087 -19433 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.A
flabel nwell 60747 -19191 60781 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.VPB
flabel pwell 61291 -19191 61325 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.VNB
flabel metal1 60747 -19191 60781 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.VPWR
flabel metal1 61291 -19191 61325 -19157 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.VGND
rlabel comment 61308 -19128 61308 -19128 4 frontAnalog_v0p0p1_4.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -19588 61356 -19128 7 frontAnalog_v0p0p1_4.RSfetsym_0.x2.VGND
rlabel metal1 60716 -19588 60812 -19128 7 frontAnalog_v0p0p1_4.RSfetsym_0.x2.VPWR
flabel metal1 57096 -23360 57296 -23160 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.VDD
flabel metal1 53056 -25350 53256 -25150 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.GND
flabel metal1 53586 -23340 53786 -23140 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.IB
flabel metal1 55576 -22840 55776 -22640 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.VIN
flabel metal1 55706 -27000 55906 -26800 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.VN
flabel metal1 57036 -24790 57236 -24590 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.CLK
flabel metal1 59956 -26510 60156 -26310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.Q
flabel metal1 56510 -23538 56710 -23338 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.VDD
flabel metal4 53070 -24788 53270 -24588 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.VSS
flabel metal1 55580 -22838 55780 -22638 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.VIP
flabel metal1 56800 -24068 57000 -23868 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.VOP
flabel metal1 56800 -25558 57000 -25358 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.VON
flabel metal1 56860 -24788 57060 -24588 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.CLK
flabel metal1 55710 -26998 55910 -26798 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.VIN
flabel metal1 53590 -23318 53790 -23118 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.class_AB_v3_sym_0.IB
flabel metal1 57127 -24223 57161 -24189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.VGND
flabel metal1 57125 -23679 57159 -23645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.VPWR
flabel locali 57125 -23679 57159 -23645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.VPWR
flabel locali 57127 -24223 57161 -24189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.VGND
flabel locali 57307 -24121 57341 -24087 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.X
flabel locali 57307 -23849 57341 -23815 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.X
flabel locali 57307 -23781 57341 -23747 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.X
flabel locali 57125 -23985 57159 -23951 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.A
flabel nwell 57125 -23679 57159 -23645 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.VPB
flabel pwell 57127 -24223 57161 -24189 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x65.VNB
rlabel comment 57096 -24206 57096 -24206 4 frontAnalog_v0p0p1_5.x65.buf_1
rlabel metal1 57096 -24254 57372 -24158 1 frontAnalog_v0p0p1_5.x65.VGND
rlabel metal1 57096 -23710 57372 -23614 1 frontAnalog_v0p0p1_5.x65.VPWR
flabel metal1 57127 -25199 57161 -25165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.VGND
flabel metal1 57125 -25743 57159 -25709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.VPWR
flabel locali 57125 -25743 57159 -25709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.VPWR
flabel locali 57127 -25199 57161 -25165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.VGND
flabel locali 57307 -25301 57341 -25267 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.X
flabel locali 57307 -25573 57341 -25539 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.X
flabel locali 57307 -25641 57341 -25607 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.X
flabel locali 57125 -25437 57159 -25403 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.A
flabel nwell 57125 -25743 57159 -25709 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.VPB
flabel pwell 57127 -25199 57161 -25165 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.x63.VNB
rlabel comment 57096 -25182 57096 -25182 2 frontAnalog_v0p0p1_5.x63.buf_1
rlabel metal1 57096 -25230 57372 -25134 5 frontAnalog_v0p0p1_5.x63.VGND
rlabel metal1 57096 -25774 57372 -25678 5 frontAnalog_v0p0p1_5.x63.VPWR
flabel metal1 58556 -24860 58756 -24660 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.VDD
flabel metal1 61166 -24310 61366 -24110 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.GND
flabel metal1 58956 -26390 59156 -26190 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.R
flabel metal1 58946 -23250 59146 -23050 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.S
flabel metal1 59956 -26510 60156 -26310 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.Q
flabel metal1 60186 -23280 60386 -23080 0 FreeSans 256 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.QN
flabel locali 60297 -24959 60331 -24925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y
flabel locali 60365 -24959 60399 -24925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y
flabel locali 60433 -24959 60467 -24925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y
flabel locali 60365 -24591 60399 -24557 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.A
flabel locali 60365 -24683 60399 -24649 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.A
flabel locali 60365 -24775 60399 -24741 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.A
flabel locali 60365 -24867 60399 -24833 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.A
flabel nwell 60671 -24591 60705 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.VPB
flabel pwell 60127 -24591 60161 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.VNB
flabel metal1 60671 -24591 60705 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.VPWR
flabel metal1 60127 -24591 60161 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.VGND
rlabel comment 60144 -24528 60144 -24528 6 frontAnalog_v0p0p1_5.RSfetsym_0.x1.inv_4
rlabel metal1 60096 -24988 60192 -24528 3 frontAnalog_v0p0p1_5.RSfetsym_0.x1.VGND
rlabel metal1 60640 -24988 60736 -24528 3 frontAnalog_v0p0p1_5.RSfetsym_0.x1.VPWR
flabel locali 61121 -24959 61155 -24925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y
flabel locali 61053 -24959 61087 -24925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y
flabel locali 60985 -24959 61019 -24925 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y
flabel locali 61053 -24591 61087 -24557 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.A
flabel locali 61053 -24683 61087 -24649 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.A
flabel locali 61053 -24775 61087 -24741 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.A
flabel locali 61053 -24867 61087 -24833 0 FreeSans 340 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.A
flabel nwell 60747 -24591 60781 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.VPB
flabel pwell 61291 -24591 61325 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.VNB
flabel metal1 60747 -24591 60781 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.VPWR
flabel metal1 61291 -24591 61325 -24557 0 FreeSans 200 0 0 0 frontAnalog_v0p0p1_5.RSfetsym_0.x2.VGND
rlabel comment 61308 -24528 61308 -24528 4 frontAnalog_v0p0p1_5.RSfetsym_0.x2.inv_4
rlabel metal1 61260 -24988 61356 -24528 7 frontAnalog_v0p0p1_5.RSfetsym_0.x2.VGND
rlabel metal1 60716 -24988 60812 -24528 7 frontAnalog_v0p0p1_5.RSfetsym_0.x2.VPWR
<< end >>
