magic
tech sky130A
magscale 1 2
timestamp 1679514808
<< nwell >>
rect -6280 3640 6340 9080
<< pwell >>
rect -10013 3327 -6817 6275
rect -4320 2860 4408 3352
rect 7047 3327 10243 6275
rect -4320 2360 4408 2852
rect -3760 1760 3750 2352
rect -3760 1140 3750 1732
rect -4320 540 4408 1132
rect -4320 -60 4408 532
<< nmos >>
rect -4110 3056 -3110 3156
rect -2892 3056 -1892 3156
rect -1674 3056 -674 3156
rect -456 3056 544 3156
rect 762 3056 1762 3156
rect 1980 3056 2980 3156
rect 3198 3056 4198 3156
rect -4110 2556 -3110 2656
rect -2892 2556 -1892 2656
rect -1674 2556 -674 2656
rect -456 2556 544 2656
rect 762 2556 1762 2656
rect 1980 2556 2980 2656
rect 3198 2556 4198 2656
rect -3550 1956 -2550 2156
rect -2332 1956 -1332 2156
rect -1114 1956 -114 2156
rect 104 1956 1104 2156
rect 1322 1956 2322 2156
rect 2540 1956 3540 2156
rect -3550 1336 -2550 1536
rect -2332 1336 -1332 1536
rect -1114 1336 -114 1536
rect 104 1336 1104 1536
rect 1322 1336 2322 1536
rect 2540 1336 3540 1536
rect -4110 736 -3110 936
rect -2892 736 -1892 936
rect -1674 736 -674 936
rect -456 736 544 936
rect 762 736 1762 936
rect 1980 736 2980 936
rect 3198 736 4198 936
rect -4110 136 -3110 336
rect -2892 136 -1892 336
rect -1674 136 -674 336
rect -456 136 544 336
rect 762 136 1762 336
rect 1980 136 2980 336
rect 3198 136 4198 336
<< pmos >>
rect -4201 8776 -3201 8876
rect -2965 8776 -1965 8876
rect -1729 8776 -729 8876
rect -493 8776 507 8876
rect 743 8776 1743 8876
rect 1979 8776 2979 8876
rect 3215 8776 4215 8876
rect -4201 8236 -3201 8336
rect -2965 8236 -1965 8336
rect -1729 8236 -729 8336
rect -493 8236 507 8336
rect 743 8236 1743 8336
rect 1979 8236 2979 8336
rect 3215 8236 4215 8336
rect -4201 7696 -3201 7796
rect -2965 7696 -1965 7796
rect -1729 7696 -729 7796
rect -493 7696 507 7796
rect 743 7696 1743 7796
rect 1979 7696 2979 7796
rect 3215 7696 4215 7796
rect -4201 7156 -3201 7256
rect -2965 7156 -1965 7256
rect -1729 7156 -729 7256
rect -493 7156 507 7256
rect 743 7156 1743 7256
rect 1979 7156 2979 7256
rect 3215 7156 4215 7256
rect -4201 6576 -3201 6676
rect -2965 6576 -1965 6676
rect -1729 6576 -729 6676
rect -493 6576 507 6676
rect 743 6576 1743 6676
rect 1979 6576 2979 6676
rect 3215 6576 4215 6676
rect -4201 5996 -3201 6096
rect -2965 5996 -1965 6096
rect -1729 5996 -729 6096
rect -493 5996 507 6096
rect 743 5996 1743 6096
rect 1979 5996 2979 6096
rect 3215 5996 4215 6096
rect -6041 5456 -5041 5556
rect -4805 5456 -3805 5556
rect -3569 5456 -2569 5556
rect -2333 5456 -1333 5556
rect -1097 5456 -97 5556
rect 139 5456 1139 5556
rect 1375 5456 2375 5556
rect 2611 5456 3611 5556
rect 3847 5456 4847 5556
rect 5083 5456 6083 5556
rect -6041 4916 -5041 5016
rect -4805 4916 -3805 5016
rect -3569 4916 -2569 5016
rect -2333 4916 -1333 5016
rect -1097 4916 -97 5016
rect 139 4916 1139 5016
rect 1375 4916 2375 5016
rect 2611 4916 3611 5016
rect 3847 4916 4847 5016
rect 5083 4916 6083 5016
rect -6041 4376 -5041 4476
rect -4805 4376 -3805 4476
rect -3569 4376 -2569 4476
rect -2333 4376 -1333 4476
rect -1097 4376 -97 4476
rect 139 4376 1139 4476
rect 1375 4376 2375 4476
rect 2611 4376 3611 4476
rect 3847 4376 4847 4476
rect 5083 4376 6083 4476
rect -6041 3836 -5041 3936
rect -4805 3836 -3805 3936
rect -3569 3836 -2569 3936
rect -2333 3836 -1333 3936
rect -1097 3836 -97 3936
rect 139 3836 1139 3936
rect 1375 3836 2375 3936
rect 2611 3836 3611 3936
rect 3847 3836 4847 3936
rect 5083 3836 6083 3936
<< ndiff >>
rect -4110 3202 -3110 3214
rect -4110 3168 -4098 3202
rect -3122 3168 -3110 3202
rect -4110 3156 -3110 3168
rect -2892 3202 -1892 3214
rect -2892 3168 -2880 3202
rect -1904 3168 -1892 3202
rect -2892 3156 -1892 3168
rect -1674 3202 -674 3214
rect -1674 3168 -1662 3202
rect -686 3168 -674 3202
rect -1674 3156 -674 3168
rect -456 3202 544 3214
rect -456 3168 -444 3202
rect 532 3168 544 3202
rect -456 3156 544 3168
rect 762 3202 1762 3214
rect 762 3168 774 3202
rect 1750 3168 1762 3202
rect 762 3156 1762 3168
rect 1980 3202 2980 3214
rect 1980 3168 1992 3202
rect 2968 3168 2980 3202
rect 1980 3156 2980 3168
rect 3198 3202 4198 3214
rect 3198 3168 3210 3202
rect 4186 3168 4198 3202
rect 3198 3156 4198 3168
rect -4110 3044 -3110 3056
rect -4110 3010 -4098 3044
rect -3122 3010 -3110 3044
rect -4110 2998 -3110 3010
rect -2892 3044 -1892 3056
rect -2892 3010 -2880 3044
rect -1904 3010 -1892 3044
rect -2892 2998 -1892 3010
rect -1674 3044 -674 3056
rect -1674 3010 -1662 3044
rect -686 3010 -674 3044
rect -1674 2998 -674 3010
rect -456 3044 544 3056
rect -456 3010 -444 3044
rect 532 3010 544 3044
rect -456 2998 544 3010
rect 762 3044 1762 3056
rect 762 3010 774 3044
rect 1750 3010 1762 3044
rect 762 2998 1762 3010
rect 1980 3044 2980 3056
rect 1980 3010 1992 3044
rect 2968 3010 2980 3044
rect 1980 2998 2980 3010
rect 3198 3044 4198 3056
rect 3198 3010 3210 3044
rect 4186 3010 4198 3044
rect 3198 2998 4198 3010
rect -4110 2702 -3110 2714
rect -4110 2668 -4098 2702
rect -3122 2668 -3110 2702
rect -4110 2656 -3110 2668
rect -2892 2702 -1892 2714
rect -2892 2668 -2880 2702
rect -1904 2668 -1892 2702
rect -2892 2656 -1892 2668
rect -1674 2702 -674 2714
rect -1674 2668 -1662 2702
rect -686 2668 -674 2702
rect -1674 2656 -674 2668
rect -456 2702 544 2714
rect -456 2668 -444 2702
rect 532 2668 544 2702
rect -456 2656 544 2668
rect 762 2702 1762 2714
rect 762 2668 774 2702
rect 1750 2668 1762 2702
rect 762 2656 1762 2668
rect 1980 2702 2980 2714
rect 1980 2668 1992 2702
rect 2968 2668 2980 2702
rect 1980 2656 2980 2668
rect 3198 2702 4198 2714
rect 3198 2668 3210 2702
rect 4186 2668 4198 2702
rect 3198 2656 4198 2668
rect -4110 2544 -3110 2556
rect -4110 2510 -4098 2544
rect -3122 2510 -3110 2544
rect -4110 2498 -3110 2510
rect -2892 2544 -1892 2556
rect -2892 2510 -2880 2544
rect -1904 2510 -1892 2544
rect -2892 2498 -1892 2510
rect -1674 2544 -674 2556
rect -1674 2510 -1662 2544
rect -686 2510 -674 2544
rect -1674 2498 -674 2510
rect -456 2544 544 2556
rect -456 2510 -444 2544
rect 532 2510 544 2544
rect -456 2498 544 2510
rect 762 2544 1762 2556
rect 762 2510 774 2544
rect 1750 2510 1762 2544
rect 762 2498 1762 2510
rect 1980 2544 2980 2556
rect 1980 2510 1992 2544
rect 2968 2510 2980 2544
rect 1980 2498 2980 2510
rect 3198 2544 4198 2556
rect 3198 2510 3210 2544
rect 4186 2510 4198 2544
rect 3198 2498 4198 2510
rect -3550 2202 -2550 2214
rect -3550 2168 -3538 2202
rect -2562 2168 -2550 2202
rect -3550 2156 -2550 2168
rect -2332 2202 -1332 2214
rect -2332 2168 -2320 2202
rect -1344 2168 -1332 2202
rect -2332 2156 -1332 2168
rect -1114 2202 -114 2214
rect -1114 2168 -1102 2202
rect -126 2168 -114 2202
rect -1114 2156 -114 2168
rect 104 2202 1104 2214
rect 104 2168 116 2202
rect 1092 2168 1104 2202
rect 104 2156 1104 2168
rect 1322 2202 2322 2214
rect 1322 2168 1334 2202
rect 2310 2168 2322 2202
rect 1322 2156 2322 2168
rect 2540 2202 3540 2214
rect 2540 2168 2552 2202
rect 3528 2168 3540 2202
rect 2540 2156 3540 2168
rect -3550 1944 -2550 1956
rect -3550 1910 -3538 1944
rect -2562 1910 -2550 1944
rect -3550 1898 -2550 1910
rect -2332 1944 -1332 1956
rect -2332 1910 -2320 1944
rect -1344 1910 -1332 1944
rect -2332 1898 -1332 1910
rect -1114 1944 -114 1956
rect -1114 1910 -1102 1944
rect -126 1910 -114 1944
rect -1114 1898 -114 1910
rect 104 1944 1104 1956
rect 104 1910 116 1944
rect 1092 1910 1104 1944
rect 104 1898 1104 1910
rect 1322 1944 2322 1956
rect 1322 1910 1334 1944
rect 2310 1910 2322 1944
rect 1322 1898 2322 1910
rect 2540 1944 3540 1956
rect 2540 1910 2552 1944
rect 3528 1910 3540 1944
rect 2540 1898 3540 1910
rect -3550 1582 -2550 1594
rect -3550 1548 -3538 1582
rect -2562 1548 -2550 1582
rect -3550 1536 -2550 1548
rect -2332 1582 -1332 1594
rect -2332 1548 -2320 1582
rect -1344 1548 -1332 1582
rect -2332 1536 -1332 1548
rect -1114 1582 -114 1594
rect -1114 1548 -1102 1582
rect -126 1548 -114 1582
rect -1114 1536 -114 1548
rect 104 1582 1104 1594
rect 104 1548 116 1582
rect 1092 1548 1104 1582
rect 104 1536 1104 1548
rect 1322 1582 2322 1594
rect 1322 1548 1334 1582
rect 2310 1548 2322 1582
rect 1322 1536 2322 1548
rect 2540 1582 3540 1594
rect 2540 1548 2552 1582
rect 3528 1548 3540 1582
rect 2540 1536 3540 1548
rect -3550 1324 -2550 1336
rect -3550 1290 -3538 1324
rect -2562 1290 -2550 1324
rect -3550 1278 -2550 1290
rect -2332 1324 -1332 1336
rect -2332 1290 -2320 1324
rect -1344 1290 -1332 1324
rect -2332 1278 -1332 1290
rect -1114 1324 -114 1336
rect -1114 1290 -1102 1324
rect -126 1290 -114 1324
rect -1114 1278 -114 1290
rect 104 1324 1104 1336
rect 104 1290 116 1324
rect 1092 1290 1104 1324
rect 104 1278 1104 1290
rect 1322 1324 2322 1336
rect 1322 1290 1334 1324
rect 2310 1290 2322 1324
rect 1322 1278 2322 1290
rect 2540 1324 3540 1336
rect 2540 1290 2552 1324
rect 3528 1290 3540 1324
rect 2540 1278 3540 1290
rect -4110 982 -3110 994
rect -4110 948 -4098 982
rect -3122 948 -3110 982
rect -4110 936 -3110 948
rect -2892 982 -1892 994
rect -2892 948 -2880 982
rect -1904 948 -1892 982
rect -2892 936 -1892 948
rect -1674 982 -674 994
rect -1674 948 -1662 982
rect -686 948 -674 982
rect -1674 936 -674 948
rect -456 982 544 994
rect -456 948 -444 982
rect 532 948 544 982
rect -456 936 544 948
rect 762 982 1762 994
rect 762 948 774 982
rect 1750 948 1762 982
rect 762 936 1762 948
rect 1980 982 2980 994
rect 1980 948 1992 982
rect 2968 948 2980 982
rect 1980 936 2980 948
rect 3198 982 4198 994
rect 3198 948 3210 982
rect 4186 948 4198 982
rect 3198 936 4198 948
rect -4110 724 -3110 736
rect -4110 690 -4098 724
rect -3122 690 -3110 724
rect -4110 678 -3110 690
rect -2892 724 -1892 736
rect -2892 690 -2880 724
rect -1904 690 -1892 724
rect -2892 678 -1892 690
rect -1674 724 -674 736
rect -1674 690 -1662 724
rect -686 690 -674 724
rect -1674 678 -674 690
rect -456 724 544 736
rect -456 690 -444 724
rect 532 690 544 724
rect -456 678 544 690
rect 762 724 1762 736
rect 762 690 774 724
rect 1750 690 1762 724
rect 762 678 1762 690
rect 1980 724 2980 736
rect 1980 690 1992 724
rect 2968 690 2980 724
rect 1980 678 2980 690
rect 3198 724 4198 736
rect 3198 690 3210 724
rect 4186 690 4198 724
rect 3198 678 4198 690
rect -4110 382 -3110 394
rect -4110 348 -4098 382
rect -3122 348 -3110 382
rect -4110 336 -3110 348
rect -2892 382 -1892 394
rect -2892 348 -2880 382
rect -1904 348 -1892 382
rect -2892 336 -1892 348
rect -1674 382 -674 394
rect -1674 348 -1662 382
rect -686 348 -674 382
rect -1674 336 -674 348
rect -456 382 544 394
rect -456 348 -444 382
rect 532 348 544 382
rect -456 336 544 348
rect 762 382 1762 394
rect 762 348 774 382
rect 1750 348 1762 382
rect 762 336 1762 348
rect 1980 382 2980 394
rect 1980 348 1992 382
rect 2968 348 2980 382
rect 1980 336 2980 348
rect 3198 382 4198 394
rect 3198 348 3210 382
rect 4186 348 4198 382
rect 3198 336 4198 348
rect -4110 124 -3110 136
rect -4110 90 -4098 124
rect -3122 90 -3110 124
rect -4110 78 -3110 90
rect -2892 124 -1892 136
rect -2892 90 -2880 124
rect -1904 90 -1892 124
rect -2892 78 -1892 90
rect -1674 124 -674 136
rect -1674 90 -1662 124
rect -686 90 -674 124
rect -1674 78 -674 90
rect -456 124 544 136
rect -456 90 -444 124
rect 532 90 544 124
rect -456 78 544 90
rect 762 124 1762 136
rect 762 90 774 124
rect 1750 90 1762 124
rect 762 78 1762 90
rect 1980 124 2980 136
rect 1980 90 1992 124
rect 2968 90 2980 124
rect 1980 78 2980 90
rect 3198 124 4198 136
rect 3198 90 3210 124
rect 4186 90 4198 124
rect 3198 78 4198 90
<< pdiff >>
rect -4201 8922 -3201 8934
rect -4201 8888 -4189 8922
rect -3213 8888 -3201 8922
rect -4201 8876 -3201 8888
rect -2965 8922 -1965 8934
rect -2965 8888 -2953 8922
rect -1977 8888 -1965 8922
rect -2965 8876 -1965 8888
rect -1729 8922 -729 8934
rect -1729 8888 -1717 8922
rect -741 8888 -729 8922
rect -1729 8876 -729 8888
rect -493 8922 507 8934
rect -493 8888 -481 8922
rect 495 8888 507 8922
rect -493 8876 507 8888
rect 743 8922 1743 8934
rect 743 8888 755 8922
rect 1731 8888 1743 8922
rect 743 8876 1743 8888
rect 1979 8922 2979 8934
rect 1979 8888 1991 8922
rect 2967 8888 2979 8922
rect 1979 8876 2979 8888
rect 3215 8922 4215 8934
rect 3215 8888 3227 8922
rect 4203 8888 4215 8922
rect 3215 8876 4215 8888
rect -4201 8764 -3201 8776
rect -4201 8730 -4189 8764
rect -3213 8730 -3201 8764
rect -4201 8718 -3201 8730
rect -2965 8764 -1965 8776
rect -2965 8730 -2953 8764
rect -1977 8730 -1965 8764
rect -2965 8718 -1965 8730
rect -1729 8764 -729 8776
rect -1729 8730 -1717 8764
rect -741 8730 -729 8764
rect -1729 8718 -729 8730
rect -493 8764 507 8776
rect -493 8730 -481 8764
rect 495 8730 507 8764
rect -493 8718 507 8730
rect 743 8764 1743 8776
rect 743 8730 755 8764
rect 1731 8730 1743 8764
rect 743 8718 1743 8730
rect 1979 8764 2979 8776
rect 1979 8730 1991 8764
rect 2967 8730 2979 8764
rect 1979 8718 2979 8730
rect 3215 8764 4215 8776
rect 3215 8730 3227 8764
rect 4203 8730 4215 8764
rect 3215 8718 4215 8730
rect -4201 8382 -3201 8394
rect -4201 8348 -4189 8382
rect -3213 8348 -3201 8382
rect -4201 8336 -3201 8348
rect -2965 8382 -1965 8394
rect -2965 8348 -2953 8382
rect -1977 8348 -1965 8382
rect -2965 8336 -1965 8348
rect -1729 8382 -729 8394
rect -1729 8348 -1717 8382
rect -741 8348 -729 8382
rect -1729 8336 -729 8348
rect -493 8382 507 8394
rect -493 8348 -481 8382
rect 495 8348 507 8382
rect -493 8336 507 8348
rect 743 8382 1743 8394
rect 743 8348 755 8382
rect 1731 8348 1743 8382
rect 743 8336 1743 8348
rect 1979 8382 2979 8394
rect 1979 8348 1991 8382
rect 2967 8348 2979 8382
rect 1979 8336 2979 8348
rect 3215 8382 4215 8394
rect 3215 8348 3227 8382
rect 4203 8348 4215 8382
rect 3215 8336 4215 8348
rect -4201 8224 -3201 8236
rect -4201 8190 -4189 8224
rect -3213 8190 -3201 8224
rect -4201 8178 -3201 8190
rect -2965 8224 -1965 8236
rect -2965 8190 -2953 8224
rect -1977 8190 -1965 8224
rect -2965 8178 -1965 8190
rect -1729 8224 -729 8236
rect -1729 8190 -1717 8224
rect -741 8190 -729 8224
rect -1729 8178 -729 8190
rect -493 8224 507 8236
rect -493 8190 -481 8224
rect 495 8190 507 8224
rect -493 8178 507 8190
rect 743 8224 1743 8236
rect 743 8190 755 8224
rect 1731 8190 1743 8224
rect 743 8178 1743 8190
rect 1979 8224 2979 8236
rect 1979 8190 1991 8224
rect 2967 8190 2979 8224
rect 1979 8178 2979 8190
rect 3215 8224 4215 8236
rect 3215 8190 3227 8224
rect 4203 8190 4215 8224
rect 3215 8178 4215 8190
rect -4201 7842 -3201 7854
rect -4201 7808 -4189 7842
rect -3213 7808 -3201 7842
rect -4201 7796 -3201 7808
rect -2965 7842 -1965 7854
rect -2965 7808 -2953 7842
rect -1977 7808 -1965 7842
rect -2965 7796 -1965 7808
rect -1729 7842 -729 7854
rect -1729 7808 -1717 7842
rect -741 7808 -729 7842
rect -1729 7796 -729 7808
rect -493 7842 507 7854
rect -493 7808 -481 7842
rect 495 7808 507 7842
rect -493 7796 507 7808
rect 743 7842 1743 7854
rect 743 7808 755 7842
rect 1731 7808 1743 7842
rect 743 7796 1743 7808
rect 1979 7842 2979 7854
rect 1979 7808 1991 7842
rect 2967 7808 2979 7842
rect 1979 7796 2979 7808
rect 3215 7842 4215 7854
rect 3215 7808 3227 7842
rect 4203 7808 4215 7842
rect 3215 7796 4215 7808
rect -4201 7684 -3201 7696
rect -4201 7650 -4189 7684
rect -3213 7650 -3201 7684
rect -4201 7638 -3201 7650
rect -2965 7684 -1965 7696
rect -2965 7650 -2953 7684
rect -1977 7650 -1965 7684
rect -2965 7638 -1965 7650
rect -1729 7684 -729 7696
rect -1729 7650 -1717 7684
rect -741 7650 -729 7684
rect -1729 7638 -729 7650
rect -493 7684 507 7696
rect -493 7650 -481 7684
rect 495 7650 507 7684
rect -493 7638 507 7650
rect 743 7684 1743 7696
rect 743 7650 755 7684
rect 1731 7650 1743 7684
rect 743 7638 1743 7650
rect 1979 7684 2979 7696
rect 1979 7650 1991 7684
rect 2967 7650 2979 7684
rect 1979 7638 2979 7650
rect 3215 7684 4215 7696
rect 3215 7650 3227 7684
rect 4203 7650 4215 7684
rect 3215 7638 4215 7650
rect -4201 7302 -3201 7314
rect -4201 7268 -4189 7302
rect -3213 7268 -3201 7302
rect -4201 7256 -3201 7268
rect -2965 7302 -1965 7314
rect -2965 7268 -2953 7302
rect -1977 7268 -1965 7302
rect -2965 7256 -1965 7268
rect -1729 7302 -729 7314
rect -1729 7268 -1717 7302
rect -741 7268 -729 7302
rect -1729 7256 -729 7268
rect -493 7302 507 7314
rect -493 7268 -481 7302
rect 495 7268 507 7302
rect -493 7256 507 7268
rect 743 7302 1743 7314
rect 743 7268 755 7302
rect 1731 7268 1743 7302
rect 743 7256 1743 7268
rect 1979 7302 2979 7314
rect 1979 7268 1991 7302
rect 2967 7268 2979 7302
rect 1979 7256 2979 7268
rect 3215 7302 4215 7314
rect 3215 7268 3227 7302
rect 4203 7268 4215 7302
rect 3215 7256 4215 7268
rect -4201 7144 -3201 7156
rect -4201 7110 -4189 7144
rect -3213 7110 -3201 7144
rect -4201 7098 -3201 7110
rect -2965 7144 -1965 7156
rect -2965 7110 -2953 7144
rect -1977 7110 -1965 7144
rect -2965 7098 -1965 7110
rect -1729 7144 -729 7156
rect -1729 7110 -1717 7144
rect -741 7110 -729 7144
rect -1729 7098 -729 7110
rect -493 7144 507 7156
rect -493 7110 -481 7144
rect 495 7110 507 7144
rect -493 7098 507 7110
rect 743 7144 1743 7156
rect 743 7110 755 7144
rect 1731 7110 1743 7144
rect 743 7098 1743 7110
rect 1979 7144 2979 7156
rect 1979 7110 1991 7144
rect 2967 7110 2979 7144
rect 1979 7098 2979 7110
rect 3215 7144 4215 7156
rect 3215 7110 3227 7144
rect 4203 7110 4215 7144
rect 3215 7098 4215 7110
rect -4201 6722 -3201 6734
rect -4201 6688 -4189 6722
rect -3213 6688 -3201 6722
rect -4201 6676 -3201 6688
rect -2965 6722 -1965 6734
rect -2965 6688 -2953 6722
rect -1977 6688 -1965 6722
rect -2965 6676 -1965 6688
rect -1729 6722 -729 6734
rect -1729 6688 -1717 6722
rect -741 6688 -729 6722
rect -1729 6676 -729 6688
rect -493 6722 507 6734
rect -493 6688 -481 6722
rect 495 6688 507 6722
rect -493 6676 507 6688
rect 743 6722 1743 6734
rect 743 6688 755 6722
rect 1731 6688 1743 6722
rect 743 6676 1743 6688
rect 1979 6722 2979 6734
rect 1979 6688 1991 6722
rect 2967 6688 2979 6722
rect 1979 6676 2979 6688
rect 3215 6722 4215 6734
rect 3215 6688 3227 6722
rect 4203 6688 4215 6722
rect 3215 6676 4215 6688
rect -4201 6564 -3201 6576
rect -4201 6530 -4189 6564
rect -3213 6530 -3201 6564
rect -4201 6518 -3201 6530
rect -2965 6564 -1965 6576
rect -2965 6530 -2953 6564
rect -1977 6530 -1965 6564
rect -2965 6518 -1965 6530
rect -1729 6564 -729 6576
rect -1729 6530 -1717 6564
rect -741 6530 -729 6564
rect -1729 6518 -729 6530
rect -493 6564 507 6576
rect -493 6530 -481 6564
rect 495 6530 507 6564
rect -493 6518 507 6530
rect 743 6564 1743 6576
rect 743 6530 755 6564
rect 1731 6530 1743 6564
rect 743 6518 1743 6530
rect 1979 6564 2979 6576
rect 1979 6530 1991 6564
rect 2967 6530 2979 6564
rect 1979 6518 2979 6530
rect 3215 6564 4215 6576
rect 3215 6530 3227 6564
rect 4203 6530 4215 6564
rect 3215 6518 4215 6530
rect -4201 6142 -3201 6154
rect -4201 6108 -4189 6142
rect -3213 6108 -3201 6142
rect -4201 6096 -3201 6108
rect -2965 6142 -1965 6154
rect -2965 6108 -2953 6142
rect -1977 6108 -1965 6142
rect -2965 6096 -1965 6108
rect -1729 6142 -729 6154
rect -1729 6108 -1717 6142
rect -741 6108 -729 6142
rect -1729 6096 -729 6108
rect -493 6142 507 6154
rect -493 6108 -481 6142
rect 495 6108 507 6142
rect -493 6096 507 6108
rect 743 6142 1743 6154
rect 743 6108 755 6142
rect 1731 6108 1743 6142
rect 743 6096 1743 6108
rect 1979 6142 2979 6154
rect 1979 6108 1991 6142
rect 2967 6108 2979 6142
rect 1979 6096 2979 6108
rect 3215 6142 4215 6154
rect 3215 6108 3227 6142
rect 4203 6108 4215 6142
rect 3215 6096 4215 6108
rect -4201 5984 -3201 5996
rect -4201 5950 -4189 5984
rect -3213 5950 -3201 5984
rect -4201 5938 -3201 5950
rect -2965 5984 -1965 5996
rect -2965 5950 -2953 5984
rect -1977 5950 -1965 5984
rect -2965 5938 -1965 5950
rect -1729 5984 -729 5996
rect -1729 5950 -1717 5984
rect -741 5950 -729 5984
rect -1729 5938 -729 5950
rect -493 5984 507 5996
rect -493 5950 -481 5984
rect 495 5950 507 5984
rect -493 5938 507 5950
rect 743 5984 1743 5996
rect 743 5950 755 5984
rect 1731 5950 1743 5984
rect 743 5938 1743 5950
rect 1979 5984 2979 5996
rect 1979 5950 1991 5984
rect 2967 5950 2979 5984
rect 1979 5938 2979 5950
rect 3215 5984 4215 5996
rect 3215 5950 3227 5984
rect 4203 5950 4215 5984
rect 3215 5938 4215 5950
rect -6041 5602 -5041 5614
rect -6041 5568 -6029 5602
rect -5053 5568 -5041 5602
rect -6041 5556 -5041 5568
rect -4805 5602 -3805 5614
rect -4805 5568 -4793 5602
rect -3817 5568 -3805 5602
rect -4805 5556 -3805 5568
rect -3569 5602 -2569 5614
rect -3569 5568 -3557 5602
rect -2581 5568 -2569 5602
rect -3569 5556 -2569 5568
rect -2333 5602 -1333 5614
rect -2333 5568 -2321 5602
rect -1345 5568 -1333 5602
rect -2333 5556 -1333 5568
rect -1097 5602 -97 5614
rect -1097 5568 -1085 5602
rect -109 5568 -97 5602
rect -1097 5556 -97 5568
rect 139 5602 1139 5614
rect 139 5568 151 5602
rect 1127 5568 1139 5602
rect 139 5556 1139 5568
rect 1375 5602 2375 5614
rect 1375 5568 1387 5602
rect 2363 5568 2375 5602
rect 1375 5556 2375 5568
rect 2611 5602 3611 5614
rect 2611 5568 2623 5602
rect 3599 5568 3611 5602
rect 2611 5556 3611 5568
rect 3847 5602 4847 5614
rect 3847 5568 3859 5602
rect 4835 5568 4847 5602
rect 3847 5556 4847 5568
rect 5083 5602 6083 5614
rect 5083 5568 5095 5602
rect 6071 5568 6083 5602
rect 5083 5556 6083 5568
rect -6041 5444 -5041 5456
rect -6041 5410 -6029 5444
rect -5053 5410 -5041 5444
rect -6041 5398 -5041 5410
rect -4805 5444 -3805 5456
rect -4805 5410 -4793 5444
rect -3817 5410 -3805 5444
rect -4805 5398 -3805 5410
rect -3569 5444 -2569 5456
rect -3569 5410 -3557 5444
rect -2581 5410 -2569 5444
rect -3569 5398 -2569 5410
rect -2333 5444 -1333 5456
rect -2333 5410 -2321 5444
rect -1345 5410 -1333 5444
rect -2333 5398 -1333 5410
rect -1097 5444 -97 5456
rect -1097 5410 -1085 5444
rect -109 5410 -97 5444
rect -1097 5398 -97 5410
rect 139 5444 1139 5456
rect 139 5410 151 5444
rect 1127 5410 1139 5444
rect 139 5398 1139 5410
rect 1375 5444 2375 5456
rect 1375 5410 1387 5444
rect 2363 5410 2375 5444
rect 1375 5398 2375 5410
rect 2611 5444 3611 5456
rect 2611 5410 2623 5444
rect 3599 5410 3611 5444
rect 2611 5398 3611 5410
rect 3847 5444 4847 5456
rect 3847 5410 3859 5444
rect 4835 5410 4847 5444
rect 3847 5398 4847 5410
rect 5083 5444 6083 5456
rect 5083 5410 5095 5444
rect 6071 5410 6083 5444
rect 5083 5398 6083 5410
rect -6041 5062 -5041 5074
rect -6041 5028 -6029 5062
rect -5053 5028 -5041 5062
rect -6041 5016 -5041 5028
rect -4805 5062 -3805 5074
rect -4805 5028 -4793 5062
rect -3817 5028 -3805 5062
rect -4805 5016 -3805 5028
rect -3569 5062 -2569 5074
rect -3569 5028 -3557 5062
rect -2581 5028 -2569 5062
rect -3569 5016 -2569 5028
rect -2333 5062 -1333 5074
rect -2333 5028 -2321 5062
rect -1345 5028 -1333 5062
rect -2333 5016 -1333 5028
rect -1097 5062 -97 5074
rect -1097 5028 -1085 5062
rect -109 5028 -97 5062
rect -1097 5016 -97 5028
rect 139 5062 1139 5074
rect 139 5028 151 5062
rect 1127 5028 1139 5062
rect 139 5016 1139 5028
rect 1375 5062 2375 5074
rect 1375 5028 1387 5062
rect 2363 5028 2375 5062
rect 1375 5016 2375 5028
rect 2611 5062 3611 5074
rect 2611 5028 2623 5062
rect 3599 5028 3611 5062
rect 2611 5016 3611 5028
rect 3847 5062 4847 5074
rect 3847 5028 3859 5062
rect 4835 5028 4847 5062
rect 3847 5016 4847 5028
rect 5083 5062 6083 5074
rect 5083 5028 5095 5062
rect 6071 5028 6083 5062
rect 5083 5016 6083 5028
rect -6041 4904 -5041 4916
rect -6041 4870 -6029 4904
rect -5053 4870 -5041 4904
rect -6041 4858 -5041 4870
rect -4805 4904 -3805 4916
rect -4805 4870 -4793 4904
rect -3817 4870 -3805 4904
rect -4805 4858 -3805 4870
rect -3569 4904 -2569 4916
rect -3569 4870 -3557 4904
rect -2581 4870 -2569 4904
rect -3569 4858 -2569 4870
rect -2333 4904 -1333 4916
rect -2333 4870 -2321 4904
rect -1345 4870 -1333 4904
rect -2333 4858 -1333 4870
rect -1097 4904 -97 4916
rect -1097 4870 -1085 4904
rect -109 4870 -97 4904
rect -1097 4858 -97 4870
rect 139 4904 1139 4916
rect 139 4870 151 4904
rect 1127 4870 1139 4904
rect 139 4858 1139 4870
rect 1375 4904 2375 4916
rect 1375 4870 1387 4904
rect 2363 4870 2375 4904
rect 1375 4858 2375 4870
rect 2611 4904 3611 4916
rect 2611 4870 2623 4904
rect 3599 4870 3611 4904
rect 2611 4858 3611 4870
rect 3847 4904 4847 4916
rect 3847 4870 3859 4904
rect 4835 4870 4847 4904
rect 3847 4858 4847 4870
rect 5083 4904 6083 4916
rect 5083 4870 5095 4904
rect 6071 4870 6083 4904
rect 5083 4858 6083 4870
rect -6041 4522 -5041 4534
rect -6041 4488 -6029 4522
rect -5053 4488 -5041 4522
rect -6041 4476 -5041 4488
rect -4805 4522 -3805 4534
rect -4805 4488 -4793 4522
rect -3817 4488 -3805 4522
rect -4805 4476 -3805 4488
rect -3569 4522 -2569 4534
rect -3569 4488 -3557 4522
rect -2581 4488 -2569 4522
rect -3569 4476 -2569 4488
rect -2333 4522 -1333 4534
rect -2333 4488 -2321 4522
rect -1345 4488 -1333 4522
rect -2333 4476 -1333 4488
rect -1097 4522 -97 4534
rect -1097 4488 -1085 4522
rect -109 4488 -97 4522
rect -1097 4476 -97 4488
rect 139 4522 1139 4534
rect 139 4488 151 4522
rect 1127 4488 1139 4522
rect 139 4476 1139 4488
rect 1375 4522 2375 4534
rect 1375 4488 1387 4522
rect 2363 4488 2375 4522
rect 1375 4476 2375 4488
rect 2611 4522 3611 4534
rect 2611 4488 2623 4522
rect 3599 4488 3611 4522
rect 2611 4476 3611 4488
rect 3847 4522 4847 4534
rect 3847 4488 3859 4522
rect 4835 4488 4847 4522
rect 3847 4476 4847 4488
rect 5083 4522 6083 4534
rect 5083 4488 5095 4522
rect 6071 4488 6083 4522
rect 5083 4476 6083 4488
rect -6041 4364 -5041 4376
rect -6041 4330 -6029 4364
rect -5053 4330 -5041 4364
rect -6041 4318 -5041 4330
rect -4805 4364 -3805 4376
rect -4805 4330 -4793 4364
rect -3817 4330 -3805 4364
rect -4805 4318 -3805 4330
rect -3569 4364 -2569 4376
rect -3569 4330 -3557 4364
rect -2581 4330 -2569 4364
rect -3569 4318 -2569 4330
rect -2333 4364 -1333 4376
rect -2333 4330 -2321 4364
rect -1345 4330 -1333 4364
rect -2333 4318 -1333 4330
rect -1097 4364 -97 4376
rect -1097 4330 -1085 4364
rect -109 4330 -97 4364
rect -1097 4318 -97 4330
rect 139 4364 1139 4376
rect 139 4330 151 4364
rect 1127 4330 1139 4364
rect 139 4318 1139 4330
rect 1375 4364 2375 4376
rect 1375 4330 1387 4364
rect 2363 4330 2375 4364
rect 1375 4318 2375 4330
rect 2611 4364 3611 4376
rect 2611 4330 2623 4364
rect 3599 4330 3611 4364
rect 2611 4318 3611 4330
rect 3847 4364 4847 4376
rect 3847 4330 3859 4364
rect 4835 4330 4847 4364
rect 3847 4318 4847 4330
rect 5083 4364 6083 4376
rect 5083 4330 5095 4364
rect 6071 4330 6083 4364
rect 5083 4318 6083 4330
rect -6041 3982 -5041 3994
rect -6041 3948 -6029 3982
rect -5053 3948 -5041 3982
rect -6041 3936 -5041 3948
rect -4805 3982 -3805 3994
rect -4805 3948 -4793 3982
rect -3817 3948 -3805 3982
rect -4805 3936 -3805 3948
rect -3569 3982 -2569 3994
rect -3569 3948 -3557 3982
rect -2581 3948 -2569 3982
rect -3569 3936 -2569 3948
rect -2333 3982 -1333 3994
rect -2333 3948 -2321 3982
rect -1345 3948 -1333 3982
rect -2333 3936 -1333 3948
rect -1097 3982 -97 3994
rect -1097 3948 -1085 3982
rect -109 3948 -97 3982
rect -1097 3936 -97 3948
rect 139 3982 1139 3994
rect 139 3948 151 3982
rect 1127 3948 1139 3982
rect 139 3936 1139 3948
rect 1375 3982 2375 3994
rect 1375 3948 1387 3982
rect 2363 3948 2375 3982
rect 1375 3936 2375 3948
rect 2611 3982 3611 3994
rect 2611 3948 2623 3982
rect 3599 3948 3611 3982
rect 2611 3936 3611 3948
rect 3847 3982 4847 3994
rect 3847 3948 3859 3982
rect 4835 3948 4847 3982
rect 3847 3936 4847 3948
rect 5083 3982 6083 3994
rect 5083 3948 5095 3982
rect 6071 3948 6083 3982
rect 5083 3936 6083 3948
rect -6041 3824 -5041 3836
rect -6041 3790 -6029 3824
rect -5053 3790 -5041 3824
rect -6041 3778 -5041 3790
rect -4805 3824 -3805 3836
rect -4805 3790 -4793 3824
rect -3817 3790 -3805 3824
rect -4805 3778 -3805 3790
rect -3569 3824 -2569 3836
rect -3569 3790 -3557 3824
rect -2581 3790 -2569 3824
rect -3569 3778 -2569 3790
rect -2333 3824 -1333 3836
rect -2333 3790 -2321 3824
rect -1345 3790 -1333 3824
rect -2333 3778 -1333 3790
rect -1097 3824 -97 3836
rect -1097 3790 -1085 3824
rect -109 3790 -97 3824
rect -1097 3778 -97 3790
rect 139 3824 1139 3836
rect 139 3790 151 3824
rect 1127 3790 1139 3824
rect 139 3778 1139 3790
rect 1375 3824 2375 3836
rect 1375 3790 1387 3824
rect 2363 3790 2375 3824
rect 1375 3778 2375 3790
rect 2611 3824 3611 3836
rect 2611 3790 2623 3824
rect 3599 3790 3611 3824
rect 2611 3778 3611 3790
rect 3847 3824 4847 3836
rect 3847 3790 3859 3824
rect 4835 3790 4847 3824
rect 3847 3778 4847 3790
rect 5083 3824 6083 3836
rect 5083 3790 5095 3824
rect 6071 3790 6083 3824
rect 5083 3778 6083 3790
<< ndiffc >>
rect -4098 3168 -3122 3202
rect -2880 3168 -1904 3202
rect -1662 3168 -686 3202
rect -444 3168 532 3202
rect 774 3168 1750 3202
rect 1992 3168 2968 3202
rect 3210 3168 4186 3202
rect -4098 3010 -3122 3044
rect -2880 3010 -1904 3044
rect -1662 3010 -686 3044
rect -444 3010 532 3044
rect 774 3010 1750 3044
rect 1992 3010 2968 3044
rect 3210 3010 4186 3044
rect -4098 2668 -3122 2702
rect -2880 2668 -1904 2702
rect -1662 2668 -686 2702
rect -444 2668 532 2702
rect 774 2668 1750 2702
rect 1992 2668 2968 2702
rect 3210 2668 4186 2702
rect -4098 2510 -3122 2544
rect -2880 2510 -1904 2544
rect -1662 2510 -686 2544
rect -444 2510 532 2544
rect 774 2510 1750 2544
rect 1992 2510 2968 2544
rect 3210 2510 4186 2544
rect -3538 2168 -2562 2202
rect -2320 2168 -1344 2202
rect -1102 2168 -126 2202
rect 116 2168 1092 2202
rect 1334 2168 2310 2202
rect 2552 2168 3528 2202
rect -3538 1910 -2562 1944
rect -2320 1910 -1344 1944
rect -1102 1910 -126 1944
rect 116 1910 1092 1944
rect 1334 1910 2310 1944
rect 2552 1910 3528 1944
rect -3538 1548 -2562 1582
rect -2320 1548 -1344 1582
rect -1102 1548 -126 1582
rect 116 1548 1092 1582
rect 1334 1548 2310 1582
rect 2552 1548 3528 1582
rect -3538 1290 -2562 1324
rect -2320 1290 -1344 1324
rect -1102 1290 -126 1324
rect 116 1290 1092 1324
rect 1334 1290 2310 1324
rect 2552 1290 3528 1324
rect -4098 948 -3122 982
rect -2880 948 -1904 982
rect -1662 948 -686 982
rect -444 948 532 982
rect 774 948 1750 982
rect 1992 948 2968 982
rect 3210 948 4186 982
rect -4098 690 -3122 724
rect -2880 690 -1904 724
rect -1662 690 -686 724
rect -444 690 532 724
rect 774 690 1750 724
rect 1992 690 2968 724
rect 3210 690 4186 724
rect -4098 348 -3122 382
rect -2880 348 -1904 382
rect -1662 348 -686 382
rect -444 348 532 382
rect 774 348 1750 382
rect 1992 348 2968 382
rect 3210 348 4186 382
rect -4098 90 -3122 124
rect -2880 90 -1904 124
rect -1662 90 -686 124
rect -444 90 532 124
rect 774 90 1750 124
rect 1992 90 2968 124
rect 3210 90 4186 124
<< pdiffc >>
rect -4189 8888 -3213 8922
rect -2953 8888 -1977 8922
rect -1717 8888 -741 8922
rect -481 8888 495 8922
rect 755 8888 1731 8922
rect 1991 8888 2967 8922
rect 3227 8888 4203 8922
rect -4189 8730 -3213 8764
rect -2953 8730 -1977 8764
rect -1717 8730 -741 8764
rect -481 8730 495 8764
rect 755 8730 1731 8764
rect 1991 8730 2967 8764
rect 3227 8730 4203 8764
rect -4189 8348 -3213 8382
rect -2953 8348 -1977 8382
rect -1717 8348 -741 8382
rect -481 8348 495 8382
rect 755 8348 1731 8382
rect 1991 8348 2967 8382
rect 3227 8348 4203 8382
rect -4189 8190 -3213 8224
rect -2953 8190 -1977 8224
rect -1717 8190 -741 8224
rect -481 8190 495 8224
rect 755 8190 1731 8224
rect 1991 8190 2967 8224
rect 3227 8190 4203 8224
rect -4189 7808 -3213 7842
rect -2953 7808 -1977 7842
rect -1717 7808 -741 7842
rect -481 7808 495 7842
rect 755 7808 1731 7842
rect 1991 7808 2967 7842
rect 3227 7808 4203 7842
rect -4189 7650 -3213 7684
rect -2953 7650 -1977 7684
rect -1717 7650 -741 7684
rect -481 7650 495 7684
rect 755 7650 1731 7684
rect 1991 7650 2967 7684
rect 3227 7650 4203 7684
rect -4189 7268 -3213 7302
rect -2953 7268 -1977 7302
rect -1717 7268 -741 7302
rect -481 7268 495 7302
rect 755 7268 1731 7302
rect 1991 7268 2967 7302
rect 3227 7268 4203 7302
rect -4189 7110 -3213 7144
rect -2953 7110 -1977 7144
rect -1717 7110 -741 7144
rect -481 7110 495 7144
rect 755 7110 1731 7144
rect 1991 7110 2967 7144
rect 3227 7110 4203 7144
rect -4189 6688 -3213 6722
rect -2953 6688 -1977 6722
rect -1717 6688 -741 6722
rect -481 6688 495 6722
rect 755 6688 1731 6722
rect 1991 6688 2967 6722
rect 3227 6688 4203 6722
rect -4189 6530 -3213 6564
rect -2953 6530 -1977 6564
rect -1717 6530 -741 6564
rect -481 6530 495 6564
rect 755 6530 1731 6564
rect 1991 6530 2967 6564
rect 3227 6530 4203 6564
rect -4189 6108 -3213 6142
rect -2953 6108 -1977 6142
rect -1717 6108 -741 6142
rect -481 6108 495 6142
rect 755 6108 1731 6142
rect 1991 6108 2967 6142
rect 3227 6108 4203 6142
rect -4189 5950 -3213 5984
rect -2953 5950 -1977 5984
rect -1717 5950 -741 5984
rect -481 5950 495 5984
rect 755 5950 1731 5984
rect 1991 5950 2967 5984
rect 3227 5950 4203 5984
rect -6029 5568 -5053 5602
rect -4793 5568 -3817 5602
rect -3557 5568 -2581 5602
rect -2321 5568 -1345 5602
rect -1085 5568 -109 5602
rect 151 5568 1127 5602
rect 1387 5568 2363 5602
rect 2623 5568 3599 5602
rect 3859 5568 4835 5602
rect 5095 5568 6071 5602
rect -6029 5410 -5053 5444
rect -4793 5410 -3817 5444
rect -3557 5410 -2581 5444
rect -2321 5410 -1345 5444
rect -1085 5410 -109 5444
rect 151 5410 1127 5444
rect 1387 5410 2363 5444
rect 2623 5410 3599 5444
rect 3859 5410 4835 5444
rect 5095 5410 6071 5444
rect -6029 5028 -5053 5062
rect -4793 5028 -3817 5062
rect -3557 5028 -2581 5062
rect -2321 5028 -1345 5062
rect -1085 5028 -109 5062
rect 151 5028 1127 5062
rect 1387 5028 2363 5062
rect 2623 5028 3599 5062
rect 3859 5028 4835 5062
rect 5095 5028 6071 5062
rect -6029 4870 -5053 4904
rect -4793 4870 -3817 4904
rect -3557 4870 -2581 4904
rect -2321 4870 -1345 4904
rect -1085 4870 -109 4904
rect 151 4870 1127 4904
rect 1387 4870 2363 4904
rect 2623 4870 3599 4904
rect 3859 4870 4835 4904
rect 5095 4870 6071 4904
rect -6029 4488 -5053 4522
rect -4793 4488 -3817 4522
rect -3557 4488 -2581 4522
rect -2321 4488 -1345 4522
rect -1085 4488 -109 4522
rect 151 4488 1127 4522
rect 1387 4488 2363 4522
rect 2623 4488 3599 4522
rect 3859 4488 4835 4522
rect 5095 4488 6071 4522
rect -6029 4330 -5053 4364
rect -4793 4330 -3817 4364
rect -3557 4330 -2581 4364
rect -2321 4330 -1345 4364
rect -1085 4330 -109 4364
rect 151 4330 1127 4364
rect 1387 4330 2363 4364
rect 2623 4330 3599 4364
rect 3859 4330 4835 4364
rect 5095 4330 6071 4364
rect -6029 3948 -5053 3982
rect -4793 3948 -3817 3982
rect -3557 3948 -2581 3982
rect -2321 3948 -1345 3982
rect -1085 3948 -109 3982
rect 151 3948 1127 3982
rect 1387 3948 2363 3982
rect 2623 3948 3599 3982
rect 3859 3948 4835 3982
rect 5095 3948 6071 3982
rect -6029 3790 -5053 3824
rect -4793 3790 -3817 3824
rect -3557 3790 -2581 3824
rect -2321 3790 -1345 3824
rect -1085 3790 -109 3824
rect 151 3790 1127 3824
rect 1387 3790 2363 3824
rect 2623 3790 3599 3824
rect 3859 3790 4835 3824
rect 5095 3790 6071 3824
<< psubdiff >>
rect -9977 6205 -9881 6239
rect -6949 6205 -6853 6239
rect -9977 6143 -9943 6205
rect -6887 6143 -6853 6205
rect -9977 4867 -9943 4929
rect 7083 6205 7179 6239
rect 10111 6205 10207 6239
rect 7083 6143 7117 6205
rect -6887 4867 -6853 4929
rect -9977 4833 -9881 4867
rect -6949 4833 -6853 4867
rect 10173 6143 10207 6205
rect 7083 4867 7117 4929
rect 10173 4867 10207 4929
rect 7083 4833 7179 4867
rect 10111 4833 10207 4867
rect -9977 4735 -9881 4769
rect -6949 4735 -6853 4769
rect -9977 4673 -9943 4735
rect -6887 4673 -6853 4735
rect -9977 3397 -9943 3459
rect 7083 4735 7179 4769
rect 10111 4735 10207 4769
rect 7083 4673 7117 4735
rect -6887 3397 -6853 3459
rect -9977 3363 -9881 3397
rect -6949 3363 -6853 3397
rect 10173 4673 10207 4735
rect 7083 3397 7117 3459
rect 10173 3397 10207 3459
rect 7083 3363 7179 3397
rect 10111 3363 10207 3397
rect -4284 3282 -4188 3316
rect 4276 3282 4372 3316
rect -4284 3220 -4250 3282
rect 4338 3220 4372 3282
rect -4284 2930 -4250 2992
rect 4338 2930 4372 2992
rect -4284 2896 -4188 2930
rect 4276 2896 4372 2930
rect -4284 2782 -4188 2816
rect 4276 2782 4372 2816
rect -4284 2720 -4250 2782
rect 4338 2720 4372 2782
rect -4284 2430 -4250 2492
rect 4338 2430 4372 2492
rect -4284 2396 -4188 2430
rect 4276 2396 4372 2430
rect -3724 2282 -3628 2316
rect 3618 2282 3714 2316
rect -3724 2220 -3690 2282
rect 3680 2220 3714 2282
rect -3724 1830 -3690 1892
rect 3680 1830 3714 1892
rect -3724 1796 -3628 1830
rect 3618 1796 3714 1830
rect -3724 1662 -3628 1696
rect 3618 1662 3714 1696
rect -3724 1600 -3690 1662
rect 3680 1600 3714 1662
rect -3724 1210 -3690 1272
rect 3680 1210 3714 1272
rect -3724 1176 -3628 1210
rect 3618 1176 3714 1210
rect -4284 1062 -4188 1096
rect 4276 1062 4372 1096
rect -4284 1000 -4250 1062
rect 4338 1000 4372 1062
rect -4284 610 -4250 672
rect 4338 610 4372 672
rect -4284 576 -4188 610
rect 4276 576 4372 610
rect -4284 462 -4188 496
rect 4276 462 4372 496
rect -4284 400 -4250 462
rect 4338 400 4372 462
rect -4284 10 -4250 72
rect 4338 10 4372 72
rect -4284 -24 -4188 10
rect 4276 -24 4372 10
<< nsubdiff >>
rect -4384 9002 -4288 9036
rect 4302 9002 4398 9036
rect -4384 8940 -4350 9002
rect 4364 8940 4398 9002
rect -4384 8650 -4350 8712
rect 4364 8650 4398 8712
rect -4384 8616 -4288 8650
rect 4302 8616 4398 8650
rect -4384 8462 -4288 8496
rect 4302 8462 4398 8496
rect -4384 8400 -4350 8462
rect 4364 8400 4398 8462
rect -4384 8110 -4350 8172
rect 4364 8110 4398 8172
rect -4384 8076 -4288 8110
rect 4302 8076 4398 8110
rect -4384 7922 -4288 7956
rect 4302 7922 4398 7956
rect -4384 7860 -4350 7922
rect 4364 7860 4398 7922
rect -4384 7570 -4350 7632
rect 4364 7570 4398 7632
rect -4384 7536 -4288 7570
rect 4302 7536 4398 7570
rect -4384 7382 -4288 7416
rect 4302 7382 4398 7416
rect -4384 7320 -4350 7382
rect 4364 7320 4398 7382
rect -4384 7030 -4350 7092
rect 4364 7030 4398 7092
rect -4384 6996 -4288 7030
rect 4302 6996 4398 7030
rect -4384 6802 -4288 6836
rect 4302 6802 4398 6836
rect -4384 6740 -4350 6802
rect 4364 6740 4398 6802
rect -4384 6450 -4350 6512
rect 4364 6450 4398 6512
rect -4384 6416 -4288 6450
rect 4302 6416 4398 6450
rect -4384 6222 -4288 6256
rect 4302 6222 4398 6256
rect -4384 6160 -4350 6222
rect 4364 6160 4398 6222
rect -4384 5870 -4350 5932
rect 4364 5870 4398 5932
rect -4384 5836 -4288 5870
rect 4302 5836 4398 5870
rect -6224 5682 -6128 5716
rect 6170 5682 6266 5716
rect -6224 5620 -6190 5682
rect 6232 5620 6266 5682
rect -6224 5330 -6190 5392
rect 6232 5330 6266 5392
rect -6224 5296 -6128 5330
rect 6170 5296 6266 5330
rect -6224 5142 -6128 5176
rect 6170 5142 6266 5176
rect -6224 5080 -6190 5142
rect 6232 5080 6266 5142
rect -6224 4790 -6190 4852
rect 6232 4790 6266 4852
rect -6224 4756 -6128 4790
rect 6170 4756 6266 4790
rect -6224 4602 -6128 4636
rect 6170 4602 6266 4636
rect -6224 4540 -6190 4602
rect 6232 4540 6266 4602
rect -6224 4250 -6190 4312
rect 6232 4250 6266 4312
rect -6224 4216 -6128 4250
rect 6170 4216 6266 4250
rect -6224 4062 -6128 4096
rect 6170 4062 6266 4096
rect -6224 4000 -6190 4062
rect 6232 4000 6266 4062
rect -6224 3710 -6190 3772
rect 6232 3710 6266 3772
rect -6224 3676 -6128 3710
rect 6170 3676 6266 3710
<< psubdiffcont >>
rect -9881 6205 -6949 6239
rect -9977 4929 -9943 6143
rect -6887 4929 -6853 6143
rect 7179 6205 10111 6239
rect -9881 4833 -6949 4867
rect 7083 4929 7117 6143
rect 10173 4929 10207 6143
rect 7179 4833 10111 4867
rect -9881 4735 -6949 4769
rect -9977 3459 -9943 4673
rect -6887 3459 -6853 4673
rect 7179 4735 10111 4769
rect -9881 3363 -6949 3397
rect 7083 3459 7117 4673
rect 10173 3459 10207 4673
rect 7179 3363 10111 3397
rect -4188 3282 4276 3316
rect -4284 2992 -4250 3220
rect 4338 2992 4372 3220
rect -4188 2896 4276 2930
rect -4188 2782 4276 2816
rect -4284 2492 -4250 2720
rect 4338 2492 4372 2720
rect -4188 2396 4276 2430
rect -3628 2282 3618 2316
rect -3724 1892 -3690 2220
rect 3680 1892 3714 2220
rect -3628 1796 3618 1830
rect -3628 1662 3618 1696
rect -3724 1272 -3690 1600
rect 3680 1272 3714 1600
rect -3628 1176 3618 1210
rect -4188 1062 4276 1096
rect -4284 672 -4250 1000
rect 4338 672 4372 1000
rect -4188 576 4276 610
rect -4188 462 4276 496
rect -4284 72 -4250 400
rect 4338 72 4372 400
rect -4188 -24 4276 10
<< nsubdiffcont >>
rect -4288 9002 4302 9036
rect -4384 8712 -4350 8940
rect 4364 8712 4398 8940
rect -4288 8616 4302 8650
rect -4288 8462 4302 8496
rect -4384 8172 -4350 8400
rect 4364 8172 4398 8400
rect -4288 8076 4302 8110
rect -4288 7922 4302 7956
rect -4384 7632 -4350 7860
rect 4364 7632 4398 7860
rect -4288 7536 4302 7570
rect -4288 7382 4302 7416
rect -4384 7092 -4350 7320
rect 4364 7092 4398 7320
rect -4288 6996 4302 7030
rect -4288 6802 4302 6836
rect -4384 6512 -4350 6740
rect 4364 6512 4398 6740
rect -4288 6416 4302 6450
rect -4288 6222 4302 6256
rect -4384 5932 -4350 6160
rect 4364 5932 4398 6160
rect -4288 5836 4302 5870
rect -6128 5682 6170 5716
rect -6224 5392 -6190 5620
rect 6232 5392 6266 5620
rect -6128 5296 6170 5330
rect -6128 5142 6170 5176
rect -6224 4852 -6190 5080
rect 6232 4852 6266 5080
rect -6128 4756 6170 4790
rect -6128 4602 6170 4636
rect -6224 4312 -6190 4540
rect 6232 4312 6266 4540
rect -6128 4216 6170 4250
rect -6128 4062 6170 4096
rect -6224 3772 -6190 4000
rect 6232 3772 6266 4000
rect -6128 3676 6170 3710
<< poly >>
rect -4298 8860 -4201 8876
rect -4298 8792 -4282 8860
rect -4248 8792 -4201 8860
rect -4298 8776 -4201 8792
rect -3201 8860 -3104 8876
rect -3201 8792 -3154 8860
rect -3120 8792 -3104 8860
rect -3201 8776 -3104 8792
rect -3062 8860 -2965 8876
rect -3062 8792 -3046 8860
rect -3012 8792 -2965 8860
rect -3062 8776 -2965 8792
rect -1965 8860 -1868 8876
rect -1965 8792 -1918 8860
rect -1884 8792 -1868 8860
rect -1965 8776 -1868 8792
rect -1826 8860 -1729 8876
rect -1826 8792 -1810 8860
rect -1776 8792 -1729 8860
rect -1826 8776 -1729 8792
rect -729 8860 -632 8876
rect -729 8792 -682 8860
rect -648 8792 -632 8860
rect -729 8776 -632 8792
rect -590 8860 -493 8876
rect -590 8792 -574 8860
rect -540 8792 -493 8860
rect -590 8776 -493 8792
rect 507 8860 604 8876
rect 507 8792 554 8860
rect 588 8792 604 8860
rect 507 8776 604 8792
rect 646 8860 743 8876
rect 646 8792 662 8860
rect 696 8792 743 8860
rect 646 8776 743 8792
rect 1743 8860 1840 8876
rect 1743 8792 1790 8860
rect 1824 8792 1840 8860
rect 1743 8776 1840 8792
rect 1882 8860 1979 8876
rect 1882 8792 1898 8860
rect 1932 8792 1979 8860
rect 1882 8776 1979 8792
rect 2979 8860 3076 8876
rect 2979 8792 3026 8860
rect 3060 8792 3076 8860
rect 2979 8776 3076 8792
rect 3118 8860 3215 8876
rect 3118 8792 3134 8860
rect 3168 8792 3215 8860
rect 3118 8776 3215 8792
rect 4215 8860 4312 8876
rect 4215 8792 4262 8860
rect 4296 8792 4312 8860
rect 4215 8776 4312 8792
rect -4298 8320 -4201 8336
rect -4298 8252 -4282 8320
rect -4248 8252 -4201 8320
rect -4298 8236 -4201 8252
rect -3201 8320 -3104 8336
rect -3201 8252 -3154 8320
rect -3120 8252 -3104 8320
rect -3201 8236 -3104 8252
rect -3062 8320 -2965 8336
rect -3062 8252 -3046 8320
rect -3012 8252 -2965 8320
rect -3062 8236 -2965 8252
rect -1965 8320 -1868 8336
rect -1965 8252 -1918 8320
rect -1884 8252 -1868 8320
rect -1965 8236 -1868 8252
rect -1826 8320 -1729 8336
rect -1826 8252 -1810 8320
rect -1776 8252 -1729 8320
rect -1826 8236 -1729 8252
rect -729 8320 -632 8336
rect -729 8252 -682 8320
rect -648 8252 -632 8320
rect -729 8236 -632 8252
rect -590 8320 -493 8336
rect -590 8252 -574 8320
rect -540 8252 -493 8320
rect -590 8236 -493 8252
rect 507 8320 604 8336
rect 507 8252 554 8320
rect 588 8252 604 8320
rect 507 8236 604 8252
rect 646 8320 743 8336
rect 646 8252 662 8320
rect 696 8252 743 8320
rect 646 8236 743 8252
rect 1743 8320 1840 8336
rect 1743 8252 1790 8320
rect 1824 8252 1840 8320
rect 1743 8236 1840 8252
rect 1882 8320 1979 8336
rect 1882 8252 1898 8320
rect 1932 8252 1979 8320
rect 1882 8236 1979 8252
rect 2979 8320 3076 8336
rect 2979 8252 3026 8320
rect 3060 8252 3076 8320
rect 2979 8236 3076 8252
rect 3118 8320 3215 8336
rect 3118 8252 3134 8320
rect 3168 8252 3215 8320
rect 3118 8236 3215 8252
rect 4215 8320 4312 8336
rect 4215 8252 4262 8320
rect 4296 8252 4312 8320
rect 4215 8236 4312 8252
rect -4298 7780 -4201 7796
rect -4298 7712 -4282 7780
rect -4248 7712 -4201 7780
rect -4298 7696 -4201 7712
rect -3201 7780 -3104 7796
rect -3201 7712 -3154 7780
rect -3120 7712 -3104 7780
rect -3201 7696 -3104 7712
rect -3062 7780 -2965 7796
rect -3062 7712 -3046 7780
rect -3012 7712 -2965 7780
rect -3062 7696 -2965 7712
rect -1965 7780 -1868 7796
rect -1965 7712 -1918 7780
rect -1884 7712 -1868 7780
rect -1965 7696 -1868 7712
rect -1826 7780 -1729 7796
rect -1826 7712 -1810 7780
rect -1776 7712 -1729 7780
rect -1826 7696 -1729 7712
rect -729 7780 -632 7796
rect -729 7712 -682 7780
rect -648 7712 -632 7780
rect -729 7696 -632 7712
rect -590 7780 -493 7796
rect -590 7712 -574 7780
rect -540 7712 -493 7780
rect -590 7696 -493 7712
rect 507 7780 604 7796
rect 507 7712 554 7780
rect 588 7712 604 7780
rect 507 7696 604 7712
rect 646 7780 743 7796
rect 646 7712 662 7780
rect 696 7712 743 7780
rect 646 7696 743 7712
rect 1743 7780 1840 7796
rect 1743 7712 1790 7780
rect 1824 7712 1840 7780
rect 1743 7696 1840 7712
rect 1882 7780 1979 7796
rect 1882 7712 1898 7780
rect 1932 7712 1979 7780
rect 1882 7696 1979 7712
rect 2979 7780 3076 7796
rect 2979 7712 3026 7780
rect 3060 7712 3076 7780
rect 2979 7696 3076 7712
rect 3118 7780 3215 7796
rect 3118 7712 3134 7780
rect 3168 7712 3215 7780
rect 3118 7696 3215 7712
rect 4215 7780 4312 7796
rect 4215 7712 4262 7780
rect 4296 7712 4312 7780
rect 4215 7696 4312 7712
rect -4298 7240 -4201 7256
rect -4298 7172 -4282 7240
rect -4248 7172 -4201 7240
rect -4298 7156 -4201 7172
rect -3201 7240 -3104 7256
rect -3201 7172 -3154 7240
rect -3120 7172 -3104 7240
rect -3201 7156 -3104 7172
rect -3062 7240 -2965 7256
rect -3062 7172 -3046 7240
rect -3012 7172 -2965 7240
rect -3062 7156 -2965 7172
rect -1965 7240 -1868 7256
rect -1965 7172 -1918 7240
rect -1884 7172 -1868 7240
rect -1965 7156 -1868 7172
rect -1826 7240 -1729 7256
rect -1826 7172 -1810 7240
rect -1776 7172 -1729 7240
rect -1826 7156 -1729 7172
rect -729 7240 -632 7256
rect -729 7172 -682 7240
rect -648 7172 -632 7240
rect -729 7156 -632 7172
rect -590 7240 -493 7256
rect -590 7172 -574 7240
rect -540 7172 -493 7240
rect -590 7156 -493 7172
rect 507 7240 604 7256
rect 507 7172 554 7240
rect 588 7172 604 7240
rect 507 7156 604 7172
rect 646 7240 743 7256
rect 646 7172 662 7240
rect 696 7172 743 7240
rect 646 7156 743 7172
rect 1743 7240 1840 7256
rect 1743 7172 1790 7240
rect 1824 7172 1840 7240
rect 1743 7156 1840 7172
rect 1882 7240 1979 7256
rect 1882 7172 1898 7240
rect 1932 7172 1979 7240
rect 1882 7156 1979 7172
rect 2979 7240 3076 7256
rect 2979 7172 3026 7240
rect 3060 7172 3076 7240
rect 2979 7156 3076 7172
rect 3118 7240 3215 7256
rect 3118 7172 3134 7240
rect 3168 7172 3215 7240
rect 3118 7156 3215 7172
rect 4215 7240 4312 7256
rect 4215 7172 4262 7240
rect 4296 7172 4312 7240
rect 4215 7156 4312 7172
rect -4298 6660 -4201 6676
rect -4298 6592 -4282 6660
rect -4248 6592 -4201 6660
rect -4298 6576 -4201 6592
rect -3201 6660 -3104 6676
rect -3201 6592 -3154 6660
rect -3120 6592 -3104 6660
rect -3201 6576 -3104 6592
rect -3062 6660 -2965 6676
rect -3062 6592 -3046 6660
rect -3012 6592 -2965 6660
rect -3062 6576 -2965 6592
rect -1965 6660 -1868 6676
rect -1965 6592 -1918 6660
rect -1884 6592 -1868 6660
rect -1965 6576 -1868 6592
rect -1826 6660 -1729 6676
rect -1826 6592 -1810 6660
rect -1776 6592 -1729 6660
rect -1826 6576 -1729 6592
rect -729 6660 -632 6676
rect -729 6592 -682 6660
rect -648 6592 -632 6660
rect -729 6576 -632 6592
rect -590 6660 -493 6676
rect -590 6592 -574 6660
rect -540 6592 -493 6660
rect -590 6576 -493 6592
rect 507 6660 604 6676
rect 507 6592 554 6660
rect 588 6592 604 6660
rect 507 6576 604 6592
rect 646 6660 743 6676
rect 646 6592 662 6660
rect 696 6592 743 6660
rect 646 6576 743 6592
rect 1743 6660 1840 6676
rect 1743 6592 1790 6660
rect 1824 6592 1840 6660
rect 1743 6576 1840 6592
rect 1882 6660 1979 6676
rect 1882 6592 1898 6660
rect 1932 6592 1979 6660
rect 1882 6576 1979 6592
rect 2979 6660 3076 6676
rect 2979 6592 3026 6660
rect 3060 6592 3076 6660
rect 2979 6576 3076 6592
rect 3118 6660 3215 6676
rect 3118 6592 3134 6660
rect 3168 6592 3215 6660
rect 3118 6576 3215 6592
rect 4215 6660 4312 6676
rect 4215 6592 4262 6660
rect 4296 6592 4312 6660
rect 4215 6576 4312 6592
rect -4298 6080 -4201 6096
rect -4298 6012 -4282 6080
rect -4248 6012 -4201 6080
rect -4298 5996 -4201 6012
rect -3201 6080 -3104 6096
rect -3201 6012 -3154 6080
rect -3120 6012 -3104 6080
rect -3201 5996 -3104 6012
rect -3062 6080 -2965 6096
rect -3062 6012 -3046 6080
rect -3012 6012 -2965 6080
rect -3062 5996 -2965 6012
rect -1965 6080 -1868 6096
rect -1965 6012 -1918 6080
rect -1884 6012 -1868 6080
rect -1965 5996 -1868 6012
rect -1826 6080 -1729 6096
rect -1826 6012 -1810 6080
rect -1776 6012 -1729 6080
rect -1826 5996 -1729 6012
rect -729 6080 -632 6096
rect -729 6012 -682 6080
rect -648 6012 -632 6080
rect -729 5996 -632 6012
rect -590 6080 -493 6096
rect -590 6012 -574 6080
rect -540 6012 -493 6080
rect -590 5996 -493 6012
rect 507 6080 604 6096
rect 507 6012 554 6080
rect 588 6012 604 6080
rect 507 5996 604 6012
rect 646 6080 743 6096
rect 646 6012 662 6080
rect 696 6012 743 6080
rect 646 5996 743 6012
rect 1743 6080 1840 6096
rect 1743 6012 1790 6080
rect 1824 6012 1840 6080
rect 1743 5996 1840 6012
rect 1882 6080 1979 6096
rect 1882 6012 1898 6080
rect 1932 6012 1979 6080
rect 1882 5996 1979 6012
rect 2979 6080 3076 6096
rect 2979 6012 3026 6080
rect 3060 6012 3076 6080
rect 2979 5996 3076 6012
rect 3118 6080 3215 6096
rect 3118 6012 3134 6080
rect 3168 6012 3215 6080
rect 3118 5996 3215 6012
rect 4215 6080 4312 6096
rect 4215 6012 4262 6080
rect 4296 6012 4312 6080
rect 4215 5996 4312 6012
rect -6138 5540 -6041 5556
rect -6138 5472 -6122 5540
rect -6088 5472 -6041 5540
rect -6138 5456 -6041 5472
rect -5041 5540 -4944 5556
rect -5041 5472 -4994 5540
rect -4960 5472 -4944 5540
rect -5041 5456 -4944 5472
rect -4902 5540 -4805 5556
rect -4902 5472 -4886 5540
rect -4852 5472 -4805 5540
rect -4902 5456 -4805 5472
rect -3805 5540 -3708 5556
rect -3805 5472 -3758 5540
rect -3724 5472 -3708 5540
rect -3805 5456 -3708 5472
rect -3666 5540 -3569 5556
rect -3666 5472 -3650 5540
rect -3616 5472 -3569 5540
rect -3666 5456 -3569 5472
rect -2569 5540 -2472 5556
rect -2569 5472 -2522 5540
rect -2488 5472 -2472 5540
rect -2569 5456 -2472 5472
rect -2430 5540 -2333 5556
rect -2430 5472 -2414 5540
rect -2380 5472 -2333 5540
rect -2430 5456 -2333 5472
rect -1333 5540 -1236 5556
rect -1333 5472 -1286 5540
rect -1252 5472 -1236 5540
rect -1333 5456 -1236 5472
rect -1194 5540 -1097 5556
rect -1194 5472 -1178 5540
rect -1144 5472 -1097 5540
rect -1194 5456 -1097 5472
rect -97 5540 0 5556
rect -97 5472 -50 5540
rect -16 5472 0 5540
rect -97 5456 0 5472
rect 42 5540 139 5556
rect 42 5472 58 5540
rect 92 5472 139 5540
rect 42 5456 139 5472
rect 1139 5540 1236 5556
rect 1139 5472 1186 5540
rect 1220 5472 1236 5540
rect 1139 5456 1236 5472
rect 1278 5540 1375 5556
rect 1278 5472 1294 5540
rect 1328 5472 1375 5540
rect 1278 5456 1375 5472
rect 2375 5540 2472 5556
rect 2375 5472 2422 5540
rect 2456 5472 2472 5540
rect 2375 5456 2472 5472
rect 2514 5540 2611 5556
rect 2514 5472 2530 5540
rect 2564 5472 2611 5540
rect 2514 5456 2611 5472
rect 3611 5540 3708 5556
rect 3611 5472 3658 5540
rect 3692 5472 3708 5540
rect 3611 5456 3708 5472
rect 3750 5540 3847 5556
rect 3750 5472 3766 5540
rect 3800 5472 3847 5540
rect 3750 5456 3847 5472
rect 4847 5540 4944 5556
rect 4847 5472 4894 5540
rect 4928 5472 4944 5540
rect 4847 5456 4944 5472
rect 4986 5540 5083 5556
rect 4986 5472 5002 5540
rect 5036 5472 5083 5540
rect 4986 5456 5083 5472
rect 6083 5540 6180 5556
rect 6083 5472 6130 5540
rect 6164 5472 6180 5540
rect 6083 5456 6180 5472
rect -6138 5000 -6041 5016
rect -6138 4932 -6122 5000
rect -6088 4932 -6041 5000
rect -6138 4916 -6041 4932
rect -5041 5000 -4944 5016
rect -5041 4932 -4994 5000
rect -4960 4932 -4944 5000
rect -5041 4916 -4944 4932
rect -4902 5000 -4805 5016
rect -4902 4932 -4886 5000
rect -4852 4932 -4805 5000
rect -4902 4916 -4805 4932
rect -3805 5000 -3708 5016
rect -3805 4932 -3758 5000
rect -3724 4932 -3708 5000
rect -3805 4916 -3708 4932
rect -3666 5000 -3569 5016
rect -3666 4932 -3650 5000
rect -3616 4932 -3569 5000
rect -3666 4916 -3569 4932
rect -2569 5000 -2472 5016
rect -2569 4932 -2522 5000
rect -2488 4932 -2472 5000
rect -2569 4916 -2472 4932
rect -2430 5000 -2333 5016
rect -2430 4932 -2414 5000
rect -2380 4932 -2333 5000
rect -2430 4916 -2333 4932
rect -1333 5000 -1236 5016
rect -1333 4932 -1286 5000
rect -1252 4932 -1236 5000
rect -1333 4916 -1236 4932
rect -1194 5000 -1097 5016
rect -1194 4932 -1178 5000
rect -1144 4932 -1097 5000
rect -1194 4916 -1097 4932
rect -97 5000 0 5016
rect -97 4932 -50 5000
rect -16 4932 0 5000
rect -97 4916 0 4932
rect 42 5000 139 5016
rect 42 4932 58 5000
rect 92 4932 139 5000
rect 42 4916 139 4932
rect 1139 5000 1236 5016
rect 1139 4932 1186 5000
rect 1220 4932 1236 5000
rect 1139 4916 1236 4932
rect 1278 5000 1375 5016
rect 1278 4932 1294 5000
rect 1328 4932 1375 5000
rect 1278 4916 1375 4932
rect 2375 5000 2472 5016
rect 2375 4932 2422 5000
rect 2456 4932 2472 5000
rect 2375 4916 2472 4932
rect 2514 5000 2611 5016
rect 2514 4932 2530 5000
rect 2564 4932 2611 5000
rect 2514 4916 2611 4932
rect 3611 5000 3708 5016
rect 3611 4932 3658 5000
rect 3692 4932 3708 5000
rect 3611 4916 3708 4932
rect 3750 5000 3847 5016
rect 3750 4932 3766 5000
rect 3800 4932 3847 5000
rect 3750 4916 3847 4932
rect 4847 5000 4944 5016
rect 4847 4932 4894 5000
rect 4928 4932 4944 5000
rect 4847 4916 4944 4932
rect 4986 5000 5083 5016
rect 4986 4932 5002 5000
rect 5036 4932 5083 5000
rect 4986 4916 5083 4932
rect 6083 5000 6180 5016
rect 6083 4932 6130 5000
rect 6164 4932 6180 5000
rect 6083 4916 6180 4932
rect -6138 4460 -6041 4476
rect -6138 4392 -6122 4460
rect -6088 4392 -6041 4460
rect -6138 4376 -6041 4392
rect -5041 4460 -4944 4476
rect -5041 4392 -4994 4460
rect -4960 4392 -4944 4460
rect -5041 4376 -4944 4392
rect -4902 4460 -4805 4476
rect -4902 4392 -4886 4460
rect -4852 4392 -4805 4460
rect -4902 4376 -4805 4392
rect -3805 4460 -3708 4476
rect -3805 4392 -3758 4460
rect -3724 4392 -3708 4460
rect -3805 4376 -3708 4392
rect -3666 4460 -3569 4476
rect -3666 4392 -3650 4460
rect -3616 4392 -3569 4460
rect -3666 4376 -3569 4392
rect -2569 4460 -2472 4476
rect -2569 4392 -2522 4460
rect -2488 4392 -2472 4460
rect -2569 4376 -2472 4392
rect -2430 4460 -2333 4476
rect -2430 4392 -2414 4460
rect -2380 4392 -2333 4460
rect -2430 4376 -2333 4392
rect -1333 4460 -1236 4476
rect -1333 4392 -1286 4460
rect -1252 4392 -1236 4460
rect -1333 4376 -1236 4392
rect -1194 4460 -1097 4476
rect -1194 4392 -1178 4460
rect -1144 4392 -1097 4460
rect -1194 4376 -1097 4392
rect -97 4460 0 4476
rect -97 4392 -50 4460
rect -16 4392 0 4460
rect -97 4376 0 4392
rect 42 4460 139 4476
rect 42 4392 58 4460
rect 92 4392 139 4460
rect 42 4376 139 4392
rect 1139 4460 1236 4476
rect 1139 4392 1186 4460
rect 1220 4392 1236 4460
rect 1139 4376 1236 4392
rect 1278 4460 1375 4476
rect 1278 4392 1294 4460
rect 1328 4392 1375 4460
rect 1278 4376 1375 4392
rect 2375 4460 2472 4476
rect 2375 4392 2422 4460
rect 2456 4392 2472 4460
rect 2375 4376 2472 4392
rect 2514 4460 2611 4476
rect 2514 4392 2530 4460
rect 2564 4392 2611 4460
rect 2514 4376 2611 4392
rect 3611 4460 3708 4476
rect 3611 4392 3658 4460
rect 3692 4392 3708 4460
rect 3611 4376 3708 4392
rect 3750 4460 3847 4476
rect 3750 4392 3766 4460
rect 3800 4392 3847 4460
rect 3750 4376 3847 4392
rect 4847 4460 4944 4476
rect 4847 4392 4894 4460
rect 4928 4392 4944 4460
rect 4847 4376 4944 4392
rect 4986 4460 5083 4476
rect 4986 4392 5002 4460
rect 5036 4392 5083 4460
rect 4986 4376 5083 4392
rect 6083 4460 6180 4476
rect 6083 4392 6130 4460
rect 6164 4392 6180 4460
rect 6083 4376 6180 4392
rect -6138 3920 -6041 3936
rect -6138 3852 -6122 3920
rect -6088 3852 -6041 3920
rect -6138 3836 -6041 3852
rect -5041 3920 -4944 3936
rect -5041 3852 -4994 3920
rect -4960 3852 -4944 3920
rect -5041 3836 -4944 3852
rect -4902 3920 -4805 3936
rect -4902 3852 -4886 3920
rect -4852 3852 -4805 3920
rect -4902 3836 -4805 3852
rect -3805 3920 -3708 3936
rect -3805 3852 -3758 3920
rect -3724 3852 -3708 3920
rect -3805 3836 -3708 3852
rect -3666 3920 -3569 3936
rect -3666 3852 -3650 3920
rect -3616 3852 -3569 3920
rect -3666 3836 -3569 3852
rect -2569 3920 -2472 3936
rect -2569 3852 -2522 3920
rect -2488 3852 -2472 3920
rect -2569 3836 -2472 3852
rect -2430 3920 -2333 3936
rect -2430 3852 -2414 3920
rect -2380 3852 -2333 3920
rect -2430 3836 -2333 3852
rect -1333 3920 -1236 3936
rect -1333 3852 -1286 3920
rect -1252 3852 -1236 3920
rect -1333 3836 -1236 3852
rect -1194 3920 -1097 3936
rect -1194 3852 -1178 3920
rect -1144 3852 -1097 3920
rect -1194 3836 -1097 3852
rect -97 3920 0 3936
rect -97 3852 -50 3920
rect -16 3852 0 3920
rect -97 3836 0 3852
rect 42 3920 139 3936
rect 42 3852 58 3920
rect 92 3852 139 3920
rect 42 3836 139 3852
rect 1139 3920 1236 3936
rect 1139 3852 1186 3920
rect 1220 3852 1236 3920
rect 1139 3836 1236 3852
rect 1278 3920 1375 3936
rect 1278 3852 1294 3920
rect 1328 3852 1375 3920
rect 1278 3836 1375 3852
rect 2375 3920 2472 3936
rect 2375 3852 2422 3920
rect 2456 3852 2472 3920
rect 2375 3836 2472 3852
rect 2514 3920 2611 3936
rect 2514 3852 2530 3920
rect 2564 3852 2611 3920
rect 2514 3836 2611 3852
rect 3611 3920 3708 3936
rect 3611 3852 3658 3920
rect 3692 3852 3708 3920
rect 3611 3836 3708 3852
rect 3750 3920 3847 3936
rect 3750 3852 3766 3920
rect 3800 3852 3847 3920
rect 3750 3836 3847 3852
rect 4847 3920 4944 3936
rect 4847 3852 4894 3920
rect 4928 3852 4944 3920
rect 4847 3836 4944 3852
rect 4986 3920 5083 3936
rect 4986 3852 5002 3920
rect 5036 3852 5083 3920
rect 4986 3836 5083 3852
rect 6083 3920 6180 3936
rect 6083 3852 6130 3920
rect 6164 3852 6180 3920
rect 6083 3836 6180 3852
rect -4198 3140 -4110 3156
rect -4198 3072 -4182 3140
rect -4148 3072 -4110 3140
rect -4198 3056 -4110 3072
rect -3110 3140 -3022 3156
rect -3110 3072 -3072 3140
rect -3038 3072 -3022 3140
rect -3110 3056 -3022 3072
rect -2980 3140 -2892 3156
rect -2980 3072 -2964 3140
rect -2930 3072 -2892 3140
rect -2980 3056 -2892 3072
rect -1892 3140 -1804 3156
rect -1892 3072 -1854 3140
rect -1820 3072 -1804 3140
rect -1892 3056 -1804 3072
rect -1762 3140 -1674 3156
rect -1762 3072 -1746 3140
rect -1712 3072 -1674 3140
rect -1762 3056 -1674 3072
rect -674 3140 -586 3156
rect -674 3072 -636 3140
rect -602 3072 -586 3140
rect -674 3056 -586 3072
rect -544 3140 -456 3156
rect -544 3072 -528 3140
rect -494 3072 -456 3140
rect -544 3056 -456 3072
rect 544 3140 632 3156
rect 544 3072 582 3140
rect 616 3072 632 3140
rect 544 3056 632 3072
rect 674 3140 762 3156
rect 674 3072 690 3140
rect 724 3072 762 3140
rect 674 3056 762 3072
rect 1762 3140 1850 3156
rect 1762 3072 1800 3140
rect 1834 3072 1850 3140
rect 1762 3056 1850 3072
rect 1892 3140 1980 3156
rect 1892 3072 1908 3140
rect 1942 3072 1980 3140
rect 1892 3056 1980 3072
rect 2980 3140 3068 3156
rect 2980 3072 3018 3140
rect 3052 3072 3068 3140
rect 2980 3056 3068 3072
rect 3110 3140 3198 3156
rect 3110 3072 3126 3140
rect 3160 3072 3198 3140
rect 3110 3056 3198 3072
rect 4198 3140 4286 3156
rect 4198 3072 4236 3140
rect 4270 3072 4286 3140
rect 4198 3056 4286 3072
rect -4198 2640 -4110 2656
rect -4198 2572 -4182 2640
rect -4148 2572 -4110 2640
rect -4198 2556 -4110 2572
rect -3110 2640 -3022 2656
rect -3110 2572 -3072 2640
rect -3038 2572 -3022 2640
rect -3110 2556 -3022 2572
rect -2980 2640 -2892 2656
rect -2980 2572 -2964 2640
rect -2930 2572 -2892 2640
rect -2980 2556 -2892 2572
rect -1892 2640 -1804 2656
rect -1892 2572 -1854 2640
rect -1820 2572 -1804 2640
rect -1892 2556 -1804 2572
rect -1762 2640 -1674 2656
rect -1762 2572 -1746 2640
rect -1712 2572 -1674 2640
rect -1762 2556 -1674 2572
rect -674 2640 -586 2656
rect -674 2572 -636 2640
rect -602 2572 -586 2640
rect -674 2556 -586 2572
rect -544 2640 -456 2656
rect -544 2572 -528 2640
rect -494 2572 -456 2640
rect -544 2556 -456 2572
rect 544 2640 632 2656
rect 544 2572 582 2640
rect 616 2572 632 2640
rect 544 2556 632 2572
rect 674 2640 762 2656
rect 674 2572 690 2640
rect 724 2572 762 2640
rect 674 2556 762 2572
rect 1762 2640 1850 2656
rect 1762 2572 1800 2640
rect 1834 2572 1850 2640
rect 1762 2556 1850 2572
rect 1892 2640 1980 2656
rect 1892 2572 1908 2640
rect 1942 2572 1980 2640
rect 1892 2556 1980 2572
rect 2980 2640 3068 2656
rect 2980 2572 3018 2640
rect 3052 2572 3068 2640
rect 2980 2556 3068 2572
rect 3110 2640 3198 2656
rect 3110 2572 3126 2640
rect 3160 2572 3198 2640
rect 3110 2556 3198 2572
rect 4198 2640 4286 2656
rect 4198 2572 4236 2640
rect 4270 2572 4286 2640
rect 4198 2556 4286 2572
rect -3638 2140 -3550 2156
rect -3638 1972 -3622 2140
rect -3588 1972 -3550 2140
rect -3638 1956 -3550 1972
rect -2550 2140 -2462 2156
rect -2550 1972 -2512 2140
rect -2478 1972 -2462 2140
rect -2550 1956 -2462 1972
rect -2420 2140 -2332 2156
rect -2420 1972 -2404 2140
rect -2370 1972 -2332 2140
rect -2420 1956 -2332 1972
rect -1332 2140 -1244 2156
rect -1332 1972 -1294 2140
rect -1260 1972 -1244 2140
rect -1332 1956 -1244 1972
rect -1202 2140 -1114 2156
rect -1202 1972 -1186 2140
rect -1152 1972 -1114 2140
rect -1202 1956 -1114 1972
rect -114 2140 -26 2156
rect -114 1972 -76 2140
rect -42 1972 -26 2140
rect -114 1956 -26 1972
rect 16 2140 104 2156
rect 16 1972 32 2140
rect 66 1972 104 2140
rect 16 1956 104 1972
rect 1104 2140 1192 2156
rect 1104 1972 1142 2140
rect 1176 1972 1192 2140
rect 1104 1956 1192 1972
rect 1234 2140 1322 2156
rect 1234 1972 1250 2140
rect 1284 1972 1322 2140
rect 1234 1956 1322 1972
rect 2322 2140 2410 2156
rect 2322 1972 2360 2140
rect 2394 1972 2410 2140
rect 2322 1956 2410 1972
rect 2452 2140 2540 2156
rect 2452 1972 2468 2140
rect 2502 1972 2540 2140
rect 2452 1956 2540 1972
rect 3540 2140 3628 2156
rect 3540 1972 3578 2140
rect 3612 1972 3628 2140
rect 3540 1956 3628 1972
rect -3638 1520 -3550 1536
rect -3638 1352 -3622 1520
rect -3588 1352 -3550 1520
rect -3638 1336 -3550 1352
rect -2550 1520 -2462 1536
rect -2550 1352 -2512 1520
rect -2478 1352 -2462 1520
rect -2550 1336 -2462 1352
rect -2420 1520 -2332 1536
rect -2420 1352 -2404 1520
rect -2370 1352 -2332 1520
rect -2420 1336 -2332 1352
rect -1332 1520 -1244 1536
rect -1332 1352 -1294 1520
rect -1260 1352 -1244 1520
rect -1332 1336 -1244 1352
rect -1202 1520 -1114 1536
rect -1202 1352 -1186 1520
rect -1152 1352 -1114 1520
rect -1202 1336 -1114 1352
rect -114 1520 -26 1536
rect -114 1352 -76 1520
rect -42 1352 -26 1520
rect -114 1336 -26 1352
rect 16 1520 104 1536
rect 16 1352 32 1520
rect 66 1352 104 1520
rect 16 1336 104 1352
rect 1104 1520 1192 1536
rect 1104 1352 1142 1520
rect 1176 1352 1192 1520
rect 1104 1336 1192 1352
rect 1234 1520 1322 1536
rect 1234 1352 1250 1520
rect 1284 1352 1322 1520
rect 1234 1336 1322 1352
rect 2322 1520 2410 1536
rect 2322 1352 2360 1520
rect 2394 1352 2410 1520
rect 2322 1336 2410 1352
rect 2452 1520 2540 1536
rect 2452 1352 2468 1520
rect 2502 1352 2540 1520
rect 2452 1336 2540 1352
rect 3540 1520 3628 1536
rect 3540 1352 3578 1520
rect 3612 1352 3628 1520
rect 3540 1336 3628 1352
rect -4198 920 -4110 936
rect -4198 752 -4182 920
rect -4148 752 -4110 920
rect -4198 736 -4110 752
rect -3110 920 -3022 936
rect -3110 752 -3072 920
rect -3038 752 -3022 920
rect -3110 736 -3022 752
rect -2980 920 -2892 936
rect -2980 752 -2964 920
rect -2930 752 -2892 920
rect -2980 736 -2892 752
rect -1892 920 -1804 936
rect -1892 752 -1854 920
rect -1820 752 -1804 920
rect -1892 736 -1804 752
rect -1762 920 -1674 936
rect -1762 752 -1746 920
rect -1712 752 -1674 920
rect -1762 736 -1674 752
rect -674 920 -586 936
rect -674 752 -636 920
rect -602 752 -586 920
rect -674 736 -586 752
rect -544 920 -456 936
rect -544 752 -528 920
rect -494 752 -456 920
rect -544 736 -456 752
rect 544 920 632 936
rect 544 752 582 920
rect 616 752 632 920
rect 544 736 632 752
rect 674 920 762 936
rect 674 752 690 920
rect 724 752 762 920
rect 674 736 762 752
rect 1762 920 1850 936
rect 1762 752 1800 920
rect 1834 752 1850 920
rect 1762 736 1850 752
rect 1892 920 1980 936
rect 1892 752 1908 920
rect 1942 752 1980 920
rect 1892 736 1980 752
rect 2980 920 3068 936
rect 2980 752 3018 920
rect 3052 752 3068 920
rect 2980 736 3068 752
rect 3110 920 3198 936
rect 3110 752 3126 920
rect 3160 752 3198 920
rect 3110 736 3198 752
rect 4198 920 4286 936
rect 4198 752 4236 920
rect 4270 752 4286 920
rect 4198 736 4286 752
rect -4198 320 -4110 336
rect -4198 152 -4182 320
rect -4148 152 -4110 320
rect -4198 136 -4110 152
rect -3110 320 -3022 336
rect -3110 152 -3072 320
rect -3038 152 -3022 320
rect -3110 136 -3022 152
rect -2980 320 -2892 336
rect -2980 152 -2964 320
rect -2930 152 -2892 320
rect -2980 136 -2892 152
rect -1892 320 -1804 336
rect -1892 152 -1854 320
rect -1820 152 -1804 320
rect -1892 136 -1804 152
rect -1762 320 -1674 336
rect -1762 152 -1746 320
rect -1712 152 -1674 320
rect -1762 136 -1674 152
rect -674 320 -586 336
rect -674 152 -636 320
rect -602 152 -586 320
rect -674 136 -586 152
rect -544 320 -456 336
rect -544 152 -528 320
rect -494 152 -456 320
rect -544 136 -456 152
rect 544 320 632 336
rect 544 152 582 320
rect 616 152 632 320
rect 544 136 632 152
rect 674 320 762 336
rect 674 152 690 320
rect 724 152 762 320
rect 674 136 762 152
rect 1762 320 1850 336
rect 1762 152 1800 320
rect 1834 152 1850 320
rect 1762 136 1850 152
rect 1892 320 1980 336
rect 1892 152 1908 320
rect 1942 152 1980 320
rect 1892 136 1980 152
rect 2980 320 3068 336
rect 2980 152 3018 320
rect 3052 152 3068 320
rect 2980 136 3068 152
rect 3110 320 3198 336
rect 3110 152 3126 320
rect 3160 152 3198 320
rect 3110 136 3198 152
rect 4198 320 4286 336
rect 4198 152 4236 320
rect 4270 152 4286 320
rect 4198 136 4286 152
<< polycont >>
rect -4282 8792 -4248 8860
rect -3154 8792 -3120 8860
rect -3046 8792 -3012 8860
rect -1918 8792 -1884 8860
rect -1810 8792 -1776 8860
rect -682 8792 -648 8860
rect -574 8792 -540 8860
rect 554 8792 588 8860
rect 662 8792 696 8860
rect 1790 8792 1824 8860
rect 1898 8792 1932 8860
rect 3026 8792 3060 8860
rect 3134 8792 3168 8860
rect 4262 8792 4296 8860
rect -4282 8252 -4248 8320
rect -3154 8252 -3120 8320
rect -3046 8252 -3012 8320
rect -1918 8252 -1884 8320
rect -1810 8252 -1776 8320
rect -682 8252 -648 8320
rect -574 8252 -540 8320
rect 554 8252 588 8320
rect 662 8252 696 8320
rect 1790 8252 1824 8320
rect 1898 8252 1932 8320
rect 3026 8252 3060 8320
rect 3134 8252 3168 8320
rect 4262 8252 4296 8320
rect -4282 7712 -4248 7780
rect -3154 7712 -3120 7780
rect -3046 7712 -3012 7780
rect -1918 7712 -1884 7780
rect -1810 7712 -1776 7780
rect -682 7712 -648 7780
rect -574 7712 -540 7780
rect 554 7712 588 7780
rect 662 7712 696 7780
rect 1790 7712 1824 7780
rect 1898 7712 1932 7780
rect 3026 7712 3060 7780
rect 3134 7712 3168 7780
rect 4262 7712 4296 7780
rect -4282 7172 -4248 7240
rect -3154 7172 -3120 7240
rect -3046 7172 -3012 7240
rect -1918 7172 -1884 7240
rect -1810 7172 -1776 7240
rect -682 7172 -648 7240
rect -574 7172 -540 7240
rect 554 7172 588 7240
rect 662 7172 696 7240
rect 1790 7172 1824 7240
rect 1898 7172 1932 7240
rect 3026 7172 3060 7240
rect 3134 7172 3168 7240
rect 4262 7172 4296 7240
rect -4282 6592 -4248 6660
rect -3154 6592 -3120 6660
rect -3046 6592 -3012 6660
rect -1918 6592 -1884 6660
rect -1810 6592 -1776 6660
rect -682 6592 -648 6660
rect -574 6592 -540 6660
rect 554 6592 588 6660
rect 662 6592 696 6660
rect 1790 6592 1824 6660
rect 1898 6592 1932 6660
rect 3026 6592 3060 6660
rect 3134 6592 3168 6660
rect 4262 6592 4296 6660
rect -4282 6012 -4248 6080
rect -3154 6012 -3120 6080
rect -3046 6012 -3012 6080
rect -1918 6012 -1884 6080
rect -1810 6012 -1776 6080
rect -682 6012 -648 6080
rect -574 6012 -540 6080
rect 554 6012 588 6080
rect 662 6012 696 6080
rect 1790 6012 1824 6080
rect 1898 6012 1932 6080
rect 3026 6012 3060 6080
rect 3134 6012 3168 6080
rect 4262 6012 4296 6080
rect -6122 5472 -6088 5540
rect -4994 5472 -4960 5540
rect -4886 5472 -4852 5540
rect -3758 5472 -3724 5540
rect -3650 5472 -3616 5540
rect -2522 5472 -2488 5540
rect -2414 5472 -2380 5540
rect -1286 5472 -1252 5540
rect -1178 5472 -1144 5540
rect -50 5472 -16 5540
rect 58 5472 92 5540
rect 1186 5472 1220 5540
rect 1294 5472 1328 5540
rect 2422 5472 2456 5540
rect 2530 5472 2564 5540
rect 3658 5472 3692 5540
rect 3766 5472 3800 5540
rect 4894 5472 4928 5540
rect 5002 5472 5036 5540
rect 6130 5472 6164 5540
rect -6122 4932 -6088 5000
rect -4994 4932 -4960 5000
rect -4886 4932 -4852 5000
rect -3758 4932 -3724 5000
rect -3650 4932 -3616 5000
rect -2522 4932 -2488 5000
rect -2414 4932 -2380 5000
rect -1286 4932 -1252 5000
rect -1178 4932 -1144 5000
rect -50 4932 -16 5000
rect 58 4932 92 5000
rect 1186 4932 1220 5000
rect 1294 4932 1328 5000
rect 2422 4932 2456 5000
rect 2530 4932 2564 5000
rect 3658 4932 3692 5000
rect 3766 4932 3800 5000
rect 4894 4932 4928 5000
rect 5002 4932 5036 5000
rect 6130 4932 6164 5000
rect -6122 4392 -6088 4460
rect -4994 4392 -4960 4460
rect -4886 4392 -4852 4460
rect -3758 4392 -3724 4460
rect -3650 4392 -3616 4460
rect -2522 4392 -2488 4460
rect -2414 4392 -2380 4460
rect -1286 4392 -1252 4460
rect -1178 4392 -1144 4460
rect -50 4392 -16 4460
rect 58 4392 92 4460
rect 1186 4392 1220 4460
rect 1294 4392 1328 4460
rect 2422 4392 2456 4460
rect 2530 4392 2564 4460
rect 3658 4392 3692 4460
rect 3766 4392 3800 4460
rect 4894 4392 4928 4460
rect 5002 4392 5036 4460
rect 6130 4392 6164 4460
rect -6122 3852 -6088 3920
rect -4994 3852 -4960 3920
rect -4886 3852 -4852 3920
rect -3758 3852 -3724 3920
rect -3650 3852 -3616 3920
rect -2522 3852 -2488 3920
rect -2414 3852 -2380 3920
rect -1286 3852 -1252 3920
rect -1178 3852 -1144 3920
rect -50 3852 -16 3920
rect 58 3852 92 3920
rect 1186 3852 1220 3920
rect 1294 3852 1328 3920
rect 2422 3852 2456 3920
rect 2530 3852 2564 3920
rect 3658 3852 3692 3920
rect 3766 3852 3800 3920
rect 4894 3852 4928 3920
rect 5002 3852 5036 3920
rect 6130 3852 6164 3920
rect -4182 3072 -4148 3140
rect -3072 3072 -3038 3140
rect -2964 3072 -2930 3140
rect -1854 3072 -1820 3140
rect -1746 3072 -1712 3140
rect -636 3072 -602 3140
rect -528 3072 -494 3140
rect 582 3072 616 3140
rect 690 3072 724 3140
rect 1800 3072 1834 3140
rect 1908 3072 1942 3140
rect 3018 3072 3052 3140
rect 3126 3072 3160 3140
rect 4236 3072 4270 3140
rect -4182 2572 -4148 2640
rect -3072 2572 -3038 2640
rect -2964 2572 -2930 2640
rect -1854 2572 -1820 2640
rect -1746 2572 -1712 2640
rect -636 2572 -602 2640
rect -528 2572 -494 2640
rect 582 2572 616 2640
rect 690 2572 724 2640
rect 1800 2572 1834 2640
rect 1908 2572 1942 2640
rect 3018 2572 3052 2640
rect 3126 2572 3160 2640
rect 4236 2572 4270 2640
rect -3622 1972 -3588 2140
rect -2512 1972 -2478 2140
rect -2404 1972 -2370 2140
rect -1294 1972 -1260 2140
rect -1186 1972 -1152 2140
rect -76 1972 -42 2140
rect 32 1972 66 2140
rect 1142 1972 1176 2140
rect 1250 1972 1284 2140
rect 2360 1972 2394 2140
rect 2468 1972 2502 2140
rect 3578 1972 3612 2140
rect -3622 1352 -3588 1520
rect -2512 1352 -2478 1520
rect -2404 1352 -2370 1520
rect -1294 1352 -1260 1520
rect -1186 1352 -1152 1520
rect -76 1352 -42 1520
rect 32 1352 66 1520
rect 1142 1352 1176 1520
rect 1250 1352 1284 1520
rect 2360 1352 2394 1520
rect 2468 1352 2502 1520
rect 3578 1352 3612 1520
rect -4182 752 -4148 920
rect -3072 752 -3038 920
rect -2964 752 -2930 920
rect -1854 752 -1820 920
rect -1746 752 -1712 920
rect -636 752 -602 920
rect -528 752 -494 920
rect 582 752 616 920
rect 690 752 724 920
rect 1800 752 1834 920
rect 1908 752 1942 920
rect 3018 752 3052 920
rect 3126 752 3160 920
rect 4236 752 4270 920
rect -4182 152 -4148 320
rect -3072 152 -3038 320
rect -2964 152 -2930 320
rect -1854 152 -1820 320
rect -1746 152 -1712 320
rect -636 152 -602 320
rect -528 152 -494 320
rect 582 152 616 320
rect 690 152 724 320
rect 1800 152 1834 320
rect 1908 152 1942 320
rect 3018 152 3052 320
rect 3126 152 3160 320
rect 4236 152 4270 320
<< xpolycontact >>
rect -9847 4963 -9415 6109
rect -7415 4963 -6983 6109
rect 7213 4963 7645 6109
rect 9645 4963 10077 6109
rect -9847 3493 -9415 4639
rect -7415 3493 -6983 4639
rect 7213 3493 7645 4639
rect 9645 3493 10077 4639
<< xpolyres >>
rect -9415 4963 -7415 6109
rect 7645 4963 9645 6109
rect -9415 3493 -7415 4639
rect 7645 3493 9645 4639
<< locali >>
rect -4384 9002 -4288 9036
rect 4302 9002 4398 9036
rect -4384 8940 -4350 9002
rect 4364 8940 4398 9002
rect -4205 8888 -4189 8922
rect -3213 8888 -3197 8922
rect -2969 8888 -2953 8922
rect -1977 8888 -1961 8922
rect -1733 8888 -1717 8922
rect -741 8888 -725 8922
rect -497 8888 -481 8922
rect 495 8888 511 8922
rect 739 8888 755 8922
rect 1731 8888 1747 8922
rect 1975 8888 1991 8922
rect 2967 8888 2983 8922
rect 3211 8888 3227 8922
rect 4203 8888 4219 8922
rect -4282 8860 -4248 8876
rect -4282 8776 -4248 8792
rect -3154 8860 -3120 8876
rect -3154 8776 -3120 8792
rect -3046 8860 -3012 8876
rect -3046 8776 -3012 8792
rect -1918 8860 -1884 8876
rect -1918 8776 -1884 8792
rect -1810 8860 -1776 8876
rect -1810 8776 -1776 8792
rect -682 8860 -648 8876
rect -682 8776 -648 8792
rect -574 8860 -540 8876
rect -574 8776 -540 8792
rect 554 8860 588 8876
rect 554 8776 588 8792
rect 662 8860 696 8876
rect 662 8776 696 8792
rect 1790 8860 1824 8876
rect 1790 8776 1824 8792
rect 1898 8860 1932 8876
rect 1898 8776 1932 8792
rect 3026 8860 3060 8876
rect 3026 8776 3060 8792
rect 3134 8860 3168 8876
rect 3134 8776 3168 8792
rect 4262 8860 4296 8876
rect 4262 8776 4296 8792
rect -4205 8730 -4189 8764
rect -3213 8730 -3197 8764
rect -2969 8730 -2953 8764
rect -1977 8730 -1961 8764
rect -1733 8730 -1717 8764
rect -741 8730 -725 8764
rect -497 8730 -481 8764
rect 495 8730 511 8764
rect 739 8730 755 8764
rect 1731 8730 1747 8764
rect 1975 8730 1991 8764
rect 2967 8730 2983 8764
rect 3211 8730 3227 8764
rect 4203 8730 4219 8764
rect -4384 8650 -4350 8712
rect 4364 8650 4398 8712
rect -4384 8616 -4288 8650
rect 4302 8616 4398 8650
rect -4384 8462 -4288 8496
rect 4302 8462 4398 8496
rect -4384 8400 -4350 8462
rect 4364 8400 4398 8462
rect -4205 8348 -4189 8382
rect -3213 8348 -3197 8382
rect -2969 8348 -2953 8382
rect -1977 8348 -1961 8382
rect -1733 8348 -1717 8382
rect -741 8348 -725 8382
rect -497 8348 -481 8382
rect 495 8348 511 8382
rect 739 8348 755 8382
rect 1731 8348 1747 8382
rect 1975 8348 1991 8382
rect 2967 8348 2983 8382
rect 3211 8348 3227 8382
rect 4203 8348 4219 8382
rect -4282 8320 -4248 8336
rect -4282 8236 -4248 8252
rect -3154 8320 -3120 8336
rect -3154 8236 -3120 8252
rect -3046 8320 -3012 8336
rect -3046 8236 -3012 8252
rect -1918 8320 -1884 8336
rect -1918 8236 -1884 8252
rect -1810 8320 -1776 8336
rect -1810 8236 -1776 8252
rect -682 8320 -648 8336
rect -682 8236 -648 8252
rect -574 8320 -540 8336
rect -574 8236 -540 8252
rect 554 8320 588 8336
rect 554 8236 588 8252
rect 662 8320 696 8336
rect 662 8236 696 8252
rect 1790 8320 1824 8336
rect 1790 8236 1824 8252
rect 1898 8320 1932 8336
rect 1898 8236 1932 8252
rect 3026 8320 3060 8336
rect 3026 8236 3060 8252
rect 3134 8320 3168 8336
rect 3134 8236 3168 8252
rect 4262 8320 4296 8336
rect 4262 8236 4296 8252
rect -4205 8190 -4189 8224
rect -3213 8190 -3197 8224
rect -2969 8190 -2953 8224
rect -1977 8190 -1961 8224
rect -1733 8190 -1717 8224
rect -741 8190 -725 8224
rect -497 8190 -481 8224
rect 495 8190 511 8224
rect 739 8190 755 8224
rect 1731 8190 1747 8224
rect 1975 8190 1991 8224
rect 2967 8190 2983 8224
rect 3211 8190 3227 8224
rect 4203 8190 4219 8224
rect -4384 8110 -4350 8172
rect 4364 8110 4398 8172
rect -4384 8076 -4288 8110
rect 4302 8076 4398 8110
rect -2600 8050 -2340 8076
rect -2600 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -2340 8050
rect -2600 7956 -2340 7980
rect -130 8060 160 8076
rect -130 8050 50 8060
rect -130 7980 -110 8050
rect -20 7990 50 8050
rect 140 7990 160 8060
rect -20 7980 160 7990
rect -130 7956 160 7980
rect 2330 8060 2620 8076
rect 2330 7990 2350 8060
rect 2430 7990 2520 8060
rect 2600 7990 2620 8060
rect 2330 7956 2620 7990
rect -4384 7922 -4288 7956
rect 4302 7922 4398 7956
rect -4384 7860 -4350 7922
rect 4364 7860 4398 7922
rect -4205 7808 -4189 7842
rect -3213 7808 -3197 7842
rect -2969 7808 -2953 7842
rect -1977 7808 -1961 7842
rect -1733 7808 -1717 7842
rect -741 7808 -725 7842
rect -497 7808 -481 7842
rect 495 7808 511 7842
rect 739 7808 755 7842
rect 1731 7808 1747 7842
rect 1975 7808 1991 7842
rect 2967 7808 2983 7842
rect 3211 7808 3227 7842
rect 4203 7808 4219 7842
rect -4282 7780 -4248 7796
rect -4282 7696 -4248 7712
rect -3154 7780 -3120 7796
rect -3154 7696 -3120 7712
rect -3046 7780 -3012 7796
rect -3046 7696 -3012 7712
rect -1918 7780 -1884 7796
rect -1918 7696 -1884 7712
rect -1810 7780 -1776 7796
rect -1810 7696 -1776 7712
rect -682 7780 -648 7796
rect -682 7696 -648 7712
rect -574 7780 -540 7796
rect -574 7696 -540 7712
rect 554 7780 588 7796
rect 554 7696 588 7712
rect 662 7780 696 7796
rect 662 7696 696 7712
rect 1790 7780 1824 7796
rect 1790 7696 1824 7712
rect 1898 7780 1932 7796
rect 1898 7696 1932 7712
rect 3026 7780 3060 7796
rect 3026 7696 3060 7712
rect 3134 7780 3168 7796
rect 3134 7696 3168 7712
rect 4262 7780 4296 7796
rect 4262 7696 4296 7712
rect -4205 7650 -4189 7684
rect -3213 7650 -3197 7684
rect -2969 7650 -2953 7684
rect -1977 7650 -1961 7684
rect -1733 7650 -1717 7684
rect -741 7650 -725 7684
rect -497 7650 -481 7684
rect 495 7650 511 7684
rect 739 7650 755 7684
rect 1731 7650 1747 7684
rect 1975 7650 1991 7684
rect 2967 7650 2983 7684
rect 3211 7650 3227 7684
rect 4203 7650 4219 7684
rect -4384 7570 -4350 7632
rect 4364 7570 4398 7632
rect -4384 7536 -4288 7570
rect 4302 7536 4398 7570
rect -2610 7520 -2320 7536
rect -2610 7440 -2590 7520
rect -2510 7440 -2420 7520
rect -2340 7440 -2320 7520
rect -2610 7416 -2320 7440
rect -130 7520 160 7536
rect -130 7440 -110 7520
rect -30 7440 60 7520
rect 140 7440 160 7520
rect -130 7416 160 7440
rect 2330 7520 2620 7536
rect 2330 7440 2350 7520
rect 2430 7440 2520 7520
rect 2600 7440 2620 7520
rect 2330 7416 2620 7440
rect -4384 7382 -4288 7416
rect 4302 7382 4398 7416
rect -4384 7320 -4350 7382
rect 4364 7320 4398 7382
rect -4205 7268 -4189 7302
rect -3213 7268 -3197 7302
rect -2969 7268 -2953 7302
rect -1977 7268 -1961 7302
rect -1733 7268 -1717 7302
rect -741 7268 -725 7302
rect -497 7268 -481 7302
rect 495 7268 511 7302
rect 739 7268 755 7302
rect 1731 7268 1747 7302
rect 1975 7268 1991 7302
rect 2967 7268 2983 7302
rect 3211 7268 3227 7302
rect 4203 7268 4219 7302
rect -4282 7240 -4248 7256
rect -4282 7156 -4248 7172
rect -3154 7240 -3120 7256
rect -3154 7156 -3120 7172
rect -3046 7240 -3012 7256
rect -3046 7156 -3012 7172
rect -1918 7240 -1884 7256
rect -1918 7156 -1884 7172
rect -1810 7240 -1776 7256
rect -1810 7156 -1776 7172
rect -682 7240 -648 7256
rect -682 7156 -648 7172
rect -574 7240 -540 7256
rect -574 7156 -540 7172
rect 554 7240 588 7256
rect 554 7156 588 7172
rect 662 7240 696 7256
rect 662 7156 696 7172
rect 1790 7240 1824 7256
rect 1790 7156 1824 7172
rect 1898 7240 1932 7256
rect 1898 7156 1932 7172
rect 3026 7240 3060 7256
rect 3026 7156 3060 7172
rect 3134 7240 3168 7256
rect 3134 7156 3168 7172
rect 4262 7240 4296 7256
rect 4262 7156 4296 7172
rect -4205 7110 -4189 7144
rect -3213 7110 -3197 7144
rect -2969 7110 -2953 7144
rect -1977 7110 -1961 7144
rect -1733 7110 -1717 7144
rect -741 7110 -725 7144
rect -497 7110 -481 7144
rect 495 7110 511 7144
rect 739 7110 755 7144
rect 1731 7110 1747 7144
rect 1975 7110 1991 7144
rect 2967 7110 2983 7144
rect 3211 7110 3227 7144
rect 4203 7110 4219 7144
rect -4384 7030 -4350 7092
rect 4364 7030 4398 7092
rect -4384 6996 -4288 7030
rect 4302 6996 4398 7030
rect -4384 6802 -4288 6836
rect 4302 6802 4398 6836
rect -4384 6740 -4350 6802
rect 4364 6740 4398 6802
rect -4205 6688 -4189 6722
rect -3213 6688 -3197 6722
rect -2969 6688 -2953 6722
rect -1977 6688 -1961 6722
rect -1733 6688 -1717 6722
rect -741 6688 -725 6722
rect -497 6688 -481 6722
rect 495 6688 511 6722
rect 739 6688 755 6722
rect 1731 6688 1747 6722
rect 1975 6688 1991 6722
rect 2967 6688 2983 6722
rect 3211 6688 3227 6722
rect 4203 6688 4219 6722
rect -4282 6660 -4248 6676
rect -4282 6576 -4248 6592
rect -3154 6660 -3120 6676
rect -3154 6576 -3120 6592
rect -3046 6660 -3012 6676
rect -3046 6576 -3012 6592
rect -1918 6660 -1884 6676
rect -1918 6576 -1884 6592
rect -1810 6660 -1776 6676
rect -1810 6576 -1776 6592
rect -682 6660 -648 6676
rect -682 6576 -648 6592
rect -574 6660 -540 6676
rect -574 6576 -540 6592
rect 554 6660 588 6676
rect 554 6576 588 6592
rect 662 6660 696 6676
rect 662 6576 696 6592
rect 1790 6660 1824 6676
rect 1790 6576 1824 6592
rect 1898 6660 1932 6676
rect 1898 6576 1932 6592
rect 3026 6660 3060 6676
rect 3026 6576 3060 6592
rect 3134 6660 3168 6676
rect 3134 6576 3168 6592
rect 4262 6660 4296 6676
rect 4262 6576 4296 6592
rect -4205 6530 -4189 6564
rect -3213 6530 -3197 6564
rect -2969 6530 -2953 6564
rect -1977 6530 -1961 6564
rect -1733 6530 -1717 6564
rect -741 6530 -725 6564
rect -497 6530 -481 6564
rect 495 6530 511 6564
rect 739 6530 755 6564
rect 1731 6530 1747 6564
rect 1975 6530 1991 6564
rect 2967 6530 2983 6564
rect 3211 6530 3227 6564
rect 4203 6530 4219 6564
rect -4384 6450 -4350 6512
rect 4364 6450 4398 6512
rect -4384 6416 -4288 6450
rect 4302 6416 4398 6450
rect -2610 6360 -2320 6416
rect -2610 6280 -2590 6360
rect -2500 6280 -2430 6360
rect -2340 6280 -2320 6360
rect -2610 6256 -2320 6280
rect -130 6350 160 6416
rect -130 6280 -110 6350
rect -30 6280 60 6350
rect 140 6280 160 6350
rect -130 6256 160 6280
rect 2330 6350 2620 6416
rect 2330 6280 2350 6350
rect 2430 6280 2520 6350
rect 2600 6280 2620 6350
rect 2330 6256 2620 6280
rect -9977 6205 -9881 6239
rect -6949 6205 -6853 6239
rect -9977 6143 -9943 6205
rect -6887 6143 -6853 6205
rect -9977 4867 -9943 4929
rect -4384 6222 -4288 6256
rect 4302 6222 4398 6256
rect -4384 6160 -4350 6222
rect 4364 6160 4398 6222
rect -4205 6108 -4189 6142
rect -3213 6108 -3197 6142
rect -2969 6108 -2953 6142
rect -1977 6108 -1961 6142
rect -1733 6108 -1717 6142
rect -741 6108 -725 6142
rect -497 6108 -481 6142
rect 495 6108 511 6142
rect 739 6108 755 6142
rect 1731 6108 1747 6142
rect 1975 6108 1991 6142
rect 2967 6108 2983 6142
rect 3211 6108 3227 6142
rect 4203 6108 4219 6142
rect -4282 6080 -4248 6096
rect -4282 5996 -4248 6012
rect -3154 6080 -3120 6096
rect -3154 5996 -3120 6012
rect -3046 6080 -3012 6096
rect -3046 5996 -3012 6012
rect -1918 6080 -1884 6096
rect -1918 5996 -1884 6012
rect -1810 6080 -1776 6096
rect -1810 5996 -1776 6012
rect -682 6080 -648 6096
rect -682 5996 -648 6012
rect -574 6080 -540 6096
rect -574 5996 -540 6012
rect 554 6080 588 6096
rect 554 5996 588 6012
rect 662 6080 696 6096
rect 662 5996 696 6012
rect 1790 6080 1824 6096
rect 1790 5996 1824 6012
rect 1898 6080 1932 6096
rect 1898 5996 1932 6012
rect 3026 6080 3060 6096
rect 3026 5996 3060 6012
rect 3134 6080 3168 6096
rect 3134 5996 3168 6012
rect 4262 6080 4296 6096
rect 4262 5996 4296 6012
rect -4205 5950 -4189 5984
rect -3213 5950 -3197 5984
rect -2969 5950 -2953 5984
rect -1977 5950 -1961 5984
rect -1733 5950 -1717 5984
rect -741 5950 -725 5984
rect -497 5950 -481 5984
rect 495 5950 511 5984
rect 739 5950 755 5984
rect 1731 5950 1747 5984
rect 1975 5950 1991 5984
rect 2967 5950 2983 5984
rect 3211 5950 3227 5984
rect 4203 5950 4219 5984
rect -4384 5870 -4350 5932
rect 4364 5870 4398 5932
rect -4384 5836 -4288 5870
rect 4302 5836 4398 5870
rect 7083 6205 7179 6239
rect 10111 6205 10207 6239
rect 7083 6143 7117 6205
rect -6224 5682 -6128 5716
rect 6170 5682 6266 5716
rect -6224 5620 -6190 5682
rect 6232 5620 6266 5682
rect -6045 5568 -6029 5602
rect -5053 5568 -5037 5602
rect -4809 5568 -4793 5602
rect -3817 5568 -3801 5602
rect -3573 5568 -3557 5602
rect -2581 5568 -2565 5602
rect -2337 5568 -2321 5602
rect -1345 5568 -1329 5602
rect -1101 5568 -1085 5602
rect -109 5568 -93 5602
rect 135 5568 151 5602
rect 1127 5568 1143 5602
rect 1371 5568 1387 5602
rect 2363 5568 2379 5602
rect 2607 5568 2623 5602
rect 3599 5568 3615 5602
rect 3843 5568 3859 5602
rect 4835 5568 4851 5602
rect 5079 5568 5095 5602
rect 6071 5568 6087 5602
rect -6122 5540 -6088 5556
rect -6122 5456 -6088 5472
rect -4994 5540 -4960 5556
rect -4994 5456 -4960 5472
rect -4886 5540 -4852 5556
rect -4886 5456 -4852 5472
rect -3758 5540 -3724 5556
rect -3758 5456 -3724 5472
rect -3650 5540 -3616 5556
rect -3650 5456 -3616 5472
rect -2522 5540 -2488 5556
rect -2522 5456 -2488 5472
rect -2414 5540 -2380 5556
rect -2414 5456 -2380 5472
rect -1286 5540 -1252 5556
rect -1286 5456 -1252 5472
rect -1178 5540 -1144 5556
rect -1178 5456 -1144 5472
rect -50 5540 -16 5556
rect -50 5456 -16 5472
rect 58 5540 92 5556
rect 58 5456 92 5472
rect 1186 5540 1220 5556
rect 1186 5456 1220 5472
rect 1294 5540 1328 5556
rect 1294 5456 1328 5472
rect 2422 5540 2456 5556
rect 2422 5456 2456 5472
rect 2530 5540 2564 5556
rect 2530 5456 2564 5472
rect 3658 5540 3692 5556
rect 3658 5456 3692 5472
rect 3766 5540 3800 5556
rect 3766 5456 3800 5472
rect 4894 5540 4928 5556
rect 4894 5456 4928 5472
rect 5002 5540 5036 5556
rect 5002 5456 5036 5472
rect 6130 5540 6164 5556
rect 6130 5456 6164 5472
rect -6045 5410 -6029 5444
rect -5053 5410 -5037 5444
rect -4809 5410 -4793 5444
rect -3817 5410 -3801 5444
rect -3573 5410 -3557 5444
rect -2581 5410 -2565 5444
rect -2337 5410 -2321 5444
rect -1345 5410 -1329 5444
rect -1101 5410 -1085 5444
rect -109 5410 -93 5444
rect 135 5410 151 5444
rect 1127 5410 1143 5444
rect 1371 5410 1387 5444
rect 2363 5410 2379 5444
rect 2607 5410 2623 5444
rect 3599 5410 3615 5444
rect 3843 5410 3859 5444
rect 4835 5410 4851 5444
rect 5079 5410 5095 5444
rect 6071 5410 6087 5444
rect -6224 5330 -6190 5392
rect 6232 5330 6266 5392
rect -6224 5296 -6128 5330
rect 6170 5296 6266 5330
rect -4470 5280 -4160 5296
rect -4470 5200 -4450 5280
rect -4360 5200 -4270 5280
rect -4180 5200 -4160 5280
rect -4470 5176 -4160 5200
rect -1940 5280 -1650 5296
rect -1940 5200 -1920 5280
rect -1830 5200 -1760 5280
rect -1670 5200 -1650 5280
rect -1940 5176 -1650 5200
rect 530 5280 820 5296
rect 530 5200 550 5280
rect 640 5200 710 5280
rect 800 5200 820 5280
rect 530 5176 820 5200
rect 2980 5280 3270 5296
rect 2980 5200 3000 5280
rect 3090 5200 3160 5280
rect 3250 5200 3270 5280
rect 2980 5176 3270 5200
rect 5480 5280 5770 5296
rect 5480 5200 5500 5280
rect 5590 5200 5660 5280
rect 5750 5200 5770 5280
rect 5480 5176 5770 5200
rect -8790 4867 -8700 4880
rect -6887 4867 -6853 4929
rect -9977 4833 -9881 4867
rect -6949 4833 -6853 4867
rect -6224 5142 -6128 5176
rect 6170 5142 6266 5176
rect -6224 5080 -6190 5142
rect 6232 5080 6266 5142
rect -6045 5028 -6029 5062
rect -5053 5028 -5037 5062
rect -4809 5028 -4793 5062
rect -3817 5028 -3801 5062
rect -3573 5028 -3557 5062
rect -2581 5028 -2565 5062
rect -2337 5028 -2321 5062
rect -1345 5028 -1329 5062
rect -1101 5028 -1085 5062
rect -109 5028 -93 5062
rect 135 5028 151 5062
rect 1127 5028 1143 5062
rect 1371 5028 1387 5062
rect 2363 5028 2379 5062
rect 2607 5028 2623 5062
rect 3599 5028 3615 5062
rect 3843 5028 3859 5062
rect 4835 5028 4851 5062
rect 5079 5028 5095 5062
rect 6071 5028 6087 5062
rect -6122 5000 -6088 5016
rect -6122 4916 -6088 4932
rect -4994 5000 -4960 5016
rect -4994 4916 -4960 4932
rect -4886 5000 -4852 5016
rect -4886 4916 -4852 4932
rect -3758 5000 -3724 5016
rect -3758 4916 -3724 4932
rect -3650 5000 -3616 5016
rect -3650 4916 -3616 4932
rect -2522 5000 -2488 5016
rect -2522 4916 -2488 4932
rect -2414 5000 -2380 5016
rect -2414 4916 -2380 4932
rect -1286 5000 -1252 5016
rect -1286 4916 -1252 4932
rect -1178 5000 -1144 5016
rect -1178 4916 -1144 4932
rect -50 5000 -16 5016
rect -50 4916 -16 4932
rect 58 5000 92 5016
rect 58 4916 92 4932
rect 1186 5000 1220 5016
rect 1186 4916 1220 4932
rect 1294 5000 1328 5016
rect 1294 4916 1328 4932
rect 2422 5000 2456 5016
rect 2422 4916 2456 4932
rect 2530 5000 2564 5016
rect 2530 4916 2564 4932
rect 3658 5000 3692 5016
rect 3658 4916 3692 4932
rect 3766 5000 3800 5016
rect 3766 4916 3800 4932
rect 4894 5000 4928 5016
rect 4894 4916 4928 4932
rect 5002 5000 5036 5016
rect 5002 4916 5036 4932
rect 6130 5000 6164 5016
rect 6130 4916 6164 4932
rect -6045 4870 -6029 4904
rect -5053 4870 -5037 4904
rect -4809 4870 -4793 4904
rect -3817 4870 -3801 4904
rect -3573 4870 -3557 4904
rect -2581 4870 -2565 4904
rect -2337 4870 -2321 4904
rect -1345 4870 -1329 4904
rect -1101 4870 -1085 4904
rect -109 4870 -93 4904
rect 135 4870 151 4904
rect 1127 4870 1143 4904
rect 1371 4870 1387 4904
rect 2363 4870 2379 4904
rect 2607 4870 2623 4904
rect 3599 4870 3615 4904
rect 3843 4870 3859 4904
rect 4835 4870 4851 4904
rect 5079 4870 5095 4904
rect 6071 4870 6087 4904
rect -8790 4769 -8700 4833
rect -6224 4790 -6190 4852
rect 6232 4790 6266 4852
rect 10173 6143 10207 6205
rect 7083 4867 7117 4929
rect 10173 4867 10207 4929
rect 7083 4833 7179 4867
rect 10111 4833 10207 4867
rect -9977 4735 -9881 4769
rect -6949 4735 -6853 4769
rect -6224 4756 -6128 4790
rect 6170 4756 6266 4790
rect 8460 4769 8600 4833
rect -9977 4673 -9943 4735
rect -6887 4673 -6853 4735
rect -9977 3397 -9943 3459
rect 7083 4735 7179 4769
rect 10111 4735 10207 4769
rect 7083 4673 7117 4735
rect -6224 4602 -6128 4636
rect 6170 4602 6266 4636
rect -6224 4540 -6190 4602
rect 6232 4540 6266 4602
rect -6045 4488 -6029 4522
rect -5053 4488 -5037 4522
rect -4809 4488 -4793 4522
rect -3817 4488 -3801 4522
rect -3573 4488 -3557 4522
rect -2581 4488 -2565 4522
rect -2337 4488 -2321 4522
rect -1345 4488 -1329 4522
rect -1101 4488 -1085 4522
rect -109 4488 -93 4522
rect 135 4488 151 4522
rect 1127 4488 1143 4522
rect 1371 4488 1387 4522
rect 2363 4488 2379 4522
rect 2607 4488 2623 4522
rect 3599 4488 3615 4522
rect 3843 4488 3859 4522
rect 4835 4488 4851 4522
rect 5079 4488 5095 4522
rect 6071 4488 6087 4522
rect -6122 4460 -6088 4476
rect -6122 4376 -6088 4392
rect -4994 4460 -4960 4476
rect -4994 4376 -4960 4392
rect -4886 4460 -4852 4476
rect -4886 4376 -4852 4392
rect -3758 4460 -3724 4476
rect -3758 4376 -3724 4392
rect -3650 4460 -3616 4476
rect -3650 4376 -3616 4392
rect -2522 4460 -2488 4476
rect -2522 4376 -2488 4392
rect -2414 4460 -2380 4476
rect -2414 4376 -2380 4392
rect -1286 4460 -1252 4476
rect -1286 4376 -1252 4392
rect -1178 4460 -1144 4476
rect -1178 4376 -1144 4392
rect -50 4460 -16 4476
rect -50 4376 -16 4392
rect 58 4460 92 4476
rect 58 4376 92 4392
rect 1186 4460 1220 4476
rect 1186 4376 1220 4392
rect 1294 4460 1328 4476
rect 1294 4376 1328 4392
rect 2422 4460 2456 4476
rect 2422 4376 2456 4392
rect 2530 4460 2564 4476
rect 2530 4376 2564 4392
rect 3658 4460 3692 4476
rect 3658 4376 3692 4392
rect 3766 4460 3800 4476
rect 3766 4376 3800 4392
rect 4894 4460 4928 4476
rect 4894 4376 4928 4392
rect 5002 4460 5036 4476
rect 5002 4376 5036 4392
rect 6130 4460 6164 4476
rect 6130 4376 6164 4392
rect -6045 4330 -6029 4364
rect -5053 4330 -5037 4364
rect -4809 4330 -4793 4364
rect -3817 4330 -3801 4364
rect -3573 4330 -3557 4364
rect -2581 4330 -2565 4364
rect -2337 4330 -2321 4364
rect -1345 4330 -1329 4364
rect -1101 4330 -1085 4364
rect -109 4330 -93 4364
rect 135 4330 151 4364
rect 1127 4330 1143 4364
rect 1371 4330 1387 4364
rect 2363 4330 2379 4364
rect 2607 4330 2623 4364
rect 3599 4330 3615 4364
rect 3843 4330 3859 4364
rect 4835 4330 4851 4364
rect 5079 4330 5095 4364
rect 6071 4330 6087 4364
rect -6224 4250 -6190 4312
rect 6232 4250 6266 4312
rect -6224 4216 -6128 4250
rect 6170 4216 6266 4250
rect -4470 4210 -4160 4216
rect -4470 4200 -4270 4210
rect -4470 4120 -4450 4200
rect -4360 4130 -4270 4200
rect -4180 4130 -4160 4210
rect -4360 4120 -4160 4130
rect -4470 4096 -4160 4120
rect -1940 4200 -1650 4216
rect -1940 4120 -1920 4200
rect -1830 4120 -1760 4200
rect -1670 4120 -1650 4200
rect -1940 4096 -1650 4120
rect 530 4200 820 4216
rect 530 4120 550 4200
rect 640 4120 710 4200
rect 800 4120 820 4200
rect 530 4096 820 4120
rect 2980 4200 3270 4216
rect 2980 4120 3000 4200
rect 3090 4120 3160 4200
rect 3250 4120 3270 4200
rect 2980 4096 3270 4120
rect 5480 4200 5770 4216
rect 5480 4120 5500 4200
rect 5590 4120 5660 4200
rect 5750 4120 5770 4200
rect 5480 4096 5770 4120
rect -6224 4062 -6128 4096
rect 6170 4062 6266 4096
rect -6224 4000 -6190 4062
rect 6232 4000 6266 4062
rect -6045 3948 -6029 3982
rect -5053 3948 -5037 3982
rect -4809 3948 -4793 3982
rect -3817 3948 -3801 3982
rect -3573 3948 -3557 3982
rect -2581 3948 -2565 3982
rect -2337 3948 -2321 3982
rect -1345 3948 -1329 3982
rect -1101 3948 -1085 3982
rect -109 3948 -93 3982
rect 135 3948 151 3982
rect 1127 3948 1143 3982
rect 1371 3948 1387 3982
rect 2363 3948 2379 3982
rect 2607 3948 2623 3982
rect 3599 3948 3615 3982
rect 3843 3948 3859 3982
rect 4835 3948 4851 3982
rect 5079 3948 5095 3982
rect 6071 3948 6087 3982
rect -6122 3920 -6088 3936
rect -6122 3836 -6088 3852
rect -4994 3920 -4960 3936
rect -4994 3836 -4960 3852
rect -4886 3920 -4852 3936
rect -4886 3836 -4852 3852
rect -3758 3920 -3724 3936
rect -3758 3836 -3724 3852
rect -3650 3920 -3616 3936
rect -3650 3836 -3616 3852
rect -2522 3920 -2488 3936
rect -2522 3836 -2488 3852
rect -2414 3920 -2380 3936
rect -2414 3836 -2380 3852
rect -1286 3920 -1252 3936
rect -1286 3836 -1252 3852
rect -1178 3920 -1144 3936
rect -1178 3836 -1144 3852
rect -50 3920 -16 3936
rect -50 3836 -16 3852
rect 58 3920 92 3936
rect 58 3836 92 3852
rect 1186 3920 1220 3936
rect 1186 3836 1220 3852
rect 1294 3920 1328 3936
rect 1294 3836 1328 3852
rect 2422 3920 2456 3936
rect 2422 3836 2456 3852
rect 2530 3920 2564 3936
rect 2530 3836 2564 3852
rect 3658 3920 3692 3936
rect 3658 3836 3692 3852
rect 3766 3920 3800 3936
rect 3766 3836 3800 3852
rect 4894 3920 4928 3936
rect 4894 3836 4928 3852
rect 5002 3920 5036 3936
rect 5002 3836 5036 3852
rect 6130 3920 6164 3936
rect 6130 3836 6164 3852
rect -6045 3790 -6029 3824
rect -5053 3790 -5037 3824
rect -4809 3790 -4793 3824
rect -3817 3790 -3801 3824
rect -3573 3790 -3557 3824
rect -2581 3790 -2565 3824
rect -2337 3790 -2321 3824
rect -1345 3790 -1329 3824
rect -1101 3790 -1085 3824
rect -109 3790 -93 3824
rect 135 3790 151 3824
rect 1127 3790 1143 3824
rect 1371 3790 1387 3824
rect 2363 3790 2379 3824
rect 2607 3790 2623 3824
rect 3599 3790 3615 3824
rect 3843 3790 3859 3824
rect 4835 3790 4851 3824
rect 5079 3790 5095 3824
rect 6071 3790 6087 3824
rect -6224 3710 -6190 3772
rect 6232 3710 6266 3772
rect -6224 3676 -6128 3710
rect 6170 3676 6266 3710
rect -6887 3397 -6853 3459
rect -9977 3363 -9881 3397
rect -6949 3363 -6853 3397
rect 10173 4673 10207 4735
rect 7083 3397 7117 3459
rect 10173 3397 10207 3459
rect 7083 3363 7179 3397
rect 10111 3363 10207 3397
rect -4284 3282 -4188 3316
rect 4276 3282 4372 3316
rect -4284 3220 -4250 3282
rect 4338 3220 4372 3282
rect -4114 3168 -4098 3202
rect -3122 3168 -3106 3202
rect -2896 3168 -2880 3202
rect -1904 3168 -1888 3202
rect -1678 3168 -1662 3202
rect -686 3168 -670 3202
rect -460 3168 -444 3202
rect 532 3168 548 3202
rect 758 3168 774 3202
rect 1750 3168 1766 3202
rect 1976 3168 1992 3202
rect 2968 3168 2984 3202
rect 3194 3168 3210 3202
rect 4186 3168 4202 3202
rect -4182 3140 -4148 3156
rect -4182 3056 -4148 3072
rect -3072 3140 -3038 3156
rect -3072 3056 -3038 3072
rect -2964 3140 -2930 3156
rect -2964 3056 -2930 3072
rect -1854 3140 -1820 3156
rect -1854 3056 -1820 3072
rect -1746 3140 -1712 3156
rect -1746 3056 -1712 3072
rect -636 3140 -602 3156
rect -636 3056 -602 3072
rect -528 3140 -494 3156
rect -528 3056 -494 3072
rect 582 3140 616 3156
rect 582 3056 616 3072
rect 690 3140 724 3156
rect 690 3056 724 3072
rect 1800 3140 1834 3156
rect 1800 3056 1834 3072
rect 1908 3140 1942 3156
rect 1908 3056 1942 3072
rect 3018 3140 3052 3156
rect 3018 3056 3052 3072
rect 3126 3140 3160 3156
rect 3126 3056 3160 3072
rect 4236 3140 4270 3156
rect 4236 3056 4270 3072
rect -4114 3010 -4098 3044
rect -3122 3010 -3106 3044
rect -2896 3010 -2880 3044
rect -1904 3010 -1888 3044
rect -1678 3010 -1662 3044
rect -686 3010 -670 3044
rect -460 3010 -444 3044
rect 532 3010 548 3044
rect 758 3010 774 3044
rect 1750 3010 1766 3044
rect 1976 3010 1992 3044
rect 2968 3010 2984 3044
rect 3194 3010 3210 3044
rect 4186 3010 4202 3044
rect -4284 2930 -4250 2992
rect 4338 2930 4372 2992
rect -4284 2896 -4188 2930
rect 4276 2896 4372 2930
rect -4284 2782 -4188 2816
rect 4276 2782 4372 2816
rect -4284 2720 -4250 2782
rect 4338 2720 4372 2782
rect -4114 2668 -4098 2702
rect -3122 2668 -3106 2702
rect -2896 2668 -2880 2702
rect -1904 2668 -1888 2702
rect -1678 2668 -1662 2702
rect -686 2668 -670 2702
rect -460 2668 -444 2702
rect 532 2668 548 2702
rect 758 2668 774 2702
rect 1750 2668 1766 2702
rect 1976 2668 1992 2702
rect 2968 2668 2984 2702
rect 3194 2668 3210 2702
rect 4186 2668 4202 2702
rect -4182 2640 -4148 2656
rect -4182 2556 -4148 2572
rect -3072 2640 -3038 2656
rect -3072 2556 -3038 2572
rect -2964 2640 -2930 2656
rect -2964 2556 -2930 2572
rect -1854 2640 -1820 2656
rect -1854 2556 -1820 2572
rect -1746 2640 -1712 2656
rect -1746 2556 -1712 2572
rect -636 2640 -602 2656
rect -636 2556 -602 2572
rect -528 2640 -494 2656
rect -528 2556 -494 2572
rect 582 2640 616 2656
rect 582 2556 616 2572
rect 690 2640 724 2656
rect 690 2556 724 2572
rect 1800 2640 1834 2656
rect 1800 2556 1834 2572
rect 1908 2640 1942 2656
rect 1908 2556 1942 2572
rect 3018 2640 3052 2656
rect 3018 2556 3052 2572
rect 3126 2640 3160 2656
rect 3126 2556 3160 2572
rect 4236 2640 4270 2656
rect 4236 2556 4270 2572
rect -4114 2510 -4098 2544
rect -3122 2510 -3106 2544
rect -2896 2510 -2880 2544
rect -1904 2510 -1888 2544
rect -1678 2510 -1662 2544
rect -686 2510 -670 2544
rect -460 2510 -444 2544
rect 532 2510 548 2544
rect 758 2510 774 2544
rect 1750 2510 1766 2544
rect 1976 2510 1992 2544
rect 2968 2510 2984 2544
rect 3194 2510 3210 2544
rect 4186 2510 4202 2544
rect -4284 2430 -4250 2492
rect 4338 2430 4372 2492
rect -4284 2396 -4188 2430
rect 4276 2396 4372 2430
rect -3724 2282 -3628 2316
rect 3618 2282 3714 2316
rect -3724 2220 -3690 2282
rect 3680 2220 3714 2282
rect -3554 2168 -3538 2202
rect -2562 2168 -2546 2202
rect -2336 2168 -2320 2202
rect -1344 2168 -1328 2202
rect -1118 2168 -1102 2202
rect -126 2168 -110 2202
rect 100 2168 116 2202
rect 1092 2168 1108 2202
rect 1318 2168 1334 2202
rect 2310 2168 2326 2202
rect 2536 2168 2552 2202
rect 3528 2168 3544 2202
rect -3622 2140 -3588 2156
rect -3622 1956 -3588 1972
rect -2512 2140 -2478 2156
rect -2512 1956 -2478 1972
rect -2404 2140 -2370 2156
rect -2404 1956 -2370 1972
rect -1294 2140 -1260 2156
rect -1294 1956 -1260 1972
rect -1186 2140 -1152 2156
rect -1186 1956 -1152 1972
rect -76 2140 -42 2156
rect -76 1956 -42 1972
rect 32 2140 66 2156
rect 32 1956 66 1972
rect 1142 2140 1176 2156
rect 1142 1956 1176 1972
rect 1250 2140 1284 2156
rect 1250 1956 1284 1972
rect 2360 2140 2394 2156
rect 2360 1956 2394 1972
rect 2468 2140 2502 2156
rect 2468 1956 2502 1972
rect 3578 2140 3612 2156
rect 3578 1956 3612 1972
rect -3554 1910 -3538 1944
rect -2562 1910 -2546 1944
rect -2336 1910 -2320 1944
rect -1344 1910 -1328 1944
rect -1118 1910 -1102 1944
rect -126 1910 -110 1944
rect 100 1910 116 1944
rect 1092 1910 1108 1944
rect 1318 1910 1334 1944
rect 2310 1910 2326 1944
rect 2536 1910 2552 1944
rect 3528 1910 3544 1944
rect -3724 1830 -3690 1892
rect 3680 1830 3714 1892
rect -3724 1796 -3628 1830
rect 3618 1796 3714 1830
rect -3030 1790 -2860 1796
rect -3030 1700 -3000 1790
rect -2890 1700 -2860 1790
rect -3030 1696 -2860 1700
rect 1880 1790 2050 1796
rect 1880 1700 1910 1790
rect 2020 1700 2050 1790
rect 1880 1696 2050 1700
rect -3724 1662 -3628 1696
rect 3618 1662 3714 1696
rect -3724 1600 -3690 1662
rect 3680 1600 3714 1662
rect -3554 1548 -3538 1582
rect -2562 1548 -2546 1582
rect -2336 1548 -2320 1582
rect -1344 1548 -1328 1582
rect -1118 1548 -1102 1582
rect -126 1548 -110 1582
rect 100 1548 116 1582
rect 1092 1548 1108 1582
rect 1318 1548 1334 1582
rect 2310 1548 2326 1582
rect 2536 1548 2552 1582
rect 3528 1548 3544 1582
rect -3622 1520 -3588 1536
rect -3622 1336 -3588 1352
rect -2512 1520 -2478 1536
rect -2512 1336 -2478 1352
rect -2404 1520 -2370 1536
rect -2404 1336 -2370 1352
rect -1294 1520 -1260 1536
rect -1294 1336 -1260 1352
rect -1186 1520 -1152 1536
rect -1186 1336 -1152 1352
rect -76 1520 -42 1536
rect -76 1336 -42 1352
rect 32 1520 66 1536
rect 32 1336 66 1352
rect 1142 1520 1176 1536
rect 1142 1336 1176 1352
rect 1250 1520 1284 1536
rect 1250 1336 1284 1352
rect 2360 1520 2394 1536
rect 2360 1336 2394 1352
rect 2468 1520 2502 1536
rect 2468 1336 2502 1352
rect 3578 1520 3612 1536
rect 3578 1336 3612 1352
rect -3554 1290 -3538 1324
rect -2562 1290 -2546 1324
rect -2336 1290 -2320 1324
rect -1344 1290 -1328 1324
rect -1118 1290 -1102 1324
rect -126 1290 -110 1324
rect 100 1290 116 1324
rect 1092 1290 1108 1324
rect 1318 1290 1334 1324
rect 2310 1290 2326 1324
rect 2536 1290 2552 1324
rect 3528 1290 3544 1324
rect -3724 1210 -3690 1272
rect 3680 1210 3714 1272
rect -3724 1176 -3628 1210
rect 3618 1176 3714 1210
rect -4284 1062 -4188 1096
rect 4276 1062 4372 1096
rect -4284 1000 -4250 1062
rect 4338 1000 4372 1062
rect -4114 948 -4098 982
rect -3122 948 -3106 982
rect -2896 948 -2880 982
rect -1904 948 -1888 982
rect -1678 948 -1662 982
rect -686 948 -670 982
rect -460 948 -444 982
rect 532 948 548 982
rect 758 948 774 982
rect 1750 948 1766 982
rect 1976 948 1992 982
rect 2968 948 2984 982
rect 3194 948 3210 982
rect 4186 948 4202 982
rect -4182 920 -4148 936
rect -4182 736 -4148 752
rect -3072 920 -3038 936
rect -3072 736 -3038 752
rect -2964 920 -2930 936
rect -2964 736 -2930 752
rect -1854 920 -1820 936
rect -1854 736 -1820 752
rect -1746 920 -1712 936
rect -1746 736 -1712 752
rect -636 920 -602 936
rect -636 736 -602 752
rect -528 920 -494 936
rect -528 736 -494 752
rect 582 920 616 936
rect 582 736 616 752
rect 690 920 724 936
rect 690 736 724 752
rect 1800 920 1834 936
rect 1800 736 1834 752
rect 1908 920 1942 936
rect 1908 736 1942 752
rect 3018 920 3052 936
rect 3018 736 3052 752
rect 3126 920 3160 936
rect 3126 736 3160 752
rect 4236 920 4270 936
rect 4236 736 4270 752
rect -4114 690 -4098 724
rect -3122 690 -3106 724
rect -2896 690 -2880 724
rect -1904 690 -1888 724
rect -1678 690 -1662 724
rect -686 690 -670 724
rect -460 690 -444 724
rect 532 690 548 724
rect 758 690 774 724
rect 1750 690 1766 724
rect 1976 690 1992 724
rect 2968 690 2984 724
rect 3194 690 3210 724
rect 4186 690 4202 724
rect -4284 610 -4250 672
rect 4338 610 4372 672
rect -4284 576 -4188 610
rect 4276 576 4372 610
rect -4284 462 -4188 496
rect 4276 462 4372 496
rect -4284 400 -4250 462
rect 4338 400 4372 462
rect -4114 348 -4098 382
rect -3122 348 -3106 382
rect -2896 348 -2880 382
rect -1904 348 -1888 382
rect -1678 348 -1662 382
rect -686 348 -670 382
rect -460 348 -444 382
rect 532 348 548 382
rect 758 348 774 382
rect 1750 348 1766 382
rect 1976 348 1992 382
rect 2968 348 2984 382
rect 3194 348 3210 382
rect 4186 348 4202 382
rect -4182 320 -4148 336
rect -4182 136 -4148 152
rect -3072 320 -3038 336
rect -3072 136 -3038 152
rect -2964 320 -2930 336
rect -2964 136 -2930 152
rect -1854 320 -1820 336
rect -1854 136 -1820 152
rect -1746 320 -1712 336
rect -1746 136 -1712 152
rect -636 320 -602 336
rect -636 136 -602 152
rect -528 320 -494 336
rect -528 136 -494 152
rect 582 320 616 336
rect 582 136 616 152
rect 690 320 724 336
rect 690 136 724 152
rect 1800 320 1834 336
rect 1800 136 1834 152
rect 1908 320 1942 336
rect 1908 136 1942 152
rect 3018 320 3052 336
rect 3018 136 3052 152
rect 3126 320 3160 336
rect 3126 136 3160 152
rect 4236 320 4270 336
rect 4236 136 4270 152
rect -4114 90 -4098 124
rect -3122 90 -3106 124
rect -2896 90 -2880 124
rect -1904 90 -1888 124
rect -1678 90 -1662 124
rect -686 90 -670 124
rect -460 90 -444 124
rect 532 90 548 124
rect 758 90 774 124
rect 1750 90 1766 124
rect 1976 90 1992 124
rect 2968 90 2984 124
rect 3194 90 3210 124
rect 4186 90 4202 124
rect -4284 10 -4250 72
rect 4338 10 4372 72
rect -4284 -24 -4188 10
rect 4276 -24 4372 10
<< viali >>
rect -2600 9036 -2510 9100
rect -2430 9036 -2340 9100
rect -110 9036 -20 9100
rect 60 9036 150 9100
rect 2350 9036 2430 9110
rect 2520 9036 2600 9110
rect -2600 9030 -2510 9036
rect -2430 9030 -2340 9036
rect -110 9030 -20 9036
rect 60 9030 150 9036
rect 2350 9030 2430 9036
rect 2520 9030 2600 9036
rect -4189 8888 -3213 8922
rect -2953 8888 -1977 8922
rect -1717 8888 -741 8922
rect -481 8888 495 8922
rect 755 8888 1731 8922
rect 1991 8888 2967 8922
rect 3227 8888 4203 8922
rect -4282 8792 -4248 8860
rect -3154 8792 -3120 8860
rect -3046 8792 -3012 8860
rect -1918 8792 -1884 8860
rect -1810 8792 -1776 8860
rect -682 8792 -648 8860
rect -574 8792 -540 8860
rect 554 8792 588 8860
rect 662 8792 696 8860
rect 1790 8792 1824 8860
rect 1898 8792 1932 8860
rect 3026 8792 3060 8860
rect 3134 8792 3168 8860
rect 4262 8792 4296 8860
rect -4189 8730 -3213 8764
rect -2953 8730 -1977 8764
rect -1717 8730 -741 8764
rect -481 8730 495 8764
rect 755 8730 1731 8764
rect 1991 8730 2967 8764
rect 3227 8730 4203 8764
rect -4189 8348 -3213 8382
rect -2953 8348 -1977 8382
rect -1717 8348 -741 8382
rect -481 8348 495 8382
rect 755 8348 1731 8382
rect 1991 8348 2967 8382
rect 3227 8348 4203 8382
rect -4282 8252 -4248 8320
rect -3154 8252 -3120 8320
rect -3046 8252 -3012 8320
rect -1918 8252 -1884 8320
rect -1810 8252 -1776 8320
rect -682 8252 -648 8320
rect -574 8252 -540 8320
rect 554 8252 588 8320
rect 662 8252 696 8320
rect 1790 8252 1824 8320
rect 1898 8252 1932 8320
rect 3026 8252 3060 8320
rect 3134 8252 3168 8320
rect 4262 8252 4296 8320
rect -4189 8190 -3213 8224
rect -2953 8190 -1977 8224
rect -1717 8190 -741 8224
rect -481 8190 495 8224
rect 755 8190 1731 8224
rect 1991 8190 2967 8224
rect 3227 8190 4203 8224
rect -2590 7980 -2500 8050
rect -2450 7980 -2360 8050
rect -110 7980 -20 8050
rect 50 7990 140 8060
rect 2350 7990 2430 8060
rect 2520 7990 2600 8060
rect -4189 7808 -3213 7842
rect -2953 7808 -1977 7842
rect -1717 7808 -741 7842
rect -481 7808 495 7842
rect 755 7808 1731 7842
rect 1991 7808 2967 7842
rect 3227 7808 4203 7842
rect -4282 7712 -4248 7780
rect -3154 7712 -3120 7780
rect -3046 7712 -3012 7780
rect -1918 7712 -1884 7780
rect -1810 7712 -1776 7780
rect -682 7712 -648 7780
rect -574 7712 -540 7780
rect 554 7712 588 7780
rect 662 7712 696 7780
rect 1790 7712 1824 7780
rect 1898 7712 1932 7780
rect 3026 7712 3060 7780
rect 3134 7712 3168 7780
rect 4262 7712 4296 7780
rect -4189 7650 -3213 7684
rect -2953 7650 -1977 7684
rect -1717 7650 -741 7684
rect -481 7650 495 7684
rect 755 7650 1731 7684
rect 1991 7650 2967 7684
rect 3227 7650 4203 7684
rect -2590 7440 -2510 7520
rect -2420 7440 -2340 7520
rect -110 7440 -30 7520
rect 60 7440 140 7520
rect 2350 7440 2430 7520
rect 2520 7440 2600 7520
rect -4189 7268 -3213 7302
rect -2953 7268 -1977 7302
rect -1717 7268 -741 7302
rect -481 7268 495 7302
rect 755 7268 1731 7302
rect 1991 7268 2967 7302
rect 3227 7268 4203 7302
rect -4282 7172 -4248 7240
rect -3154 7172 -3120 7240
rect -3046 7172 -3012 7240
rect -1918 7172 -1884 7240
rect -1810 7172 -1776 7240
rect -682 7172 -648 7240
rect -574 7172 -540 7240
rect 554 7172 588 7240
rect 662 7172 696 7240
rect 1790 7172 1824 7240
rect 1898 7172 1932 7240
rect 3026 7172 3060 7240
rect 3134 7172 3168 7240
rect 4262 7172 4296 7240
rect -4189 7110 -3213 7144
rect -2953 7110 -1977 7144
rect -1717 7110 -741 7144
rect -481 7110 495 7144
rect 755 7110 1731 7144
rect 1991 7110 2967 7144
rect 3227 7110 4203 7144
rect -4189 6688 -3213 6722
rect -2953 6688 -1977 6722
rect -1717 6688 -741 6722
rect -481 6688 495 6722
rect 755 6688 1731 6722
rect 1991 6688 2967 6722
rect 3227 6688 4203 6722
rect -4282 6592 -4248 6660
rect -3154 6592 -3120 6660
rect -3046 6592 -3012 6660
rect -1918 6592 -1884 6660
rect -1810 6592 -1776 6660
rect -682 6592 -648 6660
rect -574 6592 -540 6660
rect 554 6592 588 6660
rect 662 6592 696 6660
rect 1790 6592 1824 6660
rect 1898 6592 1932 6660
rect 3026 6592 3060 6660
rect 3134 6592 3168 6660
rect 4262 6592 4296 6660
rect -4189 6530 -3213 6564
rect -2953 6530 -1977 6564
rect -1717 6530 -741 6564
rect -481 6530 495 6564
rect 755 6530 1731 6564
rect 1991 6530 2967 6564
rect 3227 6530 4203 6564
rect -2590 6280 -2500 6360
rect -2430 6280 -2340 6360
rect -110 6280 -30 6350
rect 60 6280 140 6350
rect 2350 6280 2430 6350
rect 2520 6280 2600 6350
rect -9829 4979 -9432 6093
rect -7398 4979 -7001 6093
rect -4189 6108 -3213 6142
rect -2953 6108 -1977 6142
rect -1717 6108 -741 6142
rect -481 6108 495 6142
rect 755 6108 1731 6142
rect 1991 6108 2967 6142
rect 3227 6108 4203 6142
rect -4282 6012 -4248 6080
rect -3154 6012 -3120 6080
rect -3046 6012 -3012 6080
rect -1918 6012 -1884 6080
rect -1810 6012 -1776 6080
rect -682 6012 -648 6080
rect -574 6012 -540 6080
rect 554 6012 588 6080
rect 662 6012 696 6080
rect 1790 6012 1824 6080
rect 1898 6012 1932 6080
rect 3026 6012 3060 6080
rect 3134 6012 3168 6080
rect 4262 6012 4296 6080
rect -4189 5950 -3213 5984
rect -2953 5950 -1977 5984
rect -1717 5950 -741 5984
rect -481 5950 495 5984
rect 755 5950 1731 5984
rect 1991 5950 2967 5984
rect 3227 5950 4203 5984
rect -6029 5568 -5053 5602
rect -4793 5568 -3817 5602
rect -3557 5568 -2581 5602
rect -2321 5568 -1345 5602
rect -1085 5568 -109 5602
rect 151 5568 1127 5602
rect 1387 5568 2363 5602
rect 2623 5568 3599 5602
rect 3859 5568 4835 5602
rect 5095 5568 6071 5602
rect -6122 5472 -6088 5540
rect -4994 5472 -4960 5540
rect -4886 5472 -4852 5540
rect -3758 5472 -3724 5540
rect -3650 5472 -3616 5540
rect -2522 5472 -2488 5540
rect -2414 5472 -2380 5540
rect -1286 5472 -1252 5540
rect -1178 5472 -1144 5540
rect -50 5472 -16 5540
rect 58 5472 92 5540
rect 1186 5472 1220 5540
rect 1294 5472 1328 5540
rect 2422 5472 2456 5540
rect 2530 5472 2564 5540
rect 3658 5472 3692 5540
rect 3766 5472 3800 5540
rect 4894 5472 4928 5540
rect 5002 5472 5036 5540
rect 6130 5472 6164 5540
rect -6029 5410 -5053 5444
rect -4793 5410 -3817 5444
rect -3557 5410 -2581 5444
rect -2321 5410 -1345 5444
rect -1085 5410 -109 5444
rect 151 5410 1127 5444
rect 1387 5410 2363 5444
rect 2623 5410 3599 5444
rect 3859 5410 4835 5444
rect 5095 5410 6071 5444
rect -4450 5200 -4360 5280
rect -4270 5200 -4180 5280
rect -1920 5200 -1830 5280
rect -1760 5200 -1670 5280
rect 550 5200 640 5280
rect 710 5200 800 5280
rect 3000 5200 3090 5280
rect 3160 5200 3250 5280
rect 5500 5200 5590 5280
rect 5660 5200 5750 5280
rect -6029 5028 -5053 5062
rect -4793 5028 -3817 5062
rect -3557 5028 -2581 5062
rect -2321 5028 -1345 5062
rect -1085 5028 -109 5062
rect 151 5028 1127 5062
rect 1387 5028 2363 5062
rect 2623 5028 3599 5062
rect 3859 5028 4835 5062
rect 5095 5028 6071 5062
rect -6122 4932 -6088 5000
rect -4994 4932 -4960 5000
rect -4886 4932 -4852 5000
rect -3758 4932 -3724 5000
rect -3650 4932 -3616 5000
rect -2522 4932 -2488 5000
rect -2414 4932 -2380 5000
rect -1286 4932 -1252 5000
rect -1178 4932 -1144 5000
rect -50 4932 -16 5000
rect 58 4932 92 5000
rect 1186 4932 1220 5000
rect 1294 4932 1328 5000
rect 2422 4932 2456 5000
rect 2530 4932 2564 5000
rect 3658 4932 3692 5000
rect 3766 4932 3800 5000
rect 4894 4932 4928 5000
rect 5002 4932 5036 5000
rect 6130 4932 6164 5000
rect -6029 4870 -5053 4904
rect -4793 4870 -3817 4904
rect -3557 4870 -2581 4904
rect -2321 4870 -1345 4904
rect -1085 4870 -109 4904
rect 151 4870 1127 4904
rect 1387 4870 2363 4904
rect 2623 4870 3599 4904
rect 3859 4870 4835 4904
rect 5095 4870 6071 4904
rect 7231 4979 7628 6093
rect 9662 4979 10059 6093
rect -9829 3509 -9432 4623
rect -7398 3509 -7001 4623
rect -6029 4488 -5053 4522
rect -4793 4488 -3817 4522
rect -3557 4488 -2581 4522
rect -2321 4488 -1345 4522
rect -1085 4488 -109 4522
rect 151 4488 1127 4522
rect 1387 4488 2363 4522
rect 2623 4488 3599 4522
rect 3859 4488 4835 4522
rect 5095 4488 6071 4522
rect -6122 4392 -6088 4460
rect -4994 4392 -4960 4460
rect -4886 4392 -4852 4460
rect -3758 4392 -3724 4460
rect -3650 4392 -3616 4460
rect -2522 4392 -2488 4460
rect -2414 4392 -2380 4460
rect -1286 4392 -1252 4460
rect -1178 4392 -1144 4460
rect -50 4392 -16 4460
rect 58 4392 92 4460
rect 1186 4392 1220 4460
rect 1294 4392 1328 4460
rect 2422 4392 2456 4460
rect 2530 4392 2564 4460
rect 3658 4392 3692 4460
rect 3766 4392 3800 4460
rect 4894 4392 4928 4460
rect 5002 4392 5036 4460
rect 6130 4392 6164 4460
rect -6029 4330 -5053 4364
rect -4793 4330 -3817 4364
rect -3557 4330 -2581 4364
rect -2321 4330 -1345 4364
rect -1085 4330 -109 4364
rect 151 4330 1127 4364
rect 1387 4330 2363 4364
rect 2623 4330 3599 4364
rect 3859 4330 4835 4364
rect 5095 4330 6071 4364
rect -4450 4120 -4360 4200
rect -4270 4130 -4180 4210
rect -1920 4120 -1830 4200
rect -1760 4120 -1670 4200
rect 550 4120 640 4200
rect 710 4120 800 4200
rect 3000 4120 3090 4200
rect 3160 4120 3250 4200
rect 5500 4120 5590 4200
rect 5660 4120 5750 4200
rect -6029 3948 -5053 3982
rect -4793 3948 -3817 3982
rect -3557 3948 -2581 3982
rect -2321 3948 -1345 3982
rect -1085 3948 -109 3982
rect 151 3948 1127 3982
rect 1387 3948 2363 3982
rect 2623 3948 3599 3982
rect 3859 3948 4835 3982
rect 5095 3948 6071 3982
rect -6122 3852 -6088 3920
rect -4994 3852 -4960 3920
rect -4886 3852 -4852 3920
rect -3758 3852 -3724 3920
rect -3650 3852 -3616 3920
rect -2522 3852 -2488 3920
rect -2414 3852 -2380 3920
rect -1286 3852 -1252 3920
rect -1178 3852 -1144 3920
rect -50 3852 -16 3920
rect 58 3852 92 3920
rect 1186 3852 1220 3920
rect 1294 3852 1328 3920
rect 2422 3852 2456 3920
rect 2530 3852 2564 3920
rect 3658 3852 3692 3920
rect 3766 3852 3800 3920
rect 4894 3852 4928 3920
rect 5002 3852 5036 3920
rect 6130 3852 6164 3920
rect -6029 3790 -5053 3824
rect -4793 3790 -3817 3824
rect -3557 3790 -2581 3824
rect -2321 3790 -1345 3824
rect -1085 3790 -109 3824
rect 151 3790 1127 3824
rect 1387 3790 2363 3824
rect 2623 3790 3599 3824
rect 3859 3790 4835 3824
rect 5095 3790 6071 3824
rect -8810 3363 -8720 3390
rect -8600 3363 -8510 3390
rect 7231 3509 7628 4623
rect 9662 3509 10059 4623
rect 8500 3363 8570 3380
rect 8660 3363 8730 3380
rect -8810 3260 -8720 3363
rect -8600 3260 -8510 3363
rect 8500 3290 8570 3363
rect 8660 3290 8730 3363
rect -4098 3168 -3122 3202
rect -2880 3168 -1904 3202
rect -1662 3168 -686 3202
rect -444 3168 532 3202
rect 774 3168 1750 3202
rect 1992 3168 2968 3202
rect 3210 3168 4186 3202
rect -4182 3072 -4148 3140
rect -3072 3072 -3038 3140
rect -2964 3072 -2930 3140
rect -1854 3072 -1820 3140
rect -1746 3072 -1712 3140
rect -636 3072 -602 3140
rect -528 3072 -494 3140
rect 582 3072 616 3140
rect 690 3072 724 3140
rect 1800 3072 1834 3140
rect 1908 3072 1942 3140
rect 3018 3072 3052 3140
rect 3126 3072 3160 3140
rect 4236 3072 4270 3140
rect -4098 3010 -3122 3044
rect -2880 3010 -1904 3044
rect -1662 3010 -686 3044
rect -444 3010 532 3044
rect 774 3010 1750 3044
rect 1992 3010 2968 3044
rect 3210 3010 4186 3044
rect -2290 2896 -2180 2910
rect -1430 2896 -1320 2910
rect -220 2896 -110 2910
rect 630 2896 740 2910
rect 2200 2896 2310 2910
rect 3080 2896 3190 2910
rect -2290 2816 -2180 2896
rect -1430 2816 -1320 2896
rect -220 2816 -110 2896
rect 630 2816 740 2896
rect 2200 2816 2310 2896
rect 3080 2816 3190 2896
rect -2290 2800 -2180 2816
rect -1430 2800 -1320 2816
rect -220 2800 -110 2816
rect 630 2800 740 2816
rect 2200 2800 2310 2816
rect 3080 2800 3190 2816
rect -4098 2668 -3122 2702
rect -2880 2668 -1904 2702
rect -1662 2668 -686 2702
rect -444 2668 532 2702
rect 774 2668 1750 2702
rect 1992 2668 2968 2702
rect 3210 2668 4186 2702
rect -4182 2572 -4148 2640
rect -3072 2572 -3038 2640
rect -2964 2572 -2930 2640
rect -1854 2572 -1820 2640
rect -1746 2572 -1712 2640
rect -636 2572 -602 2640
rect -528 2572 -494 2640
rect 582 2572 616 2640
rect 690 2572 724 2640
rect 1800 2572 1834 2640
rect 1908 2572 1942 2640
rect 3018 2572 3052 2640
rect 3126 2572 3160 2640
rect 4236 2572 4270 2640
rect -4098 2510 -3122 2544
rect -2880 2510 -1904 2544
rect -1662 2510 -686 2544
rect -444 2510 532 2544
rect 774 2510 1750 2544
rect 1992 2510 2968 2544
rect 3210 2510 4186 2544
rect -3538 2168 -2562 2202
rect -2320 2168 -1344 2202
rect -1102 2168 -126 2202
rect 116 2168 1092 2202
rect 1334 2168 2310 2202
rect 2552 2168 3528 2202
rect -3622 1972 -3588 2140
rect -2512 1972 -2478 2140
rect -2404 1972 -2370 2140
rect -1294 1972 -1260 2140
rect -1186 1972 -1152 2140
rect -76 1972 -42 2140
rect 32 1972 66 2140
rect 1142 1972 1176 2140
rect 1250 1972 1284 2140
rect 2360 1972 2394 2140
rect 2468 1972 2502 2140
rect 3578 1972 3612 2140
rect -3538 1910 -2562 1944
rect -2320 1910 -1344 1944
rect -1102 1910 -126 1944
rect 116 1910 1092 1944
rect 1334 1910 2310 1944
rect 2552 1910 3528 1944
rect -3000 1700 -2890 1790
rect 1910 1700 2020 1790
rect -3538 1548 -2562 1582
rect -2320 1548 -1344 1582
rect -1102 1548 -126 1582
rect 116 1548 1092 1582
rect 1334 1548 2310 1582
rect 2552 1548 3528 1582
rect -3622 1352 -3588 1520
rect -2512 1352 -2478 1520
rect -2404 1352 -2370 1520
rect -1294 1352 -1260 1520
rect -1186 1352 -1152 1520
rect -76 1352 -42 1520
rect 32 1352 66 1520
rect 1142 1352 1176 1520
rect 1250 1352 1284 1520
rect 2360 1352 2394 1520
rect 2468 1352 2502 1520
rect 3578 1352 3612 1520
rect -3538 1290 -2562 1324
rect -2320 1290 -1344 1324
rect -1102 1290 -126 1324
rect 116 1290 1092 1324
rect 1334 1290 2310 1324
rect 2552 1290 3528 1324
rect -4098 948 -3122 982
rect -2880 948 -1904 982
rect -1662 948 -686 982
rect -444 948 532 982
rect 774 948 1750 982
rect 1992 948 2968 982
rect 3210 948 4186 982
rect -4182 752 -4148 920
rect -3072 752 -3038 920
rect -2964 752 -2930 920
rect -1854 752 -1820 920
rect -1746 752 -1712 920
rect -636 752 -602 920
rect -528 752 -494 920
rect 582 752 616 920
rect 690 752 724 920
rect 1800 752 1834 920
rect 1908 752 1942 920
rect 3018 752 3052 920
rect 3126 752 3160 920
rect 4236 752 4270 920
rect -4098 690 -3122 724
rect -2880 690 -1904 724
rect -1662 690 -686 724
rect -444 690 532 724
rect 774 690 1750 724
rect 1992 690 2968 724
rect 3210 690 4186 724
rect -3060 576 -2940 590
rect -1840 576 -1720 590
rect -630 576 -510 590
rect 590 576 710 590
rect 1820 576 1940 580
rect 3030 576 3150 590
rect -3060 496 -2940 576
rect -1840 496 -1720 576
rect -630 496 -510 576
rect 590 496 710 576
rect 1820 496 1940 576
rect 3030 496 3150 576
rect -3060 490 -2940 496
rect -1840 490 -1720 496
rect -630 490 -510 496
rect 590 490 710 496
rect 1820 480 1940 496
rect 3030 490 3150 496
rect -4098 348 -3122 382
rect -2880 348 -1904 382
rect -1662 348 -686 382
rect -444 348 532 382
rect 774 348 1750 382
rect 1992 348 2968 382
rect 3210 348 4186 382
rect -4182 152 -4148 320
rect -3072 152 -3038 320
rect -2964 152 -2930 320
rect -1854 152 -1820 320
rect -1746 152 -1712 320
rect -636 152 -602 320
rect -528 152 -494 320
rect 582 152 616 320
rect 690 152 724 320
rect 1800 152 1834 320
rect 1908 152 1942 320
rect 3018 152 3052 320
rect 3126 152 3160 320
rect 4236 152 4270 320
rect -4098 90 -3122 124
rect -2880 90 -1904 124
rect -1662 90 -686 124
rect -444 90 532 124
rect 774 90 1750 124
rect 1992 90 2968 124
rect 3210 90 4186 124
<< metal1 >>
rect 2338 9110 2442 9116
rect -2612 9100 -2498 9106
rect -2612 9030 -2600 9100
rect -2510 9030 -2498 9100
rect -2612 9024 -2498 9030
rect -2442 9100 -2328 9106
rect -2442 9030 -2430 9100
rect -2340 9030 -2328 9100
rect -2442 9024 -2328 9030
rect -122 9100 -8 9106
rect -122 9030 -110 9100
rect -20 9030 -8 9100
rect -122 9024 -8 9030
rect 48 9100 162 9106
rect 48 9030 60 9100
rect 150 9030 162 9100
rect 48 9024 162 9030
rect 2338 9030 2350 9110
rect 2430 9030 2442 9110
rect 2338 9024 2442 9030
rect 2508 9110 2612 9116
rect 2508 9030 2520 9110
rect 2600 9030 2612 9110
rect 2508 9024 2612 9030
rect -2610 8940 -2600 8990
rect -4210 8922 -2600 8940
rect -2520 8940 -2510 8990
rect -2440 8940 -2430 8990
rect -2520 8922 -2430 8940
rect -2350 8940 -2340 8990
rect -120 8940 -110 8990
rect -2350 8922 -110 8940
rect -30 8940 -20 8990
rect 50 8940 60 8990
rect -30 8922 60 8940
rect 140 8940 150 8990
rect 2340 8940 2350 8980
rect 140 8922 2350 8940
rect 2430 8940 2440 8980
rect 2510 8940 2520 8980
rect 2430 8922 2520 8940
rect 2600 8940 2610 8980
rect 2600 8922 4230 8940
rect -4210 8900 -4189 8922
rect -4201 8888 -4189 8900
rect -3213 8900 -2953 8922
rect -3213 8888 -3201 8900
rect -4201 8882 -3201 8888
rect -2965 8888 -2953 8900
rect -1977 8900 -1717 8922
rect -1977 8888 -1965 8900
rect -2965 8882 -1965 8888
rect -1729 8888 -1717 8900
rect -741 8900 -481 8922
rect -741 8888 -729 8900
rect -1729 8882 -729 8888
rect -493 8888 -481 8900
rect 495 8900 755 8922
rect 495 8888 507 8900
rect -493 8882 507 8888
rect 743 8888 755 8900
rect 1731 8900 1991 8922
rect 2967 8900 3227 8922
rect 1731 8888 1743 8900
rect 743 8882 1743 8888
rect 1979 8888 1991 8900
rect 2967 8888 2979 8900
rect 1979 8882 2979 8888
rect 3215 8888 3227 8900
rect 4203 8900 4230 8922
rect 4203 8888 4215 8900
rect 3215 8882 4215 8888
rect -4288 8860 -4242 8872
rect -4288 8810 -4282 8860
rect -4300 8792 -4282 8810
rect -4248 8850 -4242 8860
rect -3160 8860 -3114 8872
rect -3052 8860 -3006 8872
rect -3160 8850 -3154 8860
rect -4248 8820 -3154 8850
rect -4248 8792 -3480 8820
rect -4300 8764 -3480 8792
rect -3400 8764 -3330 8820
rect -3250 8792 -3154 8820
rect -3012 8850 -3006 8860
rect -1924 8860 -1878 8872
rect -1816 8860 -1770 8872
rect -688 8860 -642 8872
rect -580 8860 -534 8872
rect -1924 8850 -1918 8860
rect -3012 8792 -1918 8850
rect -1776 8850 -1770 8860
rect -690 8850 -682 8860
rect -1776 8820 -682 8850
rect -1776 8792 -990 8820
rect -3250 8790 -3150 8792
rect -3020 8790 -1910 8792
rect -1780 8790 -990 8792
rect -3250 8764 -990 8790
rect -910 8764 -840 8820
rect -760 8792 -682 8820
rect -540 8850 -534 8860
rect 548 8860 594 8872
rect 656 8860 702 8872
rect 548 8850 554 8860
rect -540 8792 554 8850
rect 696 8850 702 8860
rect 1784 8860 1830 8872
rect 1892 8860 1938 8872
rect 3020 8860 3066 8872
rect 3128 8860 3174 8872
rect 1784 8850 1790 8860
rect 696 8820 1790 8850
rect 696 8792 1490 8820
rect -760 8790 -680 8792
rect -550 8790 560 8792
rect 690 8790 1490 8792
rect -760 8764 1490 8790
rect 1570 8764 1640 8820
rect 1720 8792 1790 8820
rect 1932 8850 1940 8860
rect 3020 8850 3026 8860
rect 1932 8792 3026 8850
rect 3168 8850 3174 8860
rect 4256 8860 4302 8872
rect 4256 8850 4262 8860
rect 3168 8792 4262 8850
rect 4296 8810 4302 8860
rect 4296 8792 4310 8810
rect 1720 8790 1800 8792
rect 1930 8790 3030 8792
rect 3160 8790 4310 8792
rect 1720 8764 4310 8790
rect -4300 8730 -4189 8764
rect -3213 8730 -2953 8764
rect -1977 8730 -1717 8764
rect -741 8730 -481 8764
rect 495 8730 755 8764
rect 1731 8730 1991 8764
rect 2967 8730 3227 8764
rect 4203 8730 4310 8764
rect -4300 8710 -3870 8730
rect -3880 8670 -3870 8710
rect -3790 8710 -3700 8730
rect -3790 8670 -3780 8710
rect -3710 8670 -3700 8710
rect -3620 8710 -1350 8730
rect -3620 8670 -3610 8710
rect -1360 8670 -1350 8710
rect -1270 8710 -1180 8730
rect -1270 8670 -1260 8710
rect -1190 8670 -1180 8710
rect -1100 8710 1140 8730
rect -1100 8670 -1090 8710
rect 1130 8670 1140 8710
rect 1220 8710 1310 8730
rect 1220 8670 1230 8710
rect 1300 8670 1310 8710
rect 1390 8710 3590 8730
rect 1390 8670 1400 8710
rect 3580 8670 3590 8710
rect 3670 8710 3760 8730
rect 3670 8670 3680 8710
rect 3750 8670 3760 8710
rect 3840 8710 4310 8730
rect 3840 8670 3850 8710
rect -2610 8400 -2600 8450
rect -4210 8382 -2600 8400
rect -2520 8400 -2510 8450
rect -2440 8400 -2430 8450
rect -2520 8382 -2430 8400
rect -2350 8400 -2340 8450
rect -120 8400 -110 8450
rect -2350 8382 -110 8400
rect -30 8400 -20 8450
rect 50 8400 60 8450
rect -30 8382 60 8400
rect 140 8400 150 8450
rect 2340 8400 2350 8440
rect 140 8382 2350 8400
rect 2430 8400 2440 8440
rect 2510 8400 2520 8440
rect 2430 8382 2520 8400
rect 2600 8400 2610 8440
rect 2600 8382 4230 8400
rect -4210 8360 -4189 8382
rect -4201 8348 -4189 8360
rect -3213 8360 -2953 8382
rect -3213 8348 -3201 8360
rect -4201 8342 -3201 8348
rect -2965 8348 -2953 8360
rect -1977 8360 -1717 8382
rect -1977 8348 -1965 8360
rect -2965 8342 -1965 8348
rect -1729 8348 -1717 8360
rect -741 8360 -481 8382
rect -741 8348 -729 8360
rect -1729 8342 -729 8348
rect -493 8348 -481 8360
rect 495 8360 755 8382
rect 495 8348 507 8360
rect -493 8342 507 8348
rect 743 8348 755 8360
rect 1731 8360 1991 8382
rect 2967 8360 3227 8382
rect 1731 8348 1743 8360
rect 743 8342 1743 8348
rect 1979 8348 1991 8360
rect 2967 8348 2979 8360
rect 1979 8342 2979 8348
rect 3215 8348 3227 8360
rect 4203 8360 4230 8382
rect 4203 8348 4215 8360
rect 3215 8342 4215 8348
rect -4288 8320 -4242 8332
rect -4288 8270 -4282 8320
rect -4290 8252 -4282 8270
rect -4248 8310 -4242 8320
rect -3160 8320 -3114 8332
rect -3052 8320 -3006 8332
rect -3160 8310 -3154 8320
rect -4248 8280 -3154 8310
rect -4248 8252 -3480 8280
rect -4290 8224 -3480 8252
rect -3400 8224 -3330 8280
rect -3250 8252 -3154 8280
rect -3012 8310 -3006 8320
rect -1924 8320 -1878 8332
rect -1816 8320 -1770 8332
rect -688 8320 -642 8332
rect -580 8320 -534 8332
rect -1924 8310 -1918 8320
rect -3012 8252 -1918 8310
rect -1776 8310 -1770 8320
rect -690 8310 -682 8320
rect -1776 8280 -682 8310
rect -1776 8252 -990 8280
rect -3250 8250 -3150 8252
rect -3020 8250 -1910 8252
rect -1780 8250 -990 8252
rect -3250 8224 -990 8250
rect -910 8224 -840 8280
rect -760 8252 -682 8280
rect -540 8310 -534 8320
rect 548 8320 594 8332
rect 656 8320 702 8332
rect 548 8310 554 8320
rect -540 8252 554 8310
rect 696 8310 702 8320
rect 1784 8320 1830 8332
rect 1892 8320 1938 8332
rect 3020 8320 3066 8332
rect 3128 8320 3174 8332
rect 1784 8310 1790 8320
rect 696 8280 1790 8310
rect 696 8252 1490 8280
rect -760 8250 -680 8252
rect -550 8250 560 8252
rect 690 8250 1490 8252
rect -760 8224 1490 8250
rect 1570 8224 1640 8280
rect 1720 8252 1790 8280
rect 1932 8310 1940 8320
rect 3020 8310 3026 8320
rect 1932 8252 3026 8310
rect 3168 8310 3174 8320
rect 4256 8320 4302 8332
rect 4256 8310 4262 8320
rect 3168 8252 4262 8310
rect 4296 8252 4302 8320
rect 1720 8250 1800 8252
rect 1930 8250 3030 8252
rect 3160 8250 4302 8252
rect 1720 8240 4302 8250
rect 1720 8224 4290 8240
rect -4290 8190 -4189 8224
rect -3213 8190 -2953 8224
rect -1977 8190 -1717 8224
rect -741 8190 -481 8224
rect 495 8190 755 8224
rect 1731 8190 1991 8224
rect 2967 8190 3227 8224
rect 4203 8190 4290 8224
rect -4290 8170 -3870 8190
rect -3880 8130 -3870 8170
rect -3790 8170 -3700 8190
rect -3790 8130 -3780 8170
rect -3710 8130 -3700 8170
rect -3620 8170 -1350 8190
rect -3620 8130 -3610 8170
rect -1360 8130 -1350 8170
rect -1270 8170 -1180 8190
rect -1270 8130 -1260 8170
rect -1190 8130 -1180 8170
rect -1100 8170 1140 8190
rect -1100 8130 -1090 8170
rect 1130 8130 1140 8170
rect 1220 8170 1310 8190
rect 1220 8130 1230 8170
rect 1300 8130 1310 8170
rect 1390 8170 3590 8190
rect 1390 8130 1400 8170
rect 3580 8120 3590 8170
rect 3670 8170 3760 8190
rect 3670 8120 3680 8170
rect 3750 8120 3760 8170
rect 3840 8170 4290 8190
rect 3840 8120 3850 8170
rect -2600 8056 -2340 8090
rect 38 8060 152 8066
rect -2602 8050 -2340 8056
rect -2602 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -2340 8050
rect -2602 7974 -2340 7980
rect -122 8050 -8 8056
rect -122 7980 -110 8050
rect -20 7980 -8 8050
rect 38 7990 50 8060
rect 140 7990 152 8060
rect 38 7984 152 7990
rect 2338 8060 2442 8066
rect 2338 7990 2350 8060
rect 2430 7990 2442 8060
rect 2338 7984 2442 7990
rect 2508 8060 2612 8066
rect 2508 7990 2520 8060
rect 2600 7990 2612 8060
rect 2508 7984 2612 7990
rect -122 7974 -8 7980
rect -2600 7940 -2340 7974
rect -2610 7860 -2600 7910
rect -4210 7842 -2600 7860
rect -2520 7860 -2510 7910
rect -2440 7860 -2430 7910
rect -2520 7842 -2430 7860
rect -2350 7860 -2340 7910
rect -120 7860 -110 7920
rect -2350 7842 -110 7860
rect -30 7860 -20 7920
rect 50 7860 60 7920
rect -30 7842 60 7860
rect 140 7860 150 7920
rect 2340 7860 2350 7900
rect 140 7842 2350 7860
rect 2430 7860 2440 7900
rect 2510 7860 2520 7900
rect 2430 7842 2520 7860
rect 2600 7860 2610 7900
rect 2600 7842 4230 7860
rect -4210 7820 -4189 7842
rect -4201 7808 -4189 7820
rect -3213 7820 -2953 7842
rect -3213 7808 -3201 7820
rect -4201 7802 -3201 7808
rect -2965 7808 -2953 7820
rect -1977 7820 -1717 7842
rect -1977 7808 -1965 7820
rect -2965 7802 -1965 7808
rect -1729 7808 -1717 7820
rect -741 7820 -481 7842
rect -741 7808 -729 7820
rect -1729 7802 -729 7808
rect -493 7808 -481 7820
rect 495 7820 755 7842
rect 495 7808 507 7820
rect -493 7802 507 7808
rect 743 7808 755 7820
rect 1731 7820 1991 7842
rect 2967 7820 3227 7842
rect 1731 7808 1743 7820
rect 743 7802 1743 7808
rect 1979 7808 1991 7820
rect 2967 7808 2979 7820
rect 1979 7802 2979 7808
rect 3215 7808 3227 7820
rect 4203 7820 4230 7842
rect 4203 7808 4215 7820
rect 3215 7802 4215 7808
rect -4288 7780 -4242 7792
rect -4288 7712 -4282 7780
rect -4248 7770 -4242 7780
rect -3160 7780 -3114 7792
rect -3052 7780 -3006 7792
rect -3160 7770 -3154 7780
rect -4248 7740 -3154 7770
rect -4248 7712 -3480 7740
rect -4288 7700 -3480 7712
rect -4280 7684 -3480 7700
rect -3400 7684 -3330 7740
rect -3250 7712 -3154 7740
rect -3012 7770 -3006 7780
rect -1924 7780 -1878 7792
rect -1816 7780 -1770 7792
rect -688 7780 -642 7792
rect -580 7780 -534 7792
rect -1924 7770 -1918 7780
rect -3012 7712 -1918 7770
rect -1776 7770 -1770 7780
rect -690 7770 -682 7780
rect -1776 7740 -682 7770
rect -1776 7712 -990 7740
rect -3250 7710 -3150 7712
rect -3020 7710 -1910 7712
rect -1780 7710 -990 7712
rect -3250 7684 -990 7710
rect -910 7684 -840 7740
rect -760 7712 -682 7740
rect -540 7770 -534 7780
rect 548 7780 594 7792
rect 656 7780 702 7792
rect 548 7770 554 7780
rect -540 7712 554 7770
rect 696 7770 702 7780
rect 1784 7780 1830 7792
rect 1892 7780 1938 7792
rect 3020 7780 3066 7792
rect 3128 7780 3174 7792
rect 1784 7770 1790 7780
rect 696 7740 1790 7770
rect 696 7712 1500 7740
rect -760 7710 -680 7712
rect -550 7710 560 7712
rect 690 7710 1500 7712
rect -760 7684 1500 7710
rect 1580 7684 1640 7740
rect 1720 7712 1790 7740
rect 1932 7770 1940 7780
rect 3020 7770 3026 7780
rect 1932 7712 3026 7770
rect 3168 7770 3174 7780
rect 4256 7780 4302 7792
rect 4256 7770 4262 7780
rect 3168 7712 4262 7770
rect 4296 7712 4302 7780
rect 1720 7710 1800 7712
rect 1930 7710 3030 7712
rect 3160 7710 4302 7712
rect 1720 7700 4302 7710
rect 1720 7684 4300 7700
rect -4280 7650 -4189 7684
rect -3213 7650 -2953 7684
rect -1977 7650 -1717 7684
rect -741 7650 -481 7684
rect 495 7650 755 7684
rect 1731 7650 1991 7684
rect 2967 7650 3227 7684
rect 4203 7650 4300 7684
rect -4280 7630 -3870 7650
rect -3880 7590 -3870 7630
rect -3790 7630 -3700 7650
rect -3790 7590 -3780 7630
rect -3710 7590 -3700 7630
rect -3620 7630 -1350 7650
rect -3620 7590 -3610 7630
rect -1360 7590 -1350 7630
rect -1270 7630 -1180 7650
rect -1270 7590 -1260 7630
rect -1190 7590 -1180 7630
rect -1100 7630 1140 7650
rect -1100 7590 -1090 7630
rect 1130 7580 1140 7630
rect 1220 7630 1310 7650
rect 1220 7580 1230 7630
rect 1300 7580 1310 7630
rect 1390 7630 3590 7650
rect 1390 7580 1400 7630
rect 3580 7590 3590 7630
rect 3670 7630 3760 7650
rect 3670 7590 3680 7630
rect 3750 7590 3760 7630
rect 3840 7630 4300 7650
rect 3840 7590 3850 7630
rect -2602 7520 -2498 7526
rect -2602 7440 -2590 7520
rect -2510 7440 -2498 7520
rect -2602 7434 -2498 7440
rect -2432 7520 -2328 7526
rect -2432 7440 -2420 7520
rect -2340 7440 -2328 7520
rect -2432 7434 -2328 7440
rect -122 7520 -18 7526
rect -122 7440 -110 7520
rect -30 7440 -18 7520
rect -122 7434 -18 7440
rect 48 7520 152 7526
rect 48 7440 60 7520
rect 140 7440 152 7520
rect 48 7434 152 7440
rect 2338 7520 2442 7526
rect 2338 7440 2350 7520
rect 2430 7440 2442 7520
rect 2338 7434 2442 7440
rect 2508 7520 2612 7526
rect 2508 7440 2520 7520
rect 2600 7440 2612 7520
rect 2508 7434 2612 7440
rect -2600 7330 -2590 7390
rect -4200 7310 -2590 7330
rect -2510 7330 -2500 7390
rect -2430 7330 -2420 7390
rect -2510 7310 -2420 7330
rect -2340 7330 -2330 7390
rect -120 7330 -110 7400
rect -2340 7320 -110 7330
rect -30 7330 -20 7400
rect 50 7330 60 7400
rect -30 7320 60 7330
rect 140 7330 150 7400
rect 2340 7330 2350 7390
rect 140 7320 2350 7330
rect -2340 7310 2350 7320
rect 2430 7330 2440 7390
rect 2510 7330 2520 7390
rect 2430 7310 2520 7330
rect 2600 7330 2610 7390
rect 2600 7310 4240 7330
rect -4200 7308 4240 7310
rect -4201 7302 4240 7308
rect -4201 7268 -4189 7302
rect -3213 7290 -2953 7302
rect -3213 7268 -3201 7290
rect -4201 7262 -3201 7268
rect -2965 7268 -2953 7290
rect -1977 7290 -1717 7302
rect -1977 7268 -1965 7290
rect -2965 7262 -1965 7268
rect -1729 7268 -1717 7290
rect -741 7290 -481 7302
rect -741 7268 -729 7290
rect -1729 7262 -729 7268
rect -493 7268 -481 7290
rect 495 7290 755 7302
rect 495 7268 507 7290
rect -493 7262 507 7268
rect 743 7268 755 7290
rect 1731 7290 1991 7302
rect 1731 7268 1743 7290
rect 743 7262 1743 7268
rect 1979 7268 1991 7290
rect 2967 7290 3227 7302
rect 2967 7268 2979 7290
rect 1979 7262 2979 7268
rect 3215 7268 3227 7290
rect 4203 7290 4240 7302
rect 4203 7268 4215 7290
rect 3215 7262 4215 7268
rect -4288 7240 -4242 7252
rect -4288 7172 -4282 7240
rect -4248 7230 -4242 7240
rect -3160 7240 -3114 7252
rect -3052 7240 -3006 7252
rect -3160 7230 -3154 7240
rect -4248 7180 -3154 7230
rect -4248 7172 -4242 7180
rect -4288 7160 -4242 7172
rect -3160 7172 -3154 7180
rect -3012 7230 -3006 7240
rect -1924 7240 -1878 7252
rect -1816 7240 -1770 7252
rect -688 7240 -642 7252
rect -580 7240 -534 7252
rect -1924 7230 -1918 7240
rect -3012 7180 -1918 7230
rect -3012 7172 -3006 7180
rect -3160 7170 -3150 7172
rect -3020 7170 -3006 7172
rect -3160 7160 -3114 7170
rect -3052 7160 -3006 7170
rect -1924 7172 -1918 7180
rect -1776 7230 -1770 7240
rect -690 7230 -682 7240
rect -1776 7180 -682 7230
rect -1776 7172 -1770 7180
rect -1924 7170 -1910 7172
rect -1780 7170 -1770 7172
rect -690 7172 -682 7180
rect -540 7230 -534 7240
rect 548 7240 594 7252
rect 656 7240 702 7252
rect 1784 7240 1830 7252
rect 1892 7240 1938 7252
rect 548 7230 554 7240
rect -540 7180 554 7230
rect -540 7172 -534 7180
rect -690 7170 -680 7172
rect -550 7170 -534 7172
rect -1924 7160 -1878 7170
rect -1816 7160 -1770 7170
rect -688 7160 -642 7170
rect -580 7160 -534 7170
rect 548 7172 554 7180
rect 696 7230 702 7240
rect 1780 7230 1790 7240
rect 696 7180 1790 7230
rect 696 7172 702 7180
rect 548 7170 560 7172
rect 690 7170 702 7172
rect 1780 7170 1790 7180
rect 1932 7230 1938 7240
rect 3020 7240 3066 7252
rect 3128 7240 3174 7252
rect 3020 7230 3026 7240
rect 1932 7180 3026 7230
rect 1932 7172 1938 7180
rect 1920 7170 1938 7172
rect 548 7160 594 7170
rect 656 7160 702 7170
rect 1784 7160 1830 7170
rect 1892 7160 1938 7170
rect 3020 7172 3026 7180
rect 3168 7230 3174 7240
rect 4256 7240 4302 7252
rect 4256 7230 4262 7240
rect 3168 7180 4262 7230
rect 3168 7172 3174 7180
rect 3020 7170 3030 7172
rect 3160 7170 3174 7172
rect 3020 7160 3066 7170
rect 3128 7160 3174 7170
rect 4256 7172 4262 7180
rect 4296 7172 4302 7240
rect 4256 7160 4302 7172
rect -4201 7144 -3201 7150
rect -4201 7130 -4189 7144
rect -3213 7130 -3201 7144
rect -2965 7144 -1965 7150
rect -2965 7130 -2953 7144
rect -4210 7110 -4189 7130
rect -3213 7110 -2953 7130
rect -1977 7130 -1965 7144
rect -1729 7144 -729 7150
rect -1729 7130 -1717 7144
rect -741 7130 -729 7144
rect -493 7144 507 7150
rect -493 7130 -481 7144
rect -1977 7110 -1717 7130
rect -741 7110 -481 7130
rect 495 7130 507 7144
rect 743 7144 1743 7150
rect 743 7130 755 7144
rect 1731 7130 1743 7144
rect 1979 7144 2979 7150
rect 1979 7130 1991 7144
rect 2967 7130 2979 7144
rect 3215 7144 4215 7150
rect 3215 7130 3227 7144
rect 4203 7130 4215 7144
rect 495 7110 755 7130
rect 1731 7110 1991 7130
rect 2967 7110 3227 7130
rect 4203 7110 4230 7130
rect -4210 7090 -3870 7110
rect -3880 7050 -3870 7090
rect -3790 7090 -3700 7110
rect -3790 7050 -3780 7090
rect -3710 7050 -3700 7090
rect -3620 7090 -2190 7110
rect -3620 7050 -3610 7090
rect -2210 7060 -2190 7090
rect -2110 7060 -2080 7110
rect -2000 7090 -1360 7110
rect -2000 7060 -1980 7090
rect -2210 7030 -1980 7060
rect -1370 7050 -1360 7090
rect -1280 7090 -1190 7110
rect -1280 7050 -1270 7090
rect -1200 7050 -1190 7090
rect -1110 7090 220 7110
rect -1110 7050 -1100 7090
rect 200 7060 220 7090
rect 300 7060 330 7110
rect 410 7090 1130 7110
rect 410 7060 430 7090
rect 200 7050 430 7060
rect 1120 7050 1130 7090
rect 1210 7090 1300 7110
rect 1210 7050 1220 7090
rect 1290 7050 1300 7090
rect 1380 7090 2680 7110
rect 1380 7050 1390 7090
rect 2660 7050 2680 7090
rect 2760 7050 2790 7110
rect 2870 7090 3620 7110
rect 2870 7050 2890 7090
rect 3610 7050 3620 7090
rect 3700 7090 3790 7110
rect 3700 7050 3710 7090
rect 3780 7050 3790 7090
rect 3870 7090 4230 7110
rect 3870 7050 3880 7090
rect 2660 7030 2890 7050
rect -2600 6750 -2590 6810
rect -4210 6730 -2590 6750
rect -2510 6750 -2500 6810
rect -2430 6750 -2420 6810
rect -2510 6730 -2420 6750
rect -2340 6750 -2330 6810
rect -120 6750 -110 6820
rect -2340 6740 -110 6750
rect -30 6750 -20 6820
rect 50 6750 60 6820
rect -30 6740 60 6750
rect 140 6750 150 6820
rect 2340 6750 2350 6810
rect 140 6740 2350 6750
rect -2340 6730 2350 6740
rect 2430 6750 2440 6810
rect 2510 6750 2520 6810
rect 2430 6730 2520 6750
rect 2600 6750 2610 6810
rect 2600 6730 4230 6750
rect -4210 6722 4230 6730
rect -4210 6710 -4189 6722
rect -4201 6688 -4189 6710
rect -3213 6710 -2953 6722
rect -3213 6688 -3201 6710
rect -4201 6682 -3201 6688
rect -2965 6688 -2953 6710
rect -1977 6710 -1717 6722
rect -1977 6688 -1965 6710
rect -2965 6682 -1965 6688
rect -1729 6688 -1717 6710
rect -741 6710 -481 6722
rect -741 6688 -729 6710
rect -1729 6682 -729 6688
rect -493 6688 -481 6710
rect 495 6710 755 6722
rect 495 6688 507 6710
rect -493 6682 507 6688
rect 743 6688 755 6710
rect 1731 6710 1991 6722
rect 1731 6688 1743 6710
rect 743 6682 1743 6688
rect 1979 6688 1991 6710
rect 2967 6710 3227 6722
rect 2967 6688 2979 6710
rect 1979 6682 2979 6688
rect 3215 6688 3227 6710
rect 4203 6710 4230 6722
rect 4203 6688 4215 6710
rect 3215 6682 4215 6688
rect -4288 6660 -4242 6672
rect -4288 6592 -4282 6660
rect -4248 6650 -4242 6660
rect -3160 6660 -3114 6672
rect -3052 6660 -3006 6672
rect -3160 6650 -3154 6660
rect -4248 6600 -3154 6650
rect -4248 6592 -4242 6600
rect -4288 6580 -4242 6592
rect -3160 6592 -3154 6600
rect -3012 6650 -3006 6660
rect -1924 6660 -1878 6672
rect -1816 6660 -1770 6672
rect -1924 6650 -1918 6660
rect -3012 6600 -1918 6650
rect -3012 6592 -3006 6600
rect -3160 6590 -3150 6592
rect -3020 6590 -3006 6592
rect -3160 6580 -3114 6590
rect -3052 6580 -3006 6590
rect -1924 6592 -1918 6600
rect -1776 6650 -1770 6660
rect -688 6660 -642 6672
rect -580 6660 -534 6672
rect 548 6660 594 6672
rect 656 6660 702 6672
rect 1784 6660 1830 6672
rect 1892 6660 1938 6672
rect -688 6650 -682 6660
rect -1776 6600 -682 6650
rect -1776 6592 -1770 6600
rect -1924 6590 -1910 6592
rect -1780 6590 -1770 6592
rect -1924 6580 -1878 6590
rect -1816 6580 -1770 6590
rect -688 6592 -682 6600
rect -540 6650 -530 6660
rect 548 6650 554 6660
rect -540 6600 554 6650
rect -688 6590 -670 6592
rect -540 6590 -530 6600
rect 548 6592 554 6600
rect 696 6650 702 6660
rect 1780 6650 1790 6660
rect 696 6600 1790 6650
rect 696 6592 702 6600
rect 548 6590 560 6592
rect 690 6590 702 6592
rect 1780 6590 1790 6600
rect 1932 6650 1938 6660
rect 3020 6660 3066 6672
rect 3128 6660 3174 6672
rect 3020 6650 3026 6660
rect 1932 6600 3026 6650
rect 1932 6592 1938 6600
rect 1920 6590 1938 6592
rect -688 6580 -642 6590
rect -580 6580 -534 6590
rect 548 6580 594 6590
rect 656 6580 702 6590
rect 1784 6580 1830 6590
rect 1892 6580 1938 6590
rect 3020 6592 3026 6600
rect 3168 6650 3174 6660
rect 4256 6660 4302 6672
rect 4256 6650 4262 6660
rect 3168 6600 4262 6650
rect 3168 6592 3174 6600
rect 3020 6590 3030 6592
rect 3160 6590 3174 6592
rect 3020 6580 3066 6590
rect 3128 6580 3174 6590
rect 4256 6592 4262 6600
rect 4296 6592 4302 6660
rect 4256 6580 4302 6592
rect -4201 6564 -3201 6570
rect -4201 6550 -4189 6564
rect -3213 6550 -3201 6564
rect -2965 6564 -1965 6570
rect -2965 6550 -2953 6564
rect -4210 6530 -4189 6550
rect -3213 6530 -2953 6550
rect -1977 6550 -1965 6564
rect -1729 6564 -729 6570
rect -1729 6550 -1717 6564
rect -741 6550 -729 6564
rect -493 6564 507 6570
rect -493 6550 -481 6564
rect 495 6550 507 6564
rect 743 6564 1743 6570
rect 743 6550 755 6564
rect -1977 6530 -1717 6550
rect -741 6530 -481 6550
rect 495 6530 755 6550
rect 1731 6550 1743 6564
rect 1979 6564 2979 6570
rect 1979 6550 1991 6564
rect 2967 6550 2979 6564
rect 3215 6564 4215 6570
rect 3215 6550 3227 6564
rect 4203 6550 4215 6564
rect 1731 6530 1991 6550
rect 2967 6530 3227 6550
rect 4203 6530 4230 6550
rect -4210 6510 -3870 6530
rect -3880 6470 -3870 6510
rect -3790 6510 -3700 6530
rect -3790 6470 -3780 6510
rect -3710 6470 -3700 6510
rect -3620 6510 -2190 6530
rect -3620 6470 -3610 6510
rect -2210 6450 -2190 6510
rect -2110 6450 -2080 6530
rect -2000 6510 -1360 6530
rect -2000 6450 -1980 6510
rect -1370 6470 -1360 6510
rect -1280 6510 -1190 6530
rect -1280 6470 -1270 6510
rect -1200 6470 -1190 6510
rect -1110 6510 220 6530
rect -1110 6470 -1100 6510
rect 200 6470 220 6510
rect 300 6470 330 6530
rect 410 6510 1130 6530
rect 410 6470 430 6510
rect 200 6450 430 6470
rect 1120 6460 1130 6510
rect 1210 6510 1300 6530
rect 1210 6460 1220 6510
rect 1290 6460 1300 6510
rect 1380 6510 2680 6530
rect 1380 6460 1390 6510
rect 2660 6470 2680 6510
rect 2760 6470 2790 6530
rect 2870 6510 3620 6530
rect 2870 6470 2890 6510
rect 3610 6470 3620 6510
rect 3700 6510 3790 6530
rect 3700 6470 3710 6510
rect 3780 6470 3790 6510
rect 3870 6510 4230 6530
rect 3870 6470 3880 6510
rect 2660 6450 2890 6470
rect -2210 6440 -1980 6450
rect 9540 6440 9970 6560
rect -9960 6270 -9530 6390
rect -2602 6360 -2488 6366
rect -2602 6280 -2590 6360
rect -2500 6280 -2488 6360
rect -2602 6274 -2488 6280
rect -2442 6360 -2328 6366
rect -2442 6280 -2430 6360
rect -2340 6280 -2328 6360
rect -2442 6274 -2328 6280
rect -122 6350 -18 6356
rect -122 6280 -110 6350
rect -30 6280 -18 6350
rect -122 6274 -18 6280
rect 48 6350 152 6356
rect 48 6280 60 6350
rect 140 6280 152 6350
rect 48 6274 152 6280
rect 2338 6350 2442 6356
rect 2338 6280 2350 6350
rect 2430 6280 2442 6350
rect 2338 6274 2442 6280
rect 2508 6350 2612 6356
rect 2508 6280 2520 6350
rect 2600 6280 2612 6350
rect 2508 6274 2612 6280
rect 9540 6300 9560 6440
rect 9690 6300 9820 6440
rect 9950 6300 9970 6440
rect -9960 6130 -9940 6270
rect -9810 6130 -9690 6270
rect -9560 6130 -9530 6270
rect -2600 6170 -2590 6230
rect -4210 6150 -2590 6170
rect -2510 6170 -2500 6230
rect -2430 6170 -2420 6230
rect -2510 6150 -2420 6170
rect -2340 6170 -2330 6230
rect -120 6170 -110 6240
rect -2340 6160 -110 6170
rect -30 6170 -20 6240
rect 50 6170 60 6240
rect -30 6160 60 6170
rect 140 6170 150 6240
rect 2340 6170 2350 6230
rect 140 6160 2350 6170
rect -2340 6150 2350 6160
rect 2430 6170 2440 6230
rect 2510 6170 2520 6230
rect 2430 6150 2520 6170
rect 2600 6170 2610 6230
rect 2600 6150 4230 6170
rect -4210 6142 4230 6150
rect -4210 6130 -4189 6142
rect -9960 6105 -9530 6130
rect -4201 6108 -4189 6130
rect -3213 6130 -2953 6142
rect -3213 6108 -3201 6130
rect -9960 6093 -9426 6105
rect -9960 4979 -9829 6093
rect -9432 4979 -9426 6093
rect -7404 6093 -6995 6105
rect -4201 6102 -3201 6108
rect -2965 6108 -2953 6130
rect -1977 6130 -1717 6142
rect -1977 6108 -1965 6130
rect -2965 6102 -1965 6108
rect -1729 6108 -1717 6130
rect -741 6130 -481 6142
rect -741 6108 -729 6130
rect -1729 6102 -729 6108
rect -493 6108 -481 6130
rect 495 6130 755 6142
rect 495 6108 507 6130
rect -493 6102 507 6108
rect 743 6108 755 6130
rect 1731 6130 1991 6142
rect 1731 6108 1743 6130
rect 743 6102 1743 6108
rect 1979 6108 1991 6130
rect 2967 6130 3227 6142
rect 2967 6108 2979 6130
rect 1979 6102 2979 6108
rect 3215 6108 3227 6130
rect 4203 6130 4230 6142
rect 4203 6108 4215 6130
rect 3215 6102 4215 6108
rect 9540 6105 9970 6300
rect -7404 6000 -7398 6093
rect -9960 4967 -9426 4979
rect -7530 4979 -7398 6000
rect -7001 5560 -6995 6093
rect 7225 6093 7634 6105
rect -4288 6080 -4242 6092
rect -4288 6012 -4282 6080
rect -4248 6070 -4242 6080
rect -3160 6080 -3114 6092
rect -3052 6080 -3006 6092
rect -3160 6070 -3154 6080
rect -4248 6020 -3154 6070
rect -4248 6012 -4242 6020
rect -4288 6000 -4242 6012
rect -3160 6012 -3154 6020
rect -3012 6070 -3006 6080
rect -1924 6080 -1878 6092
rect -1816 6080 -1770 6092
rect -688 6080 -642 6092
rect -580 6080 -534 6092
rect -1924 6070 -1918 6080
rect -3012 6020 -1918 6070
rect -3012 6012 -3006 6020
rect -3160 6010 -3150 6012
rect -3020 6010 -3006 6012
rect -3160 6000 -3114 6010
rect -3052 6000 -3006 6010
rect -1924 6012 -1918 6020
rect -1884 6012 -1810 6080
rect -1776 6070 -1770 6080
rect -690 6070 -682 6080
rect -1776 6020 -682 6070
rect -1776 6012 -1770 6020
rect -1924 6010 -1770 6012
rect -690 6012 -682 6020
rect -540 6070 -534 6080
rect 548 6080 594 6092
rect 656 6080 702 6092
rect 1784 6080 1830 6092
rect 1892 6080 1938 6092
rect 548 6070 554 6080
rect -540 6020 554 6070
rect -540 6012 -534 6020
rect -690 6010 -680 6012
rect -550 6010 -534 6012
rect -1924 6000 -1878 6010
rect -1816 6000 -1770 6010
rect -688 6000 -642 6010
rect -580 6000 -534 6010
rect 548 6012 554 6020
rect 696 6070 702 6080
rect 1780 6070 1790 6080
rect 696 6020 1790 6070
rect 696 6012 702 6020
rect 548 6010 560 6012
rect 690 6010 702 6012
rect 1780 6010 1790 6020
rect 1932 6070 1938 6080
rect 3020 6080 3066 6092
rect 3128 6080 3174 6092
rect 3020 6070 3026 6080
rect 1932 6020 3026 6070
rect 1932 6012 1938 6020
rect 1920 6010 1938 6012
rect 548 6000 594 6010
rect 656 6000 702 6010
rect 1784 6000 1830 6010
rect 1892 6000 1938 6010
rect 3020 6012 3026 6020
rect 3168 6070 3174 6080
rect 4256 6080 4302 6092
rect 4256 6070 4262 6080
rect 3168 6020 4262 6070
rect 3168 6012 3174 6020
rect 3020 6010 3030 6012
rect 3160 6010 3174 6012
rect 3020 6000 3066 6010
rect 3128 6000 3174 6010
rect 4256 6012 4262 6020
rect 4296 6012 4302 6080
rect 4256 6000 4302 6012
rect 7225 6000 7231 6093
rect -4201 5984 -3201 5990
rect -4201 5960 -4189 5984
rect -4210 5950 -4189 5960
rect -3213 5960 -3201 5984
rect -2965 5984 -1965 5990
rect -2965 5960 -2953 5984
rect -3213 5950 -2953 5960
rect -1977 5960 -1965 5984
rect -1729 5984 -729 5990
rect -1729 5960 -1717 5984
rect -1977 5950 -1717 5960
rect -741 5960 -729 5984
rect -493 5984 507 5990
rect -493 5960 -481 5984
rect -741 5950 -481 5960
rect 495 5960 507 5984
rect 743 5984 1743 5990
rect 743 5960 755 5984
rect 495 5950 755 5960
rect 1731 5960 1743 5984
rect 1979 5984 2979 5990
rect 1979 5960 1991 5984
rect 1731 5950 1991 5960
rect 2967 5960 2979 5984
rect 3215 5984 4215 5990
rect 3215 5960 3227 5984
rect 2967 5950 3227 5960
rect 4203 5960 4215 5984
rect 4203 5950 4230 5960
rect -4210 5940 -1360 5950
rect -4210 5920 -3890 5940
rect -3900 5860 -3890 5920
rect -3810 5920 -3680 5940
rect -3810 5860 -3800 5920
rect -3690 5860 -3680 5920
rect -3600 5920 -1360 5940
rect -3600 5860 -3590 5920
rect -2210 5870 -1980 5920
rect -1370 5890 -1360 5920
rect -1280 5920 -1190 5950
rect -1280 5890 -1270 5920
rect -1200 5890 -1190 5920
rect -1110 5920 220 5950
rect -1110 5890 -1100 5920
rect 200 5890 220 5920
rect 300 5890 330 5950
rect 410 5920 1130 5950
rect 410 5890 430 5920
rect 1120 5890 1130 5920
rect 1210 5920 1300 5950
rect 1210 5890 1220 5920
rect 1290 5890 1300 5920
rect 1380 5920 2680 5950
rect 1380 5890 1390 5920
rect 2660 5890 2680 5920
rect 2760 5890 2790 5950
rect 2870 5920 3620 5950
rect 2870 5890 2890 5920
rect 3610 5890 3620 5920
rect 3700 5920 3790 5950
rect 3700 5890 3710 5920
rect 3780 5890 3790 5920
rect 3870 5920 4230 5950
rect 3870 5890 3880 5920
rect 200 5870 430 5890
rect 2660 5870 2890 5890
rect -4480 5630 -4470 5700
rect -6050 5620 -4470 5630
rect -4390 5630 -4380 5700
rect -4250 5630 -4240 5700
rect -4390 5620 -4240 5630
rect -4160 5630 -4150 5700
rect -1930 5630 -1920 5690
rect -4160 5620 -1920 5630
rect -6050 5610 -1920 5620
rect -1840 5630 -1830 5690
rect -1760 5630 -1750 5690
rect -1840 5610 -1750 5630
rect -1670 5630 -1660 5690
rect 530 5630 540 5690
rect -1670 5610 540 5630
rect 620 5630 630 5690
rect 720 5630 730 5690
rect 620 5610 730 5630
rect 810 5630 820 5690
rect 2980 5630 2990 5690
rect 810 5610 2990 5630
rect 3070 5630 3080 5690
rect 3170 5630 3180 5690
rect 3070 5610 3180 5630
rect 3260 5630 3270 5690
rect 5490 5630 5500 5690
rect 3260 5610 5500 5630
rect 5580 5630 5590 5690
rect 5660 5630 5670 5690
rect 5580 5610 5670 5630
rect 5750 5630 5760 5690
rect 5750 5610 6100 5630
rect -6050 5602 6100 5610
rect -6050 5580 -6029 5602
rect -6041 5568 -6029 5580
rect -5053 5580 -4793 5602
rect -5053 5568 -5041 5580
rect -6041 5562 -5041 5568
rect -4805 5568 -4793 5580
rect -3817 5580 -3557 5602
rect -3817 5568 -3805 5580
rect -4805 5562 -3805 5568
rect -3569 5568 -3557 5580
rect -2581 5580 -2321 5602
rect -2581 5568 -2569 5580
rect -3569 5562 -2569 5568
rect -2333 5568 -2321 5580
rect -1345 5580 -1085 5602
rect -1345 5568 -1333 5580
rect -2333 5562 -1333 5568
rect -1097 5568 -1085 5580
rect -109 5580 151 5602
rect -109 5568 -97 5580
rect -1097 5562 -97 5568
rect 139 5568 151 5580
rect 1127 5580 1387 5602
rect 1127 5568 1139 5580
rect 139 5562 1139 5568
rect 1375 5568 1387 5580
rect 2363 5580 2623 5602
rect 2363 5568 2375 5580
rect 1375 5562 2375 5568
rect 2611 5568 2623 5580
rect 3599 5580 3859 5602
rect 3599 5568 3611 5580
rect 2611 5562 3611 5568
rect 3847 5568 3859 5580
rect 4835 5580 5095 5602
rect 4835 5568 4847 5580
rect 3847 5562 4847 5568
rect 5083 5568 5095 5580
rect 6071 5580 6100 5602
rect 6071 5568 6083 5580
rect 5083 5562 6083 5568
rect 7100 5560 7231 6000
rect -7001 5552 -6090 5560
rect 6130 5552 7231 5560
rect -7001 5540 -6082 5552
rect -7001 5472 -6122 5540
rect -6088 5530 -6082 5540
rect -5000 5540 -4954 5552
rect -4892 5540 -4846 5552
rect -5000 5530 -4994 5540
rect -6088 5490 -4994 5530
rect -6088 5472 -6082 5490
rect -7001 5460 -6082 5472
rect -5000 5472 -4994 5490
rect -4852 5530 -4846 5540
rect -3764 5540 -3718 5552
rect -3656 5540 -3610 5552
rect -2528 5540 -2482 5552
rect -2420 5540 -2374 5552
rect -3764 5530 -3758 5540
rect -4852 5490 -3758 5530
rect -4852 5472 -4846 5490
rect -5000 5470 -4990 5472
rect -4860 5470 -4846 5472
rect -5000 5460 -4954 5470
rect -4892 5460 -4846 5470
rect -3764 5472 -3758 5490
rect -3616 5530 -3610 5540
rect -2530 5530 -2522 5540
rect -3616 5490 -2522 5530
rect -3616 5472 -3610 5490
rect -3764 5470 -3750 5472
rect -3620 5470 -3610 5472
rect -2530 5472 -2522 5490
rect -2380 5530 -2374 5540
rect -1292 5540 -1246 5552
rect -1184 5540 -1138 5552
rect -1292 5530 -1286 5540
rect -2380 5490 -1286 5530
rect -2380 5472 -2374 5490
rect -2530 5470 -2520 5472
rect -2390 5470 -2374 5472
rect -3764 5460 -3718 5470
rect -3656 5460 -3610 5470
rect -2528 5460 -2482 5470
rect -2420 5460 -2374 5470
rect -1292 5472 -1286 5490
rect -1144 5530 -1138 5540
rect -56 5540 -10 5552
rect 52 5540 98 5552
rect 1180 5540 1226 5552
rect 1288 5540 1334 5552
rect -56 5530 -50 5540
rect -1144 5490 -50 5530
rect -1144 5472 -1138 5490
rect -1292 5470 -1280 5472
rect -1150 5470 -1138 5472
rect -1292 5460 -1246 5470
rect -1184 5460 -1138 5470
rect -56 5472 -50 5490
rect 92 5530 100 5540
rect 1180 5530 1186 5540
rect 92 5490 1186 5530
rect 92 5472 100 5490
rect -56 5470 -40 5472
rect 90 5470 100 5472
rect 1180 5472 1186 5490
rect 1328 5530 1334 5540
rect 2416 5540 2462 5552
rect 2524 5540 2570 5552
rect 3652 5540 3698 5552
rect 3760 5540 3806 5552
rect 2416 5530 2422 5540
rect 1328 5490 2422 5530
rect 1328 5472 1334 5490
rect 1180 5470 1190 5472
rect 1320 5470 1334 5472
rect -56 5460 -10 5470
rect 52 5460 98 5470
rect 1180 5460 1226 5470
rect 1288 5460 1334 5470
rect 2416 5472 2422 5490
rect 2564 5530 2570 5540
rect 3650 5530 3658 5540
rect 2564 5490 3658 5530
rect 2564 5472 2570 5490
rect 2416 5470 2430 5472
rect 2560 5470 2570 5472
rect 3650 5472 3658 5490
rect 3800 5530 3806 5540
rect 4888 5540 4934 5552
rect 4996 5540 5042 5552
rect 4888 5530 4894 5540
rect 3800 5490 4894 5530
rect 3800 5472 3806 5490
rect 3650 5470 3660 5472
rect 3790 5470 3806 5472
rect 2416 5460 2462 5470
rect 2524 5460 2570 5470
rect 3652 5460 3698 5470
rect 3760 5460 3806 5470
rect 4888 5472 4894 5490
rect 5036 5530 5042 5540
rect 6124 5540 7231 5552
rect 6124 5530 6130 5540
rect 5036 5490 6130 5530
rect 5036 5472 5042 5490
rect 4888 5470 4900 5472
rect 5030 5470 5042 5472
rect 4888 5460 4934 5470
rect 4996 5460 5042 5470
rect 6124 5472 6130 5490
rect 6164 5472 7231 5540
rect 6124 5460 7231 5472
rect -7001 5020 -6995 5460
rect -6041 5444 -5041 5450
rect -6041 5430 -6029 5444
rect -6050 5410 -6029 5430
rect -5053 5430 -5041 5444
rect -4805 5444 -3805 5450
rect -4805 5430 -4793 5444
rect -5053 5410 -4793 5430
rect -3817 5430 -3805 5444
rect -3569 5444 -2569 5450
rect -3569 5430 -3557 5444
rect -3817 5410 -3557 5430
rect -2581 5430 -2569 5444
rect -2333 5444 -1333 5450
rect -2333 5430 -2321 5444
rect -2581 5410 -2321 5430
rect -1345 5430 -1333 5444
rect -1097 5444 -97 5450
rect -1097 5430 -1085 5444
rect -1345 5410 -1085 5430
rect -109 5430 -97 5444
rect 139 5444 1139 5450
rect 139 5430 151 5444
rect -109 5410 151 5430
rect 1127 5430 1139 5444
rect 1375 5444 2375 5450
rect 1375 5430 1387 5444
rect 1127 5410 1387 5430
rect 2363 5430 2375 5444
rect 2611 5444 3611 5450
rect 2611 5430 2623 5444
rect 2363 5410 2623 5430
rect 3599 5430 3611 5444
rect 3847 5444 4847 5450
rect 3847 5430 3859 5444
rect 3599 5410 3859 5430
rect 4835 5430 4847 5444
rect 5083 5444 6083 5450
rect 5083 5430 5095 5444
rect 4835 5410 5095 5430
rect 6071 5430 6083 5444
rect 6071 5410 6100 5430
rect -6050 5380 -5720 5410
rect -5730 5340 -5720 5380
rect -5640 5380 -5510 5410
rect -5640 5340 -5630 5380
rect -5520 5340 -5510 5380
rect -5430 5380 -3240 5410
rect -5430 5340 -5420 5380
rect -3250 5340 -3240 5380
rect -3160 5380 -3020 5410
rect -3160 5340 -3150 5380
rect -3030 5340 -3020 5380
rect -2940 5380 -710 5410
rect -2940 5340 -2930 5380
rect -720 5340 -710 5380
rect -630 5380 -530 5410
rect -630 5340 -620 5380
rect -540 5340 -530 5380
rect -450 5380 1750 5410
rect -450 5340 -440 5380
rect 1740 5330 1750 5380
rect 1830 5380 1930 5410
rect 1830 5330 1840 5380
rect 1920 5330 1930 5380
rect 2010 5380 4230 5410
rect 2010 5330 2020 5380
rect 4220 5330 4230 5380
rect 4310 5380 4400 5410
rect 4310 5330 4320 5380
rect 4390 5330 4400 5380
rect 4480 5380 6100 5410
rect 4480 5330 4490 5380
rect -4462 5280 -4348 5286
rect -4462 5200 -4450 5280
rect -4360 5200 -4348 5280
rect -4462 5194 -4348 5200
rect -4282 5280 -4168 5286
rect -4282 5200 -4270 5280
rect -4180 5200 -4168 5280
rect -4282 5194 -4168 5200
rect -1932 5280 -1818 5286
rect -1932 5200 -1920 5280
rect -1830 5200 -1818 5280
rect -1932 5194 -1818 5200
rect -1772 5280 -1658 5286
rect -1772 5200 -1760 5280
rect -1670 5200 -1658 5280
rect -1772 5194 -1658 5200
rect 538 5280 652 5286
rect 538 5200 550 5280
rect 640 5200 652 5280
rect 538 5194 652 5200
rect 698 5280 812 5286
rect 698 5200 710 5280
rect 800 5200 812 5280
rect 698 5194 812 5200
rect 2988 5280 3102 5286
rect 2988 5200 3000 5280
rect 3090 5200 3102 5280
rect 2988 5194 3102 5200
rect 3148 5280 3262 5286
rect 3148 5200 3160 5280
rect 3250 5200 3262 5280
rect 3148 5194 3262 5200
rect 5488 5280 5602 5286
rect 5488 5200 5500 5280
rect 5590 5200 5602 5280
rect 5488 5194 5602 5200
rect 5648 5280 5762 5286
rect 5648 5200 5660 5280
rect 5750 5200 5762 5280
rect 5648 5194 5762 5200
rect -4480 5100 -4470 5160
rect -6050 5080 -4470 5100
rect -4390 5100 -4380 5160
rect -4250 5100 -4240 5160
rect -4390 5080 -4240 5100
rect -4160 5100 -4150 5160
rect -1930 5100 -1920 5150
rect -4160 5080 -1920 5100
rect -6050 5070 -1920 5080
rect -1840 5100 -1830 5150
rect -1760 5100 -1750 5160
rect -1840 5080 -1750 5100
rect -1670 5100 -1660 5160
rect 530 5100 540 5160
rect -1670 5080 540 5100
rect 620 5100 630 5160
rect 720 5100 730 5160
rect 620 5080 730 5100
rect 810 5100 820 5160
rect 2980 5100 2990 5150
rect 810 5080 2990 5100
rect -1840 5070 2990 5080
rect 3070 5100 3080 5150
rect 3170 5100 3180 5150
rect 3070 5070 3180 5100
rect 3260 5100 3270 5150
rect 5490 5100 5500 5150
rect 3260 5070 5500 5100
rect 5580 5100 5590 5150
rect 5660 5100 5670 5150
rect 5580 5070 5670 5100
rect 5750 5100 5760 5150
rect 5750 5070 6100 5100
rect -6050 5062 6100 5070
rect -6050 5050 -6029 5062
rect -6041 5028 -6029 5050
rect -5053 5050 -4793 5062
rect -5053 5028 -5041 5050
rect -6041 5022 -5041 5028
rect -4805 5028 -4793 5050
rect -3817 5050 -3557 5062
rect -3817 5028 -3805 5050
rect -4805 5022 -3805 5028
rect -3569 5028 -3557 5050
rect -2581 5050 -2321 5062
rect -2581 5028 -2569 5050
rect -3569 5022 -2569 5028
rect -2333 5028 -2321 5050
rect -1345 5050 -1085 5062
rect -1345 5028 -1333 5050
rect -2333 5022 -1333 5028
rect -1097 5028 -1085 5050
rect -109 5050 151 5062
rect -109 5028 -97 5050
rect -1097 5022 -97 5028
rect 139 5028 151 5050
rect 1127 5050 1387 5062
rect 1127 5028 1139 5050
rect 139 5022 1139 5028
rect 1375 5028 1387 5050
rect 2363 5050 2623 5062
rect 2363 5028 2375 5050
rect 1375 5022 2375 5028
rect 2611 5028 2623 5050
rect 3599 5050 3859 5062
rect 3599 5028 3611 5050
rect 2611 5022 3611 5028
rect 3847 5028 3859 5050
rect 4835 5050 5095 5062
rect 4835 5028 4847 5050
rect 3847 5022 4847 5028
rect 5083 5028 5095 5050
rect 6071 5050 6100 5062
rect 6071 5028 6083 5050
rect 5083 5022 6083 5028
rect -7001 5012 -6090 5020
rect -7001 5000 -6082 5012
rect -7001 4979 -6122 5000
rect -9960 4635 -9530 4967
rect -7530 4932 -6122 4979
rect -6088 4990 -6082 5000
rect -5000 5010 -4954 5012
rect -4892 5010 -4846 5012
rect -5000 5000 -4990 5010
rect -4860 5000 -4846 5010
rect -5000 4990 -4994 5000
rect -6088 4950 -4994 4990
rect -6088 4932 -6082 4950
rect -7530 4920 -6082 4932
rect -5000 4932 -4994 4950
rect -4852 4990 -4846 5000
rect -3764 5000 -3718 5012
rect -3656 5000 -3610 5012
rect -2528 5000 -2482 5012
rect -2420 5000 -2374 5012
rect -3764 4990 -3758 5000
rect -4852 4950 -3758 4990
rect -4960 4932 -4954 4940
rect -5000 4920 -4954 4932
rect -4892 4932 -4886 4940
rect -4852 4932 -4846 4950
rect -4892 4920 -4846 4932
rect -3764 4932 -3758 4950
rect -3616 4990 -3610 5000
rect -2530 4990 -2522 5000
rect -3616 4950 -2522 4990
rect -3616 4932 -3610 4950
rect -3764 4930 -3750 4932
rect -3620 4930 -3610 4932
rect -2530 4932 -2522 4950
rect -2380 4990 -2374 5000
rect -1292 5000 -1246 5012
rect -1184 5000 -1138 5012
rect -1292 4990 -1286 5000
rect -2380 4950 -1286 4990
rect -2380 4932 -2374 4950
rect -2530 4930 -2520 4932
rect -2390 4930 -2374 4932
rect -3764 4920 -3718 4930
rect -3656 4920 -3610 4930
rect -2528 4920 -2482 4930
rect -2420 4920 -2374 4930
rect -1292 4932 -1286 4950
rect -1144 4990 -1138 5000
rect -56 5000 -10 5012
rect 52 5000 98 5012
rect 1180 5000 1226 5012
rect 1288 5000 1334 5012
rect -56 4990 -50 5000
rect -1144 4950 -50 4990
rect -1144 4932 -1138 4950
rect -1292 4930 -1280 4932
rect -1150 4930 -1138 4932
rect -1292 4920 -1246 4930
rect -1184 4920 -1138 4930
rect -56 4932 -50 4950
rect 92 4990 100 5000
rect 1180 4990 1186 5000
rect 92 4950 1186 4990
rect 92 4932 100 4950
rect -56 4930 -40 4932
rect 90 4930 100 4932
rect 1180 4932 1186 4950
rect 1328 4990 1334 5000
rect 2416 5000 2462 5012
rect 2524 5000 2570 5012
rect 3652 5000 3698 5012
rect 3760 5000 3806 5012
rect 2416 4990 2422 5000
rect 1328 4950 2422 4990
rect 1328 4932 1334 4950
rect 1180 4930 1190 4932
rect 1320 4930 1334 4932
rect -56 4920 -10 4930
rect 52 4920 98 4930
rect 1180 4920 1226 4930
rect 1288 4920 1334 4930
rect 2416 4932 2422 4950
rect 2564 4990 2570 5000
rect 3650 4990 3658 5000
rect 2564 4950 3658 4990
rect 2564 4932 2570 4950
rect 2416 4930 2430 4932
rect 2560 4930 2570 4932
rect 3650 4932 3658 4950
rect 3800 4990 3806 5000
rect 4888 5000 4934 5012
rect 4996 5000 5042 5012
rect 4888 4990 4894 5000
rect 3800 4950 4894 4990
rect 3800 4932 3806 4950
rect 3650 4930 3660 4932
rect 3790 4930 3806 4932
rect 2416 4920 2462 4930
rect 2524 4920 2570 4930
rect 3652 4920 3698 4930
rect 3760 4920 3806 4930
rect 4888 4932 4894 4950
rect 5036 4990 5042 5000
rect 6124 5010 6170 5012
rect 7100 5010 7231 5460
rect 6124 5000 7231 5010
rect 6124 4990 6130 5000
rect 5036 4950 6130 4990
rect 5036 4932 5042 4950
rect 4888 4930 4900 4932
rect 5030 4930 5042 4932
rect 4888 4920 4934 4930
rect 4996 4920 5042 4930
rect 6124 4932 6130 4950
rect 6164 4979 7231 5000
rect 7628 4979 7634 6093
rect 6164 4967 7634 4979
rect 9540 6093 10065 6105
rect 9540 4979 9662 6093
rect 10059 4979 10065 6093
rect 9540 4967 10065 4979
rect 6164 4932 7530 4967
rect 6124 4920 7530 4932
rect -7530 4910 -6090 4920
rect 6130 4910 7530 4920
rect -7530 4635 -7100 4910
rect -6041 4904 -5041 4910
rect -6041 4890 -6029 4904
rect -6050 4870 -6029 4890
rect -5053 4890 -5041 4904
rect -4805 4904 -3805 4910
rect -4805 4890 -4793 4904
rect -5053 4870 -4793 4890
rect -3817 4890 -3805 4904
rect -3569 4904 -2569 4910
rect -3569 4890 -3557 4904
rect -3817 4870 -3557 4890
rect -2581 4890 -2569 4904
rect -2333 4904 -1333 4910
rect -2333 4890 -2321 4904
rect -2581 4870 -2321 4890
rect -1345 4890 -1333 4904
rect -1097 4904 -97 4910
rect -1097 4890 -1085 4904
rect -1345 4870 -1085 4890
rect -109 4890 -97 4904
rect 139 4904 1139 4910
rect 139 4890 151 4904
rect -109 4870 151 4890
rect 1127 4890 1139 4904
rect 1375 4904 2375 4910
rect 1375 4890 1387 4904
rect 1127 4870 1387 4890
rect 2363 4890 2375 4904
rect 2611 4904 3611 4910
rect 2611 4890 2623 4904
rect 2363 4870 2623 4890
rect 3599 4890 3611 4904
rect 3847 4904 4847 4910
rect 3847 4890 3859 4904
rect 3599 4870 3859 4890
rect 4835 4890 4847 4904
rect 5083 4904 6083 4910
rect 5083 4890 5095 4904
rect 4835 4870 5095 4890
rect 6071 4890 6083 4904
rect 6071 4870 6100 4890
rect -6050 4840 -5720 4870
rect -5730 4800 -5720 4840
rect -5640 4840 -5510 4870
rect -5640 4800 -5630 4840
rect -5520 4800 -5510 4840
rect -5430 4840 -3240 4870
rect -5430 4800 -5420 4840
rect -3250 4800 -3240 4840
rect -3160 4840 -3020 4870
rect -3160 4800 -3150 4840
rect -3030 4800 -3020 4840
rect -2940 4840 -710 4870
rect -2940 4800 -2930 4840
rect -720 4800 -710 4840
rect -630 4840 -520 4870
rect -630 4800 -620 4840
rect -530 4800 -520 4840
rect -440 4840 1750 4870
rect -440 4800 -430 4840
rect 1740 4790 1750 4840
rect 1830 4840 1930 4870
rect 1830 4790 1840 4840
rect 1920 4790 1930 4840
rect 2010 4840 4230 4870
rect 2010 4790 2020 4840
rect 4220 4790 4230 4840
rect 4310 4840 4400 4870
rect 4310 4790 4320 4840
rect 4390 4790 4400 4840
rect 4480 4840 6100 4870
rect 4480 4790 4490 4840
rect 7100 4635 7530 4910
rect 9540 4635 9970 4967
rect -9960 4623 -9426 4635
rect -9960 3530 -9829 4623
rect -9835 3509 -9829 3530
rect -9432 3509 -9426 4623
rect -7530 4623 -6995 4635
rect -7530 3520 -7398 4623
rect -9835 3497 -9426 3509
rect -7404 3509 -7398 3520
rect -7001 4480 -6995 4623
rect 7100 4623 7634 4635
rect -4480 4560 -4470 4620
rect -6050 4540 -4470 4560
rect -4390 4560 -4380 4620
rect -4250 4560 -4240 4620
rect -4390 4540 -4240 4560
rect -4160 4560 -4150 4620
rect -1940 4560 -1930 4610
rect -4160 4540 -1930 4560
rect -6050 4530 -1930 4540
rect -1850 4560 -1840 4610
rect -1770 4560 -1760 4610
rect -1850 4530 -1760 4560
rect -1680 4560 -1670 4610
rect 530 4560 540 4610
rect -1680 4530 540 4560
rect 620 4560 630 4610
rect 710 4560 720 4610
rect 620 4530 720 4560
rect 800 4560 810 4610
rect 2980 4560 2990 4610
rect 800 4530 2990 4560
rect 3070 4560 3080 4610
rect 3170 4560 3180 4610
rect 3070 4530 3180 4560
rect 3260 4560 3270 4610
rect 5490 4560 5500 4610
rect 3260 4530 5500 4560
rect 5580 4560 5590 4610
rect 5660 4560 5670 4610
rect 5580 4530 5670 4560
rect 5750 4560 5760 4610
rect 5750 4530 6100 4560
rect -6050 4522 6100 4530
rect -6050 4510 -6029 4522
rect -6041 4488 -6029 4510
rect -5053 4510 -4793 4522
rect -5053 4488 -5041 4510
rect -6041 4482 -5041 4488
rect -4805 4488 -4793 4510
rect -3817 4510 -3557 4522
rect -3817 4488 -3805 4510
rect -4805 4482 -3805 4488
rect -3569 4488 -3557 4510
rect -2581 4510 -2321 4522
rect -2581 4488 -2569 4510
rect -3569 4482 -2569 4488
rect -2333 4488 -2321 4510
rect -1345 4510 -1085 4522
rect -1345 4488 -1333 4510
rect -2333 4482 -1333 4488
rect -1097 4488 -1085 4510
rect -109 4510 151 4522
rect -109 4488 -97 4510
rect -1097 4482 -97 4488
rect 139 4488 151 4510
rect 1127 4510 1387 4522
rect 1127 4488 1139 4510
rect 139 4482 1139 4488
rect 1375 4488 1387 4510
rect 2363 4510 2623 4522
rect 2363 4488 2375 4510
rect 1375 4482 2375 4488
rect 2611 4488 2623 4510
rect 3599 4510 3859 4522
rect 3599 4488 3611 4510
rect 2611 4482 3611 4488
rect 3847 4488 3859 4510
rect 4835 4510 5095 4522
rect 4835 4488 4847 4510
rect 3847 4482 4847 4488
rect 5083 4488 5095 4510
rect 6071 4510 6100 4522
rect 6071 4488 6083 4510
rect 5083 4482 6083 4488
rect 7100 4480 7231 4623
rect -7001 4460 -6070 4480
rect 6130 4472 7231 4480
rect -7001 4392 -6122 4460
rect -6088 4450 -6070 4460
rect -5000 4460 -4954 4472
rect -4892 4460 -4846 4472
rect -5000 4450 -4994 4460
rect -6088 4410 -4994 4450
rect -6088 4392 -6070 4410
rect -7001 4370 -6070 4392
rect -5000 4392 -4994 4410
rect -4852 4450 -4846 4460
rect -3764 4460 -3718 4472
rect -3656 4460 -3610 4472
rect -2528 4460 -2482 4472
rect -2420 4460 -2374 4472
rect -3764 4450 -3758 4460
rect -4852 4410 -3758 4450
rect -4852 4392 -4846 4410
rect -5000 4390 -4990 4392
rect -4860 4390 -4846 4392
rect -5000 4380 -4954 4390
rect -4892 4380 -4846 4390
rect -3764 4392 -3758 4410
rect -3616 4450 -3610 4460
rect -2530 4450 -2522 4460
rect -3616 4410 -2522 4450
rect -3616 4392 -3610 4410
rect -3764 4390 -3750 4392
rect -3620 4390 -3610 4392
rect -2530 4392 -2522 4410
rect -2380 4450 -2374 4460
rect -1292 4460 -1246 4472
rect -1184 4460 -1138 4472
rect -1292 4450 -1286 4460
rect -2380 4410 -1286 4450
rect -2380 4392 -2374 4410
rect -2530 4390 -2520 4392
rect -2390 4390 -2374 4392
rect -3764 4380 -3718 4390
rect -3656 4380 -3610 4390
rect -2528 4380 -2482 4390
rect -2420 4380 -2374 4390
rect -1292 4392 -1286 4410
rect -1144 4450 -1138 4460
rect -56 4460 -10 4472
rect 52 4460 98 4472
rect 1180 4460 1226 4472
rect 1288 4460 1334 4472
rect -56 4450 -50 4460
rect -1144 4410 -50 4450
rect -1144 4392 -1138 4410
rect -1292 4390 -1280 4392
rect -1150 4390 -1138 4392
rect -1292 4380 -1246 4390
rect -1184 4380 -1138 4390
rect -56 4392 -50 4410
rect 92 4450 100 4460
rect 1180 4450 1186 4460
rect 92 4410 1186 4450
rect 92 4392 100 4410
rect -56 4390 -40 4392
rect 90 4390 100 4392
rect 1180 4392 1186 4410
rect 1328 4450 1334 4460
rect 2416 4460 2462 4472
rect 2524 4460 2570 4472
rect 3652 4460 3698 4472
rect 3760 4460 3806 4472
rect 2416 4450 2422 4460
rect 1328 4410 2422 4450
rect 1328 4392 1334 4410
rect 1180 4390 1190 4392
rect 1320 4390 1334 4392
rect -56 4380 -10 4390
rect 52 4380 98 4390
rect 1180 4380 1226 4390
rect 1288 4380 1334 4390
rect 2416 4392 2422 4410
rect 2564 4450 2570 4460
rect 3650 4450 3658 4460
rect 2564 4410 3658 4450
rect 2564 4392 2570 4410
rect 2416 4390 2430 4392
rect 2560 4390 2570 4392
rect 3650 4392 3658 4410
rect 3800 4450 3806 4460
rect 4888 4460 4934 4472
rect 4996 4460 5042 4472
rect 4888 4450 4894 4460
rect 3800 4410 4894 4450
rect 3800 4392 3806 4410
rect 3650 4390 3660 4392
rect 3790 4390 3806 4392
rect 2416 4380 2462 4390
rect 2524 4380 2570 4390
rect 3652 4380 3698 4390
rect 3760 4380 3806 4390
rect 4888 4392 4894 4410
rect 5036 4450 5042 4460
rect 6124 4460 7231 4472
rect 6124 4450 6130 4460
rect 5036 4410 6130 4450
rect 5036 4392 5042 4410
rect 4888 4390 4900 4392
rect 5030 4390 5042 4392
rect 4888 4380 4934 4390
rect 4996 4380 5042 4390
rect 6124 4392 6130 4410
rect 6164 4392 7231 4460
rect 6124 4380 7231 4392
rect -7001 3940 -6995 4370
rect -6041 4364 -5041 4370
rect -6041 4350 -6029 4364
rect -6050 4330 -6029 4350
rect -5053 4350 -5041 4364
rect -4805 4364 -3805 4370
rect -4805 4350 -4793 4364
rect -5053 4330 -4793 4350
rect -3817 4350 -3805 4364
rect -3569 4364 -2569 4370
rect -3569 4350 -3557 4364
rect -3817 4330 -3557 4350
rect -2581 4350 -2569 4364
rect -2333 4364 -1333 4370
rect -2333 4350 -2321 4364
rect -2581 4330 -2321 4350
rect -1345 4350 -1333 4364
rect -1097 4364 -97 4370
rect -1097 4350 -1085 4364
rect -1345 4330 -1085 4350
rect -109 4350 -97 4364
rect 139 4364 1139 4370
rect 139 4350 151 4364
rect -109 4330 151 4350
rect 1127 4350 1139 4364
rect 1375 4364 2375 4370
rect 1375 4350 1387 4364
rect 1127 4330 1387 4350
rect 2363 4350 2375 4364
rect 2611 4364 3611 4370
rect 2611 4350 2623 4364
rect 2363 4330 2623 4350
rect 3599 4350 3611 4364
rect 3847 4364 4847 4370
rect 3847 4350 3859 4364
rect 3599 4330 3859 4350
rect 4835 4350 4847 4364
rect 5083 4364 6083 4370
rect 5083 4350 5095 4364
rect 4835 4330 5095 4350
rect 6071 4350 6083 4364
rect 6071 4330 6100 4350
rect -6050 4300 -5720 4330
rect -5730 4260 -5720 4300
rect -5640 4300 -5510 4330
rect -5640 4260 -5630 4300
rect -5520 4260 -5510 4300
rect -5430 4300 -3250 4330
rect -5430 4260 -5420 4300
rect -3260 4260 -3250 4300
rect -3170 4300 -3010 4330
rect -3170 4260 -3160 4300
rect -3020 4260 -3010 4300
rect -2930 4300 -710 4330
rect -2930 4260 -2920 4300
rect -720 4260 -710 4300
rect -630 4300 -530 4330
rect -630 4260 -620 4300
rect -540 4260 -530 4300
rect -450 4300 1760 4330
rect -450 4260 -440 4300
rect 1750 4250 1760 4300
rect 1840 4300 1930 4330
rect 1840 4250 1850 4300
rect 1920 4250 1930 4300
rect 2010 4300 4230 4330
rect 2010 4250 2020 4300
rect 4220 4250 4230 4300
rect 4310 4300 4400 4330
rect 4310 4250 4320 4300
rect 4390 4250 4400 4300
rect 4480 4300 6100 4330
rect 4480 4250 4490 4300
rect -4282 4210 -4168 4216
rect -4462 4200 -4348 4206
rect -4462 4120 -4450 4200
rect -4360 4120 -4348 4200
rect -4282 4130 -4270 4210
rect -4180 4130 -4168 4210
rect -4282 4124 -4168 4130
rect -1932 4200 -1818 4206
rect -4462 4114 -4348 4120
rect -1932 4120 -1920 4200
rect -1830 4120 -1818 4200
rect -1932 4114 -1818 4120
rect -1772 4200 -1658 4206
rect -1772 4120 -1760 4200
rect -1670 4120 -1658 4200
rect -1772 4114 -1658 4120
rect 538 4200 652 4206
rect 538 4120 550 4200
rect 640 4120 652 4200
rect 538 4114 652 4120
rect 698 4200 812 4206
rect 698 4120 710 4200
rect 800 4120 812 4200
rect 698 4114 812 4120
rect 2988 4200 3102 4206
rect 2988 4120 3000 4200
rect 3090 4120 3102 4200
rect 2988 4114 3102 4120
rect 3148 4200 3262 4206
rect 3148 4120 3160 4200
rect 3250 4120 3262 4200
rect 3148 4114 3262 4120
rect 5488 4200 5602 4206
rect 5488 4120 5500 4200
rect 5590 4120 5602 4200
rect 5488 4114 5602 4120
rect 5648 4200 5762 4206
rect 5648 4120 5660 4200
rect 5750 4120 5762 4200
rect 5648 4114 5762 4120
rect -4480 4020 -4470 4070
rect -6050 3990 -4470 4020
rect -4390 4020 -4380 4070
rect -4250 4020 -4240 4070
rect -4390 3990 -4240 4020
rect -4160 4020 -4150 4070
rect -1950 4020 -1940 4080
rect -4160 4000 -1940 4020
rect -1860 4020 -1850 4080
rect -1760 4020 -1750 4080
rect -1860 4000 -1750 4020
rect -1670 4020 -1660 4080
rect 530 4020 540 4070
rect -1670 4000 540 4020
rect -4160 3990 540 4000
rect 620 4020 630 4070
rect 720 4020 730 4070
rect 620 3990 730 4020
rect 810 4020 820 4070
rect 2980 4020 2990 4070
rect 810 3990 2990 4020
rect 3070 4020 3080 4070
rect 3170 4020 3180 4070
rect 3070 3990 3180 4020
rect 3260 4020 3270 4070
rect 5490 4020 5500 4060
rect 3260 3990 5500 4020
rect -6050 3982 5500 3990
rect 5580 4020 5590 4060
rect 5660 4020 5670 4060
rect 5580 3982 5670 4020
rect 5750 4020 5760 4060
rect 5750 3982 6100 4020
rect -6050 3970 -6029 3982
rect -6041 3948 -6029 3970
rect -5053 3970 -4793 3982
rect -5053 3948 -5041 3970
rect -6041 3942 -5041 3948
rect -4805 3948 -4793 3970
rect -3817 3970 -3557 3982
rect -3817 3948 -3805 3970
rect -4805 3942 -3805 3948
rect -3569 3948 -3557 3970
rect -2581 3970 -2321 3982
rect -2581 3948 -2569 3970
rect -3569 3942 -2569 3948
rect -2333 3948 -2321 3970
rect -1345 3970 -1085 3982
rect -1345 3948 -1333 3970
rect -2333 3942 -1333 3948
rect -1097 3948 -1085 3970
rect -109 3970 151 3982
rect -109 3948 -97 3970
rect -1097 3942 -97 3948
rect 139 3948 151 3970
rect 1127 3970 1387 3982
rect 1127 3948 1139 3970
rect 139 3942 1139 3948
rect 1375 3948 1387 3970
rect 2363 3970 2623 3982
rect 2363 3948 2375 3970
rect 1375 3942 2375 3948
rect 2611 3948 2623 3970
rect 3599 3970 3859 3982
rect 3599 3948 3611 3970
rect 2611 3942 3611 3948
rect 3847 3948 3859 3970
rect 4835 3970 5095 3982
rect 4835 3948 4847 3970
rect 3847 3942 4847 3948
rect 5083 3948 5095 3970
rect 6071 3970 6100 3982
rect 6071 3948 6083 3970
rect 5083 3942 6083 3948
rect 7100 3940 7231 4380
rect -7001 3920 -6080 3940
rect 6130 3932 7231 3940
rect -7001 3852 -6122 3920
rect -6088 3910 -6080 3920
rect -5000 3920 -4954 3932
rect -4892 3920 -4846 3932
rect -5000 3910 -4994 3920
rect -6088 3870 -4994 3910
rect -6088 3852 -6080 3870
rect -7001 3830 -6080 3852
rect -5000 3852 -4994 3870
rect -4852 3910 -4846 3920
rect -3764 3920 -3718 3932
rect -3656 3920 -3610 3932
rect -2528 3920 -2482 3932
rect -2420 3920 -2374 3932
rect -3764 3910 -3758 3920
rect -4852 3870 -3758 3910
rect -4852 3852 -4846 3870
rect -5000 3850 -4990 3852
rect -4860 3850 -4846 3852
rect -5000 3840 -4954 3850
rect -4892 3840 -4846 3850
rect -3764 3852 -3758 3870
rect -3616 3910 -3610 3920
rect -2530 3910 -2522 3920
rect -3616 3870 -2522 3910
rect -3616 3852 -3610 3870
rect -3764 3850 -3750 3852
rect -3620 3850 -3610 3852
rect -2530 3852 -2522 3870
rect -2380 3910 -2374 3920
rect -1292 3920 -1246 3932
rect -1184 3920 -1138 3932
rect -1292 3910 -1286 3920
rect -2380 3870 -1286 3910
rect -2380 3852 -2374 3870
rect -2530 3850 -2520 3852
rect -2390 3850 -2374 3852
rect -3764 3840 -3718 3850
rect -3656 3840 -3610 3850
rect -2528 3840 -2482 3850
rect -2420 3840 -2374 3850
rect -1292 3852 -1286 3870
rect -1144 3910 -1138 3920
rect -56 3920 -10 3932
rect 52 3920 98 3932
rect 1180 3920 1226 3932
rect 1288 3920 1334 3932
rect -56 3910 -50 3920
rect -1144 3870 -50 3910
rect -1144 3852 -1138 3870
rect -1292 3850 -1280 3852
rect -1150 3850 -1138 3852
rect -1292 3840 -1246 3850
rect -1184 3840 -1138 3850
rect -56 3852 -50 3870
rect 92 3910 100 3920
rect 1180 3910 1186 3920
rect 92 3870 1186 3910
rect 92 3852 100 3870
rect -56 3850 -40 3852
rect 90 3850 100 3852
rect 1180 3852 1186 3870
rect 1328 3910 1334 3920
rect 2416 3920 2462 3932
rect 2524 3920 2570 3932
rect 3652 3920 3698 3932
rect 3760 3920 3806 3932
rect 2416 3910 2422 3920
rect 1328 3870 2422 3910
rect 1328 3852 1334 3870
rect 1180 3850 1190 3852
rect 1320 3850 1334 3852
rect -56 3840 -10 3850
rect 52 3840 98 3850
rect 1180 3840 1226 3850
rect 1288 3840 1334 3850
rect 2416 3852 2422 3870
rect 2564 3910 2570 3920
rect 3650 3910 3658 3920
rect 2564 3870 3658 3910
rect 2564 3852 2570 3870
rect 2416 3850 2430 3852
rect 2560 3850 2570 3852
rect 3650 3852 3658 3870
rect 3800 3910 3806 3920
rect 4888 3920 4934 3932
rect 4996 3920 5042 3932
rect 4888 3910 4894 3920
rect 3800 3870 4894 3910
rect 3800 3852 3806 3870
rect 3650 3850 3660 3852
rect 3790 3850 3806 3852
rect 2416 3840 2462 3850
rect 2524 3840 2570 3850
rect 3652 3840 3698 3850
rect 3760 3840 3806 3850
rect 4888 3852 4894 3870
rect 5036 3910 5042 3920
rect 6124 3920 7231 3932
rect 6124 3910 6130 3920
rect 5036 3870 6130 3910
rect 5036 3852 5042 3870
rect 4888 3850 4900 3852
rect 5030 3850 5042 3852
rect 4888 3840 4934 3850
rect 4996 3840 5042 3850
rect 6124 3852 6130 3870
rect 6164 3852 7231 3920
rect 6124 3840 7231 3852
rect -7001 3509 -6995 3830
rect -6041 3824 -5041 3830
rect -6041 3810 -6029 3824
rect -6050 3790 -6029 3810
rect -5053 3810 -5041 3824
rect -4805 3824 -3805 3830
rect -4805 3810 -4793 3824
rect -5053 3790 -4793 3810
rect -3817 3810 -3805 3824
rect -3569 3824 -2569 3830
rect -3569 3810 -3557 3824
rect -3817 3790 -3557 3810
rect -2581 3810 -2569 3824
rect -2333 3824 -1333 3830
rect -2333 3810 -2321 3824
rect -2581 3790 -2321 3810
rect -1345 3810 -1333 3824
rect -1097 3824 -97 3830
rect -1097 3810 -1085 3824
rect -1345 3790 -1085 3810
rect -109 3810 -97 3824
rect 139 3824 1139 3830
rect 139 3810 151 3824
rect -109 3790 151 3810
rect 1127 3810 1139 3824
rect 1375 3824 2375 3830
rect 1375 3810 1387 3824
rect 1127 3790 1387 3810
rect 2363 3810 2375 3824
rect 2611 3824 3611 3830
rect 2611 3810 2623 3824
rect 2363 3790 2623 3810
rect 3599 3810 3611 3824
rect 3847 3824 4847 3830
rect 3847 3810 3859 3824
rect 3599 3790 3859 3810
rect 4835 3810 4847 3824
rect 5083 3824 6083 3830
rect 5083 3810 5095 3824
rect 4835 3790 5095 3810
rect 6071 3810 6083 3824
rect 6071 3790 6100 3810
rect -6050 3760 -5720 3790
rect -5730 3720 -5720 3760
rect -5640 3760 -5510 3790
rect -5640 3720 -5630 3760
rect -5520 3720 -5510 3760
rect -5430 3760 -3250 3790
rect -5430 3720 -5420 3760
rect -3260 3710 -3250 3760
rect -3170 3760 -3010 3790
rect -3170 3710 -3160 3760
rect -3020 3710 -3010 3760
rect -2930 3760 -710 3790
rect -2930 3710 -2920 3760
rect -720 3720 -710 3760
rect -630 3760 -520 3790
rect -630 3720 -620 3760
rect -530 3720 -520 3760
rect -440 3760 1750 3790
rect -440 3720 -430 3760
rect 1740 3710 1750 3760
rect 1830 3760 1940 3790
rect 1830 3710 1840 3760
rect 1930 3710 1940 3760
rect 2020 3780 6100 3790
rect 2020 3760 4230 3780
rect 2020 3710 2030 3760
rect 4220 3700 4230 3760
rect 4310 3760 4400 3780
rect 4310 3700 4320 3760
rect 4390 3700 4400 3760
rect 4480 3760 6100 3780
rect 4480 3700 4490 3760
rect 7100 3520 7231 3840
rect -7404 3497 -6995 3509
rect 7225 3509 7231 3520
rect 7628 3509 7634 4623
rect 7225 3497 7634 3509
rect 9540 4623 10065 4635
rect 9540 3509 9662 4623
rect 10059 3509 10065 4623
rect 9540 3500 10065 3509
rect 9656 3497 10065 3500
rect -8816 3390 -8714 3402
rect -8606 3390 -8504 3402
rect -8820 3260 -8810 3390
rect -8720 3260 -8710 3390
rect -8610 3260 -8600 3390
rect -8510 3260 -8500 3390
rect 8494 3380 8576 3392
rect 8654 3380 8736 3392
rect 8490 3290 8500 3380
rect 8570 3290 8580 3380
rect 8650 3290 8660 3380
rect 8730 3290 8740 3380
rect -2210 3270 -1980 3280
rect -8816 3248 -8714 3260
rect -8606 3248 -8504 3260
rect -3760 3220 -3750 3270
rect -4120 3202 -3750 3220
rect -3620 3220 -3610 3270
rect -2440 3260 -2340 3270
rect -2530 3220 -2520 3260
rect -3620 3202 -2520 3220
rect -2390 3220 -2340 3260
rect -2210 3220 -2190 3270
rect -2390 3202 -2190 3220
rect -2110 3202 -2080 3270
rect -2000 3220 -1980 3270
rect -20 3260 80 3290
rect 200 3270 430 3290
rect 2660 3280 2890 3290
rect -1290 3220 -1280 3260
rect -2000 3202 -1280 3220
rect -1150 3220 -1140 3260
rect -50 3220 -40 3260
rect -1150 3202 -40 3220
rect 90 3220 100 3260
rect 200 3220 220 3270
rect 90 3202 220 3220
rect 300 3202 330 3270
rect 410 3220 430 3270
rect 1180 3220 1190 3260
rect 410 3202 1190 3220
rect 1320 3220 1330 3260
rect 2410 3220 2430 3280
rect 1320 3210 2430 3220
rect 2560 3220 2570 3280
rect 2660 3220 2680 3280
rect 2560 3210 2680 3220
rect 1320 3202 2680 3210
rect 2760 3202 2790 3280
rect 2870 3220 2890 3280
rect 8494 3278 8576 3290
rect 8654 3278 8736 3290
rect 3650 3220 3660 3260
rect 2870 3202 3660 3220
rect 3790 3220 3800 3260
rect 3790 3202 4210 3220
rect -4120 3180 -4098 3202
rect -4110 3168 -4098 3180
rect -3122 3180 -2880 3202
rect -3122 3168 -3110 3180
rect -4110 3162 -3110 3168
rect -2892 3168 -2880 3180
rect -1904 3180 -1662 3202
rect -1904 3168 -1892 3180
rect -2892 3162 -1892 3168
rect -1674 3168 -1662 3180
rect -686 3180 -444 3202
rect -686 3168 -674 3180
rect -1674 3162 -674 3168
rect -456 3168 -444 3180
rect 532 3180 774 3202
rect 532 3168 544 3180
rect -456 3162 544 3168
rect 762 3168 774 3180
rect 1750 3180 1992 3202
rect 1750 3168 1762 3180
rect 762 3162 1762 3168
rect 1980 3168 1992 3180
rect 2968 3180 3210 3202
rect 2968 3168 2980 3180
rect 1980 3162 2980 3168
rect 3198 3168 3210 3180
rect 4186 3180 4210 3202
rect 4186 3168 4198 3180
rect 3198 3162 4198 3168
rect -4188 3140 -4142 3152
rect -4188 3130 -4182 3140
rect -4190 3090 -4182 3130
rect -4188 3072 -4182 3090
rect -4148 3130 -4142 3140
rect -3078 3140 -3032 3152
rect -3078 3130 -3072 3140
rect -4148 3090 -3072 3130
rect -4148 3072 -4142 3090
rect -4188 3060 -4142 3072
rect -3078 3072 -3072 3090
rect -3038 3130 -3032 3140
rect -2970 3140 -2924 3152
rect -2970 3130 -2964 3140
rect -3038 3090 -2964 3130
rect -3038 3072 -3032 3090
rect -3078 3060 -3032 3072
rect -2970 3072 -2964 3090
rect -2930 3130 -2924 3140
rect -1860 3140 -1814 3152
rect -1752 3140 -1706 3152
rect -1860 3130 -1854 3140
rect -2930 3090 -1854 3130
rect -2930 3072 -2924 3090
rect -2970 3060 -2924 3072
rect -1860 3072 -1854 3090
rect -1820 3072 -1746 3140
rect -1712 3130 -1706 3140
rect -642 3140 -596 3152
rect -534 3140 -488 3152
rect -642 3130 -636 3140
rect -1712 3090 -636 3130
rect -1712 3072 -1706 3090
rect -1860 3070 -1706 3072
rect -1860 3060 -1814 3070
rect -1752 3060 -1706 3070
rect -642 3072 -636 3090
rect -602 3072 -528 3140
rect -494 3130 -488 3140
rect 576 3140 622 3152
rect 684 3140 730 3152
rect 576 3130 582 3140
rect -494 3090 582 3130
rect -494 3072 -488 3090
rect -642 3070 -488 3072
rect -642 3060 -596 3070
rect -534 3060 -488 3070
rect 576 3072 582 3090
rect 616 3072 690 3140
rect 724 3130 730 3140
rect 1794 3140 1840 3152
rect 1902 3140 1948 3152
rect 3012 3140 3058 3152
rect 3120 3140 3166 3152
rect 1794 3130 1800 3140
rect 724 3090 1800 3130
rect 724 3072 730 3090
rect 576 3070 730 3072
rect 576 3060 622 3070
rect 684 3060 730 3070
rect 1794 3072 1800 3090
rect 1834 3072 1908 3140
rect 1942 3130 1950 3140
rect 3010 3130 3018 3140
rect 1942 3090 3018 3130
rect 1942 3072 1950 3090
rect 1794 3070 1950 3072
rect 3010 3072 3018 3090
rect 3052 3072 3126 3140
rect 3160 3130 3166 3140
rect 4230 3140 4276 3152
rect 4230 3130 4236 3140
rect 3160 3090 4236 3130
rect 3160 3072 3166 3090
rect 3010 3070 3166 3072
rect 1794 3060 1840 3070
rect 1902 3060 1948 3070
rect 3012 3060 3058 3070
rect 3120 3060 3166 3070
rect 4230 3072 4236 3090
rect 4270 3072 4276 3140
rect 4230 3060 4276 3072
rect -4110 3044 -3110 3050
rect -4110 3030 -4098 3044
rect -4120 3010 -4098 3030
rect -3122 3030 -3110 3044
rect -2892 3044 -1892 3050
rect -2892 3030 -2880 3044
rect -3122 3010 -2880 3030
rect -1904 3030 -1892 3044
rect -1674 3044 -674 3050
rect -1674 3030 -1662 3044
rect -1904 3010 -1662 3030
rect -686 3030 -674 3044
rect -456 3044 544 3050
rect -456 3030 -444 3044
rect -686 3010 -444 3030
rect 532 3030 544 3044
rect 762 3044 1762 3050
rect 762 3030 774 3044
rect 532 3010 774 3030
rect 1750 3030 1762 3044
rect 1980 3044 2980 3050
rect 1980 3030 1992 3044
rect 1750 3010 1992 3030
rect 2968 3030 2980 3044
rect 3198 3044 4198 3050
rect 3198 3030 3210 3044
rect 2968 3010 3210 3030
rect 4186 3030 4198 3044
rect 4186 3010 4210 3030
rect -4120 3000 1200 3010
rect -4120 2990 -3810 3000
rect -3820 2920 -3810 2990
rect -3720 2920 -3670 3000
rect -3580 2990 1200 3000
rect -3580 2920 -3570 2990
rect -1230 2940 -1130 2990
rect 1190 2940 1200 2990
rect 1290 2940 1340 3010
rect 1430 2990 4210 3010
rect 1430 2940 1440 2990
rect -3810 2770 -3580 2920
rect -2302 2910 -2168 2916
rect -2302 2800 -2290 2910
rect -2180 2800 -2168 2910
rect -2302 2794 -2168 2800
rect -1442 2910 -1308 2916
rect -1442 2800 -1430 2910
rect -1320 2800 -1308 2910
rect -1442 2794 -1308 2800
rect -232 2910 -98 2916
rect -232 2800 -220 2910
rect -110 2800 -98 2910
rect -232 2794 -98 2800
rect 618 2910 752 2916
rect 618 2800 630 2910
rect 740 2800 752 2910
rect 618 2794 752 2800
rect -3820 2720 -3810 2770
rect -4120 2702 -3810 2720
rect -3720 2702 -3670 2770
rect -3580 2720 -3570 2770
rect -2440 2720 -2340 2770
rect -20 2720 80 2790
rect 1200 2760 1430 2940
rect 3650 2930 3750 2990
rect 2188 2910 2322 2916
rect 2188 2800 2200 2910
rect 2310 2800 2322 2910
rect 2188 2794 2322 2800
rect 3068 2910 3202 2916
rect 3068 2800 3080 2910
rect 3190 2800 3202 2910
rect 3068 2794 3202 2800
rect 1190 2720 1200 2760
rect -3580 2702 1200 2720
rect 1290 2702 1340 2760
rect 1430 2720 1440 2760
rect 2410 2720 2510 2780
rect 1430 2702 4210 2720
rect -4120 2680 -4098 2702
rect -4110 2668 -4098 2680
rect -3122 2680 -2880 2702
rect -3122 2668 -3110 2680
rect -4110 2662 -3110 2668
rect -2892 2668 -2880 2680
rect -1904 2680 -1662 2702
rect -1904 2668 -1892 2680
rect -2892 2662 -1892 2668
rect -1674 2668 -1662 2680
rect -686 2680 -444 2702
rect -686 2668 -674 2680
rect -1674 2662 -674 2668
rect -456 2668 -444 2680
rect 532 2680 774 2702
rect 1750 2680 1992 2702
rect 532 2668 544 2680
rect -456 2662 544 2668
rect 762 2668 774 2680
rect 1750 2668 1762 2680
rect 762 2662 1762 2668
rect 1980 2668 1992 2680
rect 2968 2680 3210 2702
rect 2968 2668 2980 2680
rect 1980 2662 2980 2668
rect 3198 2668 3210 2680
rect 4186 2680 4210 2702
rect 4186 2668 4198 2680
rect 3198 2662 4198 2668
rect -4188 2640 -4142 2652
rect -4188 2572 -4182 2640
rect -4148 2630 -4142 2640
rect -3078 2640 -3032 2652
rect -3078 2630 -3072 2640
rect -4148 2590 -3072 2630
rect -4148 2572 -4142 2590
rect -4188 2560 -4142 2572
rect -3078 2572 -3072 2590
rect -3038 2630 -3032 2640
rect -2970 2640 -2924 2652
rect -2970 2630 -2964 2640
rect -3038 2590 -2964 2630
rect -3038 2572 -3032 2590
rect -3078 2560 -3032 2572
rect -2970 2572 -2964 2590
rect -2930 2630 -2924 2640
rect -1860 2640 -1814 2652
rect -1752 2640 -1706 2652
rect -1860 2630 -1854 2640
rect -2930 2590 -1854 2630
rect -2930 2572 -2924 2590
rect -2970 2560 -2924 2572
rect -1860 2572 -1854 2590
rect -1820 2572 -1746 2640
rect -1712 2630 -1706 2640
rect -642 2640 -596 2652
rect -534 2640 -488 2652
rect -642 2630 -636 2640
rect -1712 2590 -636 2630
rect -1712 2572 -1706 2590
rect -1860 2570 -1706 2572
rect -1860 2560 -1814 2570
rect -1752 2560 -1706 2570
rect -642 2572 -636 2590
rect -602 2572 -528 2640
rect -494 2630 -488 2640
rect 576 2640 622 2652
rect 684 2640 730 2652
rect 576 2630 582 2640
rect -494 2590 582 2630
rect -494 2572 -488 2590
rect -642 2570 -488 2572
rect -642 2560 -596 2570
rect -534 2560 -488 2570
rect 576 2572 582 2590
rect 616 2572 690 2640
rect 724 2630 730 2640
rect 1794 2640 1840 2652
rect 1902 2640 1948 2652
rect 3012 2640 3058 2652
rect 3120 2640 3166 2652
rect 1794 2630 1800 2640
rect 724 2590 1800 2630
rect 724 2572 730 2590
rect 576 2570 730 2572
rect 576 2560 622 2570
rect 684 2560 730 2570
rect 1794 2572 1800 2590
rect 1834 2572 1908 2640
rect 1942 2630 1950 2640
rect 3010 2630 3018 2640
rect 1942 2590 3018 2630
rect 1942 2572 1950 2590
rect 1794 2570 1950 2572
rect 3010 2572 3018 2590
rect 3052 2572 3126 2640
rect 3160 2630 3166 2640
rect 4230 2640 4276 2652
rect 4230 2630 4236 2640
rect 3160 2590 4236 2630
rect 3160 2572 3166 2590
rect 3010 2570 3166 2572
rect 1794 2560 1840 2570
rect 1902 2560 1948 2570
rect 3012 2560 3058 2570
rect 3120 2560 3166 2570
rect 4230 2572 4236 2590
rect 4270 2630 4276 2640
rect 4270 2590 4280 2630
rect 4270 2572 4276 2590
rect 4230 2560 4276 2572
rect -4110 2544 -3110 2550
rect -4110 2530 -4098 2544
rect -4120 2510 -4098 2530
rect -3122 2530 -3110 2544
rect -2892 2544 -1892 2550
rect -2892 2530 -2880 2544
rect -3122 2510 -2880 2530
rect -1904 2530 -1892 2544
rect -1674 2544 -674 2550
rect -1674 2530 -1662 2544
rect -686 2530 -674 2544
rect -456 2544 544 2550
rect -456 2530 -444 2544
rect -1904 2510 -1662 2530
rect -686 2510 -444 2530
rect 532 2530 544 2544
rect 762 2544 1762 2550
rect 762 2530 774 2544
rect 1750 2530 1762 2544
rect 1980 2544 2980 2550
rect 1980 2530 1992 2544
rect 532 2510 774 2530
rect 1750 2510 1992 2530
rect 2968 2530 2980 2544
rect 3198 2544 4198 2550
rect 3198 2530 3210 2544
rect 2968 2510 3210 2530
rect 4186 2530 4198 2544
rect 4186 2510 4210 2530
rect -4120 2490 -3480 2510
rect -3680 2440 -3580 2490
rect -3490 2430 -3480 2490
rect -3400 2490 -3330 2510
rect -3400 2430 -3390 2490
rect -3340 2430 -3330 2490
rect -3250 2490 -990 2510
rect -3250 2430 -3240 2490
rect -2530 2470 -2380 2490
rect -1290 2460 -1130 2490
rect -1230 2440 -1130 2460
rect -1000 2450 -990 2490
rect -910 2490 -840 2510
rect -910 2450 -900 2490
rect -850 2450 -840 2490
rect -760 2490 1490 2510
rect -760 2450 -750 2490
rect -50 2460 100 2490
rect 1210 2430 1310 2490
rect 1480 2450 1490 2490
rect 1570 2490 1630 2510
rect 1570 2450 1580 2490
rect 1620 2450 1630 2490
rect 1710 2490 4210 2510
rect 1710 2450 1720 2490
rect 2420 2460 2570 2490
rect 3650 2460 3800 2490
rect 3650 2430 3750 2460
rect -3120 2280 -2810 2310
rect -3240 2220 -3030 2280
rect -3560 2202 -3030 2220
rect -2950 2202 -2920 2280
rect -2840 2220 -2810 2280
rect 1820 2270 2040 2280
rect -630 2220 -620 2250
rect -2840 2202 -620 2220
rect -540 2220 -530 2250
rect 1820 2220 1830 2270
rect -540 2202 1830 2220
rect 1910 2202 1950 2270
rect 2030 2220 2040 2270
rect 3020 2220 3030 2260
rect 2030 2202 3030 2220
rect 3110 2220 3120 2260
rect 3110 2202 3560 2220
rect -3560 2180 -3538 2202
rect -3550 2168 -3538 2180
rect -2562 2180 -2320 2202
rect -2562 2168 -2550 2180
rect -3550 2162 -2550 2168
rect -2332 2168 -2320 2180
rect -1344 2180 -1102 2202
rect -1344 2168 -1332 2180
rect -2332 2162 -1332 2168
rect -1114 2168 -1102 2180
rect -126 2180 116 2202
rect -126 2168 -114 2180
rect -1114 2162 -114 2168
rect 104 2168 116 2180
rect 1092 2180 1334 2202
rect 1092 2168 1104 2180
rect 104 2162 1104 2168
rect 1322 2168 1334 2180
rect 2310 2180 2552 2202
rect 3528 2180 3560 2202
rect 2310 2168 2322 2180
rect 1322 2162 2322 2168
rect 2540 2168 2552 2180
rect 3528 2168 3540 2180
rect 2540 2162 3540 2168
rect -3628 2140 -3582 2152
rect -3628 2120 -3622 2140
rect -3640 2000 -3622 2120
rect -3628 1972 -3622 2000
rect -3588 2120 -3582 2140
rect -2518 2140 -2472 2152
rect -2518 2120 -2512 2140
rect -3588 2000 -2512 2120
rect -3588 1972 -3582 2000
rect -3628 1960 -3582 1972
rect -2518 1972 -2512 2000
rect -2478 2120 -2472 2140
rect -2410 2140 -2364 2152
rect -2410 2120 -2404 2140
rect -2478 2000 -2404 2120
rect -2478 1972 -2472 2000
rect -2518 1960 -2472 1972
rect -2410 1972 -2404 2000
rect -2370 2120 -2364 2140
rect -1300 2140 -1254 2152
rect -1300 2120 -1294 2140
rect -2370 2100 -1294 2120
rect -2370 2020 -1850 2100
rect -1770 2020 -1294 2100
rect -2370 2000 -1294 2020
rect -2370 1972 -2364 2000
rect -2410 1960 -2364 1972
rect -1300 1972 -1294 2000
rect -1260 2120 -1254 2140
rect -1192 2140 -1146 2152
rect -1192 2120 -1186 2140
rect -1260 2000 -1186 2120
rect -1260 1972 -1254 2000
rect -1300 1960 -1254 1972
rect -1192 1972 -1186 2000
rect -1152 2120 -1146 2140
rect -82 2140 -36 2152
rect -82 2120 -76 2140
rect -1152 2000 -76 2120
rect -1152 1972 -1146 2000
rect -1192 1960 -1146 1972
rect -82 1972 -76 2000
rect -42 2120 -36 2140
rect 26 2140 72 2152
rect 26 2120 32 2140
rect -42 2000 32 2120
rect -42 1972 -36 2000
rect -82 1960 -36 1972
rect 26 1972 32 2000
rect 66 2120 72 2140
rect 1136 2140 1182 2152
rect 1136 2120 1142 2140
rect 66 2100 1142 2120
rect 66 2020 560 2100
rect 640 2020 1142 2100
rect 66 2000 1142 2020
rect 66 1972 72 2000
rect 26 1960 72 1972
rect 1136 1972 1142 2000
rect 1176 2120 1182 2140
rect 1244 2140 1290 2152
rect 1244 2120 1250 2140
rect 1176 2000 1250 2120
rect 1176 1972 1182 2000
rect 1136 1960 1182 1972
rect 1244 1972 1250 2000
rect 1284 2120 1290 2140
rect 2354 2140 2400 2152
rect 2354 2120 2360 2140
rect 1284 2000 2360 2120
rect 1284 1972 1290 2000
rect 1244 1960 1290 1972
rect 2354 1972 2360 2000
rect 2394 2120 2400 2140
rect 2462 2140 2508 2152
rect 2462 2120 2468 2140
rect 2394 2000 2468 2120
rect 2394 1972 2400 2000
rect 2354 1960 2400 1972
rect 2462 1972 2468 2000
rect 2502 2120 2508 2140
rect 3572 2140 3618 2152
rect 3572 2120 3578 2140
rect 2502 2000 3578 2120
rect 2502 1972 2508 2000
rect 2462 1960 2508 1972
rect 3572 1972 3578 2000
rect 3612 1972 3618 2140
rect 3572 1960 3618 1972
rect -3550 1944 -2550 1950
rect -3550 1920 -3538 1944
rect -2562 1920 -2550 1944
rect -2332 1944 -1332 1950
rect -2332 1920 -2320 1944
rect -3560 1910 -3538 1920
rect -2562 1910 -2320 1920
rect -1344 1920 -1332 1944
rect -1114 1944 -114 1950
rect -1114 1920 -1102 1944
rect -1344 1910 -1102 1920
rect -126 1920 -114 1944
rect 104 1944 1104 1950
rect 104 1920 116 1944
rect -126 1910 116 1920
rect 1092 1920 1104 1944
rect 1322 1944 2322 1950
rect 1322 1920 1334 1944
rect 2310 1920 2322 1944
rect 2540 1944 3540 1950
rect 2540 1920 2552 1944
rect 1092 1910 1334 1920
rect 2310 1910 2552 1920
rect 3528 1920 3540 1944
rect 3528 1910 3560 1920
rect -3560 1880 -3110 1910
rect -3120 1840 -3110 1880
rect -3030 1880 1780 1910
rect -3030 1840 -3020 1880
rect 1770 1840 1780 1880
rect 1860 1880 3560 1910
rect 1860 1840 1870 1880
rect -3012 1790 -2878 1796
rect -3012 1700 -3000 1790
rect -2890 1700 -2878 1790
rect -3012 1694 -2878 1700
rect 1898 1790 2032 1796
rect 1898 1700 1910 1790
rect 2020 1700 2032 1790
rect 1898 1694 2032 1700
rect -630 1600 -620 1630
rect -3560 1582 -620 1600
rect -540 1600 -530 1630
rect 3020 1600 3030 1640
rect -540 1582 3030 1600
rect 3110 1600 3120 1640
rect 3110 1582 3560 1600
rect -3560 1560 -3538 1582
rect -3550 1548 -3538 1560
rect -2562 1560 -2320 1582
rect -2562 1548 -2550 1560
rect -3550 1542 -2550 1548
rect -2332 1548 -2320 1560
rect -1344 1560 -1102 1582
rect -1344 1548 -1332 1560
rect -2332 1542 -1332 1548
rect -1114 1548 -1102 1560
rect -126 1560 116 1582
rect -126 1548 -114 1560
rect -1114 1542 -114 1548
rect 104 1548 116 1560
rect 1092 1560 1334 1582
rect 1092 1548 1104 1560
rect 104 1542 1104 1548
rect 1322 1548 1334 1560
rect 2310 1560 2552 1582
rect 3528 1560 3560 1582
rect 2310 1548 2322 1560
rect 1322 1542 2322 1548
rect 2540 1548 2552 1560
rect 3528 1548 3540 1560
rect 2540 1542 3540 1548
rect -3628 1520 -3582 1532
rect -3628 1490 -3622 1520
rect -3660 1390 -3622 1490
rect -3628 1352 -3622 1390
rect -3588 1500 -3582 1520
rect -2518 1520 -2472 1532
rect -2518 1500 -2512 1520
rect -3588 1380 -2512 1500
rect -3588 1352 -3582 1380
rect -3628 1340 -3582 1352
rect -2518 1352 -2512 1380
rect -2478 1500 -2472 1520
rect -2410 1520 -2364 1532
rect -2410 1500 -2404 1520
rect -2478 1480 -2404 1500
rect -2370 1500 -2364 1520
rect -1300 1520 -1254 1532
rect -1300 1500 -1294 1520
rect -2370 1480 -1294 1500
rect -2478 1400 -2460 1480
rect -2370 1400 -2340 1480
rect -2250 1400 -1850 1480
rect -1770 1400 -1294 1480
rect -2478 1380 -2404 1400
rect -2478 1352 -2472 1380
rect -2518 1340 -2472 1352
rect -2410 1352 -2404 1380
rect -2370 1380 -1294 1400
rect -2370 1352 -2364 1380
rect -2410 1340 -2364 1352
rect -1300 1352 -1294 1380
rect -1260 1500 -1254 1520
rect -1192 1520 -1146 1532
rect -1192 1500 -1186 1520
rect -1260 1380 -1186 1500
rect -1260 1352 -1254 1380
rect -1300 1340 -1254 1352
rect -1192 1352 -1186 1380
rect -1152 1500 -1146 1520
rect -82 1520 -36 1532
rect -82 1500 -76 1520
rect -1152 1380 -76 1500
rect -1152 1352 -1146 1380
rect -1192 1340 -1146 1352
rect -82 1352 -76 1380
rect -42 1500 -36 1520
rect 26 1520 72 1532
rect 26 1500 32 1520
rect -42 1480 32 1500
rect 66 1500 72 1520
rect 1136 1520 1182 1532
rect 1136 1500 1142 1520
rect 66 1480 1142 1500
rect -42 1400 -10 1480
rect 80 1400 110 1480
rect 200 1400 560 1480
rect 640 1400 1142 1480
rect -42 1380 32 1400
rect -42 1352 -36 1380
rect -82 1340 -36 1352
rect 26 1352 32 1380
rect 66 1380 1142 1400
rect 66 1352 72 1380
rect 26 1340 72 1352
rect 1136 1352 1142 1380
rect 1176 1500 1182 1520
rect 1244 1520 1290 1532
rect 1244 1500 1250 1520
rect 1176 1380 1250 1500
rect 1176 1352 1182 1380
rect 1136 1340 1182 1352
rect 1244 1352 1250 1380
rect 1284 1500 1290 1520
rect 2354 1520 2400 1532
rect 2354 1500 2360 1520
rect 1284 1380 2360 1500
rect 1284 1352 1290 1380
rect 1244 1340 1290 1352
rect 2354 1352 2360 1380
rect 2394 1500 2400 1520
rect 2462 1520 2508 1532
rect 2462 1500 2468 1520
rect 2394 1490 2468 1500
rect 2502 1500 2508 1520
rect 3572 1520 3618 1532
rect 3572 1500 3578 1520
rect 2502 1490 3578 1500
rect 2394 1400 2420 1490
rect 2630 1400 3578 1490
rect 2394 1380 2468 1400
rect 2394 1352 2400 1380
rect 2354 1340 2400 1352
rect 2462 1352 2468 1380
rect 2502 1380 3578 1400
rect 2502 1352 2508 1380
rect 2462 1340 2508 1352
rect 3572 1352 3578 1380
rect 3612 1500 3618 1520
rect 3612 1380 3620 1500
rect 3612 1352 3618 1380
rect 3572 1340 3618 1352
rect -3550 1324 -2550 1330
rect -3550 1300 -3538 1324
rect -2562 1300 -2550 1324
rect -2332 1324 -1332 1330
rect -2332 1300 -2320 1324
rect -3560 1290 -3538 1300
rect -2562 1290 -2320 1300
rect -1344 1300 -1332 1324
rect -1114 1324 -114 1330
rect -1114 1300 -1102 1324
rect -1344 1290 -1102 1300
rect -126 1300 -114 1324
rect 104 1324 1104 1330
rect 104 1300 116 1324
rect -126 1290 116 1300
rect 1092 1300 1104 1324
rect 1322 1324 2322 1330
rect 1322 1300 1334 1324
rect 2310 1300 2322 1324
rect 2540 1324 3540 1330
rect 2540 1300 2552 1324
rect 1092 1290 1334 1300
rect 2310 1290 2552 1300
rect 3528 1300 3540 1324
rect 3528 1290 3560 1300
rect -3560 1260 -3110 1290
rect -3120 1220 -3110 1260
rect -3030 1260 1780 1290
rect -3030 1220 -3020 1260
rect 1770 1220 1780 1260
rect 1860 1260 3560 1290
rect 1860 1220 1870 1260
rect -1240 1020 -1230 1050
rect -4120 982 -1230 1020
rect -1140 1020 -1130 1050
rect 3640 1020 3650 1070
rect -1140 990 3650 1020
rect 3740 1020 3750 1070
rect 3740 990 4200 1020
rect -1140 982 4200 990
rect -4120 980 -4098 982
rect -4110 948 -4098 980
rect -3122 980 -2880 982
rect -3122 948 -3110 980
rect -4110 942 -3110 948
rect -2892 948 -2880 980
rect -1904 980 -1662 982
rect -1904 948 -1892 980
rect -2892 942 -1892 948
rect -1674 948 -1662 980
rect -686 980 -444 982
rect -686 948 -674 980
rect -1674 942 -674 948
rect -456 948 -444 980
rect 532 980 774 982
rect 532 948 544 980
rect -456 942 544 948
rect 762 948 774 980
rect 1750 980 1992 982
rect 1750 948 1762 980
rect 762 942 1762 948
rect 1980 948 1992 980
rect 2968 980 3210 982
rect 2968 948 2980 980
rect 1980 942 2980 948
rect 3198 948 3210 980
rect 4186 980 4200 982
rect 4186 948 4198 980
rect 3198 942 4198 948
rect -4188 920 -4142 932
rect -4188 900 -4182 920
rect -4200 780 -4182 900
rect -4188 752 -4182 780
rect -4148 900 -4142 920
rect -3078 920 -3032 932
rect -3078 900 -3072 920
rect -4148 780 -3072 900
rect -4148 752 -4142 780
rect -4188 740 -4142 752
rect -3078 752 -3072 780
rect -3038 900 -3032 920
rect -2970 920 -2924 932
rect -2970 900 -2964 920
rect -3038 780 -2964 900
rect -3038 752 -3032 780
rect -3078 740 -3032 752
rect -2970 752 -2964 780
rect -2930 900 -2924 920
rect -1860 920 -1814 932
rect -1860 900 -1854 920
rect -2930 880 -1854 900
rect -2930 800 -2460 880
rect -2370 800 -2340 880
rect -2250 800 -1854 880
rect -2930 780 -1854 800
rect -2930 752 -2924 780
rect -2970 740 -2924 752
rect -1860 752 -1854 780
rect -1820 900 -1814 920
rect -1752 920 -1706 932
rect -1752 900 -1746 920
rect -1820 780 -1746 900
rect -1820 752 -1814 780
rect -1860 740 -1814 752
rect -1752 752 -1746 780
rect -1712 900 -1706 920
rect -642 920 -596 932
rect -642 900 -636 920
rect -1712 780 -636 900
rect -1712 752 -1706 780
rect -1752 740 -1706 752
rect -642 752 -636 780
rect -602 900 -596 920
rect -534 920 -488 932
rect -534 900 -528 920
rect -602 780 -528 900
rect -602 752 -596 780
rect -642 740 -596 752
rect -534 752 -528 780
rect -494 900 -488 920
rect 576 920 622 932
rect 576 900 582 920
rect -494 880 582 900
rect -494 800 -10 880
rect 80 800 110 880
rect 200 800 582 880
rect -494 780 582 800
rect -494 752 -488 780
rect -534 740 -488 752
rect 576 752 582 780
rect 616 900 622 920
rect 684 920 730 932
rect 684 900 690 920
rect 616 780 690 900
rect 616 752 622 780
rect 576 740 622 752
rect 684 752 690 780
rect 724 900 730 920
rect 1794 920 1840 932
rect 1794 900 1800 920
rect 724 780 1800 900
rect 724 752 730 780
rect 684 740 730 752
rect 1794 752 1800 780
rect 1834 900 1840 920
rect 1902 920 1948 932
rect 1902 900 1908 920
rect 1834 780 1908 900
rect 1834 752 1840 780
rect 1794 740 1840 752
rect 1902 752 1908 780
rect 1942 900 1948 920
rect 3012 920 3058 932
rect 3012 900 3018 920
rect 1942 880 3018 900
rect 1942 800 2420 880
rect 2510 800 2540 880
rect 2630 800 3018 880
rect 1942 780 3018 800
rect 1942 752 1948 780
rect 1902 740 1948 752
rect 3012 752 3018 780
rect 3052 900 3058 920
rect 3120 920 3166 932
rect 3120 900 3126 920
rect 3052 780 3126 900
rect 3052 752 3058 780
rect 3012 740 3058 752
rect 3120 752 3126 780
rect 3160 900 3166 920
rect 4230 920 4276 932
rect 4230 900 4236 920
rect 3160 780 4236 900
rect 3160 752 3166 780
rect 3120 740 3166 752
rect 4230 752 4236 780
rect 4270 900 4276 920
rect 4270 780 4280 900
rect 4270 752 4276 780
rect 4230 740 4276 752
rect -4110 724 -3110 730
rect -4110 700 -4098 724
rect -4120 690 -4098 700
rect -3122 700 -3110 724
rect -2892 724 -1892 730
rect -2892 700 -2880 724
rect -3122 690 -2880 700
rect -1904 700 -1892 724
rect -1674 724 -674 730
rect -1674 700 -1662 724
rect -1904 690 -1662 700
rect -686 700 -674 724
rect -456 724 544 730
rect -456 700 -444 724
rect -686 690 -444 700
rect 532 700 544 724
rect 762 724 1762 730
rect 762 700 774 724
rect 532 690 774 700
rect 1750 700 1762 724
rect 1980 724 2980 730
rect 1980 700 1992 724
rect 1750 690 1992 700
rect 2968 700 2980 724
rect 3198 724 4198 730
rect 3198 700 3210 724
rect 2968 690 3210 700
rect 4186 700 4198 724
rect 4186 690 4200 700
rect -4120 660 -3810 690
rect -3820 640 -3810 660
rect -3720 660 -3670 690
rect -3720 640 -3710 660
rect -3680 640 -3670 660
rect -3580 660 1200 690
rect -3580 640 -3570 660
rect 1190 640 1200 660
rect 1290 660 1340 690
rect 1290 640 1300 660
rect 1330 640 1340 660
rect 1430 660 4200 690
rect 1430 640 1440 660
rect -3080 590 -2920 600
rect -3080 490 -3060 590
rect -2940 490 -2920 590
rect -3080 420 -2920 490
rect -1860 590 -1700 600
rect -1860 490 -1840 590
rect -1720 490 -1700 590
rect -1860 420 -1700 490
rect -650 590 -490 600
rect 578 590 722 596
rect 3018 590 3162 596
rect -650 490 -630 590
rect -510 490 -490 590
rect -1240 420 -1230 450
rect -4120 382 -1230 420
rect -1140 420 -1130 450
rect -650 420 -490 490
rect 570 490 590 590
rect 710 490 730 590
rect 1808 580 1952 586
rect 570 420 730 490
rect 1800 480 1820 580
rect 1940 480 1960 580
rect 1800 420 1960 480
rect 3010 490 3030 590
rect 3150 490 3170 590
rect 3010 420 3170 490
rect 3640 420 3650 470
rect -1140 390 3650 420
rect 3740 420 3750 470
rect 3740 390 4200 420
rect -1140 382 4200 390
rect -4120 380 -4098 382
rect -4110 348 -4098 380
rect -3122 380 -2880 382
rect -3122 348 -3110 380
rect -4110 342 -3110 348
rect -2892 348 -2880 380
rect -1904 380 -1662 382
rect -1904 348 -1892 380
rect -2892 342 -1892 348
rect -1674 348 -1662 380
rect -686 380 -444 382
rect -686 348 -674 380
rect -1674 342 -674 348
rect -456 348 -444 380
rect 532 380 774 382
rect 532 348 544 380
rect -456 342 544 348
rect 762 348 774 380
rect 1750 380 1992 382
rect 1750 348 1762 380
rect 762 342 1762 348
rect 1980 348 1992 380
rect 2968 380 3210 382
rect 2968 348 2980 380
rect 1980 342 2980 348
rect 3198 348 3210 380
rect 4186 380 4200 382
rect 4186 348 4198 380
rect 3198 342 4198 348
rect -4188 320 -4142 332
rect -4188 152 -4182 320
rect -4148 300 -4142 320
rect -3078 320 -3032 332
rect -3078 300 -3072 320
rect -4148 180 -3072 300
rect -4148 152 -4142 180
rect -4188 140 -4142 152
rect -3078 152 -3072 180
rect -3038 300 -3032 320
rect -2970 320 -2924 332
rect -2970 300 -2964 320
rect -3038 180 -2964 300
rect -3038 152 -3032 180
rect -3078 140 -3032 152
rect -2970 152 -2964 180
rect -2930 300 -2924 320
rect -1860 320 -1814 332
rect -1860 300 -1854 320
rect -2930 280 -1854 300
rect -2930 200 -2460 280
rect -2370 200 -2340 280
rect -2250 200 -1854 280
rect -2930 180 -1854 200
rect -2930 152 -2924 180
rect -2970 140 -2924 152
rect -1860 152 -1854 180
rect -1820 300 -1814 320
rect -1752 320 -1706 332
rect -1752 300 -1746 320
rect -1820 180 -1746 300
rect -1820 152 -1814 180
rect -1860 140 -1814 152
rect -1752 152 -1746 180
rect -1712 300 -1706 320
rect -642 320 -596 332
rect -642 300 -636 320
rect -1712 180 -636 300
rect -1712 152 -1706 180
rect -1752 140 -1706 152
rect -642 152 -636 180
rect -602 300 -596 320
rect -534 320 -488 332
rect -534 300 -528 320
rect -602 180 -528 300
rect -602 152 -596 180
rect -642 140 -596 152
rect -534 152 -528 180
rect -494 300 -488 320
rect 576 320 622 332
rect 576 300 582 320
rect -494 280 582 300
rect -494 200 -10 280
rect 80 200 110 280
rect 200 200 582 280
rect -494 180 582 200
rect -494 152 -488 180
rect -534 140 -488 152
rect 576 152 582 180
rect 616 300 622 320
rect 684 320 730 332
rect 684 300 690 320
rect 616 180 690 300
rect 616 152 622 180
rect 576 140 622 152
rect 684 152 690 180
rect 724 300 730 320
rect 1794 320 1840 332
rect 1794 300 1800 320
rect 724 180 1800 300
rect 724 152 730 180
rect 684 140 730 152
rect 1794 152 1800 180
rect 1834 300 1840 320
rect 1902 320 1948 332
rect 1902 300 1908 320
rect 1834 180 1908 300
rect 1834 152 1840 180
rect 1794 140 1840 152
rect 1902 152 1908 180
rect 1942 300 1948 320
rect 3012 320 3058 332
rect 3012 300 3018 320
rect 1942 280 3018 300
rect 1942 200 2420 280
rect 2510 200 2540 280
rect 2630 200 3018 280
rect 1942 180 3018 200
rect 1942 152 1948 180
rect 1902 140 1948 152
rect 3012 152 3018 180
rect 3052 300 3058 320
rect 3120 320 3166 332
rect 3120 300 3126 320
rect 3052 180 3126 300
rect 3052 152 3058 180
rect 3012 140 3058 152
rect 3120 152 3126 180
rect 3160 300 3166 320
rect 4230 320 4276 332
rect 4230 300 4236 320
rect 3160 180 4236 300
rect 3160 152 3166 180
rect 3120 140 3166 152
rect 4230 152 4236 180
rect 4270 300 4276 320
rect 4270 180 4280 300
rect 4270 152 4276 180
rect 4230 140 4276 152
rect -4110 124 -3110 130
rect -4110 100 -4098 124
rect -3122 100 -3110 124
rect -2892 124 -1892 130
rect -2892 100 -2880 124
rect -4120 90 -4098 100
rect -3122 90 -2880 100
rect -1904 100 -1892 124
rect -1674 124 -674 130
rect -1674 100 -1662 124
rect -1904 90 -1662 100
rect -686 100 -674 124
rect -456 124 544 130
rect -456 100 -444 124
rect -686 90 -444 100
rect 532 100 544 124
rect 762 124 1762 130
rect 762 100 774 124
rect 532 90 774 100
rect 1750 100 1762 124
rect 1980 124 2980 130
rect 1980 100 1992 124
rect 1750 90 1992 100
rect 2968 100 2980 124
rect 3198 124 4198 130
rect 3198 100 3210 124
rect 2968 90 3210 100
rect 4186 100 4198 124
rect 4186 90 4200 100
rect -4120 60 -3810 90
rect -3820 20 -3810 60
rect -3720 60 -3670 90
rect -3720 20 -3710 60
rect -3680 20 -3670 60
rect -3580 60 1200 90
rect -3580 20 -3570 60
rect 1190 40 1200 60
rect 1290 60 1340 90
rect 1290 40 1300 60
rect 1330 40 1340 60
rect 1430 60 4200 90
rect 1430 40 1440 60
<< via1 >>
rect -2600 9030 -2510 9100
rect -2430 9030 -2340 9100
rect -110 9030 -20 9100
rect 60 9030 150 9100
rect 2350 9030 2430 9110
rect 2520 9030 2600 9110
rect -2600 8922 -2520 8990
rect -2430 8922 -2350 8990
rect -110 8922 -30 8990
rect 60 8922 140 8990
rect 2350 8922 2430 8980
rect 2520 8922 2600 8980
rect -2600 8910 -2520 8922
rect -2430 8910 -2350 8922
rect -110 8910 -30 8922
rect 60 8910 140 8922
rect 2350 8900 2430 8922
rect 2520 8900 2600 8922
rect -3480 8764 -3400 8820
rect -3330 8764 -3250 8820
rect -3150 8792 -3120 8860
rect -3120 8792 -3046 8860
rect -3046 8792 -3020 8860
rect -1910 8792 -1884 8860
rect -1884 8792 -1810 8860
rect -1810 8792 -1780 8860
rect -3150 8790 -3020 8792
rect -1910 8790 -1780 8792
rect -990 8764 -910 8820
rect -840 8764 -760 8820
rect -680 8792 -648 8860
rect -648 8792 -574 8860
rect -574 8792 -550 8860
rect 560 8792 588 8860
rect 588 8792 662 8860
rect 662 8792 690 8860
rect -680 8790 -550 8792
rect 560 8790 690 8792
rect 1490 8764 1570 8820
rect 1640 8764 1720 8820
rect 1800 8792 1824 8860
rect 1824 8792 1898 8860
rect 1898 8792 1930 8860
rect 3030 8792 3060 8860
rect 3060 8792 3134 8860
rect 3134 8792 3160 8860
rect 1800 8790 1930 8792
rect 3030 8790 3160 8792
rect -3870 8730 -3790 8750
rect -3700 8730 -3620 8750
rect -3480 8740 -3400 8764
rect -3330 8740 -3250 8764
rect -1350 8730 -1270 8750
rect -1180 8730 -1100 8750
rect -990 8740 -910 8764
rect -840 8740 -760 8764
rect 1140 8730 1220 8750
rect 1310 8730 1390 8750
rect 1490 8740 1570 8764
rect 1640 8740 1720 8764
rect 3590 8730 3670 8750
rect 3760 8730 3840 8750
rect -3870 8670 -3790 8730
rect -3700 8670 -3620 8730
rect -1350 8670 -1270 8730
rect -1180 8670 -1100 8730
rect 1140 8670 1220 8730
rect 1310 8670 1390 8730
rect 3590 8670 3670 8730
rect 3760 8670 3840 8730
rect -2600 8382 -2520 8450
rect -2430 8382 -2350 8450
rect -110 8382 -30 8450
rect 60 8382 140 8450
rect 2350 8382 2430 8440
rect 2520 8382 2600 8440
rect -2600 8370 -2520 8382
rect -2430 8370 -2350 8382
rect -110 8370 -30 8382
rect 60 8370 140 8382
rect 2350 8360 2430 8382
rect 2520 8360 2600 8382
rect -3480 8224 -3400 8280
rect -3330 8224 -3250 8280
rect -3150 8252 -3120 8320
rect -3120 8252 -3046 8320
rect -3046 8252 -3020 8320
rect -1910 8252 -1884 8320
rect -1884 8252 -1810 8320
rect -1810 8252 -1780 8320
rect -3150 8250 -3020 8252
rect -1910 8250 -1780 8252
rect -990 8224 -910 8280
rect -840 8224 -760 8280
rect -680 8252 -648 8320
rect -648 8252 -574 8320
rect -574 8252 -550 8320
rect 560 8252 588 8320
rect 588 8252 662 8320
rect 662 8252 690 8320
rect -680 8250 -550 8252
rect 560 8250 690 8252
rect 1490 8224 1570 8280
rect 1640 8224 1720 8280
rect 1800 8252 1824 8320
rect 1824 8252 1898 8320
rect 1898 8252 1930 8320
rect 3030 8252 3060 8320
rect 3060 8252 3134 8320
rect 3134 8252 3160 8320
rect 1800 8250 1930 8252
rect 3030 8250 3160 8252
rect -3870 8190 -3790 8210
rect -3700 8190 -3620 8210
rect -3480 8200 -3400 8224
rect -3330 8200 -3250 8224
rect -1350 8190 -1270 8210
rect -1180 8190 -1100 8210
rect -990 8200 -910 8224
rect -840 8200 -760 8224
rect 1140 8190 1220 8210
rect 1310 8190 1390 8210
rect 1490 8200 1570 8224
rect 1640 8200 1720 8224
rect 3590 8190 3670 8200
rect 3760 8190 3840 8200
rect -3870 8130 -3790 8190
rect -3700 8130 -3620 8190
rect -1350 8130 -1270 8190
rect -1180 8130 -1100 8190
rect 1140 8130 1220 8190
rect 1310 8130 1390 8190
rect 3590 8120 3670 8190
rect 3760 8120 3840 8190
rect -2590 7980 -2500 8050
rect -2450 7980 -2360 8050
rect -110 7980 -20 8050
rect 50 7990 140 8060
rect 2350 7990 2430 8060
rect 2520 7990 2600 8060
rect -2600 7842 -2520 7910
rect -2430 7842 -2350 7910
rect -110 7842 -30 7920
rect 60 7842 140 7920
rect 2350 7842 2430 7900
rect 2520 7842 2600 7900
rect -2600 7830 -2520 7842
rect -2430 7830 -2350 7842
rect -110 7840 -30 7842
rect 60 7840 140 7842
rect 2350 7820 2430 7842
rect 2520 7820 2600 7842
rect -3480 7684 -3400 7740
rect -3330 7684 -3250 7740
rect -3150 7712 -3120 7780
rect -3120 7712 -3046 7780
rect -3046 7712 -3020 7780
rect -1910 7712 -1884 7780
rect -1884 7712 -1810 7780
rect -1810 7712 -1780 7780
rect -3150 7710 -3020 7712
rect -1910 7710 -1780 7712
rect -990 7684 -910 7740
rect -840 7684 -760 7740
rect -680 7712 -648 7780
rect -648 7712 -574 7780
rect -574 7712 -550 7780
rect 560 7712 588 7780
rect 588 7712 662 7780
rect 662 7712 690 7780
rect -680 7710 -550 7712
rect 560 7710 690 7712
rect 1500 7684 1580 7740
rect 1640 7684 1720 7740
rect 1800 7712 1824 7780
rect 1824 7712 1898 7780
rect 1898 7712 1930 7780
rect 3030 7712 3060 7780
rect 3060 7712 3134 7780
rect 3134 7712 3160 7780
rect 1800 7710 1930 7712
rect 3030 7710 3160 7712
rect -3870 7650 -3790 7670
rect -3700 7650 -3620 7670
rect -3480 7660 -3400 7684
rect -3330 7660 -3250 7684
rect -1350 7650 -1270 7670
rect -1180 7650 -1100 7670
rect -990 7660 -910 7684
rect -840 7660 -760 7684
rect 1500 7660 1580 7684
rect 1640 7660 1720 7684
rect 1140 7650 1220 7660
rect 1310 7650 1390 7660
rect 3590 7650 3670 7670
rect 3760 7650 3840 7670
rect -3870 7590 -3790 7650
rect -3700 7590 -3620 7650
rect -1350 7590 -1270 7650
rect -1180 7590 -1100 7650
rect 1140 7580 1220 7650
rect 1310 7580 1390 7650
rect 3590 7590 3670 7650
rect 3760 7590 3840 7650
rect -2590 7440 -2510 7520
rect -2420 7440 -2340 7520
rect -110 7440 -30 7520
rect 60 7440 140 7520
rect 2350 7440 2430 7520
rect 2520 7440 2600 7520
rect -2590 7310 -2510 7390
rect -2420 7310 -2340 7390
rect -110 7320 -30 7400
rect 60 7320 140 7400
rect 2350 7310 2430 7390
rect 2520 7310 2600 7390
rect -3150 7172 -3120 7240
rect -3120 7172 -3046 7240
rect -3046 7172 -3020 7240
rect -3150 7170 -3020 7172
rect -1910 7172 -1884 7240
rect -1884 7172 -1810 7240
rect -1810 7172 -1780 7240
rect -1910 7170 -1780 7172
rect -680 7172 -648 7240
rect -648 7172 -574 7240
rect -574 7172 -550 7240
rect -680 7170 -550 7172
rect 560 7172 588 7240
rect 588 7172 662 7240
rect 662 7172 690 7240
rect 560 7170 690 7172
rect 1790 7172 1824 7240
rect 1824 7172 1898 7240
rect 1898 7172 1920 7240
rect 1790 7170 1920 7172
rect 3030 7172 3060 7240
rect 3060 7172 3134 7240
rect 3134 7172 3160 7240
rect 3030 7170 3160 7172
rect -3870 7110 -3790 7130
rect -3700 7110 -3620 7130
rect -2190 7110 -2110 7140
rect -2080 7110 -2000 7140
rect -1360 7110 -1280 7130
rect -1190 7110 -1110 7130
rect 220 7110 300 7140
rect 330 7110 410 7140
rect 1130 7110 1210 7130
rect 1300 7110 1380 7130
rect 2680 7110 2760 7130
rect 2790 7110 2870 7130
rect 3620 7110 3700 7130
rect 3790 7110 3870 7130
rect -3870 7050 -3790 7110
rect -3700 7050 -3620 7110
rect -2190 7060 -2110 7110
rect -2080 7060 -2000 7110
rect -1360 7050 -1280 7110
rect -1190 7050 -1110 7110
rect 220 7060 300 7110
rect 330 7060 410 7110
rect 1130 7050 1210 7110
rect 1300 7050 1380 7110
rect 2680 7050 2760 7110
rect 2790 7050 2870 7110
rect 3620 7050 3700 7110
rect 3790 7050 3870 7110
rect -2590 6730 -2510 6810
rect -2420 6730 -2340 6810
rect -110 6740 -30 6820
rect 60 6740 140 6820
rect 2350 6730 2430 6810
rect 2520 6730 2600 6810
rect -3150 6592 -3120 6660
rect -3120 6592 -3046 6660
rect -3046 6592 -3020 6660
rect -3150 6590 -3020 6592
rect -1910 6592 -1884 6660
rect -1884 6592 -1810 6660
rect -1810 6592 -1780 6660
rect -1910 6590 -1780 6592
rect -670 6592 -648 6660
rect -648 6592 -574 6660
rect -574 6592 -540 6660
rect -670 6590 -540 6592
rect 560 6592 588 6660
rect 588 6592 662 6660
rect 662 6592 690 6660
rect 560 6590 690 6592
rect 1790 6592 1824 6660
rect 1824 6592 1898 6660
rect 1898 6592 1920 6660
rect 1790 6590 1920 6592
rect 3030 6592 3060 6660
rect 3060 6592 3134 6660
rect 3134 6592 3160 6660
rect 3030 6590 3160 6592
rect -3870 6530 -3790 6550
rect -3700 6530 -3620 6550
rect -1360 6530 -1280 6550
rect -1190 6530 -1110 6550
rect 220 6530 300 6550
rect 330 6530 410 6550
rect 1130 6530 1210 6540
rect 1300 6530 1380 6540
rect 2680 6530 2760 6550
rect 2790 6530 2870 6550
rect 3620 6530 3700 6550
rect 3790 6530 3870 6550
rect -3870 6470 -3790 6530
rect -3700 6470 -3620 6530
rect -2190 6450 -2110 6530
rect -2080 6450 -2000 6530
rect -1360 6470 -1280 6530
rect -1190 6470 -1110 6530
rect 220 6470 300 6530
rect 330 6470 410 6530
rect 1130 6460 1210 6530
rect 1300 6460 1380 6530
rect 2680 6470 2760 6530
rect 2790 6470 2870 6530
rect 3620 6470 3700 6530
rect 3790 6470 3870 6530
rect -2590 6280 -2500 6360
rect -2430 6280 -2340 6360
rect -110 6280 -30 6350
rect 60 6280 140 6350
rect 2350 6280 2430 6350
rect 2520 6280 2600 6350
rect 9560 6300 9690 6440
rect 9820 6300 9950 6440
rect -9940 6130 -9810 6270
rect -9690 6130 -9560 6270
rect -2590 6150 -2510 6230
rect -2420 6150 -2340 6230
rect -110 6160 -30 6240
rect 60 6160 140 6240
rect 2350 6150 2430 6230
rect 2520 6150 2600 6230
rect -3150 6012 -3120 6080
rect -3120 6012 -3046 6080
rect -3046 6012 -3020 6080
rect -3150 6010 -3020 6012
rect -680 6012 -648 6080
rect -648 6012 -574 6080
rect -574 6012 -550 6080
rect -680 6010 -550 6012
rect 560 6012 588 6080
rect 588 6012 662 6080
rect 662 6012 690 6080
rect 560 6010 690 6012
rect 1790 6012 1824 6080
rect 1824 6012 1898 6080
rect 1898 6012 1920 6080
rect 1790 6010 1920 6012
rect 3030 6012 3060 6080
rect 3060 6012 3134 6080
rect 3134 6012 3160 6080
rect 3030 6010 3160 6012
rect -1360 5950 -1280 5970
rect -1190 5950 -1110 5970
rect 220 5950 300 5970
rect 330 5950 410 5970
rect 1130 5950 1210 5970
rect 1300 5950 1380 5970
rect 2680 5950 2760 5970
rect 2790 5950 2870 5970
rect 3620 5950 3700 5970
rect 3790 5950 3870 5970
rect -3890 5860 -3810 5940
rect -3680 5860 -3600 5940
rect -1360 5890 -1280 5950
rect -1190 5890 -1110 5950
rect 220 5890 300 5950
rect 330 5890 410 5950
rect 1130 5890 1210 5950
rect 1300 5890 1380 5950
rect 2680 5890 2760 5950
rect 2790 5890 2870 5950
rect 3620 5890 3700 5950
rect 3790 5890 3870 5950
rect -4470 5620 -4390 5700
rect -4240 5620 -4160 5700
rect -1920 5610 -1840 5690
rect -1750 5610 -1670 5690
rect 540 5610 620 5690
rect 730 5610 810 5690
rect 2990 5610 3070 5690
rect 3180 5610 3260 5690
rect 5500 5610 5580 5690
rect 5670 5610 5750 5690
rect -4990 5472 -4960 5540
rect -4960 5472 -4886 5540
rect -4886 5472 -4860 5540
rect -4990 5470 -4860 5472
rect -3750 5472 -3724 5540
rect -3724 5472 -3650 5540
rect -3650 5472 -3620 5540
rect -3750 5470 -3620 5472
rect -2520 5472 -2488 5540
rect -2488 5472 -2414 5540
rect -2414 5472 -2390 5540
rect -2520 5470 -2390 5472
rect -1280 5472 -1252 5540
rect -1252 5472 -1178 5540
rect -1178 5472 -1150 5540
rect -1280 5470 -1150 5472
rect -40 5472 -16 5540
rect -16 5472 58 5540
rect 58 5472 90 5540
rect -40 5470 90 5472
rect 1190 5472 1220 5540
rect 1220 5472 1294 5540
rect 1294 5472 1320 5540
rect 1190 5470 1320 5472
rect 2430 5472 2456 5540
rect 2456 5472 2530 5540
rect 2530 5472 2560 5540
rect 2430 5470 2560 5472
rect 3660 5472 3692 5540
rect 3692 5472 3766 5540
rect 3766 5472 3790 5540
rect 3660 5470 3790 5472
rect 4900 5472 4928 5540
rect 4928 5472 5002 5540
rect 5002 5472 5030 5540
rect 4900 5470 5030 5472
rect -5720 5410 -5640 5420
rect -5510 5410 -5430 5420
rect -3240 5410 -3160 5420
rect -3020 5410 -2940 5420
rect -710 5410 -630 5420
rect -530 5410 -450 5420
rect -5720 5340 -5640 5410
rect -5510 5340 -5430 5410
rect -3240 5340 -3160 5410
rect -3020 5340 -2940 5410
rect -710 5340 -630 5410
rect -530 5340 -450 5410
rect 1750 5330 1830 5410
rect 1930 5330 2010 5410
rect 4230 5330 4310 5410
rect 4400 5330 4480 5410
rect -4450 5200 -4360 5280
rect -4270 5200 -4180 5280
rect -1920 5200 -1830 5280
rect -1760 5200 -1670 5280
rect 550 5200 640 5280
rect 710 5200 800 5280
rect 3000 5200 3090 5280
rect 3160 5200 3250 5280
rect 5500 5200 5590 5280
rect 5660 5200 5750 5280
rect -4470 5080 -4390 5160
rect -4240 5080 -4160 5160
rect -1920 5070 -1840 5150
rect -1750 5080 -1670 5160
rect 540 5080 620 5160
rect 730 5080 810 5160
rect 2990 5070 3070 5150
rect 3180 5070 3260 5150
rect 5500 5070 5580 5150
rect 5670 5070 5750 5150
rect -4990 5000 -4860 5010
rect -4990 4940 -4960 5000
rect -4960 4940 -4886 5000
rect -4886 4940 -4860 5000
rect -3750 4932 -3724 5000
rect -3724 4932 -3650 5000
rect -3650 4932 -3620 5000
rect -3750 4930 -3620 4932
rect -2520 4932 -2488 5000
rect -2488 4932 -2414 5000
rect -2414 4932 -2390 5000
rect -2520 4930 -2390 4932
rect -1280 4932 -1252 5000
rect -1252 4932 -1178 5000
rect -1178 4932 -1150 5000
rect -1280 4930 -1150 4932
rect -40 4932 -16 5000
rect -16 4932 58 5000
rect 58 4932 90 5000
rect -40 4930 90 4932
rect 1190 4932 1220 5000
rect 1220 4932 1294 5000
rect 1294 4932 1320 5000
rect 1190 4930 1320 4932
rect 2430 4932 2456 5000
rect 2456 4932 2530 5000
rect 2530 4932 2560 5000
rect 2430 4930 2560 4932
rect 3660 4932 3692 5000
rect 3692 4932 3766 5000
rect 3766 4932 3790 5000
rect 3660 4930 3790 4932
rect 4900 4932 4928 5000
rect 4928 4932 5002 5000
rect 5002 4932 5030 5000
rect 4900 4930 5030 4932
rect -5720 4870 -5640 4880
rect -5510 4870 -5430 4880
rect -3240 4870 -3160 4880
rect -3020 4870 -2940 4880
rect -710 4870 -630 4880
rect -520 4870 -440 4880
rect -5720 4800 -5640 4870
rect -5510 4800 -5430 4870
rect -3240 4800 -3160 4870
rect -3020 4800 -2940 4870
rect -710 4800 -630 4870
rect -520 4800 -440 4870
rect 1750 4790 1830 4870
rect 1930 4790 2010 4870
rect 4230 4790 4310 4870
rect 4400 4790 4480 4870
rect -4470 4540 -4390 4620
rect -4240 4540 -4160 4620
rect -1930 4530 -1850 4610
rect -1760 4530 -1680 4610
rect 540 4530 620 4610
rect 720 4530 800 4610
rect 2990 4530 3070 4610
rect 3180 4530 3260 4610
rect 5500 4530 5580 4610
rect 5670 4530 5750 4610
rect -4990 4392 -4960 4460
rect -4960 4392 -4886 4460
rect -4886 4392 -4860 4460
rect -4990 4390 -4860 4392
rect -3750 4392 -3724 4460
rect -3724 4392 -3650 4460
rect -3650 4392 -3620 4460
rect -3750 4390 -3620 4392
rect -2520 4392 -2488 4460
rect -2488 4392 -2414 4460
rect -2414 4392 -2390 4460
rect -2520 4390 -2390 4392
rect -1280 4392 -1252 4460
rect -1252 4392 -1178 4460
rect -1178 4392 -1150 4460
rect -1280 4390 -1150 4392
rect -40 4392 -16 4460
rect -16 4392 58 4460
rect 58 4392 90 4460
rect -40 4390 90 4392
rect 1190 4392 1220 4460
rect 1220 4392 1294 4460
rect 1294 4392 1320 4460
rect 1190 4390 1320 4392
rect 2430 4392 2456 4460
rect 2456 4392 2530 4460
rect 2530 4392 2560 4460
rect 2430 4390 2560 4392
rect 3660 4392 3692 4460
rect 3692 4392 3766 4460
rect 3766 4392 3790 4460
rect 3660 4390 3790 4392
rect 4900 4392 4928 4460
rect 4928 4392 5002 4460
rect 5002 4392 5030 4460
rect 4900 4390 5030 4392
rect -5720 4330 -5640 4340
rect -5510 4330 -5430 4340
rect -3250 4330 -3170 4340
rect -3010 4330 -2930 4340
rect -710 4330 -630 4340
rect -530 4330 -450 4340
rect -5720 4260 -5640 4330
rect -5510 4260 -5430 4330
rect -3250 4260 -3170 4330
rect -3010 4260 -2930 4330
rect -710 4260 -630 4330
rect -530 4260 -450 4330
rect 1760 4250 1840 4330
rect 1930 4250 2010 4330
rect 4230 4250 4310 4330
rect 4400 4250 4480 4330
rect -4450 4120 -4360 4200
rect -4270 4130 -4180 4210
rect -1920 4120 -1830 4200
rect -1760 4120 -1670 4200
rect 550 4120 640 4200
rect 710 4120 800 4200
rect 3000 4120 3090 4200
rect 3160 4120 3250 4200
rect 5500 4120 5590 4200
rect 5660 4120 5750 4200
rect -4470 3990 -4390 4070
rect -4240 3990 -4160 4070
rect -1940 4000 -1860 4080
rect -1750 4000 -1670 4080
rect 540 3990 620 4070
rect 730 3990 810 4070
rect 2990 3990 3070 4070
rect 3180 3990 3260 4070
rect 5500 3982 5580 4060
rect 5670 3982 5750 4060
rect 5500 3980 5580 3982
rect 5670 3980 5750 3982
rect -4990 3852 -4960 3920
rect -4960 3852 -4886 3920
rect -4886 3852 -4860 3920
rect -4990 3850 -4860 3852
rect -3750 3852 -3724 3920
rect -3724 3852 -3650 3920
rect -3650 3852 -3620 3920
rect -3750 3850 -3620 3852
rect -2520 3852 -2488 3920
rect -2488 3852 -2414 3920
rect -2414 3852 -2390 3920
rect -2520 3850 -2390 3852
rect -1280 3852 -1252 3920
rect -1252 3852 -1178 3920
rect -1178 3852 -1150 3920
rect -1280 3850 -1150 3852
rect -40 3852 -16 3920
rect -16 3852 58 3920
rect 58 3852 90 3920
rect -40 3850 90 3852
rect 1190 3852 1220 3920
rect 1220 3852 1294 3920
rect 1294 3852 1320 3920
rect 1190 3850 1320 3852
rect 2430 3852 2456 3920
rect 2456 3852 2530 3920
rect 2530 3852 2560 3920
rect 2430 3850 2560 3852
rect 3660 3852 3692 3920
rect 3692 3852 3766 3920
rect 3766 3852 3790 3920
rect 3660 3850 3790 3852
rect 4900 3852 4928 3920
rect 4928 3852 5002 3920
rect 5002 3852 5030 3920
rect 4900 3850 5030 3852
rect -5720 3790 -5640 3800
rect -5510 3790 -5430 3800
rect -710 3790 -630 3800
rect -520 3790 -440 3800
rect -5720 3720 -5640 3790
rect -5510 3720 -5430 3790
rect -3250 3710 -3170 3790
rect -3010 3710 -2930 3790
rect -710 3720 -630 3790
rect -520 3720 -440 3790
rect 1750 3710 1830 3790
rect 1940 3710 2020 3790
rect 4230 3700 4310 3780
rect 4400 3700 4480 3780
rect -8810 3260 -8720 3390
rect -8600 3260 -8510 3390
rect 8500 3290 8570 3380
rect 8660 3290 8730 3380
rect -3750 3202 -3620 3270
rect -2520 3202 -2390 3260
rect -2190 3202 -2110 3270
rect -2080 3202 -2000 3270
rect -1280 3202 -1150 3260
rect -40 3202 90 3260
rect 220 3202 300 3270
rect 330 3202 410 3270
rect 1190 3202 1320 3260
rect 2430 3210 2560 3280
rect 2680 3202 2760 3280
rect 2790 3202 2870 3280
rect 3660 3202 3790 3260
rect -3750 3200 -3620 3202
rect -2520 3190 -2390 3202
rect -2190 3190 -2110 3202
rect -2080 3190 -2000 3202
rect -1280 3190 -1150 3202
rect -40 3190 90 3202
rect 220 3190 300 3202
rect 330 3190 410 3202
rect 1190 3190 1320 3202
rect 2680 3200 2760 3202
rect 2790 3200 2870 3202
rect 3660 3190 3790 3202
rect 1200 3010 1290 3020
rect 1340 3010 1430 3020
rect -3810 2920 -3720 3000
rect -3670 2920 -3580 3000
rect 1200 2940 1290 3010
rect 1340 2940 1430 3010
rect -2290 2800 -2180 2910
rect -1430 2800 -1320 2910
rect -220 2800 -110 2910
rect 630 2800 740 2910
rect -3810 2702 -3720 2770
rect -3670 2702 -3580 2770
rect 2200 2800 2310 2910
rect 3080 2800 3190 2910
rect 1200 2702 1290 2760
rect 1340 2702 1430 2760
rect -3810 2690 -3720 2702
rect -3670 2690 -3580 2702
rect 1200 2680 1290 2702
rect 1340 2680 1430 2702
rect -990 2510 -910 2530
rect -840 2510 -760 2530
rect 1490 2510 1570 2530
rect 1630 2510 1710 2530
rect -3480 2430 -3400 2510
rect -3330 2430 -3250 2510
rect -990 2450 -910 2510
rect -840 2450 -760 2510
rect 1490 2450 1570 2510
rect 1630 2450 1710 2510
rect -3030 2202 -2950 2280
rect -2920 2202 -2840 2280
rect -620 2202 -540 2250
rect 1830 2202 1910 2270
rect 1950 2202 2030 2270
rect 3030 2202 3110 2260
rect -3030 2200 -2950 2202
rect -2920 2200 -2840 2202
rect -620 2170 -540 2202
rect 1830 2190 1910 2202
rect 1950 2190 2030 2202
rect 3030 2180 3110 2202
rect -1850 2020 -1770 2100
rect 560 2020 640 2100
rect -3110 1910 -3030 1920
rect 1780 1910 1860 1920
rect -3110 1840 -3030 1910
rect 1780 1840 1860 1910
rect -3000 1700 -2890 1790
rect 1910 1700 2020 1790
rect -620 1582 -540 1630
rect 3030 1582 3110 1640
rect -620 1550 -540 1582
rect 3030 1560 3110 1582
rect -2460 1400 -2404 1480
rect -2404 1400 -2370 1480
rect -2340 1400 -2250 1480
rect -1850 1400 -1770 1480
rect -10 1400 32 1480
rect 32 1400 66 1480
rect 66 1400 80 1480
rect 110 1400 200 1480
rect 560 1400 640 1480
rect 2420 1400 2468 1490
rect 2468 1400 2502 1490
rect 2502 1400 2630 1490
rect -3110 1290 -3030 1300
rect 1780 1290 1860 1300
rect -3110 1220 -3030 1290
rect 1780 1220 1860 1290
rect -1230 982 -1140 1050
rect 3650 990 3740 1070
rect -1230 970 -1140 982
rect -2460 800 -2370 880
rect -2340 800 -2250 880
rect -10 800 80 880
rect 110 800 200 880
rect 2420 800 2510 880
rect 2540 800 2630 880
rect -3810 690 -3720 720
rect -3670 690 -3580 720
rect 1200 690 1290 720
rect 1340 690 1430 720
rect -3810 640 -3720 690
rect -3670 640 -3580 690
rect 1200 640 1290 690
rect 1340 640 1430 690
rect -3060 490 -2940 590
rect -1840 490 -1720 590
rect -630 490 -510 590
rect -1230 382 -1140 450
rect 590 490 710 590
rect 1820 480 1940 580
rect 3030 490 3150 590
rect 3650 390 3740 470
rect -1230 370 -1140 382
rect -2460 200 -2370 280
rect -2340 200 -2250 280
rect -10 200 80 280
rect 110 200 200 280
rect 2420 200 2510 280
rect 2540 200 2630 280
rect -3810 90 -3720 100
rect -3670 90 -3580 100
rect 1200 90 1290 120
rect 1340 90 1430 120
rect -3810 20 -3720 90
rect -3670 20 -3580 90
rect 1200 40 1290 90
rect 1340 40 1430 90
<< metal2 >>
rect -2620 9100 -2330 9120
rect -2620 9030 -2600 9100
rect -2510 9030 -2430 9100
rect -2340 9030 -2330 9100
rect -2620 8990 -2330 9030
rect -2620 8910 -2600 8990
rect -2520 8910 -2430 8990
rect -2350 8910 -2330 8990
rect -130 9100 160 9120
rect -130 9030 -110 9100
rect -20 9030 60 9100
rect 150 9030 160 9100
rect -130 8990 160 9030
rect -3890 8750 -3600 8870
rect -3160 8860 -3010 8910
rect -3890 8670 -3870 8750
rect -3790 8670 -3700 8750
rect -3620 8670 -3600 8750
rect -3480 8820 -3400 8830
rect -3480 8730 -3400 8740
rect -3330 8820 -3250 8830
rect -3330 8730 -3250 8740
rect -3160 8790 -3150 8860
rect -3020 8790 -3010 8860
rect -3890 8210 -3600 8670
rect -3160 8320 -3010 8790
rect -3890 8130 -3870 8210
rect -3790 8130 -3700 8210
rect -3620 8130 -3600 8210
rect -3480 8280 -3400 8290
rect -3480 8190 -3400 8200
rect -3330 8280 -3250 8290
rect -3330 8190 -3250 8200
rect -3160 8250 -3150 8320
rect -3020 8250 -3010 8320
rect -3890 7670 -3600 8130
rect -3160 7780 -3010 8250
rect -2620 8450 -2330 8910
rect -2620 8370 -2600 8450
rect -2520 8370 -2430 8450
rect -2350 8370 -2330 8450
rect -2620 8050 -2330 8370
rect -2620 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -2330 8050
rect -2620 7910 -2330 7980
rect -2620 7830 -2600 7910
rect -2520 7830 -2430 7910
rect -2350 7830 -2330 7910
rect -2620 7820 -2330 7830
rect -1920 8860 -1770 8920
rect -1920 8790 -1910 8860
rect -1780 8790 -1770 8860
rect -1920 8320 -1770 8790
rect -1920 8250 -1910 8320
rect -1780 8250 -1770 8320
rect -3890 7590 -3870 7670
rect -3790 7590 -3700 7670
rect -3620 7590 -3600 7670
rect -3480 7740 -3400 7750
rect -3480 7650 -3400 7660
rect -3330 7740 -3250 7750
rect -3330 7650 -3250 7660
rect -3160 7710 -3150 7780
rect -3020 7710 -3010 7780
rect -3890 7570 -3600 7590
rect -3160 7240 -3010 7710
rect -1920 7780 -1770 8250
rect -1920 7710 -1910 7780
rect -1780 7710 -1770 7780
rect -2590 7520 -2510 7530
rect -2590 7430 -2510 7440
rect -2420 7520 -2340 7530
rect -2420 7430 -2340 7440
rect -3160 7170 -3150 7240
rect -3020 7170 -3010 7240
rect -3890 7130 -3600 7160
rect -3890 7050 -3870 7130
rect -3790 7050 -3700 7130
rect -3620 7050 -3600 7130
rect -3890 6550 -3600 7050
rect -3890 6470 -3870 6550
rect -3790 6470 -3700 6550
rect -3620 6470 -3600 6550
rect -9940 6270 -9810 6280
rect -9940 6120 -9810 6130
rect -9690 6270 -9560 6280
rect -9690 6120 -9560 6130
rect -3890 5940 -3600 6470
rect -3160 6660 -3010 7170
rect -3160 6590 -3150 6660
rect -3020 6590 -3010 6660
rect -3160 6080 -3010 6590
rect -2610 7390 -2320 7430
rect -2610 7310 -2590 7390
rect -2510 7310 -2420 7390
rect -2340 7310 -2320 7390
rect -2610 6810 -2320 7310
rect -1920 7240 -1770 7710
rect -1370 8750 -1080 8950
rect -130 8910 -110 8990
rect -30 8910 60 8990
rect 140 8910 160 8990
rect 2330 9110 2620 9150
rect 2330 9030 2350 9110
rect 2430 9030 2520 9110
rect 2600 9030 2620 9110
rect 2330 8980 2620 9030
rect -690 8860 -540 8910
rect -1370 8670 -1350 8750
rect -1270 8670 -1180 8750
rect -1100 8670 -1080 8750
rect -990 8820 -910 8830
rect -990 8730 -910 8740
rect -840 8820 -760 8830
rect -840 8730 -760 8740
rect -690 8790 -680 8860
rect -550 8790 -540 8860
rect -1370 8210 -1080 8670
rect -690 8320 -540 8790
rect -1370 8130 -1350 8210
rect -1270 8130 -1180 8210
rect -1100 8130 -1080 8210
rect -990 8280 -910 8290
rect -990 8190 -910 8200
rect -840 8280 -760 8290
rect -840 8190 -760 8200
rect -690 8250 -680 8320
rect -550 8250 -540 8320
rect -1370 7670 -1080 8130
rect -690 7780 -540 8250
rect -130 8450 160 8910
rect -130 8370 -110 8450
rect -30 8370 60 8450
rect 140 8370 160 8450
rect -130 8060 160 8370
rect -130 8050 50 8060
rect -130 7980 -110 8050
rect -20 7990 50 8050
rect 140 7990 160 8060
rect -20 7980 160 7990
rect -130 7920 160 7980
rect -130 7840 -110 7920
rect -30 7840 60 7920
rect 140 7840 160 7920
rect -130 7820 160 7840
rect 550 8860 700 8910
rect 550 8790 560 8860
rect 690 8790 700 8860
rect 550 8320 700 8790
rect 550 8250 560 8320
rect 690 8250 700 8320
rect -1370 7590 -1350 7670
rect -1270 7590 -1180 7670
rect -1100 7590 -1080 7670
rect -990 7740 -910 7750
rect -990 7650 -910 7660
rect -840 7740 -760 7750
rect -840 7650 -760 7660
rect -690 7710 -680 7780
rect -550 7710 -540 7780
rect -1370 7560 -1080 7590
rect -1920 7170 -1910 7240
rect -1780 7170 -1770 7240
rect -690 7240 -540 7710
rect 550 7780 700 8250
rect 550 7710 560 7780
rect 690 7710 700 7780
rect -110 7520 -30 7530
rect 60 7520 140 7530
rect -2190 7140 -2110 7150
rect -2190 7050 -2110 7060
rect -2080 7140 -2000 7150
rect -2080 7050 -2000 7060
rect -2610 6730 -2590 6810
rect -2510 6730 -2420 6810
rect -2340 6730 -2320 6810
rect -2610 6360 -2320 6730
rect -1920 6660 -1770 7170
rect -1920 6590 -1910 6660
rect -1780 6590 -1770 6660
rect -2190 6530 -2110 6540
rect -2190 6440 -2110 6450
rect -2080 6530 -2000 6540
rect -2080 6440 -2000 6450
rect -2610 6280 -2590 6360
rect -2500 6280 -2430 6360
rect -2340 6280 -2320 6360
rect -2610 6230 -2320 6280
rect -2610 6150 -2590 6230
rect -2510 6150 -2420 6230
rect -2340 6150 -2320 6230
rect -1920 6170 -1770 6590
rect -1388 7130 -1056 7180
rect -1388 7050 -1360 7130
rect -1280 7050 -1190 7130
rect -1110 7050 -1056 7130
rect -1388 6550 -1056 7050
rect -1388 6470 -1360 6550
rect -1280 6470 -1190 6550
rect -1110 6470 -1056 6550
rect -2610 6130 -2320 6150
rect -3160 6010 -3150 6080
rect -3020 6010 -3010 6080
rect -3160 5970 -3010 6010
rect -1388 5970 -1056 6470
rect -690 7170 -680 7240
rect -550 7170 -540 7240
rect -690 6660 -540 7170
rect -690 6590 -670 6660
rect -690 6080 -540 6590
rect -130 7400 160 7440
rect -130 7320 -110 7400
rect -30 7320 60 7400
rect 140 7320 160 7400
rect -130 6820 160 7320
rect 550 7240 700 7710
rect 1120 8750 1410 8950
rect 2330 8900 2350 8980
rect 2430 8900 2520 8980
rect 2600 8900 2620 8980
rect 1790 8860 1940 8900
rect 1120 8670 1140 8750
rect 1220 8670 1310 8750
rect 1390 8670 1410 8750
rect 1490 8820 1570 8830
rect 1490 8730 1570 8740
rect 1640 8820 1720 8830
rect 1640 8730 1720 8740
rect 1790 8790 1800 8860
rect 1930 8790 1940 8860
rect 1120 8210 1410 8670
rect 1790 8570 1940 8790
rect 1780 8320 1940 8570
rect 1120 8130 1140 8210
rect 1220 8130 1310 8210
rect 1390 8130 1410 8210
rect 1490 8280 1570 8290
rect 1490 8190 1570 8200
rect 1640 8280 1720 8290
rect 1640 8190 1720 8200
rect 1780 8250 1800 8320
rect 1930 8250 1940 8320
rect 1120 7660 1410 8130
rect 1780 7780 1940 8250
rect 1120 7580 1140 7660
rect 1220 7580 1310 7660
rect 1390 7580 1410 7660
rect 1500 7740 1580 7750
rect 1500 7650 1580 7660
rect 1640 7740 1720 7750
rect 1640 7650 1720 7660
rect 1780 7710 1800 7780
rect 1930 7710 1940 7780
rect 1780 7670 1940 7710
rect 2330 8440 2620 8900
rect 2330 8360 2350 8440
rect 2430 8360 2520 8440
rect 2600 8360 2620 8440
rect 2330 8060 2620 8360
rect 2330 7990 2350 8060
rect 2430 7990 2520 8060
rect 2600 7990 2620 8060
rect 2330 7900 2620 7990
rect 2330 7820 2350 7900
rect 2430 7820 2520 7900
rect 2600 7820 2620 7900
rect 1120 7560 1410 7580
rect 550 7170 560 7240
rect 690 7170 700 7240
rect 1780 7240 1930 7670
rect 2330 7570 2620 7820
rect 3020 8860 3170 8890
rect 3020 8790 3030 8860
rect 3160 8790 3170 8860
rect 3020 8320 3170 8790
rect 3020 8250 3030 8320
rect 3160 8250 3170 8320
rect 3020 7780 3170 8250
rect 3020 7710 3030 7780
rect 3160 7710 3170 7780
rect 2350 7520 2430 7530
rect 2520 7520 2600 7530
rect 1780 7170 1790 7240
rect 1920 7170 1930 7240
rect 220 7140 300 7150
rect 220 7050 300 7060
rect 330 7140 410 7150
rect 330 7050 410 7060
rect -130 6740 -110 6820
rect -30 6740 60 6820
rect 140 6740 160 6820
rect -130 6350 160 6740
rect 550 6660 700 7170
rect 550 6590 560 6660
rect 690 6590 700 6660
rect 220 6550 300 6560
rect 220 6460 300 6470
rect 330 6550 410 6560
rect 330 6460 410 6470
rect -130 6280 -110 6350
rect -30 6280 60 6350
rect 140 6280 160 6350
rect -130 6240 160 6280
rect -130 6160 -110 6240
rect -30 6160 60 6240
rect 140 6160 160 6240
rect -130 6140 160 6160
rect -690 6010 -680 6080
rect -550 6010 -540 6080
rect -690 5980 -540 6010
rect 550 6080 700 6590
rect 550 6010 560 6080
rect 690 6010 700 6080
rect 550 5980 700 6010
rect 1110 7130 1400 7170
rect 1110 7050 1130 7130
rect 1210 7050 1300 7130
rect 1380 7050 1400 7130
rect 1110 6540 1400 7050
rect 1110 6460 1130 6540
rect 1210 6460 1300 6540
rect 1380 6460 1400 6540
rect -5720 5790 -5430 5870
rect -3810 5860 -3680 5940
rect -3890 5850 -3810 5860
rect -3680 5850 -3600 5860
rect -1388 5890 -1360 5970
rect -1280 5890 -1190 5970
rect -1110 5890 -1056 5970
rect -1388 5832 -1056 5890
rect 220 5970 300 5980
rect 220 5880 300 5890
rect 330 5970 410 5980
rect 330 5880 410 5890
rect 1110 5970 1400 6460
rect 1780 6660 1930 7170
rect 1780 6590 1790 6660
rect 1920 6590 1930 6660
rect 1780 6080 1930 6590
rect 2330 7390 2620 7440
rect 2330 7310 2350 7390
rect 2430 7310 2520 7390
rect 2600 7310 2620 7390
rect 2330 6810 2620 7310
rect 3020 7240 3170 7710
rect 3570 8750 3860 9020
rect 3570 8670 3590 8750
rect 3670 8670 3760 8750
rect 3840 8670 3860 8750
rect 3570 8200 3860 8670
rect 3570 8120 3590 8200
rect 3670 8120 3760 8200
rect 3840 8120 3860 8200
rect 3570 7670 3860 8120
rect 3570 7590 3590 7670
rect 3670 7590 3760 7670
rect 3840 7590 3860 7670
rect 3570 7580 3860 7590
rect 3020 7170 3030 7240
rect 3160 7170 3170 7240
rect 2680 7130 2760 7140
rect 2680 7040 2760 7050
rect 2790 7130 2870 7140
rect 2790 7040 2870 7050
rect 2330 6730 2350 6810
rect 2430 6730 2520 6810
rect 2600 6730 2620 6810
rect 2330 6350 2620 6730
rect 3020 6660 3170 7170
rect 3020 6590 3030 6660
rect 3160 6590 3170 6660
rect 2680 6550 2760 6560
rect 2680 6460 2760 6470
rect 2790 6550 2870 6560
rect 2790 6460 2870 6470
rect 2330 6280 2350 6350
rect 2430 6280 2520 6350
rect 2600 6280 2620 6350
rect 2330 6230 2620 6280
rect 2330 6150 2350 6230
rect 2430 6150 2520 6230
rect 2600 6150 2620 6230
rect 2330 6140 2620 6150
rect 1780 6010 1790 6080
rect 1920 6010 1930 6080
rect 1780 5970 1930 6010
rect 3020 6080 3170 6590
rect 3020 6010 3030 6080
rect 3160 6010 3170 6080
rect 3020 5980 3170 6010
rect 3600 7130 3890 7220
rect 3600 7050 3620 7130
rect 3700 7050 3790 7130
rect 3870 7050 3890 7130
rect 3600 6550 3890 7050
rect 3600 6470 3620 6550
rect 3700 6470 3790 6550
rect 3870 6470 3890 6550
rect 2680 5970 2760 5980
rect 1110 5890 1130 5970
rect 1210 5890 1300 5970
rect 1380 5890 1400 5970
rect 1110 5870 1400 5890
rect 2680 5880 2760 5890
rect 2790 5970 2870 5980
rect 2790 5880 2870 5890
rect 3600 5970 3890 6470
rect 9560 6440 9690 6450
rect 9560 6290 9690 6300
rect 9820 6440 9950 6450
rect 9820 6290 9950 6300
rect 3600 5890 3620 5970
rect 3700 5890 3790 5970
rect 3870 5890 3890 5970
rect 3600 5870 3890 5890
rect -5720 5680 -5700 5790
rect -5610 5680 -5540 5790
rect -5450 5680 -5430 5790
rect 4210 5740 4500 5780
rect -5720 5420 -5430 5680
rect -4470 5700 -4160 5720
rect -4390 5620 -4240 5700
rect -5640 5340 -5510 5420
rect -5720 4880 -5430 5340
rect -5640 4800 -5510 4880
rect -5720 4340 -5430 4800
rect -5640 4260 -5510 4340
rect -5720 3800 -5430 4260
rect -5000 5540 -4850 5570
rect -5000 5470 -4990 5540
rect -4860 5470 -4850 5540
rect -5000 5010 -4850 5470
rect -5000 4940 -4990 5010
rect -4860 4940 -4850 5010
rect -5000 4460 -4850 4940
rect -5000 4390 -4990 4460
rect -4860 4390 -4850 4460
rect -5000 3920 -4850 4390
rect -4470 5280 -4160 5620
rect -1940 5690 -1650 5720
rect -1940 5610 -1920 5690
rect -1840 5610 -1750 5690
rect -1670 5610 -1650 5690
rect -4470 5200 -4450 5280
rect -4360 5200 -4270 5280
rect -4180 5200 -4160 5280
rect -4470 5160 -4160 5200
rect -4390 5080 -4240 5160
rect -4470 4620 -4160 5080
rect -4390 4540 -4240 4620
rect -4470 4210 -4160 4540
rect -4470 4200 -4270 4210
rect -4470 4120 -4450 4200
rect -4360 4130 -4270 4200
rect -4180 4130 -4160 4210
rect -4360 4120 -4160 4130
rect -4470 4070 -4160 4120
rect -4390 3990 -4240 4070
rect -4470 3980 -4160 3990
rect -3760 5540 -3610 5580
rect -3760 5470 -3750 5540
rect -3620 5470 -3610 5540
rect -3760 5000 -3610 5470
rect -2530 5540 -2380 5570
rect -2530 5470 -2520 5540
rect -2390 5470 -2380 5540
rect -3760 4930 -3750 5000
rect -3620 4930 -3610 5000
rect -3760 4460 -3610 4930
rect -3760 4390 -3750 4460
rect -3620 4390 -3610 4460
rect -5000 3850 -4990 3920
rect -4860 3850 -4850 3920
rect -5000 3810 -4850 3850
rect -3760 3920 -3610 4390
rect -3760 3850 -3750 3920
rect -3620 3850 -3610 3920
rect -5640 3720 -5510 3800
rect -5720 3710 -5430 3720
rect -8810 3390 -8720 3400
rect -8810 3250 -8720 3260
rect -8600 3390 -8510 3400
rect -8600 3250 -8510 3260
rect -3760 3270 -3610 3850
rect -3250 5420 -2930 5450
rect -3250 5340 -3240 5420
rect -3160 5340 -3020 5420
rect -2940 5340 -2930 5420
rect -3250 4880 -2930 5340
rect -3250 4800 -3240 4880
rect -3160 4800 -3020 4880
rect -2940 4800 -2930 4880
rect -3250 4340 -2930 4800
rect -3170 4260 -3010 4340
rect -3250 3870 -2930 4260
rect -2530 5000 -2380 5470
rect -2530 4930 -2520 5000
rect -2390 4930 -2380 5000
rect -2530 4460 -2380 4930
rect -2530 4390 -2520 4460
rect -2390 4390 -2380 4460
rect -2530 3920 -2380 4390
rect -1940 5280 -1650 5610
rect 530 5690 820 5730
rect 530 5610 540 5690
rect 620 5610 730 5690
rect 810 5610 820 5690
rect -1940 5200 -1920 5280
rect -1830 5200 -1760 5280
rect -1670 5200 -1650 5280
rect -1940 5160 -1650 5200
rect -1940 5150 -1750 5160
rect -1940 5070 -1920 5150
rect -1840 5080 -1750 5150
rect -1670 5080 -1650 5160
rect -1840 5070 -1650 5080
rect -1940 4610 -1650 5070
rect -1940 4530 -1930 4610
rect -1850 4530 -1760 4610
rect -1680 4530 -1650 4610
rect -1940 4200 -1650 4530
rect -1940 4120 -1920 4200
rect -1830 4120 -1760 4200
rect -1670 4120 -1650 4200
rect -1940 4080 -1650 4120
rect -1860 4000 -1750 4080
rect -1670 4000 -1650 4080
rect -1940 3970 -1650 4000
rect -1290 5540 -1140 5570
rect -1290 5470 -1280 5540
rect -1150 5470 -1140 5540
rect -50 5540 100 5560
rect -1290 5000 -1140 5470
rect -1290 4930 -1280 5000
rect -1150 4930 -1140 5000
rect -1290 4460 -1140 4930
rect -1290 4390 -1280 4460
rect -1150 4390 -1140 4460
rect -3250 3790 -2840 3870
rect -3170 3710 -3010 3790
rect -2930 3710 -2840 3790
rect -3250 3610 -2840 3710
rect -3760 3200 -3750 3270
rect -3620 3200 -3610 3270
rect -3760 3190 -3610 3200
rect -3810 3000 -3720 3010
rect -3670 3000 -3580 3010
rect -3720 2920 -3670 2990
rect -3810 2770 -3580 2920
rect -3720 2690 -3670 2770
rect -3810 720 -3580 2690
rect -3500 2510 -3230 2520
rect -3500 2430 -3480 2510
rect -3400 2430 -3330 2510
rect -3250 2430 -3230 2510
rect -3480 2420 -3400 2430
rect -3330 2420 -3250 2430
rect -3030 2310 -2840 3610
rect -2530 3850 -2520 3920
rect -2390 3850 -2380 3920
rect -2530 3260 -2380 3850
rect -1290 3920 -1140 4390
rect -1290 3850 -1280 3920
rect -1150 3850 -1140 3920
rect -2530 3190 -2520 3260
rect -2390 3190 -2380 3260
rect -2530 3140 -2380 3190
rect -2190 3270 -2110 3280
rect -2190 3180 -2110 3190
rect -2080 3270 -2000 3280
rect -2080 3180 -2000 3190
rect -1290 3260 -1140 3850
rect -1290 3190 -1280 3260
rect -1150 3190 -1140 3260
rect -1290 3100 -1140 3190
rect -720 5420 -430 5510
rect -720 5340 -710 5420
rect -630 5340 -530 5420
rect -450 5340 -430 5420
rect -720 4880 -430 5340
rect -720 4800 -710 4880
rect -630 4800 -520 4880
rect -440 4800 -430 4880
rect -720 4340 -430 4800
rect -720 4260 -710 4340
rect -630 4260 -530 4340
rect -450 4260 -430 4340
rect -720 3800 -430 4260
rect -720 3720 -710 3800
rect -630 3720 -520 3800
rect -440 3720 -430 3800
rect -2290 2910 -2180 2920
rect -2290 2790 -2180 2800
rect -1430 2910 -1320 2920
rect -1430 2790 -1320 2800
rect -990 2530 -910 2540
rect -990 2440 -910 2450
rect -840 2530 -760 2540
rect -840 2440 -760 2450
rect -3120 2280 -2810 2310
rect -3120 2200 -3030 2280
rect -2950 2200 -2920 2280
rect -2840 2200 -2810 2280
rect -720 2250 -430 3720
rect -50 5470 -40 5540
rect 90 5470 100 5540
rect -50 5000 100 5470
rect -50 4930 -40 5000
rect 90 4930 100 5000
rect -50 4460 100 4930
rect -50 4390 -40 4460
rect 90 4390 100 4460
rect -50 3920 100 4390
rect 530 5280 820 5610
rect 2980 5690 3270 5720
rect 2980 5610 2990 5690
rect 3070 5610 3180 5690
rect 3260 5610 3270 5690
rect 530 5200 550 5280
rect 640 5200 710 5280
rect 800 5200 820 5280
rect 530 5160 820 5200
rect 530 5080 540 5160
rect 620 5080 730 5160
rect 810 5080 820 5160
rect 530 4610 820 5080
rect 530 4530 540 4610
rect 620 4530 720 4610
rect 800 4530 820 4610
rect 530 4200 820 4530
rect 530 4120 550 4200
rect 640 4120 710 4200
rect 800 4120 820 4200
rect 530 4070 820 4120
rect 530 3990 540 4070
rect 620 3990 730 4070
rect 810 3990 820 4070
rect 530 3980 820 3990
rect 1180 5540 1330 5570
rect 1180 5470 1190 5540
rect 1320 5470 1330 5540
rect 2420 5540 2570 5590
rect 1180 5000 1330 5470
rect 1180 4930 1190 5000
rect 1320 4930 1330 5000
rect 1180 4460 1330 4930
rect 1180 4390 1190 4460
rect 1320 4390 1330 4460
rect -50 3850 -40 3920
rect 90 3850 100 3920
rect -50 3260 100 3850
rect 1180 3920 1330 4390
rect 1180 3850 1190 3920
rect 1320 3850 1330 3920
rect -50 3190 -40 3260
rect 90 3190 100 3260
rect -50 3120 100 3190
rect 220 3270 300 3280
rect 220 3180 300 3190
rect 330 3270 410 3280
rect 330 3180 410 3190
rect 1180 3260 1330 3850
rect 1740 5410 2030 5510
rect 1740 5330 1750 5410
rect 1830 5330 1930 5410
rect 2010 5330 2030 5410
rect 1740 4870 2030 5330
rect 1740 4790 1750 4870
rect 1830 4790 1930 4870
rect 2010 4790 2030 4870
rect 1740 4330 2030 4790
rect 1740 4250 1760 4330
rect 1840 4250 1930 4330
rect 2010 4250 2030 4330
rect 1740 3890 2030 4250
rect 2420 5470 2430 5540
rect 2560 5470 2570 5540
rect 2420 5000 2570 5470
rect 2420 4930 2430 5000
rect 2560 4930 2570 5000
rect 2420 4460 2570 4930
rect 2420 4390 2430 4460
rect 2560 4390 2570 4460
rect 2420 3920 2570 4390
rect 1740 3790 2040 3890
rect 1740 3710 1750 3790
rect 1830 3710 1940 3790
rect 2020 3710 2040 3790
rect 1740 3690 2040 3710
rect 1180 3190 1190 3260
rect 1320 3190 1330 3260
rect 1180 3180 1330 3190
rect 1200 3020 1290 3030
rect 1340 3020 1430 3030
rect 1290 2940 1340 3020
rect -220 2910 -110 2920
rect -220 2790 -110 2800
rect 630 2910 740 2920
rect 630 2790 740 2800
rect -720 2200 -620 2250
rect -3120 2180 -2810 2200
rect -540 2200 -430 2250
rect 1200 2760 1430 2940
rect 1290 2680 1340 2760
rect -1850 2100 -1770 2130
rect -3110 1920 -3030 1950
rect -3110 1830 -3030 1840
rect -3110 1790 -2850 1830
rect -3110 1700 -3000 1790
rect -2890 1700 -2850 1790
rect -3110 1660 -2850 1700
rect -3110 1300 -3030 1660
rect -3110 1210 -3030 1220
rect -2460 1480 -2250 1500
rect -2370 1400 -2340 1480
rect -3720 640 -3670 720
rect -3810 100 -3580 640
rect -2460 880 -2250 1400
rect -1850 1480 -1770 2020
rect -620 1630 -540 2170
rect -620 1540 -540 1550
rect 560 2100 640 2130
rect -1850 1390 -1770 1400
rect -10 1480 200 1500
rect 80 1400 110 1480
rect -2370 800 -2340 880
rect -3060 590 -2940 600
rect -3060 480 -2940 490
rect -2460 280 -2250 800
rect -1230 1050 -1140 1080
rect -1840 590 -1720 600
rect -1840 480 -1720 490
rect -1230 450 -1140 970
rect -10 880 200 1400
rect 560 1480 640 2020
rect 560 1390 640 1400
rect 80 800 110 880
rect -630 590 -510 600
rect -630 480 -510 490
rect -1230 360 -1140 370
rect -2370 200 -2340 280
rect -2460 190 -2250 200
rect -10 280 200 800
rect 1200 720 1430 2680
rect 1490 2530 1570 2540
rect 1490 2440 1570 2450
rect 1630 2530 1710 2540
rect 1630 2440 1710 2450
rect 1820 2270 2040 3690
rect 2420 3850 2430 3920
rect 2560 3850 2570 3920
rect 2420 3280 2570 3850
rect 2980 5280 3270 5610
rect 4210 5660 4230 5740
rect 4310 5660 4400 5740
rect 4480 5660 4500 5740
rect 2980 5200 3000 5280
rect 3090 5200 3160 5280
rect 3250 5200 3270 5280
rect 2980 5150 3270 5200
rect 2980 5070 2990 5150
rect 3070 5070 3180 5150
rect 3260 5070 3270 5150
rect 2980 4610 3270 5070
rect 2980 4530 2990 4610
rect 3070 4530 3180 4610
rect 3260 4530 3270 4610
rect 2980 4200 3270 4530
rect 2980 4120 3000 4200
rect 3090 4120 3160 4200
rect 3250 4120 3270 4200
rect 2980 4070 3270 4120
rect 2980 3990 2990 4070
rect 3070 3990 3180 4070
rect 3260 3990 3270 4070
rect 2980 3740 3270 3990
rect 3650 5540 3800 5580
rect 3650 5470 3660 5540
rect 3790 5470 3800 5540
rect 3650 5000 3800 5470
rect 3650 4930 3660 5000
rect 3790 4930 3800 5000
rect 3650 4460 3800 4930
rect 3650 4390 3660 4460
rect 3790 4390 3800 4460
rect 3650 3920 3800 4390
rect 3650 3850 3660 3920
rect 3790 3850 3800 3920
rect 2420 3210 2430 3280
rect 2560 3210 2570 3280
rect 2420 3150 2570 3210
rect 2680 3280 2760 3290
rect 2680 3190 2760 3200
rect 2790 3280 2870 3290
rect 2790 3190 2870 3200
rect 3650 3260 3800 3850
rect 4210 5410 4500 5660
rect 5480 5690 5770 5710
rect 5480 5610 5500 5690
rect 5580 5610 5670 5690
rect 5750 5610 5770 5690
rect 4210 5330 4230 5410
rect 4310 5330 4400 5410
rect 4480 5330 4500 5410
rect 4210 4870 4500 5330
rect 4210 4790 4230 4870
rect 4310 4790 4400 4870
rect 4480 4790 4500 4870
rect 4210 4330 4500 4790
rect 4210 4250 4230 4330
rect 4310 4250 4400 4330
rect 4480 4250 4500 4330
rect 4210 3780 4500 4250
rect 4890 5540 5040 5580
rect 4890 5470 4900 5540
rect 5030 5470 5040 5540
rect 4890 5000 5040 5470
rect 4890 4930 4900 5000
rect 5030 4930 5040 5000
rect 4890 4460 5040 4930
rect 4890 4390 4900 4460
rect 5030 4390 5040 4460
rect 4890 3920 5040 4390
rect 5480 5280 5770 5610
rect 5480 5200 5500 5280
rect 5590 5200 5660 5280
rect 5750 5200 5770 5280
rect 5480 5150 5770 5200
rect 5480 5070 5500 5150
rect 5580 5070 5670 5150
rect 5750 5070 5770 5150
rect 5480 4610 5770 5070
rect 5480 4530 5500 4610
rect 5580 4530 5670 4610
rect 5750 4530 5770 4610
rect 5480 4200 5770 4530
rect 5480 4120 5500 4200
rect 5590 4120 5660 4200
rect 5750 4120 5770 4200
rect 5480 4060 5770 4120
rect 5480 3980 5500 4060
rect 5580 3980 5670 4060
rect 5750 3980 5770 4060
rect 5480 3960 5770 3980
rect 4890 3850 4900 3920
rect 5030 3850 5040 3920
rect 4890 3820 5040 3850
rect 4210 3700 4230 3780
rect 4310 3700 4400 3780
rect 4480 3700 4500 3780
rect 4210 3690 4500 3700
rect 8500 3380 8570 3390
rect 8500 3280 8570 3290
rect 8660 3380 8730 3390
rect 8660 3280 8730 3290
rect 3650 3190 3660 3260
rect 3790 3190 3800 3260
rect 3650 3150 3800 3190
rect 2200 2910 2310 2920
rect 2200 2790 2310 2800
rect 3080 2910 3190 2920
rect 3080 2790 3190 2800
rect 1820 2190 1830 2270
rect 1910 2190 1950 2270
rect 2030 2190 2040 2270
rect 2980 2260 3270 2270
rect 2980 2220 3030 2260
rect 1820 2180 2040 2190
rect 3110 2220 3270 2260
rect 1780 1920 1860 1950
rect 1780 1830 1860 1840
rect 1780 1790 2050 1830
rect 1780 1700 1910 1790
rect 2020 1700 2050 1790
rect 1780 1660 2050 1700
rect 1780 1300 1860 1660
rect 3030 1640 3110 2180
rect 3030 1550 3110 1560
rect 2410 1490 2640 1500
rect 2410 1400 2420 1490
rect 2630 1400 2640 1490
rect 2410 1390 2640 1400
rect 1780 1210 1860 1220
rect 1290 640 1340 720
rect 590 590 710 600
rect 590 480 710 490
rect 80 200 110 280
rect -10 190 200 200
rect -3720 20 -3670 100
rect 1200 120 1430 640
rect 2420 880 2630 1390
rect 2510 800 2540 880
rect 1820 580 1940 590
rect 1820 470 1940 480
rect 2420 280 2630 800
rect 3650 1070 3740 1100
rect 3030 590 3150 600
rect 3030 480 3150 490
rect 3650 470 3740 990
rect 3650 380 3740 390
rect 2510 200 2540 280
rect 2420 190 2630 200
rect 1290 40 1340 120
rect 1200 30 1430 40
rect -3810 10 -3580 20
<< via2 >>
rect -2600 9030 -2510 9100
rect -2430 9030 -2340 9100
rect -110 9030 -20 9100
rect 60 9030 150 9100
rect -3480 8740 -3400 8820
rect -3330 8740 -3250 8820
rect -3480 8200 -3400 8280
rect -3330 8200 -3250 8280
rect -2590 7980 -2500 8050
rect -2450 7980 -2360 8050
rect -3480 7660 -3400 7740
rect -3330 7660 -3250 7740
rect -2590 7440 -2510 7520
rect -2420 7440 -2340 7520
rect -9940 6130 -9810 6270
rect -9690 6130 -9560 6270
rect 2350 9030 2430 9110
rect 2520 9030 2600 9110
rect -990 8740 -910 8820
rect -840 8740 -760 8820
rect -990 8200 -910 8280
rect -840 8200 -760 8280
rect -110 7980 -20 8050
rect 50 7990 140 8060
rect -990 7660 -910 7740
rect -840 7660 -760 7740
rect -110 7440 -30 7520
rect 60 7440 140 7520
rect -2190 7060 -2110 7140
rect -2080 7060 -2000 7140
rect -2190 6450 -2110 6530
rect -2080 6450 -2000 6530
rect -2590 6280 -2500 6360
rect -2430 6280 -2340 6360
rect 1490 8740 1570 8820
rect 1640 8740 1720 8820
rect 1490 8200 1570 8280
rect 1640 8200 1720 8280
rect 1500 7660 1580 7740
rect 1640 7660 1720 7740
rect 2350 7990 2430 8060
rect 2520 7990 2600 8060
rect 2350 7440 2430 7520
rect 2520 7440 2600 7520
rect 220 7060 300 7140
rect 330 7060 410 7140
rect 220 6470 300 6550
rect 330 6470 410 6550
rect -110 6280 -30 6350
rect 60 6280 140 6350
rect 220 5890 300 5970
rect 330 5890 410 5970
rect 2680 7050 2760 7130
rect 2790 7050 2870 7130
rect 2680 6470 2760 6550
rect 2790 6470 2870 6550
rect 2350 6280 2430 6350
rect 2520 6280 2600 6350
rect 2680 5890 2760 5970
rect 2790 5890 2870 5970
rect 9560 6300 9690 6440
rect 9820 6300 9950 6440
rect -5700 5680 -5610 5790
rect -5540 5680 -5450 5790
rect -4450 5200 -4360 5280
rect -4270 5200 -4180 5280
rect -4450 4120 -4360 4200
rect -4270 4130 -4180 4210
rect -8810 3260 -8720 3390
rect -8600 3260 -8510 3390
rect -1920 5200 -1830 5280
rect -1760 5200 -1670 5280
rect -1920 4120 -1830 4200
rect -1760 4120 -1670 4200
rect -3480 2430 -3400 2510
rect -3330 2430 -3250 2510
rect -2190 3190 -2110 3270
rect -2080 3190 -2000 3270
rect -2290 2800 -2180 2910
rect -1430 2800 -1320 2910
rect -990 2450 -910 2530
rect -840 2450 -760 2530
rect 550 5200 640 5280
rect 710 5200 800 5280
rect 550 4120 640 4200
rect 710 4120 800 4200
rect 220 3190 300 3270
rect 330 3190 410 3270
rect -220 2800 -110 2910
rect 630 2800 740 2910
rect -3000 1700 -2890 1790
rect -3060 490 -2940 590
rect -1840 490 -1720 590
rect -630 490 -510 590
rect 1490 2450 1570 2530
rect 1630 2450 1710 2530
rect 4230 5660 4310 5740
rect 4400 5660 4480 5740
rect 3000 5200 3090 5280
rect 3160 5200 3250 5280
rect 3000 4120 3090 4200
rect 3160 4120 3250 4200
rect 2680 3200 2760 3280
rect 2790 3200 2870 3280
rect 5500 5200 5590 5280
rect 5660 5200 5750 5280
rect 5500 4120 5590 4200
rect 5660 4120 5750 4200
rect 8500 3290 8570 3380
rect 8660 3290 8730 3380
rect 2200 2800 2310 2910
rect 3080 2800 3190 2910
rect 1910 1700 2020 1790
rect 590 490 710 590
rect 3030 490 3150 590
<< metal3 >>
rect -9960 13130 -9520 13180
rect -9960 13000 -9930 13130
rect -9830 13000 -9670 13130
rect -9570 13000 -9520 13130
rect 9540 13130 9970 13190
rect -9960 6270 -9520 13000
rect -7400 13059 -4000 13079
rect -7400 12995 -7372 13059
rect -4028 12995 -4000 13059
rect -7400 9580 -4000 12995
rect -3600 13059 -200 13079
rect -3600 12995 -3572 13059
rect -228 12995 -200 13059
rect -3600 9580 -200 12995
rect 200 13059 3600 13079
rect 200 12995 228 13059
rect 3572 12995 3600 13059
rect 200 9580 3600 12995
rect 4000 13059 7400 13079
rect 4000 12995 4028 13059
rect 7372 12995 7400 13059
rect 4000 9580 7400 12995
rect 9540 13000 9560 13130
rect 9670 13000 9820 13130
rect 9930 13000 9970 13130
rect -4650 9110 6930 9350
rect -4650 9100 2350 9110
rect -4650 9030 -2600 9100
rect -2510 9030 -2430 9100
rect -2340 9030 -110 9100
rect -20 9030 60 9100
rect 150 9030 2350 9100
rect 2430 9030 2520 9110
rect 2600 9030 6930 9110
rect -4650 8990 6930 9030
rect -3500 8820 -3230 8840
rect -3500 8740 -3480 8820
rect -3400 8740 -3330 8820
rect -3250 8740 -3230 8820
rect -3500 8720 -3230 8740
rect -1010 8820 -740 8830
rect -1010 8740 -990 8820
rect -910 8740 -840 8820
rect -760 8740 -740 8820
rect -1010 8720 -740 8740
rect 1470 8820 1740 8840
rect 1470 8740 1490 8820
rect 1570 8740 1640 8820
rect 1720 8740 1740 8820
rect 1470 8720 1740 8740
rect -3500 8280 -3230 8300
rect -3500 8200 -3480 8280
rect -3400 8200 -3330 8280
rect -3250 8200 -3230 8280
rect -3500 8180 -3230 8200
rect -1010 8280 -740 8290
rect -1010 8200 -990 8280
rect -910 8200 -840 8280
rect -760 8200 -740 8280
rect -1010 8180 -740 8200
rect 1470 8280 1740 8300
rect 1470 8200 1490 8280
rect 1570 8200 1640 8280
rect 1720 8200 1740 8280
rect 1470 8180 1740 8200
rect 6520 8120 6930 8990
rect -4890 8060 6930 8120
rect -4890 8050 50 8060
rect -4890 7980 -2590 8050
rect -2500 7980 -2450 8050
rect -2360 7980 -110 8050
rect -20 7990 50 8050
rect 140 7990 2350 8060
rect 2430 7990 2520 8060
rect 2600 7990 6930 8060
rect -20 7980 6930 7990
rect -4890 7890 6930 7980
rect -3500 7740 -3230 7770
rect -3500 7660 -3480 7740
rect -3400 7660 -3330 7740
rect -3250 7660 -3230 7740
rect -3500 7640 -3230 7660
rect -1010 7740 -740 7750
rect -1010 7660 -990 7740
rect -910 7660 -840 7740
rect -760 7660 -740 7740
rect -1010 7640 -740 7660
rect 1470 7740 1740 7770
rect 1470 7660 1500 7740
rect 1580 7660 1640 7740
rect 1720 7660 1740 7740
rect 1470 7640 1740 7660
rect 6520 7530 6930 7890
rect -4500 7520 6930 7530
rect -4500 7440 -2590 7520
rect -2510 7440 -2420 7520
rect -2340 7440 -110 7520
rect -30 7440 60 7520
rect 140 7440 2350 7520
rect 2430 7440 2520 7520
rect 2600 7440 6930 7520
rect -4500 7310 6930 7440
rect -2210 7140 -1980 7160
rect -2210 7060 -2190 7140
rect -2110 7060 -2080 7140
rect -2000 7060 -1980 7140
rect -2210 7030 -1980 7060
rect 200 7140 430 7160
rect 200 7060 220 7140
rect 300 7060 330 7140
rect 410 7060 430 7140
rect 200 7050 430 7060
rect 2660 7130 2890 7140
rect 2660 7050 2680 7130
rect 2760 7050 2790 7130
rect 2870 7050 2890 7130
rect 2660 7030 2890 7050
rect 200 6550 430 6560
rect -2210 6530 -1980 6540
rect -2210 6450 -2190 6530
rect -2110 6450 -2080 6530
rect -2000 6450 -1980 6530
rect 200 6470 220 6550
rect 300 6470 330 6550
rect 410 6470 430 6550
rect 200 6450 430 6470
rect 2660 6550 2890 6560
rect 2660 6470 2680 6550
rect 2760 6470 2790 6550
rect 2870 6470 2890 6550
rect 2660 6450 2890 6470
rect -2210 6440 -1980 6450
rect 6520 6370 6930 7310
rect -9960 6130 -9940 6270
rect -9810 6130 -9690 6270
rect -9560 6130 -9520 6270
rect -4580 6360 6930 6370
rect -4580 6280 -2590 6360
rect -2500 6280 -2430 6360
rect -2340 6350 6930 6360
rect -2340 6280 -110 6350
rect -30 6280 60 6350
rect 140 6280 2350 6350
rect 2430 6280 2520 6350
rect 2600 6280 6930 6350
rect 9540 6440 9970 13000
rect 9540 6300 9560 6440
rect 9690 6300 9820 6440
rect 9950 6300 9970 6440
rect 9540 6290 9970 6300
rect -4580 6190 6930 6280
rect -9960 6110 -9520 6130
rect -2210 5970 -1980 5990
rect -2210 5890 -2190 5970
rect -2110 5890 -2080 5970
rect -2000 5890 -1980 5970
rect -2210 5870 -1980 5890
rect 200 5970 430 5980
rect 200 5890 220 5970
rect 300 5890 330 5970
rect 410 5890 430 5970
rect 200 5870 430 5890
rect 2660 5970 2890 5980
rect 2660 5890 2680 5970
rect 2760 5890 2790 5970
rect 2870 5890 2890 5970
rect 2660 5870 2890 5890
rect -5720 5790 -5430 5810
rect -5720 5680 -5700 5790
rect -5610 5680 -5540 5790
rect -5450 5680 -5430 5790
rect -5720 5670 -5430 5680
rect 4210 5740 4502 5750
rect 4210 5660 4230 5740
rect 4310 5660 4400 5740
rect 4480 5660 4502 5740
rect 4210 5652 4502 5660
rect 6520 5460 6930 6190
rect -6730 5280 6930 5460
rect -6730 5200 -4450 5280
rect -4360 5200 -4270 5280
rect -4180 5200 -1920 5280
rect -1830 5200 -1760 5280
rect -1670 5200 550 5280
rect 640 5200 710 5280
rect 800 5200 3000 5280
rect 3090 5200 3160 5280
rect 3250 5200 5500 5280
rect 5590 5200 5660 5280
rect 5750 5200 6930 5280
rect -6730 5100 6930 5200
rect 6520 4330 6930 5100
rect -6360 4210 6930 4330
rect -6360 4200 -4270 4210
rect -6360 4120 -4450 4200
rect -4360 4130 -4270 4200
rect -4180 4200 6930 4210
rect -4180 4130 -1920 4200
rect -4360 4120 -1920 4130
rect -1830 4120 -1760 4200
rect -1670 4120 550 4200
rect 640 4120 710 4200
rect 800 4120 3000 4200
rect 3090 4120 3160 4200
rect 3250 4120 5500 4200
rect 5590 4120 5660 4200
rect 5750 4120 6930 4200
rect -6360 3990 6930 4120
rect -8830 3390 -8480 3400
rect -8830 3260 -8810 3390
rect -8720 3260 -8600 3390
rect -8510 3260 -8480 3390
rect 8490 3380 8750 3390
rect 8490 3290 8500 3380
rect 8570 3290 8660 3380
rect 8730 3290 8750 3380
rect -8830 3060 -8480 3260
rect -2210 3270 -1980 3280
rect -2210 3190 -2190 3270
rect -2110 3190 -2080 3270
rect -2000 3190 -1980 3270
rect -2210 3180 -1980 3190
rect 200 3270 430 3290
rect 200 3190 220 3270
rect 300 3190 330 3270
rect 410 3190 430 3270
rect 2660 3280 2890 3290
rect 2660 3200 2680 3280
rect 2760 3200 2790 3280
rect 2870 3200 2890 3280
rect 2660 3190 2890 3200
rect 200 3180 430 3190
rect -9330 3050 -4660 3060
rect 8490 3050 8750 3290
rect -9330 2910 9880 3050
rect -9330 2830 -2290 2910
rect -4940 2800 -2290 2830
rect -2180 2800 -1430 2910
rect -1320 2800 -220 2910
rect -110 2800 630 2910
rect 740 2800 2200 2910
rect 2310 2800 3080 2910
rect 3190 2800 9880 2910
rect -4940 2690 9880 2800
rect -4940 1990 -4660 2690
rect 4830 2680 9880 2690
rect -1010 2530 -740 2540
rect -3500 2510 -3230 2530
rect -3500 2430 -3480 2510
rect -3400 2430 -3330 2510
rect -3250 2430 -3230 2510
rect -1010 2450 -990 2530
rect -910 2450 -840 2530
rect -760 2450 -740 2530
rect -1010 2430 -740 2450
rect 1470 2530 1740 2540
rect 1470 2450 1490 2530
rect 1570 2450 1630 2530
rect 1710 2450 1740 2530
rect 1470 2430 1740 2450
rect -3500 2400 -3230 2430
rect 4900 1990 5120 2680
rect -4940 1790 5120 1990
rect -4940 1700 -3000 1790
rect -2890 1700 1910 1790
rect 2020 1700 5120 1790
rect -4940 1530 5120 1700
rect -4940 810 -4660 1530
rect 4900 810 5120 1530
rect -4940 590 5120 810
rect -4940 490 -3060 590
rect -2940 490 -1840 590
rect -1720 490 -630 590
rect -510 490 590 590
rect 710 580 3030 590
rect 710 490 1820 580
rect -4940 480 1820 490
rect 1940 490 3030 580
rect 3150 490 5120 590
rect 1940 480 5120 490
rect -4940 350 5120 480
<< via3 >>
rect -9930 13000 -9830 13130
rect -9670 13000 -9570 13130
rect -7372 12995 -4028 13059
rect -3572 12995 -228 13059
rect 228 12995 3572 13059
rect 4028 12995 7372 13059
rect 9560 13000 9670 13130
rect 9820 13000 9930 13130
rect -3480 8740 -3400 8820
rect -3330 8740 -3250 8820
rect -990 8740 -910 8820
rect -840 8740 -760 8820
rect 1490 8740 1570 8820
rect 1640 8740 1720 8820
rect -3480 8200 -3400 8280
rect -3330 8200 -3250 8280
rect -990 8200 -910 8280
rect -840 8200 -760 8280
rect 1490 8200 1570 8280
rect 1640 8200 1720 8280
rect -3480 7660 -3400 7740
rect -3330 7660 -3250 7740
rect -990 7660 -910 7740
rect -840 7660 -760 7740
rect 1500 7660 1580 7740
rect 1640 7660 1720 7740
rect -2190 7060 -2110 7140
rect -2080 7060 -2000 7140
rect 220 7060 300 7140
rect 330 7060 410 7140
rect 2680 7050 2760 7130
rect 2790 7050 2870 7130
rect -2190 6450 -2110 6530
rect -2080 6450 -2000 6530
rect 220 6470 300 6550
rect 330 6470 410 6550
rect 2680 6470 2760 6550
rect 2790 6470 2870 6550
rect -2190 5890 -2110 5970
rect -2080 5890 -2000 5970
rect 220 5890 300 5970
rect 330 5890 410 5970
rect 2680 5890 2760 5970
rect 2790 5890 2870 5970
rect -5700 5680 -5610 5790
rect -5540 5680 -5450 5790
rect 4230 5660 4310 5740
rect 4400 5660 4480 5740
rect -2190 3190 -2110 3270
rect -2080 3190 -2000 3270
rect 220 3190 300 3270
rect 330 3190 410 3270
rect 2680 3200 2760 3280
rect 2790 3200 2870 3280
rect -3480 2430 -3400 2510
rect -3330 2430 -3250 2510
rect -990 2450 -910 2530
rect -840 2450 -760 2530
rect 1490 2450 1570 2530
rect 1630 2450 1710 2530
rect 1820 480 1940 580
<< mimcap >>
rect -7300 12840 -4100 12880
rect -7300 9720 -7260 12840
rect -4140 9720 -4100 12840
rect -7300 9680 -4100 9720
rect -3500 12840 -300 12880
rect -3500 9720 -3460 12840
rect -340 9720 -300 12840
rect -3500 9680 -300 9720
rect 300 12840 3500 12880
rect 300 9720 340 12840
rect 3460 9720 3500 12840
rect 300 9680 3500 9720
rect 4100 12840 7300 12880
rect 4100 9720 4140 12840
rect 7260 9720 7300 12840
rect 4100 9680 7300 9720
<< mimcapcontact >>
rect -7260 9720 -4140 12840
rect -3460 9720 -340 12840
rect 340 9720 3460 12840
rect 4140 9720 7260 12840
<< metal4 >>
rect -9970 13130 9970 13190
rect -9970 13000 -9930 13130
rect -9830 13000 -9670 13130
rect -9570 13059 9560 13130
rect -9570 13000 -7372 13059
rect -9970 12995 -7372 13000
rect -4028 12995 -3572 13059
rect -228 12995 228 13059
rect 3572 12995 4028 13059
rect 7372 13000 9560 13059
rect 9670 13000 9820 13130
rect 9930 13000 9970 13130
rect 7372 12995 9970 13000
rect -9970 12950 9970 12995
rect -7261 12840 -4139 12841
rect -7261 9720 -7260 12840
rect -4140 11690 -4139 12840
rect -3461 12840 -339 12841
rect -3461 11690 -3460 12840
rect -4140 11330 -3460 11690
rect -4140 9720 -4139 11330
rect -7261 9719 -4139 9720
rect -3920 9510 -3750 11330
rect -3461 9720 -3460 11330
rect -340 11690 -339 12840
rect 339 12840 3461 12841
rect 339 11690 340 12840
rect -340 11330 340 11690
rect -340 9720 -339 11330
rect -3461 9719 -339 9720
rect 339 9720 340 11330
rect 3460 11690 3461 12840
rect 4139 12840 7261 12841
rect 4139 11690 4140 12840
rect 3460 11330 4140 11690
rect 3460 9720 3461 11330
rect 339 9719 3461 9720
rect -5720 9320 -3750 9510
rect 3720 9530 3880 11330
rect 4139 9720 4140 11330
rect 7260 9720 7261 12840
rect 4139 9719 7261 9720
rect 3720 9400 4500 9530
rect -5720 5790 -5430 9320
rect -5720 5680 -5700 5790
rect -5610 5680 -5540 5790
rect -5450 5680 -5430 5790
rect -5720 5460 -5430 5680
rect -3500 8820 -3230 8950
rect -3500 8740 -3480 8820
rect -3400 8740 -3330 8820
rect -3250 8740 -3230 8820
rect -3500 8280 -3230 8740
rect -3500 8200 -3480 8280
rect -3400 8200 -3330 8280
rect -3250 8200 -3230 8280
rect -3500 7740 -3230 8200
rect -3500 7660 -3480 7740
rect -3400 7660 -3330 7740
rect -3250 7660 -3230 7740
rect -3500 2510 -3230 7660
rect -1010 8820 -740 9000
rect -1010 8740 -990 8820
rect -910 8740 -840 8820
rect -760 8740 -740 8820
rect -1010 8280 -740 8740
rect -1010 8200 -990 8280
rect -910 8200 -840 8280
rect -760 8200 -740 8280
rect -1010 7740 -740 8200
rect -1010 7660 -990 7740
rect -910 7660 -840 7740
rect -760 7660 -740 7740
rect -2210 7140 -1980 7160
rect -2210 7060 -2190 7140
rect -2110 7060 -2080 7140
rect -2000 7060 -1980 7140
rect -2210 6530 -1980 7060
rect -2210 6450 -2190 6530
rect -2110 6450 -2080 6530
rect -2000 6450 -1980 6530
rect -2210 5970 -1980 6450
rect -2210 5890 -2190 5970
rect -2110 5890 -2080 5970
rect -2000 5890 -1980 5970
rect -2210 3270 -1980 5890
rect -2210 3190 -2190 3270
rect -2110 3190 -2080 3270
rect -2000 3190 -1980 3270
rect -2210 3170 -1980 3190
rect -3500 2430 -3480 2510
rect -3400 2430 -3330 2510
rect -3250 2430 -3230 2510
rect -1010 2530 -740 7660
rect 1470 8820 1740 9010
rect 1470 8740 1490 8820
rect 1570 8740 1640 8820
rect 1720 8740 1740 8820
rect 1470 8280 1740 8740
rect 1470 8200 1490 8280
rect 1570 8200 1640 8280
rect 1720 8200 1740 8280
rect 1470 7740 1740 8200
rect 1470 7660 1500 7740
rect 1580 7660 1640 7740
rect 1720 7660 1740 7740
rect 200 7140 430 7160
rect 200 7060 220 7140
rect 300 7060 330 7140
rect 410 7060 430 7140
rect 200 6550 430 7060
rect 200 6470 220 6550
rect 300 6470 330 6550
rect 410 6470 430 6550
rect 200 5970 430 6470
rect 200 5890 220 5970
rect 300 5890 330 5970
rect 410 5890 430 5970
rect 200 3270 430 5890
rect 200 3190 220 3270
rect 300 3190 330 3270
rect 410 3190 430 3270
rect 200 3170 430 3190
rect -1010 2450 -990 2530
rect -910 2450 -840 2530
rect -760 2450 -740 2530
rect -1010 2430 -740 2450
rect 1470 2530 1740 7660
rect 2660 7130 2890 7170
rect 2660 7050 2680 7130
rect 2760 7050 2790 7130
rect 2870 7050 2890 7130
rect 2660 6550 2890 7050
rect 2660 6470 2680 6550
rect 2760 6470 2790 6550
rect 2870 6470 2890 6550
rect 2660 5970 2890 6470
rect 2660 5890 2680 5970
rect 2760 5890 2790 5970
rect 2870 5890 2890 5970
rect 2660 3280 2890 5890
rect 4210 5740 4500 9400
rect 4210 5660 4230 5740
rect 4310 5660 4400 5740
rect 4480 5660 4500 5740
rect 4210 5250 4500 5660
rect 2660 3200 2680 3280
rect 2760 3200 2790 3280
rect 2870 3200 2890 3280
rect 2660 3180 2890 3200
rect 1470 2450 1490 2530
rect 1570 2450 1630 2530
rect 1710 2450 1740 2530
rect 1470 2430 1740 2450
rect -3500 2400 -3230 2430
rect 1819 580 1941 581
rect 1819 480 1820 580
rect 1940 480 1941 580
rect 1819 479 1941 480
<< res5p73 >>
rect -9417 4961 -7413 6111
rect 7643 4961 9647 6111
rect -9417 3491 -7413 4641
rect 7643 3491 9647 4641
<< labels >>
rlabel metal3 5110 1800 5110 1800 1 VSS
port 4 n
rlabel metal3 6920 7930 6920 7930 1 VDD
port 3 n
rlabel metal2 -440 3590 -440 3590 1 Vout
port 2 n
rlabel metal1 -1780 200 -1780 200 1 Vin
port 1 n
rlabel space -300 3530 -160 3590 1 find
rlabel metal1 -1784 2574 -1784 2574 1 Vn_OR
port 5 n
rlabel metal1 -1784 3086 -1784 3086 1 Vp_OR
port 6 n
rlabel metal1 6364 5554 6364 5554 1 Vmid
port 7 n
<< end >>
