magic
tech sky130A
timestamp 1709390584
<< pwell >>
rect -360 -355 360 355
<< nmos >>
rect -262 -250 -212 250
rect -183 -250 -133 250
rect -104 -250 -54 250
rect -25 -250 25 250
rect 54 -250 104 250
rect 133 -250 183 250
rect 212 -250 262 250
<< ndiff >>
rect -291 244 -262 250
rect -291 -244 -285 244
rect -268 -244 -262 244
rect -291 -250 -262 -244
rect -212 244 -183 250
rect -212 -244 -206 244
rect -189 -244 -183 244
rect -212 -250 -183 -244
rect -133 244 -104 250
rect -133 -244 -127 244
rect -110 -244 -104 244
rect -133 -250 -104 -244
rect -54 244 -25 250
rect -54 -244 -48 244
rect -31 -244 -25 244
rect -54 -250 -25 -244
rect 25 244 54 250
rect 25 -244 31 244
rect 48 -244 54 244
rect 25 -250 54 -244
rect 104 244 133 250
rect 104 -244 110 244
rect 127 -244 133 244
rect 104 -250 133 -244
rect 183 244 212 250
rect 183 -244 189 244
rect 206 -244 212 244
rect 183 -250 212 -244
rect 262 244 291 250
rect 262 -244 268 244
rect 285 -244 291 244
rect 262 -250 291 -244
<< ndiffc >>
rect -285 -244 -268 244
rect -206 -244 -189 244
rect -127 -244 -110 244
rect -48 -244 -31 244
rect 31 -244 48 244
rect 110 -244 127 244
rect 189 -244 206 244
rect 268 -244 285 244
<< psubdiff >>
rect -342 320 -294 337
rect 294 320 342 337
rect -342 289 -325 320
rect 325 289 342 320
rect -342 -320 -325 -289
rect 325 -320 342 -289
rect -342 -337 -294 -320
rect 294 -337 342 -320
<< psubdiffcont >>
rect -294 320 294 337
rect -342 -289 -325 289
rect 325 -289 342 289
rect -294 -337 294 -320
<< poly >>
rect -262 286 -212 294
rect -262 269 -254 286
rect -220 269 -212 286
rect -262 250 -212 269
rect -183 286 -133 294
rect -183 269 -175 286
rect -141 269 -133 286
rect -183 250 -133 269
rect -104 286 -54 294
rect -104 269 -96 286
rect -62 269 -54 286
rect -104 250 -54 269
rect -25 286 25 294
rect -25 269 -17 286
rect 17 269 25 286
rect -25 250 25 269
rect 54 286 104 294
rect 54 269 62 286
rect 96 269 104 286
rect 54 250 104 269
rect 133 286 183 294
rect 133 269 141 286
rect 175 269 183 286
rect 133 250 183 269
rect 212 286 262 294
rect 212 269 220 286
rect 254 269 262 286
rect 212 250 262 269
rect -262 -269 -212 -250
rect -262 -286 -254 -269
rect -220 -286 -212 -269
rect -262 -294 -212 -286
rect -183 -269 -133 -250
rect -183 -286 -175 -269
rect -141 -286 -133 -269
rect -183 -294 -133 -286
rect -104 -269 -54 -250
rect -104 -286 -96 -269
rect -62 -286 -54 -269
rect -104 -294 -54 -286
rect -25 -269 25 -250
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect -25 -294 25 -286
rect 54 -269 104 -250
rect 54 -286 62 -269
rect 96 -286 104 -269
rect 54 -294 104 -286
rect 133 -269 183 -250
rect 133 -286 141 -269
rect 175 -286 183 -269
rect 133 -294 183 -286
rect 212 -269 262 -250
rect 212 -286 220 -269
rect 254 -286 262 -269
rect 212 -294 262 -286
<< polycont >>
rect -254 269 -220 286
rect -175 269 -141 286
rect -96 269 -62 286
rect -17 269 17 286
rect 62 269 96 286
rect 141 269 175 286
rect 220 269 254 286
rect -254 -286 -220 -269
rect -175 -286 -141 -269
rect -96 -286 -62 -269
rect -17 -286 17 -269
rect 62 -286 96 -269
rect 141 -286 175 -269
rect 220 -286 254 -269
<< locali >>
rect -342 320 -294 337
rect 294 320 342 337
rect -342 289 -325 320
rect 325 289 342 320
rect -262 269 -254 286
rect -220 269 -212 286
rect -183 269 -175 286
rect -141 269 -133 286
rect -104 269 -96 286
rect -62 269 -54 286
rect -25 269 -17 286
rect 17 269 25 286
rect 54 269 62 286
rect 96 269 104 286
rect 133 269 141 286
rect 175 269 183 286
rect 212 269 220 286
rect 254 269 262 286
rect -285 244 -268 252
rect -285 -252 -268 -244
rect -206 244 -189 252
rect -206 -252 -189 -244
rect -127 244 -110 252
rect -127 -252 -110 -244
rect -48 244 -31 252
rect -48 -252 -31 -244
rect 31 244 48 252
rect 31 -252 48 -244
rect 110 244 127 252
rect 110 -252 127 -244
rect 189 244 206 252
rect 189 -252 206 -244
rect 268 244 285 252
rect 268 -252 285 -244
rect -262 -286 -254 -269
rect -220 -286 -212 -269
rect -183 -286 -175 -269
rect -141 -286 -133 -269
rect -104 -286 -96 -269
rect -62 -286 -54 -269
rect -25 -286 -17 -269
rect 17 -286 25 -269
rect 54 -286 62 -269
rect 96 -286 104 -269
rect 133 -286 141 -269
rect 175 -286 183 -269
rect 212 -286 220 -269
rect 254 -286 262 -269
rect -342 -320 -325 -289
rect 325 -320 342 -289
rect -342 -337 -294 -320
rect 294 -337 342 -320
<< viali >>
rect -254 269 -220 286
rect -175 269 -141 286
rect -96 269 -62 286
rect -17 269 17 286
rect 62 269 96 286
rect 141 269 175 286
rect 220 269 254 286
rect -285 -244 -268 244
rect -206 -244 -189 244
rect -127 -244 -110 244
rect -48 -244 -31 244
rect 31 -244 48 244
rect 110 -244 127 244
rect 189 -244 206 244
rect 268 -244 285 244
rect -254 -286 -220 -269
rect -175 -286 -141 -269
rect -96 -286 -62 -269
rect -17 -286 17 -269
rect 62 -286 96 -269
rect 141 -286 175 -269
rect 220 -286 254 -269
<< metal1 >>
rect -260 286 -214 289
rect -260 269 -254 286
rect -220 269 -214 286
rect -260 266 -214 269
rect -181 286 -135 289
rect -181 269 -175 286
rect -141 269 -135 286
rect -181 266 -135 269
rect -102 286 -56 289
rect -102 269 -96 286
rect -62 269 -56 286
rect -102 266 -56 269
rect -23 286 23 289
rect -23 269 -17 286
rect 17 269 23 286
rect -23 266 23 269
rect 56 286 102 289
rect 56 269 62 286
rect 96 269 102 286
rect 56 266 102 269
rect 135 286 181 289
rect 135 269 141 286
rect 175 269 181 286
rect 135 266 181 269
rect 214 286 260 289
rect 214 269 220 286
rect 254 269 260 286
rect 214 266 260 269
rect -288 244 -265 250
rect -288 -244 -285 244
rect -268 -244 -265 244
rect -288 -250 -265 -244
rect -209 244 -186 250
rect -209 -244 -206 244
rect -189 -244 -186 244
rect -209 -250 -186 -244
rect -130 244 -107 250
rect -130 -244 -127 244
rect -110 -244 -107 244
rect -130 -250 -107 -244
rect -51 244 -28 250
rect -51 -244 -48 244
rect -31 -244 -28 244
rect -51 -250 -28 -244
rect 28 244 51 250
rect 28 -244 31 244
rect 48 -244 51 244
rect 28 -250 51 -244
rect 107 244 130 250
rect 107 -244 110 244
rect 127 -244 130 244
rect 107 -250 130 -244
rect 186 244 209 250
rect 186 -244 189 244
rect 206 -244 209 244
rect 186 -250 209 -244
rect 265 244 288 250
rect 265 -244 268 244
rect 285 -244 288 244
rect 265 -250 288 -244
rect -260 -269 -214 -266
rect -260 -286 -254 -269
rect -220 -286 -214 -269
rect -260 -289 -214 -286
rect -181 -269 -135 -266
rect -181 -286 -175 -269
rect -141 -286 -135 -269
rect -181 -289 -135 -286
rect -102 -269 -56 -266
rect -102 -286 -96 -269
rect -62 -286 -56 -269
rect -102 -289 -56 -286
rect -23 -269 23 -266
rect -23 -286 -17 -269
rect 17 -286 23 -269
rect -23 -289 23 -286
rect 56 -269 102 -266
rect 56 -286 62 -269
rect 96 -286 102 -269
rect 56 -289 102 -286
rect 135 -269 181 -266
rect 135 -286 141 -269
rect 175 -286 181 -269
rect 135 -289 181 -286
rect 214 -269 260 -266
rect 214 -286 220 -269
rect 254 -286 260 -269
rect 214 -289 260 -286
<< properties >>
string FIXED_BBOX -333 -328 333 328
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
