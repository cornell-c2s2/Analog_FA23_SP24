magic
tech sky130A
timestamp 1716869746
<< pwell >>
rect -128 -305 128 305
<< nmoslvt >>
rect -30 -200 30 200
<< ndiff >>
rect -59 194 -30 200
rect -59 -194 -53 194
rect -36 -194 -30 194
rect -59 -200 -30 -194
rect 30 194 59 200
rect 30 -194 36 194
rect 53 -194 59 194
rect 30 -200 59 -194
<< ndiffc >>
rect -53 -194 -36 194
rect 36 -194 53 194
<< psubdiff >>
rect -110 270 -62 287
rect 62 270 110 287
rect -110 239 -93 270
rect 93 239 110 270
rect -110 -270 -93 -239
rect 93 -270 110 -239
rect -110 -287 -62 -270
rect 62 -287 110 -270
<< psubdiffcont >>
rect -62 270 62 287
rect -110 -239 -93 239
rect 93 -239 110 239
rect -62 -287 62 -270
<< poly >>
rect -30 236 30 244
rect -30 219 -22 236
rect 22 219 30 236
rect -30 200 30 219
rect -30 -219 30 -200
rect -30 -236 -22 -219
rect 22 -236 30 -219
rect -30 -244 30 -236
<< polycont >>
rect -22 219 22 236
rect -22 -236 22 -219
<< locali >>
rect -110 270 -62 287
rect 62 270 110 287
rect -110 239 -93 270
rect 93 239 110 270
rect -30 219 -22 236
rect 22 219 30 236
rect -53 194 -36 202
rect -53 -202 -36 -194
rect 36 194 53 202
rect 36 -202 53 -194
rect -30 -236 -22 -219
rect 22 -236 30 -219
rect -110 -270 -93 -239
rect 93 -270 110 -239
rect -110 -287 -62 -270
rect 62 -287 110 -270
<< viali >>
rect -22 219 22 236
rect -53 -194 -36 194
rect 36 -194 53 194
rect -22 -236 22 -219
<< metal1 >>
rect -28 236 28 239
rect -28 219 -22 236
rect 22 219 28 236
rect -28 216 28 219
rect -56 194 -33 200
rect -56 -194 -53 194
rect -36 -194 -33 194
rect -56 -200 -33 -194
rect 33 194 56 200
rect 33 -194 36 194
rect 53 -194 56 194
rect 33 -200 56 -194
rect -28 -219 28 -216
rect -28 -236 -22 -219
rect 22 -236 28 -219
rect -28 -239 28 -236
<< properties >>
string FIXED_BBOX -101 -278 101 278
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
