magic
tech sky130A
timestamp 1708718592
<< checkpaint >>
rect -649 1202 1063 1226
rect -649 1178 1496 1202
rect -649 1154 1929 1178
rect -649 1130 2362 1154
rect -649 1106 2611 1130
rect -649 1082 3044 1106
rect -649 1058 3477 1082
rect -649 1034 3910 1058
rect -649 1010 4343 1034
rect -649 986 4500 1010
rect -649 -354 4749 986
rect -630 -426 4749 -354
rect -630 -1630 730 -426
rect 1083 -450 4749 -426
rect 1332 -474 4749 -450
rect 1765 -498 4749 -474
rect 2198 -522 4749 -498
rect 2631 -546 4749 -522
rect 3064 -570 4749 -546
rect 3221 -594 4749 -570
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
use sky130_fd_sc_hd__nand2_4  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 0 0 1 300
box -19 -24 433 296
use sky130_fd_sc_hd__nand2_4  x4
timestamp 1701704242
transform 1 0 433 0 1 276
box -19 -24 433 296
use sky130_fd_sc_hd__nand2_4  x5
timestamp 1701704242
transform 1 0 866 0 1 252
box -19 -24 433 296
use sky130_fd_sc_hd__nand2_4  x6
timestamp 1701704242
transform 1 0 1299 0 1 228
box -19 -24 433 296
use sky130_fd_sc_hd__inv_4  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1732 0 1 204
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_4  x9
timestamp 1701704242
transform 1 0 1981 0 1 180
box -19 -24 433 296
use sky130_fd_sc_hd__nand2_4  x10
timestamp 1701704242
transform 1 0 2414 0 1 156
box -19 -24 433 296
use sky130_fd_sc_hd__nand2_4  x11
timestamp 1701704242
transform 1 0 2847 0 1 132
box -19 -24 433 296
use sky130_fd_sc_hd__nand2_4  x12
timestamp 1701704242
transform 1 0 3280 0 1 108
box -19 -24 433 296
use sky130_fd_sc_hd__inv_4  x13
timestamp 1701704242
transform 1 0 3870 0 1 60
box -19 -24 249 296
use sky130_fd_sc_hd__clkinv_1  x14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3713 0 1 84
box -19 -24 157 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 VDD
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 SIG
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 OUT
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 CLK
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 VSS
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 VMID
port 5 nsew
<< end >>
