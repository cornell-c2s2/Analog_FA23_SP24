magic
tech sky130A
magscale 1 2
timestamp 1713027377
<< error_s >>
rect -1678 5424 -1142 5472
rect -1678 5376 -828 5424
rect -1678 5328 -330 5376
rect -1678 5280 1180 5328
rect -1678 5232 1494 5280
rect -1678 5184 1992 5232
rect -1678 5151 3502 5184
rect -1180 5136 3502 5151
rect -1180 5103 3816 5136
rect -866 5088 3816 5103
rect -1403 5021 -1351 5067
rect -1584 4937 -1532 5021
rect -1502 4937 -1448 5021
rect -1418 4937 -1351 5021
rect -1321 4937 -1269 5067
rect -866 5055 4314 5088
rect -368 5040 4314 5055
rect -1074 4889 -1022 5019
rect -992 4889 -940 5019
rect -368 5007 5824 5040
rect -791 4841 -739 4971
rect -709 4841 -655 4971
rect -625 4841 -571 4971
rect -541 4841 -487 4971
rect -457 4841 -405 4971
rect 1142 4959 5824 5007
rect -290 4793 -238 4923
rect -208 4793 -154 4923
rect -124 4793 -70 4923
rect -40 4793 14 4923
rect 44 4793 98 4923
rect 128 4793 182 4923
rect 212 4793 266 4923
rect 296 4793 350 4923
rect 380 4793 434 4923
rect 464 4793 518 4923
rect 548 4793 602 4923
rect 632 4793 686 4923
rect 716 4793 770 4923
rect 800 4793 854 4923
rect 884 4793 938 4923
rect 968 4793 1022 4923
rect 1052 4793 1104 4923
rect 1456 4911 5824 4959
rect 1248 4745 1300 4875
rect 1330 4745 1382 4875
rect 1954 4863 5824 4911
rect 1531 4697 1583 4827
rect 1613 4697 1667 4827
rect 1697 4697 1751 4827
rect 1781 4697 1835 4827
rect 1865 4697 1917 4827
rect 3464 4815 5824 4863
rect 2032 4649 2084 4779
rect 2114 4649 2168 4779
rect 2198 4649 2252 4779
rect 2282 4649 2336 4779
rect 2366 4649 2420 4779
rect 2450 4649 2504 4779
rect 2534 4649 2588 4779
rect 2618 4649 2672 4779
rect 2702 4649 2756 4779
rect 2786 4649 2840 4779
rect 2870 4649 2924 4779
rect 2954 4649 3008 4779
rect 3038 4649 3092 4779
rect 3122 4649 3176 4779
rect 3206 4649 3260 4779
rect 3290 4649 3344 4779
rect 3374 4649 3426 4779
rect 3778 4767 5824 4815
rect 3570 4601 3622 4731
rect 3652 4601 3704 4731
rect 4276 4719 5824 4767
rect 8108 4800 8460 4848
rect 8108 4752 8958 4800
rect 3853 4553 3905 4683
rect 3935 4553 3989 4683
rect 4019 4553 4073 4683
rect 4103 4553 4157 4683
rect 4187 4553 4239 4683
rect 4354 4505 4406 4635
rect 4436 4505 4490 4635
rect 4520 4505 4574 4635
rect 4604 4505 4658 4635
rect 4688 4505 4742 4635
rect 4772 4505 4826 4635
rect 4856 4505 4910 4635
rect 4940 4505 4994 4635
rect 5024 4505 5078 4635
rect 5108 4505 5162 4635
rect 5192 4505 5246 4635
rect 5276 4505 5330 4635
rect 5360 4505 5414 4635
rect 5444 4505 5498 4635
rect 5528 4505 5582 4635
rect 5612 4505 5666 4635
rect 5696 4505 5748 4635
rect 8108 4527 9456 4752
rect 8422 4479 9456 4527
rect 8214 4313 8266 4443
rect 8296 4313 8348 4443
rect 8920 4431 9456 4479
rect 16748 4464 18296 4512
rect 20798 4488 22346 4536
rect 8697 4349 8749 4395
rect 8516 4265 8568 4349
rect 8598 4265 8652 4349
rect 8682 4265 8749 4349
rect 8779 4265 8831 4395
rect 9195 4301 9247 4347
rect 9014 4217 9066 4301
rect 9096 4217 9150 4301
rect 9180 4217 9247 4301
rect 9277 4217 9329 4347
rect 16748 4191 19806 4464
rect 20798 4440 23856 4488
rect 20798 4392 25366 4440
rect 20798 4344 26876 4392
rect 20798 4296 28386 4344
rect 20798 4248 29896 4296
rect 20798 4215 31406 4248
rect 18258 4143 19806 4191
rect 22308 4200 31406 4215
rect 22308 4167 32916 4200
rect 23818 4152 32916 4167
rect 16826 3977 16878 4107
rect 16908 3977 16962 4107
rect 16992 3977 17046 4107
rect 17076 3977 17130 4107
rect 17160 3977 17214 4107
rect 17244 3977 17298 4107
rect 17328 3977 17382 4107
rect 17412 3977 17466 4107
rect 17496 3977 17550 4107
rect 17580 3977 17634 4107
rect 17664 3977 17718 4107
rect 17748 3977 17802 4107
rect 17832 3977 17886 4107
rect 17916 3977 17970 4107
rect 18000 3977 18054 4107
rect 18084 3977 18138 4107
rect 18168 3977 18220 4107
rect 18336 3929 18388 4059
rect 18418 3929 18472 4059
rect 18502 3929 18556 4059
rect 18586 3929 18640 4059
rect 18670 3929 18724 4059
rect 18754 3929 18808 4059
rect 18838 3929 18892 4059
rect 18922 3929 18976 4059
rect 19006 3929 19060 4059
rect 19090 3929 19144 4059
rect 19174 3929 19228 4059
rect 19258 3929 19312 4059
rect 19342 3929 19396 4059
rect 19426 3929 19480 4059
rect 19510 3929 19564 4059
rect 19594 3929 19648 4059
rect 19678 3929 19730 4059
rect 20876 4001 20928 4131
rect 20958 4001 21012 4131
rect 21042 4001 21096 4131
rect 21126 4001 21180 4131
rect 21210 4001 21264 4131
rect 21294 4001 21348 4131
rect 21378 4001 21432 4131
rect 21462 4001 21516 4131
rect 21546 4001 21600 4131
rect 21630 4001 21684 4131
rect 21714 4001 21768 4131
rect 21798 4001 21852 4131
rect 21882 4001 21936 4131
rect 21966 4001 22020 4131
rect 22050 4001 22104 4131
rect 22134 4001 22188 4131
rect 22218 4001 22270 4131
rect 23818 4119 34426 4152
rect 25328 4104 34426 4119
rect 22386 3953 22438 4083
rect 22468 3953 22522 4083
rect 22552 3953 22606 4083
rect 22636 3953 22690 4083
rect 22720 3953 22774 4083
rect 22804 3953 22858 4083
rect 22888 3953 22942 4083
rect 22972 3953 23026 4083
rect 23056 3953 23110 4083
rect 23140 3953 23194 4083
rect 23224 3953 23278 4083
rect 23308 3953 23362 4083
rect 23392 3953 23446 4083
rect 23476 3953 23530 4083
rect 23560 3953 23614 4083
rect 23644 3953 23698 4083
rect 23728 3953 23780 4083
rect 25328 4071 35936 4104
rect 23896 3905 23948 4035
rect 23978 3905 24032 4035
rect 24062 3905 24116 4035
rect 24146 3905 24200 4035
rect 24230 3905 24284 4035
rect 24314 3905 24368 4035
rect 24398 3905 24452 4035
rect 24482 3905 24536 4035
rect 24566 3905 24620 4035
rect 24650 3905 24704 4035
rect 24734 3905 24788 4035
rect 24818 3905 24872 4035
rect 24902 3905 24956 4035
rect 24986 3905 25040 4035
rect 25070 3905 25124 4035
rect 25154 3905 25208 4035
rect 25238 3905 25290 4035
rect 26838 4023 35936 4071
rect 25406 3857 25458 3987
rect 25488 3857 25542 3987
rect 25572 3857 25626 3987
rect 25656 3857 25710 3987
rect 25740 3857 25794 3987
rect 25824 3857 25878 3987
rect 25908 3857 25962 3987
rect 25992 3857 26046 3987
rect 26076 3857 26130 3987
rect 26160 3857 26214 3987
rect 26244 3857 26298 3987
rect 26328 3857 26382 3987
rect 26412 3857 26466 3987
rect 26496 3857 26550 3987
rect 26580 3857 26634 3987
rect 26664 3857 26718 3987
rect 26748 3857 26800 3987
rect 28348 3975 35936 4023
rect 26916 3809 26968 3939
rect 26998 3809 27052 3939
rect 27082 3809 27136 3939
rect 27166 3809 27220 3939
rect 27250 3809 27304 3939
rect 27334 3809 27388 3939
rect 27418 3809 27472 3939
rect 27502 3809 27556 3939
rect 27586 3809 27640 3939
rect 27670 3809 27724 3939
rect 27754 3809 27808 3939
rect 27838 3809 27892 3939
rect 27922 3809 27976 3939
rect 28006 3809 28060 3939
rect 28090 3809 28144 3939
rect 28174 3809 28228 3939
rect 28258 3809 28310 3939
rect 29858 3927 35936 3975
rect 28426 3761 28478 3891
rect 28508 3761 28562 3891
rect 28592 3761 28646 3891
rect 28676 3761 28730 3891
rect 28760 3761 28814 3891
rect 28844 3761 28898 3891
rect 28928 3761 28982 3891
rect 29012 3761 29066 3891
rect 29096 3761 29150 3891
rect 29180 3761 29234 3891
rect 29264 3761 29318 3891
rect 29348 3761 29402 3891
rect 29432 3761 29486 3891
rect 29516 3761 29570 3891
rect 29600 3761 29654 3891
rect 29684 3761 29738 3891
rect 29768 3761 29820 3891
rect 31368 3879 35936 3927
rect 29936 3713 29988 3843
rect 30018 3713 30072 3843
rect 30102 3713 30156 3843
rect 30186 3713 30240 3843
rect 30270 3713 30324 3843
rect 30354 3713 30408 3843
rect 30438 3713 30492 3843
rect 30522 3713 30576 3843
rect 30606 3713 30660 3843
rect 30690 3713 30744 3843
rect 30774 3713 30828 3843
rect 30858 3713 30912 3843
rect 30942 3713 30996 3843
rect 31026 3713 31080 3843
rect 31110 3713 31164 3843
rect 31194 3713 31248 3843
rect 31278 3713 31330 3843
rect 32878 3831 35936 3879
rect 31446 3665 31498 3795
rect 31528 3665 31582 3795
rect 31612 3665 31666 3795
rect 31696 3665 31750 3795
rect 31780 3665 31834 3795
rect 31864 3665 31918 3795
rect 31948 3665 32002 3795
rect 32032 3665 32086 3795
rect 32116 3665 32170 3795
rect 32200 3665 32254 3795
rect 32284 3665 32338 3795
rect 32368 3665 32422 3795
rect 32452 3665 32506 3795
rect 32536 3665 32590 3795
rect 32620 3665 32674 3795
rect 32704 3665 32758 3795
rect 32788 3665 32840 3795
rect 34388 3783 35936 3831
rect 32956 3617 33008 3747
rect 33038 3617 33092 3747
rect 33122 3617 33176 3747
rect 33206 3617 33260 3747
rect 33290 3617 33344 3747
rect 33374 3617 33428 3747
rect 33458 3617 33512 3747
rect 33542 3617 33596 3747
rect 33626 3617 33680 3747
rect 33710 3617 33764 3747
rect 33794 3617 33848 3747
rect 33878 3617 33932 3747
rect 33962 3617 34016 3747
rect 34046 3617 34100 3747
rect 34130 3617 34184 3747
rect 34214 3617 34268 3747
rect 34298 3617 34350 3747
rect 34466 3569 34518 3699
rect 34548 3569 34602 3699
rect 34632 3569 34686 3699
rect 34716 3569 34770 3699
rect 34800 3569 34854 3699
rect 34884 3569 34938 3699
rect 34968 3569 35022 3699
rect 35052 3569 35106 3699
rect 35136 3569 35190 3699
rect 35220 3569 35274 3699
rect 35304 3569 35358 3699
rect 35388 3569 35442 3699
rect 35472 3569 35526 3699
rect 35556 3569 35610 3699
rect 35640 3569 35694 3699
rect 35724 3569 35778 3699
rect 35808 3569 35860 3699
rect 8790 -690 8814 -666
rect 8876 -690 8900 -666
rect 8766 -714 8790 -690
rect 8900 -714 8924 -690
rect 8766 -800 8790 -776
rect 8900 -800 8924 -776
rect 8790 -824 8814 -800
rect 8876 -824 8900 -800
rect 10650 -1140 10690 -1132
rect 10650 -1178 10690 -1170
rect 8910 -1223 8963 -1216
rect 8997 -1223 9014 -1216
rect 9384 -1225 9426 -1216
rect 11883 -1225 11916 -1025
rect 11946 -1225 12000 -1025
rect 12030 -1225 12084 -1025
rect 12114 -1225 12168 -1025
rect 12198 -1225 12250 -1025
rect 12328 -1225 12380 -1025
rect 12410 -1225 12464 -1025
rect 12494 -1225 12548 -1025
rect 12578 -1225 12632 -1025
rect 12662 -1225 12716 -1025
rect 12746 -1225 12800 -1025
rect 12830 -1225 12884 -1025
rect 12914 -1225 12968 -1025
rect 12998 -1225 13052 -1025
rect 13082 -1225 13136 -1025
rect 13166 -1225 13220 -1025
rect 13250 -1225 13304 -1025
rect 13334 -1225 13388 -1025
rect 13418 -1225 13472 -1025
rect 13502 -1225 13556 -1025
rect 13586 -1225 13640 -1025
rect 13670 -1225 13722 -1025
rect 13800 -1225 13852 -1025
rect 13882 -1225 13936 -1025
rect 13966 -1225 14020 -1025
rect 14050 -1225 14104 -1025
rect 14134 -1225 14188 -1025
rect 14218 -1225 14272 -1025
rect 14302 -1225 14356 -1025
rect 14386 -1225 14440 -1025
rect 14470 -1225 14524 -1025
rect 14554 -1225 14608 -1025
rect 14638 -1225 14692 -1025
rect 14722 -1225 14776 -1025
rect 14806 -1225 14860 -1025
rect 14890 -1225 14944 -1025
rect 14974 -1225 15028 -1025
rect 15058 -1225 15112 -1025
rect 15142 -1225 15194 -1025
rect 15272 -1225 15324 -1025
rect 15354 -1225 15408 -1025
rect 15438 -1225 15492 -1025
rect 15522 -1225 15576 -1025
rect 15606 -1225 15660 -1025
rect 15690 -1225 15744 -1025
rect 15774 -1225 15828 -1025
rect 15858 -1225 15912 -1025
rect 15942 -1225 15996 -1025
rect 16026 -1225 16080 -1025
rect 16110 -1225 16164 -1025
rect 16194 -1225 16248 -1025
rect 16278 -1225 16332 -1025
rect 16362 -1225 16416 -1025
rect 16446 -1225 16500 -1025
rect 16530 -1225 16584 -1025
rect 16614 -1225 16666 -1025
rect 8876 -1257 8980 -1250
rect 9350 -1259 9430 -1250
rect 8676 -1475 8728 -1345
rect 8758 -1475 8810 -1345
rect 8921 -1475 8973 -1345
rect 9003 -1475 9057 -1345
rect 9087 -1475 9141 -1345
rect 9171 -1475 9225 -1345
rect 9255 -1475 9307 -1345
rect 9384 -1475 9436 -1345
rect 9466 -1475 9520 -1345
rect 9550 -1475 9604 -1345
rect 9634 -1475 9688 -1345
rect 9718 -1475 9772 -1345
rect 9802 -1475 9856 -1345
rect 9886 -1475 9940 -1345
rect 9970 -1475 10024 -1345
rect 10054 -1475 10108 -1345
rect 10138 -1475 10192 -1345
rect 10222 -1475 10276 -1345
rect 10306 -1475 10360 -1345
rect 10390 -1475 10444 -1345
rect 10474 -1475 10528 -1345
rect 10558 -1475 10612 -1345
rect 10642 -1475 10696 -1345
rect 10726 -1475 10778 -1345
rect 10856 -1475 10908 -1345
rect 10938 -1475 10992 -1345
rect 11022 -1475 11076 -1345
rect 11106 -1475 11160 -1345
rect 11190 -1475 11244 -1345
rect 11274 -1475 11328 -1345
rect 11358 -1475 11412 -1345
rect 11442 -1475 11496 -1345
rect 11526 -1475 11580 -1345
rect 11610 -1475 11664 -1345
rect 11694 -1475 11748 -1345
rect 11778 -1475 11832 -1345
rect 11862 -1475 11916 -1345
rect 11946 -1475 12000 -1345
rect 12030 -1475 12084 -1345
rect 12114 -1475 12168 -1345
rect 12198 -1475 12250 -1345
rect 12328 -1475 12380 -1345
rect 12410 -1475 12464 -1345
rect 12494 -1475 12548 -1345
rect 12578 -1475 12632 -1345
rect 12662 -1475 12716 -1345
rect 12746 -1475 12800 -1345
rect 12830 -1475 12884 -1345
rect 12914 -1475 12968 -1345
rect 12998 -1475 13052 -1345
rect 13082 -1475 13136 -1345
rect 13166 -1475 13220 -1345
rect 13250 -1475 13304 -1345
rect 13334 -1475 13388 -1345
rect 13418 -1475 13472 -1345
rect 13502 -1475 13556 -1345
rect 13586 -1475 13640 -1345
rect 13670 -1475 13722 -1345
rect 13800 -1475 13852 -1345
rect 13882 -1475 13936 -1345
rect 13966 -1475 14020 -1345
rect 14050 -1475 14104 -1345
rect 14134 -1475 14188 -1345
rect 14218 -1475 14272 -1345
rect 14302 -1475 14356 -1345
rect 14386 -1475 14440 -1345
rect 14470 -1475 14524 -1345
rect 14554 -1475 14608 -1345
rect 14638 -1475 14692 -1345
rect 14722 -1475 14776 -1345
rect 14806 -1475 14860 -1345
rect 14890 -1475 14944 -1345
rect 14974 -1475 15028 -1345
rect 15058 -1475 15112 -1345
rect 15142 -1475 15194 -1345
rect 15272 -1475 15324 -1345
rect 15354 -1475 15408 -1345
rect 15438 -1475 15492 -1345
rect 15522 -1475 15576 -1345
rect 15606 -1475 15660 -1345
rect 15690 -1475 15744 -1345
rect 15774 -1475 15828 -1345
rect 15858 -1475 15912 -1345
rect 15942 -1475 15996 -1345
rect 16026 -1475 16080 -1345
rect 16110 -1475 16164 -1345
rect 16194 -1475 16248 -1345
rect 16278 -1475 16332 -1345
rect 16362 -1475 16416 -1345
rect 16446 -1475 16500 -1345
rect 16530 -1475 16584 -1345
rect 16614 -1475 16666 -1345
rect 2340 -10090 2460 -9890
<< nwell >>
rect 8560 -1270 16750 -540
<< pwell >>
rect 8560 -1510 16750 -1310
<< nsubdiffcont >>
rect 8790 -800 8900 -690
<< locali >>
rect 8780 -1310 8980 -1250
rect 9270 -1310 9430 -1250
<< viali >>
rect 10650 -1140 10690 -1100
rect 10650 -1210 10690 -1170
rect 10650 -1310 10690 -1270
rect 10650 -1400 10690 -1360
<< metal1 >>
rect 480 -610 920 -600
rect 480 -790 690 -610
rect 910 -790 920 -610
rect 480 -800 920 -790
rect 480 -940 920 -930
rect -4260 -1260 -4060 -1060
rect -3710 -1210 -3510 -1010
rect -3130 -1150 -2930 -950
rect -2670 -1190 -2470 -990
rect 480 -1120 690 -940
rect 910 -1120 920 -940
rect 8600 -1030 16710 -920
rect 480 -1130 920 -1120
rect 10630 -1100 10710 -1090
rect 10630 -1140 10650 -1100
rect 10690 -1140 10710 -1100
rect 10630 -1170 10710 -1140
rect 10630 -1210 10650 -1170
rect 10690 -1210 10710 -1170
rect 10630 -1270 10710 -1210
rect 10630 -1310 10650 -1270
rect 10690 -1310 10710 -1270
rect 10630 -1360 10710 -1310
rect 10630 -1400 10650 -1360
rect 10690 -1400 10710 -1360
rect 480 -1430 920 -1420
rect 10630 -1430 10710 -1400
rect 480 -1610 690 -1430
rect 910 -1610 920 -1430
rect 8600 -1580 16710 -1470
rect 480 -1620 920 -1610
rect 480 -1710 920 -1700
rect 480 -1890 690 -1710
rect 910 -1890 920 -1710
rect 480 -1900 920 -1890
rect 480 -2170 920 -2160
rect 480 -2350 690 -2170
rect 910 -2350 920 -2170
rect 480 -2360 920 -2350
rect 480 -2530 920 -2520
rect 480 -2710 690 -2530
rect 910 -2710 920 -2530
rect 480 -2720 920 -2710
rect 480 -2930 920 -2920
rect 480 -3110 690 -2930
rect 910 -3110 920 -2930
rect 480 -3120 920 -3110
rect 480 -3380 920 -3370
rect 480 -3560 690 -3380
rect 910 -3560 920 -3380
rect 480 -3570 920 -3560
rect 480 -3750 920 -3740
rect 480 -3930 690 -3750
rect 910 -3930 920 -3750
rect 480 -3940 920 -3930
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8950 920 -8770
rect 680 -8960 920 -8950
rect 470 -9100 920 -9090
rect 470 -9280 690 -9100
rect 910 -9280 920 -9100
rect 470 -9290 920 -9280
rect 470 -9590 920 -9580
rect 470 -9770 690 -9590
rect 910 -9770 920 -9590
rect 470 -9780 920 -9770
rect 470 -9870 920 -9860
rect 470 -10050 690 -9870
rect 910 -10050 920 -9870
rect 470 -10060 920 -10050
rect 470 -10330 920 -10320
rect 470 -10510 690 -10330
rect 910 -10510 920 -10330
rect 470 -10520 920 -10510
rect 470 -10690 920 -10680
rect 470 -10870 690 -10690
rect 910 -10870 920 -10690
rect 470 -10880 920 -10870
rect 470 -11090 920 -11080
rect 470 -11270 690 -11090
rect 910 -11270 920 -11090
rect 470 -11280 920 -11270
rect 470 -11540 920 -11530
rect 470 -11720 690 -11540
rect 910 -11720 920 -11540
rect 470 -11730 920 -11720
rect 480 -11910 920 -11900
rect 480 -12090 690 -11910
rect 910 -12090 920 -11910
rect 480 -12100 920 -12090
<< via1 >>
rect 690 -790 910 -610
rect 690 -1120 910 -940
rect 690 -1610 910 -1430
rect 690 -1890 910 -1710
rect 690 -2350 910 -2170
rect 690 -2710 910 -2530
rect 690 -3110 910 -2930
rect 690 -3560 910 -3380
rect 690 -3930 910 -3750
rect 690 -8950 910 -8770
rect 690 -9280 910 -9100
rect 690 -9770 910 -9590
rect 690 -10050 910 -9870
rect 690 -10510 910 -10330
rect 690 -10870 910 -10690
rect 690 -11270 910 -11090
rect 690 -11720 910 -11540
rect 690 -12090 910 -11910
<< metal2 >>
rect 680 -610 920 -600
rect 680 -790 690 -610
rect 910 -790 920 -610
rect 680 -800 920 -790
rect 680 -940 920 -930
rect 680 -1120 690 -940
rect 910 -1120 920 -940
rect 680 -1130 920 -1120
rect 680 -1430 920 -1420
rect 680 -1610 690 -1430
rect 910 -1610 920 -1430
rect 680 -1620 920 -1610
rect 680 -1710 920 -1700
rect 680 -1890 690 -1710
rect 910 -1890 920 -1710
rect 680 -1900 920 -1890
rect 680 -2170 920 -2160
rect 680 -2350 690 -2170
rect 910 -2350 920 -2170
rect 680 -2360 920 -2350
rect 680 -2530 920 -2520
rect 680 -2710 690 -2530
rect 910 -2710 920 -2530
rect 680 -2720 920 -2710
rect 680 -2930 920 -2920
rect 680 -3110 690 -2930
rect 910 -3110 920 -2930
rect 680 -3120 920 -3110
rect 680 -3380 920 -3370
rect 680 -3560 690 -3380
rect 910 -3560 920 -3380
rect 680 -3570 920 -3560
rect 680 -3750 920 -3740
rect 680 -3930 690 -3750
rect 910 -3930 920 -3750
rect 680 -3940 920 -3930
rect 1080 -3770 1220 -1150
rect 1080 -3910 1090 -3770
rect 1210 -3910 1220 -3770
rect 1080 -3940 1220 -3910
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8950 920 -8770
rect 680 -8960 920 -8950
rect 680 -9100 920 -9090
rect 680 -9280 690 -9100
rect 910 -9280 920 -9100
rect 680 -9290 920 -9280
rect 680 -9590 920 -9580
rect 680 -9770 690 -9590
rect 910 -9770 920 -9590
rect 680 -9780 920 -9770
rect 680 -9870 920 -9860
rect 680 -10050 690 -9870
rect 910 -10050 920 -9870
rect 680 -10060 920 -10050
rect 680 -10330 920 -10320
rect 680 -10510 690 -10330
rect 910 -10510 920 -10330
rect 680 -10520 920 -10510
rect 680 -10690 920 -10680
rect 680 -10870 690 -10690
rect 910 -10870 920 -10690
rect 680 -10880 920 -10870
rect 680 -11090 920 -11080
rect 680 -11270 690 -11090
rect 910 -11270 920 -11090
rect 680 -11280 920 -11270
rect 680 -11540 920 -11530
rect 680 -11720 690 -11540
rect 910 -11720 920 -11540
rect 680 -11730 920 -11720
rect 680 -11910 920 -11900
rect 680 -12090 690 -11910
rect 910 -12090 920 -11910
rect 680 -12100 920 -12090
rect 1080 -11930 1220 -9310
rect 1080 -12070 1090 -11930
rect 1210 -12070 1220 -11930
rect 1080 -12100 1220 -12070
<< via2 >>
rect 690 -790 910 -610
rect 3090 -890 3210 -790
rect 690 -1120 910 -940
rect 2840 -1090 2960 -970
rect 690 -1610 910 -1430
rect 690 -1890 910 -1710
rect 690 -2350 910 -2170
rect 690 -2710 910 -2530
rect 690 -3110 910 -2930
rect 690 -3560 910 -3380
rect 690 -3930 910 -3750
rect 2590 -1590 2710 -1450
rect 2340 -1870 2460 -1730
rect 1840 -2690 1960 -2550
rect 1590 -3090 1710 -2960
rect 1340 -3540 1460 -3400
rect 1090 -3910 1210 -3770
rect 690 -8950 910 -8770
rect 3090 -9050 3210 -8950
rect 690 -9280 910 -9100
rect 2840 -9250 2960 -9130
rect 690 -9770 910 -9590
rect 690 -10050 910 -9870
rect 690 -10510 910 -10330
rect 690 -10870 910 -10690
rect 690 -11270 910 -11090
rect 690 -11720 910 -11540
rect 690 -12090 910 -11910
rect 2590 -9750 2710 -9610
rect 2340 -10030 2460 -9890
rect 1840 -10850 1960 -10710
rect 1590 -11250 1710 -11110
rect 1340 -11700 1460 -11560
rect 1090 -12070 1210 -11930
<< metal3 >>
rect 680 -610 920 -600
rect 680 -790 690 -610
rect 910 -620 920 -610
rect 910 -780 1240 -620
rect 910 -790 920 -780
rect 680 -800 920 -790
rect 1080 -790 3220 -780
rect 1080 -890 3090 -790
rect 3210 -890 3220 -790
rect 1080 -900 3220 -890
rect 680 -940 920 -930
rect 680 -1120 690 -940
rect 910 -960 920 -940
rect 910 -970 2970 -960
rect 910 -1090 2840 -970
rect 2960 -1090 2970 -970
rect 910 -1100 2970 -1090
rect 910 -1120 920 -1100
rect 680 -1130 920 -1120
rect 680 -1430 920 -1420
rect 680 -1610 690 -1430
rect 910 -1440 920 -1430
rect 910 -1450 2720 -1440
rect 910 -1590 2590 -1450
rect 2710 -1590 2720 -1450
rect 910 -1600 2720 -1590
rect 910 -1610 920 -1600
rect 680 -1620 920 -1610
rect 680 -1710 920 -1700
rect 680 -1890 690 -1710
rect 910 -1720 920 -1710
rect 910 -1730 2470 -1720
rect 910 -1870 2340 -1730
rect 2460 -1870 2470 -1730
rect 910 -1880 2470 -1870
rect 910 -1890 920 -1880
rect 680 -1900 920 -1890
rect 680 -2170 920 -2160
rect 680 -2350 690 -2170
rect 910 -2180 920 -2170
rect 910 -2340 2220 -2180
rect 910 -2350 920 -2340
rect 680 -2360 920 -2350
rect 680 -2530 920 -2520
rect 680 -2710 690 -2530
rect 910 -2540 920 -2530
rect 910 -2550 1970 -2540
rect 910 -2690 1840 -2550
rect 1960 -2690 1970 -2550
rect 910 -2700 1970 -2690
rect 910 -2710 920 -2700
rect 680 -2720 920 -2710
rect 680 -2930 920 -2920
rect 680 -3110 690 -2930
rect 910 -2950 920 -2930
rect 910 -2960 1720 -2950
rect 910 -3090 1590 -2960
rect 1710 -3090 1720 -2960
rect 910 -3100 1720 -3090
rect 910 -3110 920 -3100
rect 680 -3120 920 -3110
rect 680 -3380 920 -3370
rect 680 -3560 690 -3380
rect 910 -3390 920 -3380
rect 910 -3400 1470 -3390
rect 910 -3540 1340 -3400
rect 1460 -3540 1470 -3400
rect 910 -3550 1470 -3540
rect 910 -3560 920 -3550
rect 680 -3570 920 -3560
rect 680 -3750 920 -3740
rect 680 -3930 690 -3750
rect 910 -3760 920 -3750
rect 910 -3770 1220 -3760
rect 910 -3910 1090 -3770
rect 1210 -3910 1220 -3770
rect 910 -3920 1220 -3910
rect 910 -3930 920 -3920
rect 680 -3940 920 -3930
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8780 920 -8770
rect 910 -8940 1240 -8780
rect 910 -8950 920 -8940
rect 680 -8960 920 -8950
rect 1080 -8950 3220 -8940
rect 1080 -9050 3090 -8950
rect 3210 -9050 3220 -8950
rect 1080 -9060 3220 -9050
rect 680 -9100 920 -9090
rect 680 -9280 690 -9100
rect 910 -9120 920 -9100
rect 910 -9130 2970 -9120
rect 910 -9250 2840 -9130
rect 2960 -9250 2970 -9130
rect 910 -9260 2970 -9250
rect 910 -9280 920 -9260
rect 680 -9290 920 -9280
rect 680 -9590 920 -9580
rect 680 -9770 690 -9590
rect 910 -9600 920 -9590
rect 910 -9610 2720 -9600
rect 910 -9750 2590 -9610
rect 2710 -9750 2720 -9610
rect 910 -9760 2720 -9750
rect 910 -9770 920 -9760
rect 680 -9780 920 -9770
rect 680 -9870 920 -9860
rect 680 -10050 690 -9870
rect 910 -9880 920 -9870
rect 910 -9890 2470 -9880
rect 910 -10030 2340 -9890
rect 2460 -10030 2470 -9890
rect 910 -10040 2470 -10030
rect 910 -10050 920 -10040
rect 680 -10060 920 -10050
rect 680 -10330 920 -10320
rect 680 -10510 690 -10330
rect 910 -10340 920 -10330
rect 910 -10500 2220 -10340
rect 910 -10510 920 -10500
rect 680 -10520 920 -10510
rect 680 -10690 920 -10680
rect 680 -10870 690 -10690
rect 910 -10700 920 -10690
rect 910 -10710 1970 -10700
rect 910 -10850 1840 -10710
rect 1960 -10850 1970 -10710
rect 910 -10860 1970 -10850
rect 910 -10870 920 -10860
rect 680 -10880 920 -10870
rect 680 -11090 920 -11080
rect 680 -11270 690 -11090
rect 910 -11100 920 -11090
rect 910 -11110 1720 -11100
rect 910 -11250 1590 -11110
rect 1710 -11250 1720 -11110
rect 910 -11260 1720 -11250
rect 910 -11270 920 -11260
rect 680 -11280 920 -11270
rect 680 -11540 920 -11530
rect 680 -11720 690 -11540
rect 910 -11550 920 -11540
rect 910 -11560 1470 -11550
rect 910 -11700 1340 -11560
rect 1460 -11700 1470 -11560
rect 910 -11710 1470 -11700
rect 910 -11720 920 -11710
rect 680 -11730 920 -11720
rect 680 -11910 920 -11900
rect 680 -12090 690 -11910
rect 910 -11920 920 -11910
rect 910 -11930 1220 -11920
rect 910 -12070 1090 -11930
rect 1210 -12070 1220 -11930
rect 910 -12080 1220 -12070
rect 910 -12090 920 -12080
rect 680 -12100 920 -12090
<< metal4 >>
rect 4140 -500 8390 300
rect 4140 -15670 4950 -500
rect 7640 -15750 8390 -500
<< metal5 >>
rect 5330 -15300 17310 10
use sky130_fd_sc_hd__or2_1  x1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8460 0 1 4218
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  x2
timestamp 1701704242
transform 1 0 8958 0 1 4170
box -38 -48 498 592
use 8to3_Priority_Encoder_v0p2p0  x3
timestamp 1713021466
transform 1 0 4960 0 1 -8740
box -3910 -7130 3570 700
use sky130_fd_sc_hd__inv_16  x4 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12288 0 1 -1522
box -38 -48 1510 592
use 8to3_Priority_Encoder_v0p2p0  x5
timestamp 1713021466
transform 1 0 4960 0 1 -700
box -3910 -7130 3570 700
use sky130_fd_sc_hd__inv_16  x6
timestamp 1701704242
transform 1 0 10816 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8146 0 1 4266
box -38 -48 314 592
use sky130_fd_sc_hd__inv_16  x8
timestamp 1701704242
transform 1 0 13760 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x9
timestamp 1701704242
transform 1 0 15232 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x10
timestamp 1701704242
transform 1 0 16786 0 1 3930
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  x11
timestamp 1701704242
transform 1 0 -1640 0 1 4890
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x12
timestamp 1701704242
transform 1 0 18296 0 1 3882
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x13
timestamp 1701704242
transform 1 0 20836 0 1 3954
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x14
timestamp 1701704242
transform 1 0 22346 0 1 3906
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x15
timestamp 1701704242
transform 1 0 23856 0 1 3858
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x16
timestamp 1701704242
transform 1 0 25366 0 1 3810
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x17
timestamp 1701704242
transform 1 0 26876 0 1 3762
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x18
timestamp 1701704242
transform 1 0 28386 0 1 3714
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x19
timestamp 1701704242
transform 1 0 29896 0 1 3666
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x20
timestamp 1701704242
transform 1 0 -1142 0 1 4842
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x21 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 -828 0 1 4794
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x22
timestamp 1701704242
transform 1 0 -330 0 1 4746
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x23
timestamp 1701704242
transform 1 0 31406 0 1 3618
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x24
timestamp 1701704242
transform 1 0 32916 0 1 3570
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x25
timestamp 1701704242
transform 1 0 34426 0 1 3522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x27
timestamp 1701704242
transform 1 0 1180 0 1 4698
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x28
timestamp 1701704242
transform 1 0 1494 0 1 4650
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x29
timestamp 1701704242
transform 1 0 1992 0 1 4602
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x34
timestamp 1701704242
transform 1 0 3502 0 1 4554
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x35
timestamp 1701704242
transform 1 0 3816 0 1 4506
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x36
timestamp 1701704242
transform 1 0 4314 0 1 4458
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x41
timestamp 1701704242
transform 1 0 8608 0 1 -1522
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x42
timestamp 1701704242
transform 1 0 8884 0 1 -1522
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x43
timestamp 1701704242
transform 1 0 9344 0 1 -1522
box -38 -48 1510 592
<< labels >>
flabel metal1 480 -1130 680 -930 0 FreeSans 256 0 0 0 I15
port 2 nsew
flabel metal1 480 -800 680 -600 0 FreeSans 256 0 0 0 EI
port 1 nsew
flabel metal1 480 -1620 680 -1420 0 FreeSans 256 0 0 0 I14
port 3 nsew
flabel metal1 480 -1900 680 -1700 0 FreeSans 256 0 0 0 I13
port 4 nsew
flabel metal1 480 -2360 680 -2160 0 FreeSans 256 0 0 0 I12
port 5 nsew
flabel metal1 480 -2720 680 -2520 0 FreeSans 256 0 0 0 I11
port 6 nsew
flabel metal1 480 -3120 680 -2920 0 FreeSans 256 0 0 0 I10
port 7 nsew
flabel metal1 480 -3570 680 -3370 0 FreeSans 256 0 0 0 I9
port 9 nsew
flabel metal1 480 -3940 680 -3740 0 FreeSans 256 0 0 0 I8
port 10 nsew
flabel metal1 480 -12100 680 -11900 0 FreeSans 256 0 0 0 I0
port 19 nsew
flabel metal1 470 -11730 670 -11530 0 FreeSans 256 0 0 0 I1
port 18 nsew
flabel metal1 470 -11280 670 -11080 0 FreeSans 256 0 0 0 I2
port 17 nsew
flabel metal1 470 -10880 670 -10680 0 FreeSans 256 0 0 0 I3
port 16 nsew
flabel metal1 470 -10520 670 -10320 0 FreeSans 256 0 0 0 I4
port 14 nsew
flabel metal1 470 -10060 670 -9860 0 FreeSans 256 0 0 0 I5
port 13 nsew
flabel metal1 470 -9780 670 -9580 0 FreeSans 256 0 0 0 I6
port 12 nsew
flabel metal1 470 -9290 670 -9090 0 FreeSans 256 0 0 0 I7
port 11 nsew
flabel metal1 -4260 -1260 -4060 -1060 0 FreeSans 256 0 0 0 A3
port 0 nsew
flabel metal1 -3710 -1210 -3510 -1010 0 FreeSans 256 0 0 0 A2
port 8 nsew
flabel metal1 -3130 -1150 -2930 -950 0 FreeSans 256 0 0 0 A1
port 15 nsew
flabel metal1 -2670 -1190 -2470 -990 0 FreeSans 256 0 0 0 A0
port 20 nsew
<< end >>
